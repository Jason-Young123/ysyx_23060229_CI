//Generate the verilog at 2025-09-29T17:20:45 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_B ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ;
wire \myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__A_B ;
wire \mylsu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[6]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

AND3_X4 _08922_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01414_ ) );
AND3_X4 _08923_ ( .A1(_01414_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01415_ ) );
AND3_X4 _08924_ ( .A1(_01415_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01416_ ) );
AND3_X4 _08925_ ( .A1(_01416_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01417_ ) );
AND3_X4 _08926_ ( .A1(_01417_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01418_ ) );
AND3_X4 _08927_ ( .A1(_01418_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01419_ ) );
AND3_X4 _08928_ ( .A1(_01419_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01420_ ) );
AND3_X4 _08929_ ( .A1(_01420_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01421_ ) );
AND3_X4 _08930_ ( .A1(_01421_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01422_ ) );
AND3_X4 _08931_ ( .A1(_01422_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01423_ ) );
AND3_X4 _08932_ ( .A1(_01423_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01424_ ) );
AND3_X4 _08933_ ( .A1(_01424_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01425_ ) );
AND3_X4 _08934_ ( .A1(_01425_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01426_ ) );
AND2_X2 _08935_ ( .A1(_01426_ ), .A2(\myclint.mtime [27] ), .ZN(_01427_ ) );
AND2_X1 _08936_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01428_ ) );
AND2_X2 _08937_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01429_ ) );
AND4_X4 _08938_ ( .A1(\myclint.mtime [33] ), .A2(_01427_ ), .A3(_01428_ ), .A4(_01429_ ), .ZN(_01430_ ) );
AND3_X2 _08939_ ( .A1(_01430_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01431_ ) );
AND3_X4 _08940_ ( .A1(_01431_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [35] ), .ZN(_01432_ ) );
AND3_X2 _08941_ ( .A1(_01432_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [37] ), .ZN(_01433_ ) );
AND2_X2 _08942_ ( .A1(_01433_ ), .A2(\myclint.mtime [39] ), .ZN(_01434_ ) );
AND2_X1 _08943_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01435_ ) );
AND2_X2 _08944_ ( .A1(_01434_ ), .A2(_01435_ ), .ZN(_01436_ ) );
AND2_X1 _08945_ ( .A1(\myclint.mtime [42] ), .A2(\myclint.mtime [43] ), .ZN(_01437_ ) );
AND2_X4 _08946_ ( .A1(_01436_ ), .A2(_01437_ ), .ZN(_01438_ ) );
AND2_X1 _08947_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01439_ ) );
AND3_X1 _08948_ ( .A1(_01439_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01440_ ) );
AND2_X1 _08949_ ( .A1(_01438_ ), .A2(_01440_ ), .ZN(_01441_ ) );
AND2_X1 _08950_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01442_ ) );
AND2_X1 _08951_ ( .A1(_01441_ ), .A2(_01442_ ), .ZN(_01443_ ) );
AND2_X1 _08952_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01444_ ) );
AND2_X1 _08953_ ( .A1(_01443_ ), .A2(_01444_ ), .ZN(_01445_ ) );
AND2_X1 _08954_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01446_ ) );
AND2_X1 _08955_ ( .A1(_01445_ ), .A2(_01446_ ), .ZN(_01447_ ) );
AND2_X1 _08956_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01448_ ) );
AND2_X1 _08957_ ( .A1(_01447_ ), .A2(_01448_ ), .ZN(_01449_ ) );
AND2_X1 _08958_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01450_ ) );
AND2_X1 _08959_ ( .A1(_01449_ ), .A2(_01450_ ), .ZN(_01451_ ) );
AND2_X1 _08960_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01452_ ) );
AND2_X2 _08961_ ( .A1(_01451_ ), .A2(_01452_ ), .ZN(_01453_ ) );
INV_X1 _08962_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01454_ ) );
AND2_X1 _08963_ ( .A1(\myclint.mtime [60] ), .A2(\myclint.mtime [61] ), .ZN(_01455_ ) );
AND3_X2 _08964_ ( .A1(_01453_ ), .A2(_01454_ ), .A3(_01455_ ), .ZN(_01456_ ) );
AND2_X1 _08965_ ( .A1(_01456_ ), .A2(\myclint.mtime [63] ), .ZN(_01457_ ) );
INV_X1 _08966_ ( .A(fanout_net_1 ), .ZN(_01458_ ) );
BUF_X4 _08967_ ( .A(_01458_ ), .Z(_01459_ ) );
BUF_X4 _08968_ ( .A(_01459_ ), .Z(_01460_ ) );
OAI21_X1 _08969_ ( .A(_01460_ ), .B1(_01456_ ), .B2(\myclint.mtime [63] ), .ZN(_01461_ ) );
NOR2_X1 _08970_ ( .A1(_01457_ ), .A2(_01461_ ), .ZN(_00000_ ) );
AND2_X1 _08971_ ( .A1(_01414_ ), .A2(\myclint.mtime [3] ), .ZN(_01462_ ) );
AND4_X1 _08972_ ( .A1(\myclint.mtime [6] ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [5] ), .A4(\myclint.mtime [7] ), .ZN(_01463_ ) );
AND2_X1 _08973_ ( .A1(_01462_ ), .A2(_01463_ ), .ZN(_01464_ ) );
AND4_X1 _08974_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01465_ ) );
AND2_X1 _08975_ ( .A1(\myclint.mtime [8] ), .A2(\myclint.mtime [9] ), .ZN(_01466_ ) );
AND4_X1 _08976_ ( .A1(\myclint.mtime [10] ), .A2(_01465_ ), .A3(\myclint.mtime [11] ), .A4(_01466_ ), .ZN(_01467_ ) );
AND2_X1 _08977_ ( .A1(_01464_ ), .A2(_01467_ ), .ZN(_01468_ ) );
AND2_X1 _08978_ ( .A1(\myclint.mtime [16] ), .A2(\myclint.mtime [17] ), .ZN(_01469_ ) );
NAND3_X1 _08979_ ( .A1(_01469_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [19] ), .ZN(_01470_ ) );
NAND4_X1 _08980_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01471_ ) );
NOR2_X1 _08981_ ( .A1(_01470_ ), .A2(_01471_ ), .ZN(_01472_ ) );
AND2_X1 _08982_ ( .A1(\myclint.mtime [24] ), .A2(\myclint.mtime [25] ), .ZN(_01473_ ) );
AND3_X1 _08983_ ( .A1(_01473_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [27] ), .ZN(_01474_ ) );
AND4_X1 _08984_ ( .A1(_01428_ ), .A2(_01472_ ), .A3(_01429_ ), .A4(_01474_ ), .ZN(_01475_ ) );
NAND2_X1 _08985_ ( .A1(_01468_ ), .A2(_01475_ ), .ZN(_01476_ ) );
AND2_X1 _08986_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01477_ ) );
NAND3_X1 _08987_ ( .A1(_01477_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01478_ ) );
NAND4_X1 _08988_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01479_ ) );
NOR2_X1 _08989_ ( .A1(_01478_ ), .A2(_01479_ ), .ZN(_01480_ ) );
AND2_X1 _08990_ ( .A1(_01437_ ), .A2(_01435_ ), .ZN(_01481_ ) );
AND3_X1 _08991_ ( .A1(_01480_ ), .A2(_01440_ ), .A3(_01481_ ), .ZN(_01482_ ) );
INV_X1 _08992_ ( .A(_01482_ ), .ZN(_01483_ ) );
NOR2_X1 _08993_ ( .A1(_01476_ ), .A2(_01483_ ), .ZN(_01484_ ) );
AND4_X1 _08994_ ( .A1(_01448_ ), .A2(_01446_ ), .A3(_01444_ ), .A4(_01442_ ), .ZN(_01485_ ) );
AND2_X1 _08995_ ( .A1(_01484_ ), .A2(_01485_ ), .ZN(_01486_ ) );
AND4_X1 _08996_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01487_ ) );
NAND3_X1 _08997_ ( .A1(_01486_ ), .A2(_01455_ ), .A3(_01487_ ), .ZN(_01488_ ) );
OR2_X1 _08998_ ( .A1(_01488_ ), .A2(\myclint.mtime [62] ), .ZN(_01489_ ) );
NAND2_X1 _08999_ ( .A1(_01488_ ), .A2(\myclint.mtime [62] ), .ZN(_01490_ ) );
AOI21_X1 _09000_ ( .A(fanout_net_1 ), .B1(_01489_ ), .B2(_01490_ ), .ZN(_00001_ ) );
AND2_X1 _09001_ ( .A1(_01444_ ), .A2(_01442_ ), .ZN(_01491_ ) );
NAND2_X1 _09002_ ( .A1(_01484_ ), .A2(_01491_ ), .ZN(_01492_ ) );
OR3_X1 _09003_ ( .A1(_01492_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [53] ), .ZN(_01493_ ) );
OAI21_X1 _09004_ ( .A(\myclint.mtime [53] ), .B1(_01492_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01494_ ) );
AOI21_X1 _09005_ ( .A(fanout_net_1 ), .B1(_01493_ ), .B2(_01494_ ), .ZN(_00002_ ) );
OR2_X1 _09006_ ( .A1(_01492_ ), .A2(\myclint.mtime [52] ), .ZN(_01495_ ) );
NAND2_X1 _09007_ ( .A1(_01492_ ), .A2(\myclint.mtime [52] ), .ZN(_01496_ ) );
AOI21_X1 _09008_ ( .A(fanout_net_1 ), .B1(_01495_ ), .B2(_01496_ ), .ZN(_00003_ ) );
INV_X1 _09009_ ( .A(_01476_ ), .ZN(_01497_ ) );
NAND3_X1 _09010_ ( .A1(_01497_ ), .A2(_01442_ ), .A3(_01482_ ), .ZN(_01498_ ) );
OR3_X1 _09011_ ( .A1(_01498_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [51] ), .ZN(_01499_ ) );
OAI21_X1 _09012_ ( .A(\myclint.mtime [51] ), .B1(_01498_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01500_ ) );
AOI21_X1 _09013_ ( .A(fanout_net_1 ), .B1(_01499_ ), .B2(_01500_ ), .ZN(_00004_ ) );
OR2_X1 _09014_ ( .A1(_01498_ ), .A2(\myclint.mtime [50] ), .ZN(_01501_ ) );
NAND2_X1 _09015_ ( .A1(_01498_ ), .A2(\myclint.mtime [50] ), .ZN(_01502_ ) );
AOI21_X1 _09016_ ( .A(fanout_net_1 ), .B1(_01501_ ), .B2(_01502_ ), .ZN(_00005_ ) );
INV_X1 _09017_ ( .A(_01438_ ), .ZN(_01503_ ) );
INV_X1 _09018_ ( .A(_01440_ ), .ZN(_01504_ ) );
NOR3_X1 _09019_ ( .A1(_01503_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01504_ ), .ZN(_01505_ ) );
AND2_X1 _09020_ ( .A1(_01505_ ), .A2(\myclint.mtime [49] ), .ZN(_01506_ ) );
OAI21_X1 _09021_ ( .A(_01460_ ), .B1(_01505_ ), .B2(\myclint.mtime [49] ), .ZN(_01507_ ) );
NOR2_X1 _09022_ ( .A1(_01506_ ), .A2(_01507_ ), .ZN(_00006_ ) );
NAND2_X1 _09023_ ( .A1(_01464_ ), .A2(_01467_ ), .ZN(_01508_ ) );
NAND4_X1 _09024_ ( .A1(_01472_ ), .A2(_01428_ ), .A3(_01429_ ), .A4(_01474_ ), .ZN(_01509_ ) );
OR4_X1 _09025_ ( .A1(\myclint.mtime [48] ), .A2(_01483_ ), .A3(_01508_ ), .A4(_01509_ ), .ZN(_01510_ ) );
OAI21_X1 _09026_ ( .A(\myclint.mtime [48] ), .B1(_01476_ ), .B2(_01483_ ), .ZN(_01511_ ) );
AOI21_X1 _09027_ ( .A(fanout_net_1 ), .B1(_01510_ ), .B2(_01511_ ), .ZN(_00007_ ) );
NAND3_X1 _09028_ ( .A1(_01436_ ), .A2(\myclint.mtime [44] ), .A3(_01437_ ), .ZN(_01512_ ) );
INV_X1 _09029_ ( .A(\myclint.mtime [45] ), .ZN(_01513_ ) );
NOR3_X1 _09030_ ( .A1(_01512_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01513_ ), .ZN(_01514_ ) );
AND2_X1 _09031_ ( .A1(_01514_ ), .A2(\myclint.mtime [47] ), .ZN(_01515_ ) );
BUF_X4 _09032_ ( .A(_01459_ ), .Z(_01516_ ) );
NAND3_X1 _09033_ ( .A1(_01436_ ), .A2(_01439_ ), .A3(_01437_ ), .ZN(_01517_ ) );
NOR2_X1 _09034_ ( .A1(_01517_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01518_ ) );
OAI21_X1 _09035_ ( .A(_01516_ ), .B1(_01518_ ), .B2(\myclint.mtime [47] ), .ZN(_01519_ ) );
NOR2_X1 _09036_ ( .A1(_01515_ ), .A2(_01519_ ), .ZN(_00008_ ) );
AND2_X1 _09037_ ( .A1(_01497_ ), .A2(_01480_ ), .ZN(_01520_ ) );
AND3_X1 _09038_ ( .A1(_01520_ ), .A2(_01439_ ), .A3(_01481_ ), .ZN(_01521_ ) );
XNOR2_X1 _09039_ ( .A(_01521_ ), .B(\myclint.mtime [46] ), .ZN(_01522_ ) );
NOR2_X1 _09040_ ( .A1(_01522_ ), .A2(fanout_net_1 ), .ZN(_00009_ ) );
INV_X1 _09041_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01523_ ) );
AND3_X1 _09042_ ( .A1(_01436_ ), .A2(_01523_ ), .A3(_01437_ ), .ZN(_01524_ ) );
AND2_X1 _09043_ ( .A1(_01524_ ), .A2(\myclint.mtime [45] ), .ZN(_01525_ ) );
OAI21_X1 _09044_ ( .A(_01516_ ), .B1(_01524_ ), .B2(\myclint.mtime [45] ), .ZN(_01526_ ) );
NOR2_X1 _09045_ ( .A1(_01525_ ), .A2(_01526_ ), .ZN(_00010_ ) );
AND2_X1 _09046_ ( .A1(_01520_ ), .A2(_01481_ ), .ZN(_01527_ ) );
XNOR2_X1 _09047_ ( .A(_01527_ ), .B(\myclint.mtime [44] ), .ZN(_01528_ ) );
NOR2_X1 _09048_ ( .A1(_01528_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
AND2_X1 _09049_ ( .A1(_01486_ ), .A2(_01487_ ), .ZN(_01529_ ) );
INV_X1 _09050_ ( .A(_01529_ ), .ZN(_01530_ ) );
OR3_X1 _09051_ ( .A1(_01530_ ), .A2(\myclint.mtime [61] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01531_ ) );
OAI21_X1 _09052_ ( .A(\myclint.mtime [61] ), .B1(_01530_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01532_ ) );
AOI21_X1 _09053_ ( .A(fanout_net_1 ), .B1(_01531_ ), .B2(_01532_ ), .ZN(_00012_ ) );
NAND3_X1 _09054_ ( .A1(_01497_ ), .A2(_01435_ ), .A3(_01480_ ), .ZN(_01533_ ) );
OR3_X1 _09055_ ( .A1(_01533_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [43] ), .ZN(_01534_ ) );
OAI21_X1 _09056_ ( .A(\myclint.mtime [43] ), .B1(_01533_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01535_ ) );
AOI21_X1 _09057_ ( .A(fanout_net_1 ), .B1(_01534_ ), .B2(_01535_ ), .ZN(_00013_ ) );
OR2_X1 _09058_ ( .A1(_01533_ ), .A2(\myclint.mtime [42] ), .ZN(_01536_ ) );
NAND2_X1 _09059_ ( .A1(_01533_ ), .A2(\myclint.mtime [42] ), .ZN(_01537_ ) );
AOI21_X1 _09060_ ( .A(fanout_net_1 ), .B1(_01536_ ), .B2(_01537_ ), .ZN(_00014_ ) );
INV_X1 _09061_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01538_ ) );
AND3_X1 _09062_ ( .A1(_01433_ ), .A2(_01538_ ), .A3(\myclint.mtime [39] ), .ZN(_01539_ ) );
AND2_X1 _09063_ ( .A1(_01539_ ), .A2(\myclint.mtime [41] ), .ZN(_01540_ ) );
OAI21_X1 _09064_ ( .A(_01516_ ), .B1(_01539_ ), .B2(\myclint.mtime [41] ), .ZN(_01541_ ) );
NOR2_X1 _09065_ ( .A1(_01540_ ), .A2(_01541_ ), .ZN(_00015_ ) );
INV_X1 _09066_ ( .A(_01520_ ), .ZN(_01542_ ) );
NAND2_X1 _09067_ ( .A1(_01542_ ), .A2(\myclint.mtime [40] ), .ZN(_01543_ ) );
OR4_X1 _09068_ ( .A1(\myclint.mtime [40] ), .A2(_01476_ ), .A3(_01479_ ), .A4(_01478_ ), .ZN(_01544_ ) );
AOI21_X1 _09069_ ( .A(fanout_net_1 ), .B1(_01543_ ), .B2(_01544_ ), .ZN(_00016_ ) );
BUF_X2 _09070_ ( .A(_01459_ ), .Z(_01545_ ) );
INV_X1 _09071_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01546_ ) );
AND3_X1 _09072_ ( .A1(_01432_ ), .A2(_01546_ ), .A3(\myclint.mtime [37] ), .ZN(_01547_ ) );
OAI21_X1 _09073_ ( .A(_01545_ ), .B1(_01547_ ), .B2(\myclint.mtime [39] ), .ZN(_01548_ ) );
NAND4_X1 _09074_ ( .A1(_01427_ ), .A2(\myclint.mtime [33] ), .A3(_01428_ ), .A4(_01429_ ), .ZN(_01549_ ) );
INV_X1 _09075_ ( .A(\myclint.mtime [32] ), .ZN(_01550_ ) );
NOR2_X1 _09076_ ( .A1(_01549_ ), .A2(_01550_ ), .ZN(_01551_ ) );
AND3_X1 _09077_ ( .A1(_01551_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01552_ ) );
AND3_X1 _09078_ ( .A1(_01552_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .ZN(_01553_ ) );
AND3_X1 _09079_ ( .A1(_01553_ ), .A2(_01546_ ), .A3(\myclint.mtime [39] ), .ZN(_01554_ ) );
NOR2_X1 _09080_ ( .A1(_01548_ ), .A2(_01554_ ), .ZN(_00017_ ) );
BUF_X4 _09081_ ( .A(_01459_ ), .Z(_01555_ ) );
OAI21_X1 _09082_ ( .A(_01555_ ), .B1(_01553_ ), .B2(\myclint.mtime [38] ), .ZN(_01556_ ) );
NOR2_X1 _09083_ ( .A1(_01556_ ), .A2(_01433_ ), .ZN(_00018_ ) );
INV_X1 _09084_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01557_ ) );
AND3_X1 _09085_ ( .A1(_01431_ ), .A2(_01557_ ), .A3(\myclint.mtime [35] ), .ZN(_01558_ ) );
OAI21_X1 _09086_ ( .A(_01555_ ), .B1(_01558_ ), .B2(\myclint.mtime [37] ), .ZN(_01559_ ) );
AND3_X1 _09087_ ( .A1(_01552_ ), .A2(\myclint.mtime [37] ), .A3(_01557_ ), .ZN(_01560_ ) );
NOR2_X1 _09088_ ( .A1(_01559_ ), .A2(_01560_ ), .ZN(_00019_ ) );
OAI21_X1 _09089_ ( .A(_01555_ ), .B1(_01552_ ), .B2(\myclint.mtime [36] ), .ZN(_01561_ ) );
NOR2_X1 _09090_ ( .A1(_01561_ ), .A2(_01432_ ), .ZN(_00020_ ) );
NOR3_X1 _09091_ ( .A1(_01549_ ), .A2(_01550_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01562_ ) );
OAI21_X1 _09092_ ( .A(_01555_ ), .B1(_01562_ ), .B2(\myclint.mtime [35] ), .ZN(_01563_ ) );
INV_X1 _09093_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01564_ ) );
AND3_X1 _09094_ ( .A1(_01551_ ), .A2(_01564_ ), .A3(\myclint.mtime [35] ), .ZN(_01565_ ) );
NOR2_X1 _09095_ ( .A1(_01563_ ), .A2(_01565_ ), .ZN(_00021_ ) );
OAI21_X1 _09096_ ( .A(_01555_ ), .B1(_01551_ ), .B2(\myclint.mtime [34] ), .ZN(_01566_ ) );
NOR2_X1 _09097_ ( .A1(_01566_ ), .A2(_01431_ ), .ZN(_00022_ ) );
XNOR2_X1 _09098_ ( .A(_01529_ ), .B(\myclint.mtime [60] ), .ZN(_01567_ ) );
NOR2_X1 _09099_ ( .A1(_01567_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
AND2_X1 _09100_ ( .A1(_01427_ ), .A2(_01429_ ), .ZN(_01568_ ) );
INV_X1 _09101_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01569_ ) );
AND3_X1 _09102_ ( .A1(_01568_ ), .A2(_01569_ ), .A3(_01428_ ), .ZN(_01570_ ) );
AND2_X1 _09103_ ( .A1(_01570_ ), .A2(\myclint.mtime [33] ), .ZN(_01571_ ) );
OAI21_X1 _09104_ ( .A(_01516_ ), .B1(_01570_ ), .B2(\myclint.mtime [33] ), .ZN(_01572_ ) );
NOR2_X1 _09105_ ( .A1(_01571_ ), .A2(_01572_ ), .ZN(_00024_ ) );
NAND4_X1 _09106_ ( .A1(_01475_ ), .A2(_01550_ ), .A3(_01464_ ), .A4(_01467_ ), .ZN(_01573_ ) );
OAI21_X1 _09107_ ( .A(\myclint.mtime [32] ), .B1(_01508_ ), .B2(_01509_ ), .ZN(_01574_ ) );
AOI21_X1 _09108_ ( .A(fanout_net_1 ), .B1(_01573_ ), .B2(_01574_ ), .ZN(_00025_ ) );
INV_X1 _09109_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01575_ ) );
AND3_X1 _09110_ ( .A1(_01427_ ), .A2(_01575_ ), .A3(_01429_ ), .ZN(_01576_ ) );
AND2_X1 _09111_ ( .A1(_01576_ ), .A2(\myclint.mtime [31] ), .ZN(_01577_ ) );
OAI21_X1 _09112_ ( .A(_01516_ ), .B1(_01576_ ), .B2(\myclint.mtime [31] ), .ZN(_01578_ ) );
NOR2_X1 _09113_ ( .A1(_01577_ ), .A2(_01578_ ), .ZN(_00026_ ) );
AND2_X1 _09114_ ( .A1(_01468_ ), .A2(_01472_ ), .ZN(_01579_ ) );
NAND3_X1 _09115_ ( .A1(_01579_ ), .A2(_01429_ ), .A3(_01474_ ), .ZN(_01580_ ) );
OR2_X1 _09116_ ( .A1(_01580_ ), .A2(\myclint.mtime [30] ), .ZN(_01581_ ) );
NAND2_X1 _09117_ ( .A1(_01580_ ), .A2(\myclint.mtime [30] ), .ZN(_01582_ ) );
AOI21_X1 _09118_ ( .A(fanout_net_1 ), .B1(_01581_ ), .B2(_01582_ ), .ZN(_00027_ ) );
INV_X1 _09119_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01583_ ) );
AND3_X1 _09120_ ( .A1(_01426_ ), .A2(_01583_ ), .A3(\myclint.mtime [27] ), .ZN(_01584_ ) );
AND2_X1 _09121_ ( .A1(_01584_ ), .A2(\myclint.mtime [29] ), .ZN(_01585_ ) );
OAI21_X1 _09122_ ( .A(_01516_ ), .B1(_01584_ ), .B2(\myclint.mtime [29] ), .ZN(_01586_ ) );
NOR2_X1 _09123_ ( .A1(_01585_ ), .A2(_01586_ ), .ZN(_00028_ ) );
NAND2_X1 _09124_ ( .A1(_01579_ ), .A2(_01474_ ), .ZN(_01587_ ) );
OR2_X1 _09125_ ( .A1(_01587_ ), .A2(\myclint.mtime [28] ), .ZN(_01588_ ) );
NAND2_X1 _09126_ ( .A1(_01587_ ), .A2(\myclint.mtime [28] ), .ZN(_01589_ ) );
AOI21_X1 _09127_ ( .A(fanout_net_1 ), .B1(_01588_ ), .B2(_01589_ ), .ZN(_00029_ ) );
NAND3_X1 _09128_ ( .A1(_01468_ ), .A2(_01473_ ), .A3(_01472_ ), .ZN(_01590_ ) );
OR3_X1 _09129_ ( .A1(_01590_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01591_ ) );
OAI21_X1 _09130_ ( .A(\myclint.mtime [27] ), .B1(_01590_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01592_ ) );
AOI21_X1 _09131_ ( .A(fanout_net_1 ), .B1(_01591_ ), .B2(_01592_ ), .ZN(_00030_ ) );
AND2_X1 _09132_ ( .A1(_01425_ ), .A2(\myclint.mtime [25] ), .ZN(_01593_ ) );
OAI21_X1 _09133_ ( .A(_01555_ ), .B1(_01593_ ), .B2(\myclint.mtime [26] ), .ZN(_01594_ ) );
NOR2_X1 _09134_ ( .A1(_01594_ ), .A2(_01426_ ), .ZN(_00031_ ) );
INV_X1 _09135_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01595_ ) );
AND3_X1 _09136_ ( .A1(_01424_ ), .A2(_01595_ ), .A3(\myclint.mtime [23] ), .ZN(_01596_ ) );
AND2_X1 _09137_ ( .A1(_01596_ ), .A2(\myclint.mtime [25] ), .ZN(_01597_ ) );
OAI21_X1 _09138_ ( .A(_01516_ ), .B1(_01596_ ), .B2(\myclint.mtime [25] ), .ZN(_01598_ ) );
NOR2_X1 _09139_ ( .A1(_01597_ ), .A2(_01598_ ), .ZN(_00032_ ) );
AND2_X1 _09140_ ( .A1(_01424_ ), .A2(\myclint.mtime [23] ), .ZN(_01599_ ) );
OAI21_X1 _09141_ ( .A(_01555_ ), .B1(_01599_ ), .B2(\myclint.mtime [24] ), .ZN(_01600_ ) );
NOR2_X1 _09142_ ( .A1(_01600_ ), .A2(_01425_ ), .ZN(_00033_ ) );
NAND3_X1 _09143_ ( .A1(_01484_ ), .A2(_01450_ ), .A3(_01485_ ), .ZN(_01601_ ) );
OR3_X1 _09144_ ( .A1(_01601_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [59] ), .ZN(_01602_ ) );
OAI21_X1 _09145_ ( .A(\myclint.mtime [59] ), .B1(_01601_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01603_ ) );
AOI21_X1 _09146_ ( .A(fanout_net_1 ), .B1(_01602_ ), .B2(_01603_ ), .ZN(_00034_ ) );
NOR2_X1 _09147_ ( .A1(_01508_ ), .A2(_01470_ ), .ZN(_01604_ ) );
NAND3_X1 _09148_ ( .A1(_01604_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01605_ ) );
OR3_X1 _09149_ ( .A1(_01605_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01606_ ) );
OAI21_X1 _09150_ ( .A(\myclint.mtime [23] ), .B1(_01605_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01607_ ) );
AOI21_X1 _09151_ ( .A(fanout_net_1 ), .B1(_01606_ ), .B2(_01607_ ), .ZN(_00035_ ) );
AND2_X1 _09152_ ( .A1(_01423_ ), .A2(\myclint.mtime [21] ), .ZN(_01608_ ) );
OAI21_X1 _09153_ ( .A(_01555_ ), .B1(_01608_ ), .B2(\myclint.mtime [22] ), .ZN(_01609_ ) );
NOR2_X1 _09154_ ( .A1(_01609_ ), .A2(_01424_ ), .ZN(_00036_ ) );
OR3_X1 _09155_ ( .A1(_01508_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01470_ ), .ZN(_01610_ ) );
NAND2_X1 _09156_ ( .A1(_01610_ ), .A2(\myclint.mtime [21] ), .ZN(_01611_ ) );
OR4_X1 _09157_ ( .A1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01508_ ), .A3(\myclint.mtime [21] ), .A4(_01470_ ), .ZN(_01612_ ) );
AOI21_X1 _09158_ ( .A(fanout_net_1 ), .B1(_01611_ ), .B2(_01612_ ), .ZN(_00037_ ) );
AND2_X1 _09159_ ( .A1(_01422_ ), .A2(\myclint.mtime [19] ), .ZN(_01613_ ) );
OAI21_X1 _09160_ ( .A(_01555_ ), .B1(_01613_ ), .B2(\myclint.mtime [20] ), .ZN(_01614_ ) );
NOR2_X1 _09161_ ( .A1(_01614_ ), .A2(_01423_ ), .ZN(_00038_ ) );
NAND3_X1 _09162_ ( .A1(_01464_ ), .A2(_01467_ ), .A3(_01469_ ), .ZN(_01615_ ) );
OR3_X1 _09163_ ( .A1(_01615_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01616_ ) );
OAI21_X1 _09164_ ( .A(\myclint.mtime [19] ), .B1(_01615_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01617_ ) );
AOI21_X1 _09165_ ( .A(fanout_net_1 ), .B1(_01616_ ), .B2(_01617_ ), .ZN(_00039_ ) );
AND2_X1 _09166_ ( .A1(_01421_ ), .A2(\myclint.mtime [17] ), .ZN(_01618_ ) );
OAI21_X1 _09167_ ( .A(_01555_ ), .B1(_01618_ ), .B2(\myclint.mtime [18] ), .ZN(_01619_ ) );
NOR2_X1 _09168_ ( .A1(_01619_ ), .A2(_01422_ ), .ZN(_00040_ ) );
INV_X1 _09169_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01620_ ) );
AND3_X1 _09170_ ( .A1(_01420_ ), .A2(_01620_ ), .A3(\myclint.mtime [15] ), .ZN(_01621_ ) );
AND2_X1 _09171_ ( .A1(_01621_ ), .A2(\myclint.mtime [17] ), .ZN(_01622_ ) );
OAI21_X1 _09172_ ( .A(_01516_ ), .B1(_01621_ ), .B2(\myclint.mtime [17] ), .ZN(_01623_ ) );
NOR2_X1 _09173_ ( .A1(_01622_ ), .A2(_01623_ ), .ZN(_00041_ ) );
AND2_X1 _09174_ ( .A1(_01420_ ), .A2(\myclint.mtime [15] ), .ZN(_01624_ ) );
OAI21_X1 _09175_ ( .A(_01460_ ), .B1(_01624_ ), .B2(\myclint.mtime [16] ), .ZN(_01625_ ) );
NOR2_X1 _09176_ ( .A1(_01625_ ), .A2(_01421_ ), .ZN(_00042_ ) );
AND3_X1 _09177_ ( .A1(_01466_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [11] ), .ZN(_01626_ ) );
AND2_X1 _09178_ ( .A1(_01464_ ), .A2(_01626_ ), .ZN(_01627_ ) );
NAND3_X1 _09179_ ( .A1(_01627_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01628_ ) );
OR3_X1 _09180_ ( .A1(_01628_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01629_ ) );
OAI21_X1 _09181_ ( .A(\myclint.mtime [15] ), .B1(_01628_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01630_ ) );
AOI21_X1 _09182_ ( .A(fanout_net_1 ), .B1(_01629_ ), .B2(_01630_ ), .ZN(_00043_ ) );
AND2_X1 _09183_ ( .A1(_01419_ ), .A2(\myclint.mtime [13] ), .ZN(_01631_ ) );
OAI21_X1 _09184_ ( .A(_01460_ ), .B1(_01631_ ), .B2(\myclint.mtime [14] ), .ZN(_01632_ ) );
NOR2_X1 _09185_ ( .A1(_01632_ ), .A2(_01420_ ), .ZN(_00044_ ) );
OR2_X1 _09186_ ( .A1(_01601_ ), .A2(\myclint.mtime [58] ), .ZN(_01633_ ) );
NAND2_X1 _09187_ ( .A1(_01601_ ), .A2(\myclint.mtime [58] ), .ZN(_01634_ ) );
AOI21_X1 _09188_ ( .A(fanout_net_1 ), .B1(_01633_ ), .B2(_01634_ ), .ZN(_00045_ ) );
INV_X1 _09189_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01635_ ) );
AND3_X1 _09190_ ( .A1(_01418_ ), .A2(_01635_ ), .A3(\myclint.mtime [11] ), .ZN(_01636_ ) );
AND2_X1 _09191_ ( .A1(_01636_ ), .A2(\myclint.mtime [13] ), .ZN(_01637_ ) );
OAI21_X1 _09192_ ( .A(_01516_ ), .B1(_01636_ ), .B2(\myclint.mtime [13] ), .ZN(_01638_ ) );
NOR2_X1 _09193_ ( .A1(_01637_ ), .A2(_01638_ ), .ZN(_00046_ ) );
AND2_X1 _09194_ ( .A1(_01418_ ), .A2(\myclint.mtime [11] ), .ZN(_01639_ ) );
OAI21_X1 _09195_ ( .A(_01460_ ), .B1(_01639_ ), .B2(\myclint.mtime [12] ), .ZN(_01640_ ) );
NOR2_X1 _09196_ ( .A1(_01640_ ), .A2(_01419_ ), .ZN(_00047_ ) );
NAND3_X1 _09197_ ( .A1(_01462_ ), .A2(_01463_ ), .A3(_01466_ ), .ZN(_01641_ ) );
OR3_X1 _09198_ ( .A1(_01641_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_01642_ ) );
OAI21_X1 _09199_ ( .A(\myclint.mtime [11] ), .B1(_01641_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01643_ ) );
AOI21_X1 _09200_ ( .A(fanout_net_1 ), .B1(_01642_ ), .B2(_01643_ ), .ZN(_00048_ ) );
AND2_X1 _09201_ ( .A1(_01417_ ), .A2(\myclint.mtime [9] ), .ZN(_01644_ ) );
OAI21_X1 _09202_ ( .A(_01460_ ), .B1(_01644_ ), .B2(\myclint.mtime [10] ), .ZN(_01645_ ) );
NOR2_X1 _09203_ ( .A1(_01645_ ), .A2(_01418_ ), .ZN(_00049_ ) );
AND2_X1 _09204_ ( .A1(_01416_ ), .A2(\myclint.mtime [7] ), .ZN(_01646_ ) );
INV_X1 _09205_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01647_ ) );
AND3_X1 _09206_ ( .A1(_01646_ ), .A2(\myclint.mtime [9] ), .A3(_01647_ ), .ZN(_01648_ ) );
AOI21_X1 _09207_ ( .A(\myclint.mtime [9] ), .B1(_01646_ ), .B2(_01647_ ), .ZN(_01649_ ) );
NOR3_X1 _09208_ ( .A1(_01648_ ), .A2(_01649_ ), .A3(fanout_net_1 ), .ZN(_00050_ ) );
OAI21_X1 _09209_ ( .A(_01460_ ), .B1(_01646_ ), .B2(\myclint.mtime [8] ), .ZN(_01650_ ) );
NOR2_X1 _09210_ ( .A1(_01650_ ), .A2(_01417_ ), .ZN(_00051_ ) );
AND2_X1 _09211_ ( .A1(_01415_ ), .A2(\myclint.mtime [5] ), .ZN(_01651_ ) );
INV_X1 _09212_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01652_ ) );
AND3_X1 _09213_ ( .A1(_01651_ ), .A2(_01652_ ), .A3(\myclint.mtime [7] ), .ZN(_01653_ ) );
AOI21_X1 _09214_ ( .A(\myclint.mtime [7] ), .B1(_01651_ ), .B2(_01652_ ), .ZN(_01654_ ) );
NOR3_X1 _09215_ ( .A1(_01653_ ), .A2(_01654_ ), .A3(fanout_net_1 ), .ZN(_00052_ ) );
OAI21_X1 _09216_ ( .A(_01460_ ), .B1(_01651_ ), .B2(\myclint.mtime [6] ), .ZN(_01655_ ) );
NOR2_X1 _09217_ ( .A1(_01655_ ), .A2(_01416_ ), .ZN(_00053_ ) );
INV_X1 _09218_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01656_ ) );
AND3_X1 _09219_ ( .A1(_01462_ ), .A2(\myclint.mtime [5] ), .A3(_01656_ ), .ZN(_01657_ ) );
AOI21_X1 _09220_ ( .A(\myclint.mtime [5] ), .B1(_01462_ ), .B2(_01656_ ), .ZN(_01658_ ) );
NOR3_X1 _09221_ ( .A1(_01657_ ), .A2(_01658_ ), .A3(fanout_net_1 ), .ZN(_00054_ ) );
OAI21_X1 _09222_ ( .A(_01460_ ), .B1(_01462_ ), .B2(\myclint.mtime [4] ), .ZN(_01659_ ) );
NOR2_X1 _09223_ ( .A1(_01659_ ), .A2(_01415_ ), .ZN(_00055_ ) );
INV_X1 _09224_ ( .A(_01486_ ), .ZN(_01660_ ) );
OR3_X1 _09225_ ( .A1(_01660_ ), .A2(\myclint.mtime [57] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01661_ ) );
OAI21_X1 _09226_ ( .A(\myclint.mtime [57] ), .B1(_01660_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01662_ ) );
AOI21_X1 _09227_ ( .A(fanout_net_1 ), .B1(_01661_ ), .B2(_01662_ ), .ZN(_00056_ ) );
AND2_X1 _09228_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01663_ ) );
INV_X1 _09229_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01664_ ) );
AND3_X1 _09230_ ( .A1(_01663_ ), .A2(_01664_ ), .A3(\myclint.mtime [3] ), .ZN(_01665_ ) );
AOI21_X1 _09231_ ( .A(\myclint.mtime [3] ), .B1(_01663_ ), .B2(_01664_ ), .ZN(_01666_ ) );
NOR3_X1 _09232_ ( .A1(_01665_ ), .A2(_01666_ ), .A3(fanout_net_1 ), .ZN(_00057_ ) );
AOI21_X1 _09233_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01667_ ) );
NOR3_X1 _09234_ ( .A1(_01414_ ), .A2(_01667_ ), .A3(fanout_net_2 ), .ZN(_00058_ ) );
NOR2_X1 _09235_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01668_ ) );
NOR3_X1 _09236_ ( .A1(_01663_ ), .A2(_01668_ ), .A3(fanout_net_2 ), .ZN(_00059_ ) );
INV_X1 _09237_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_01669_ ) );
NOR2_X1 _09238_ ( .A1(_01669_ ), .A2(fanout_net_2 ), .ZN(_00060_ ) );
XNOR2_X1 _09239_ ( .A(_01486_ ), .B(\myclint.mtime [56] ), .ZN(_01670_ ) );
NOR2_X1 _09240_ ( .A1(_01670_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
NAND3_X1 _09241_ ( .A1(_01484_ ), .A2(_01446_ ), .A3(_01491_ ), .ZN(_01671_ ) );
OR3_X1 _09242_ ( .A1(_01671_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01672_ ) );
OAI21_X1 _09243_ ( .A(\myclint.mtime [55] ), .B1(_01671_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01673_ ) );
AOI21_X1 _09244_ ( .A(fanout_net_2 ), .B1(_01672_ ), .B2(_01673_ ), .ZN(_00062_ ) );
OR2_X1 _09245_ ( .A1(_01671_ ), .A2(\myclint.mtime [54] ), .ZN(_01674_ ) );
NAND2_X1 _09246_ ( .A1(_01671_ ), .A2(\myclint.mtime [54] ), .ZN(_01675_ ) );
AOI21_X1 _09247_ ( .A(fanout_net_2 ), .B1(_01674_ ), .B2(_01675_ ), .ZN(_00063_ ) );
INV_X32 _09248_ ( .A(fanout_net_42 ), .ZN(_01676_ ) );
CLKBUF_X2 _09249_ ( .A(_01676_ ), .Z(_01677_ ) );
OR2_X1 _09250_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[1][4] ), .ZN(_01678_ ) );
INV_X32 _09251_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01679_ ) );
BUF_X4 _09252_ ( .A(_01679_ ), .Z(_01680_ ) );
BUF_X4 _09253_ ( .A(_01680_ ), .Z(_01681_ ) );
OAI211_X1 _09254_ ( .A(_01678_ ), .B(_01681_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][4] ), .ZN(_01682_ ) );
OR2_X1 _09255_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[3][4] ), .ZN(_01683_ ) );
OAI211_X1 _09256_ ( .A(_01683_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[2][4] ), .ZN(_01684_ ) );
NAND2_X1 _09257_ ( .A1(_01682_ ), .A2(_01684_ ), .ZN(_01685_ ) );
INV_X1 _09258_ ( .A(\IF_ID_pc [9] ), .ZN(_01686_ ) );
XNOR2_X1 _09259_ ( .A(_01685_ ), .B(_01686_ ), .ZN(_01687_ ) );
BUF_X32 _09260_ ( .A(_01676_ ), .Z(_01688_ ) );
OR2_X4 _09261_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[1][13] ), .ZN(_01689_ ) );
OAI211_X2 _09262_ ( .A(_01689_ ), .B(_01680_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][13] ), .ZN(_01690_ ) );
OR2_X4 _09263_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[3][13] ), .ZN(_01691_ ) );
OAI211_X2 _09264_ ( .A(_01691_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[2][13] ), .ZN(_01692_ ) );
AOI21_X2 _09265_ ( .A(\IF_ID_pc [18] ), .B1(_01690_ ), .B2(_01692_ ), .ZN(_01693_ ) );
OR2_X4 _09266_ ( .A1(_01676_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01694_ ) );
OAI211_X2 _09267_ ( .A(_01694_ ), .B(_01679_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01695_ ) );
OR2_X4 _09268_ ( .A1(_01676_ ), .A2(\myifu.myicache.tag[3][12] ), .ZN(_01696_ ) );
OAI211_X4 _09269_ ( .A(_01696_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[2][12] ), .ZN(_01697_ ) );
NAND2_X2 _09270_ ( .A1(_01695_ ), .A2(_01697_ ), .ZN(_01698_ ) );
INV_X1 _09271_ ( .A(\IF_ID_pc [17] ), .ZN(_01699_ ) );
XNOR2_X2 _09272_ ( .A(_01698_ ), .B(_01699_ ), .ZN(_01700_ ) );
MUX2_X1 _09273_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_42 ), .Z(_01701_ ) );
OR2_X1 _09274_ ( .A1(_01701_ ), .A2(_01680_ ), .ZN(_01702_ ) );
MUX2_X1 _09275_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_42 ), .Z(_01703_ ) );
OAI21_X1 _09276_ ( .A(_01702_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01703_ ), .ZN(_01704_ ) );
AOI211_X2 _09277_ ( .A(_01693_ ), .B(_01700_ ), .C1(\IF_ID_pc [16] ), .C2(_01704_ ), .ZN(_01705_ ) );
MUX2_X1 _09278_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(fanout_net_42 ), .Z(_01706_ ) );
OR2_X1 _09279_ ( .A1(_01706_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01707_ ) );
MUX2_X1 _09280_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(fanout_net_42 ), .Z(_01708_ ) );
OAI21_X1 _09281_ ( .A(_01707_ ), .B1(_01681_ ), .B2(_01708_ ), .ZN(_01709_ ) );
OR2_X1 _09282_ ( .A1(_01709_ ), .A2(\IF_ID_pc [20] ), .ZN(_01710_ ) );
NAND3_X1 _09283_ ( .A1(_01690_ ), .A2(_01692_ ), .A3(\IF_ID_pc [18] ), .ZN(_01711_ ) );
MUX2_X1 _09284_ ( .A(\myifu.myicache.tag[2][14] ), .B(\myifu.myicache.tag[3][14] ), .S(fanout_net_42 ), .Z(_01712_ ) );
OR2_X2 _09285_ ( .A1(_01712_ ), .A2(_01679_ ), .ZN(_01713_ ) );
MUX2_X1 _09286_ ( .A(\myifu.myicache.tag[0][14] ), .B(\myifu.myicache.tag[1][14] ), .S(fanout_net_42 ), .Z(_01714_ ) );
OR2_X2 _09287_ ( .A1(_01714_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01715_ ) );
AND2_X2 _09288_ ( .A1(_01713_ ), .A2(_01715_ ), .ZN(_01716_ ) );
XNOR2_X1 _09289_ ( .A(_01716_ ), .B(\IF_ID_pc [19] ), .ZN(_01717_ ) );
NAND4_X1 _09290_ ( .A1(_01705_ ), .A2(_01710_ ), .A3(_01711_ ), .A4(_01717_ ), .ZN(_01718_ ) );
MUX2_X1 _09291_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(fanout_net_42 ), .Z(_01719_ ) );
AND2_X1 _09292_ ( .A1(_01719_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01720_ ) );
MUX2_X1 _09293_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(fanout_net_42 ), .Z(_01721_ ) );
AOI21_X1 _09294_ ( .A(_01720_ ), .B1(_01681_ ), .B2(_01721_ ), .ZN(_01722_ ) );
NAND2_X1 _09295_ ( .A1(_01722_ ), .A2(\IF_ID_pc [12] ), .ZN(_01723_ ) );
MUX2_X1 _09296_ ( .A(\myifu.myicache.tag[2][3] ), .B(\myifu.myicache.tag[3][3] ), .S(fanout_net_42 ), .Z(_01724_ ) );
OR2_X1 _09297_ ( .A1(_01724_ ), .A2(_01680_ ), .ZN(_01725_ ) );
MUX2_X1 _09298_ ( .A(\myifu.myicache.tag[0][3] ), .B(\myifu.myicache.tag[1][3] ), .S(fanout_net_42 ), .Z(_01726_ ) );
OAI21_X1 _09299_ ( .A(_01725_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01726_ ), .ZN(_01727_ ) );
INV_X1 _09300_ ( .A(\IF_ID_pc [21] ), .ZN(_01728_ ) );
OR2_X4 _09301_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[1][16] ), .ZN(_01729_ ) );
OAI211_X1 _09302_ ( .A(_01729_ ), .B(_01680_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][16] ), .ZN(_01730_ ) );
OR2_X4 _09303_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[3][16] ), .ZN(_01731_ ) );
OAI211_X2 _09304_ ( .A(_01731_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[2][16] ), .ZN(_01732_ ) );
NAND2_X1 _09305_ ( .A1(_01730_ ), .A2(_01732_ ), .ZN(_01733_ ) );
AOI22_X1 _09306_ ( .A1(_01727_ ), .A2(\IF_ID_pc [8] ), .B1(_01728_ ), .B2(_01733_ ), .ZN(_01734_ ) );
OAI211_X1 _09307_ ( .A(_01723_ ), .B(_01734_ ), .C1(\IF_ID_pc [8] ), .C2(_01727_ ), .ZN(_01735_ ) );
OR2_X1 _09308_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_01736_ ) );
OAI211_X1 _09309_ ( .A(_01736_ ), .B(_01680_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_01737_ ) );
OR2_X1 _09310_ ( .A1(fanout_net_42 ), .A2(\myifu.myicache.tag[2][6] ), .ZN(_01738_ ) );
OAI211_X1 _09311_ ( .A(_01738_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01677_ ), .C2(\myifu.myicache.tag[3][6] ), .ZN(_01739_ ) );
NAND2_X1 _09312_ ( .A1(_01737_ ), .A2(_01739_ ), .ZN(_01740_ ) );
INV_X1 _09313_ ( .A(\IF_ID_pc [11] ), .ZN(_01741_ ) );
XNOR2_X1 _09314_ ( .A(_01740_ ), .B(_01741_ ), .ZN(_01742_ ) );
OR4_X4 _09315_ ( .A1(_01687_ ), .A2(_01718_ ), .A3(_01735_ ), .A4(_01742_ ), .ZN(_01743_ ) );
MUX2_X1 _09316_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(fanout_net_42 ), .Z(_01744_ ) );
MUX2_X1 _09317_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(fanout_net_42 ), .Z(_01745_ ) );
MUX2_X1 _09318_ ( .A(_01744_ ), .B(_01745_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01746_ ) );
OR2_X4 _09319_ ( .A1(_01676_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_01747_ ) );
OAI211_X2 _09320_ ( .A(_01747_ ), .B(_01679_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_01748_ ) );
OR2_X4 _09321_ ( .A1(_01676_ ), .A2(\myifu.myicache.tag[3][25] ), .ZN(_01749_ ) );
OAI211_X2 _09322_ ( .A(_01749_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[2][25] ), .ZN(_01750_ ) );
NAND2_X2 _09323_ ( .A1(_01748_ ), .A2(_01750_ ), .ZN(_01751_ ) );
XOR2_X1 _09324_ ( .A(_01751_ ), .B(\IF_ID_pc [30] ), .Z(_01752_ ) );
INV_X1 _09325_ ( .A(\IF_ID_pc [31] ), .ZN(_01753_ ) );
MUX2_X1 _09326_ ( .A(\myifu.myicache.tag[0][26] ), .B(\myifu.myicache.tag[1][26] ), .S(fanout_net_42 ), .Z(_01754_ ) );
MUX2_X1 _09327_ ( .A(\myifu.myicache.tag[2][26] ), .B(\myifu.myicache.tag[3][26] ), .S(fanout_net_42 ), .Z(_01755_ ) );
MUX2_X1 _09328_ ( .A(_01754_ ), .B(_01755_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01756_ ) );
MUX2_X1 _09329_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(fanout_net_42 ), .Z(_01757_ ) );
OR2_X1 _09330_ ( .A1(_01757_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01758_ ) );
MUX2_X1 _09331_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(fanout_net_42 ), .Z(_01759_ ) );
OAI21_X1 _09332_ ( .A(_01758_ ), .B1(_01680_ ), .B2(_01759_ ), .ZN(_01760_ ) );
AOI221_X2 _09333_ ( .A(_01752_ ), .B1(_01753_ ), .B2(_01756_ ), .C1(\IF_ID_pc [29] ), .C2(_01760_ ), .ZN(_01761_ ) );
OR2_X1 _09334_ ( .A1(_01756_ ), .A2(_01753_ ), .ZN(_01762_ ) );
OR2_X1 _09335_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[1][0] ), .ZN(_01763_ ) );
OAI211_X1 _09336_ ( .A(_01763_ ), .B(_01680_ ), .C1(fanout_net_42 ), .C2(\myifu.myicache.tag[0][0] ), .ZN(_01764_ ) );
OR2_X1 _09337_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[3][0] ), .ZN(_01765_ ) );
OAI211_X1 _09338_ ( .A(_01765_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][0] ), .ZN(_01766_ ) );
NAND2_X1 _09339_ ( .A1(_01764_ ), .A2(_01766_ ), .ZN(_01767_ ) );
XOR2_X1 _09340_ ( .A(_01767_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .Z(_01768_ ) );
AND4_X2 _09341_ ( .A1(_01746_ ), .A2(_01761_ ), .A3(_01762_ ), .A4(_01768_ ), .ZN(_01769_ ) );
OR2_X1 _09342_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[1][21] ), .ZN(_01770_ ) );
OAI211_X1 _09343_ ( .A(_01770_ ), .B(_01681_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][21] ), .ZN(_01771_ ) );
OR2_X1 _09344_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[3][21] ), .ZN(_01772_ ) );
OAI211_X1 _09345_ ( .A(_01772_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][21] ), .ZN(_01773_ ) );
NAND2_X1 _09346_ ( .A1(_01771_ ), .A2(_01773_ ), .ZN(_01774_ ) );
INV_X1 _09347_ ( .A(\IF_ID_pc [26] ), .ZN(_01775_ ) );
XNOR2_X1 _09348_ ( .A(_01774_ ), .B(_01775_ ), .ZN(_01776_ ) );
INV_X1 _09349_ ( .A(_01776_ ), .ZN(_01777_ ) );
MUX2_X1 _09350_ ( .A(\myifu.myicache.tag[0][23] ), .B(\myifu.myicache.tag[1][23] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01778_ ) );
NAND2_X1 _09351_ ( .A1(_01778_ ), .A2(_01681_ ), .ZN(_01779_ ) );
MUX2_X1 _09352_ ( .A(\myifu.myicache.tag[2][23] ), .B(\myifu.myicache.tag[3][23] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01780_ ) );
NAND2_X1 _09353_ ( .A1(_01780_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01781_ ) );
NAND2_X1 _09354_ ( .A1(_01779_ ), .A2(_01781_ ), .ZN(_01782_ ) );
XNOR2_X1 _09355_ ( .A(_01782_ ), .B(\IF_ID_pc [28] ), .ZN(_01783_ ) );
AND3_X1 _09356_ ( .A1(_01730_ ), .A2(_01732_ ), .A3(\IF_ID_pc [21] ), .ZN(_01784_ ) );
MUX2_X1 _09357_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01785_ ) );
MUX2_X1 _09358_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01786_ ) );
MUX2_X2 _09359_ ( .A(_01785_ ), .B(_01786_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01787_ ) );
INV_X1 _09360_ ( .A(\IF_ID_pc [25] ), .ZN(_01788_ ) );
NAND2_X1 _09361_ ( .A1(_01787_ ), .A2(_01788_ ), .ZN(_01789_ ) );
INV_X1 _09362_ ( .A(\IF_ID_pc [23] ), .ZN(_01790_ ) );
MUX2_X1 _09363_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01791_ ) );
MUX2_X1 _09364_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01792_ ) );
MUX2_X1 _09365_ ( .A(_01791_ ), .B(_01792_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01793_ ) );
OAI21_X1 _09366_ ( .A(_01789_ ), .B1(_01790_ ), .B2(_01793_ ), .ZN(_01794_ ) );
AOI211_X1 _09367_ ( .A(_01784_ ), .B(_01794_ ), .C1(_01790_ ), .C2(_01793_ ), .ZN(_01795_ ) );
NAND4_X4 _09368_ ( .A1(_01769_ ), .A2(_01777_ ), .A3(_01783_ ), .A4(_01795_ ), .ZN(_01796_ ) );
NOR2_X4 _09369_ ( .A1(_01743_ ), .A2(_01796_ ), .ZN(_01797_ ) );
MUX2_X1 _09370_ ( .A(\myifu.myicache.tag[2][2] ), .B(\myifu.myicache.tag[3][2] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01798_ ) );
OR2_X1 _09371_ ( .A1(_01798_ ), .A2(_01680_ ), .ZN(_01799_ ) );
MUX2_X1 _09372_ ( .A(\myifu.myicache.tag[0][2] ), .B(\myifu.myicache.tag[1][2] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01800_ ) );
OR2_X1 _09373_ ( .A1(_01800_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01801_ ) );
AND3_X1 _09374_ ( .A1(_01799_ ), .A2(_01801_ ), .A3(\IF_ID_pc [7] ), .ZN(_01802_ ) );
AOI21_X1 _09375_ ( .A(\IF_ID_pc [7] ), .B1(_01799_ ), .B2(_01801_ ), .ZN(_01803_ ) );
OR2_X1 _09376_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[1][1] ), .ZN(_01804_ ) );
OAI211_X1 _09377_ ( .A(_01804_ ), .B(_01680_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][1] ), .ZN(_01805_ ) );
OR2_X1 _09378_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[3][1] ), .ZN(_01806_ ) );
OAI211_X1 _09379_ ( .A(_01806_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][1] ), .ZN(_01807_ ) );
INV_X1 _09380_ ( .A(\IF_ID_pc [6] ), .ZN(_01808_ ) );
AND3_X1 _09381_ ( .A1(_01805_ ), .A2(_01807_ ), .A3(_01808_ ), .ZN(_01809_ ) );
AOI21_X1 _09382_ ( .A(_01808_ ), .B1(_01805_ ), .B2(_01807_ ), .ZN(_01810_ ) );
OAI22_X1 _09383_ ( .A1(_01802_ ), .A2(_01803_ ), .B1(_01809_ ), .B2(_01810_ ), .ZN(_01811_ ) );
NOR2_X1 _09384_ ( .A1(_01722_ ), .A2(\IF_ID_pc [12] ), .ZN(_01812_ ) );
MUX2_X1 _09385_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01813_ ) );
AND2_X2 _09386_ ( .A1(_01813_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01814_ ) );
MUX2_X1 _09387_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01815_ ) );
AOI21_X4 _09388_ ( .A(_01814_ ), .B1(_01681_ ), .B2(_01815_ ), .ZN(_01816_ ) );
AND2_X1 _09389_ ( .A1(_01816_ ), .A2(\IF_ID_pc [10] ), .ZN(_01817_ ) );
NAND2_X1 _09390_ ( .A1(_01709_ ), .A2(\IF_ID_pc [20] ), .ZN(_01818_ ) );
OAI21_X2 _09391_ ( .A(_01818_ ), .B1(\IF_ID_pc [10] ), .B2(_01816_ ), .ZN(_01819_ ) );
NOR4_X2 _09392_ ( .A1(_01811_ ), .A2(_01812_ ), .A3(_01817_ ), .A4(_01819_ ), .ZN(_01820_ ) );
OR2_X1 _09393_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[1][10] ), .ZN(_01821_ ) );
OAI211_X1 _09394_ ( .A(_01821_ ), .B(_01681_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][10] ), .ZN(_01822_ ) );
OR2_X1 _09395_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[3][10] ), .ZN(_01823_ ) );
OAI211_X1 _09396_ ( .A(_01823_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][10] ), .ZN(_01824_ ) );
NAND2_X1 _09397_ ( .A1(_01822_ ), .A2(_01824_ ), .ZN(_01825_ ) );
XNOR2_X1 _09398_ ( .A(_01825_ ), .B(\IF_ID_pc [15] ), .ZN(_01826_ ) );
MUX2_X1 _09399_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01827_ ) );
MUX2_X1 _09400_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01828_ ) );
MUX2_X1 _09401_ ( .A(_01827_ ), .B(_01828_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01829_ ) );
INV_X1 _09402_ ( .A(\IF_ID_pc [14] ), .ZN(_01830_ ) );
NAND2_X1 _09403_ ( .A1(_01829_ ), .A2(_01830_ ), .ZN(_01831_ ) );
OAI22_X1 _09404_ ( .A1(_01704_ ), .A2(\IF_ID_pc [16] ), .B1(_01830_ ), .B2(_01829_ ), .ZN(_01832_ ) );
OR2_X1 _09405_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[1][8] ), .ZN(_01833_ ) );
OAI211_X1 _09406_ ( .A(_01833_ ), .B(_01681_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][8] ), .ZN(_01834_ ) );
OR2_X1 _09407_ ( .A1(_01688_ ), .A2(\myifu.myicache.tag[3][8] ), .ZN(_01835_ ) );
OAI211_X1 _09408_ ( .A(_01835_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][8] ), .ZN(_01836_ ) );
NAND2_X1 _09409_ ( .A1(_01834_ ), .A2(_01836_ ), .ZN(_01837_ ) );
INV_X1 _09410_ ( .A(\IF_ID_pc [13] ), .ZN(_01838_ ) );
XNOR2_X1 _09411_ ( .A(_01837_ ), .B(_01838_ ), .ZN(_01839_ ) );
NOR2_X1 _09412_ ( .A1(_01832_ ), .A2(_01839_ ), .ZN(_01840_ ) );
NAND4_X1 _09413_ ( .A1(_01820_ ), .A2(_01826_ ), .A3(_01831_ ), .A4(_01840_ ), .ZN(_01841_ ) );
OR2_X1 _09414_ ( .A1(_01677_ ), .A2(\myifu.myicache.tag[1][17] ), .ZN(_01842_ ) );
OAI211_X1 _09415_ ( .A(_01842_ ), .B(_01681_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][17] ), .ZN(_01843_ ) );
OR2_X1 _09416_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][17] ), .ZN(_01844_ ) );
OAI211_X1 _09417_ ( .A(_01844_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01677_ ), .C2(\myifu.myicache.tag[3][17] ), .ZN(_01845_ ) );
NAND2_X1 _09418_ ( .A1(_01843_ ), .A2(_01845_ ), .ZN(_01846_ ) );
INV_X1 _09419_ ( .A(\IF_ID_pc [22] ), .ZN(_01847_ ) );
XNOR2_X1 _09420_ ( .A(_01846_ ), .B(_01847_ ), .ZN(_01848_ ) );
NOR2_X1 _09421_ ( .A1(_01787_ ), .A2(_01788_ ), .ZN(_01849_ ) );
INV_X1 _09422_ ( .A(\IF_ID_pc [27] ), .ZN(_01850_ ) );
MUX2_X1 _09423_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01851_ ) );
MUX2_X1 _09424_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01852_ ) );
MUX2_X1 _09425_ ( .A(_01851_ ), .B(_01852_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01853_ ) );
AOI21_X1 _09426_ ( .A(_01849_ ), .B1(_01850_ ), .B2(_01853_ ), .ZN(_01854_ ) );
OAI221_X1 _09427_ ( .A(_01854_ ), .B1(\IF_ID_pc [29] ), .B2(_01760_ ), .C1(_01850_ ), .C2(_01853_ ), .ZN(_01855_ ) );
MUX2_X1 _09428_ ( .A(\myifu.myicache.tag[2][19] ), .B(\myifu.myicache.tag[3][19] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01856_ ) );
NOR2_X1 _09429_ ( .A1(_01856_ ), .A2(_01681_ ), .ZN(_01857_ ) );
MUX2_X1 _09430_ ( .A(\myifu.myicache.tag[0][19] ), .B(\myifu.myicache.tag[1][19] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01858_ ) );
NOR2_X1 _09431_ ( .A1(_01858_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01859_ ) );
NOR2_X1 _09432_ ( .A1(_01857_ ), .A2(_01859_ ), .ZN(_01860_ ) );
INV_X1 _09433_ ( .A(\IF_ID_pc [24] ), .ZN(_01861_ ) );
XNOR2_X1 _09434_ ( .A(_01860_ ), .B(_01861_ ), .ZN(_01862_ ) );
NOR4_X4 _09435_ ( .A1(_01841_ ), .A2(_01848_ ), .A3(_01855_ ), .A4(_01862_ ), .ZN(_01863_ ) );
NAND2_X4 _09436_ ( .A1(_01797_ ), .A2(_01863_ ), .ZN(_01864_ ) );
AND2_X4 _09437_ ( .A1(_01864_ ), .A2(\myifu.state [0] ), .ZN(_01865_ ) );
INV_X1 _09438_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01866_ ) );
NOR2_X4 _09439_ ( .A1(_01865_ ), .A2(_01866_ ), .ZN(_01867_ ) );
NOR2_X1 _09440_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01868_ ) );
NOR2_X4 _09441_ ( .A1(_01867_ ), .A2(_01868_ ), .ZN(_01869_ ) );
INV_X32 _09442_ ( .A(\EX_LS_flag [1] ), .ZN(_01870_ ) );
INV_X1 _09443_ ( .A(\EX_LS_flag [0] ), .ZN(_01871_ ) );
OR4_X1 _09444_ ( .A1(\EX_LS_flag [2] ), .A2(_01870_ ), .A3(_01871_ ), .A4(\mylsu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__A_B ), .ZN(_01872_ ) );
INV_X1 _09445_ ( .A(EXU_valid_LSU ), .ZN(_01873_ ) );
NOR2_X1 _09446_ ( .A1(_01872_ ), .A2(_01873_ ), .ZN(_01874_ ) );
INV_X1 _09447_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01875_ ) );
NOR2_X1 _09448_ ( .A1(_01874_ ), .A2(_01875_ ), .ZN(_01876_ ) );
NOR2_X4 _09449_ ( .A1(_01869_ ), .A2(_01876_ ), .ZN(_01877_ ) );
BUF_X4 _09450_ ( .A(_01877_ ), .Z(_01878_ ) );
CLKBUF_X2 _09451_ ( .A(_01872_ ), .Z(_01879_ ) );
OR3_X1 _09452_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(_01873_ ), .ZN(_01880_ ) );
BUF_X4 _09453_ ( .A(_01874_ ), .Z(_01881_ ) );
OAI211_X1 _09454_ ( .A(_01878_ ), .B(_01880_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01881_ ), .ZN(_01882_ ) );
INV_X4 _09455_ ( .A(_01869_ ), .ZN(_01883_ ) );
OAI21_X1 _09456_ ( .A(_01882_ ), .B1(_01790_ ), .B2(_01883_ ), .ZN(\io_master_araddr [23] ) );
BUF_X8 _09457_ ( .A(_01877_ ), .Z(_01884_ ) );
CLKBUF_X2 _09458_ ( .A(_01872_ ), .Z(_01885_ ) );
CLKBUF_X2 _09459_ ( .A(_01873_ ), .Z(_01886_ ) );
OR3_X1 _09460_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(_01886_ ), .ZN(_01887_ ) );
BUF_X4 _09461_ ( .A(_01874_ ), .Z(_01888_ ) );
OAI211_X1 _09462_ ( .A(_01884_ ), .B(_01887_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01888_ ), .ZN(_01889_ ) );
BUF_X2 _09463_ ( .A(_01865_ ), .Z(_01890_ ) );
BUF_X4 _09464_ ( .A(_01866_ ), .Z(_01891_ ) );
OAI221_X1 _09465_ ( .A(\IF_ID_pc [30] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01890_ ), .C2(_01891_ ), .ZN(_01892_ ) );
AND2_X1 _09466_ ( .A1(_01889_ ), .A2(_01892_ ), .ZN(_01893_ ) );
OR3_X1 _09467_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(_01886_ ), .ZN(_01894_ ) );
OAI211_X1 _09468_ ( .A(_01878_ ), .B(_01894_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01888_ ), .ZN(_01895_ ) );
OAI221_X1 _09469_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01890_ ), .C2(_01891_ ), .ZN(_01896_ ) );
AND2_X1 _09470_ ( .A1(_01895_ ), .A2(_01896_ ), .ZN(_01897_ ) );
OR3_X1 _09471_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(_01886_ ), .ZN(_01898_ ) );
OAI211_X1 _09472_ ( .A(_01878_ ), .B(_01898_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01881_ ), .ZN(_01899_ ) );
OAI221_X1 _09473_ ( .A(\IF_ID_pc [24] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01890_ ), .C2(_01891_ ), .ZN(_01900_ ) );
AND2_X1 _09474_ ( .A1(_01899_ ), .A2(_01900_ ), .ZN(_01901_ ) );
OR3_X1 _09475_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [25] ), .A3(_01886_ ), .ZN(_01902_ ) );
OAI211_X4 _09476_ ( .A(_01884_ ), .B(_01902_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_01888_ ), .ZN(_01903_ ) );
OAI21_X4 _09477_ ( .A(_01903_ ), .B1(_01788_ ), .B2(_01883_ ), .ZN(\io_master_araddr [25] ) );
NAND4_X1 _09478_ ( .A1(_01893_ ), .A2(_01897_ ), .A3(_01901_ ), .A4(\io_master_araddr [25] ), .ZN(_01904_ ) );
OR3_X1 _09479_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(_01886_ ), .ZN(_01905_ ) );
OAI211_X1 _09480_ ( .A(_01878_ ), .B(_01905_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01881_ ), .ZN(_01906_ ) );
OAI21_X1 _09481_ ( .A(_01906_ ), .B1(_01699_ ), .B2(_01883_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09482_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(_01873_ ), .ZN(_01907_ ) );
OAI211_X1 _09483_ ( .A(_01878_ ), .B(_01907_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01881_ ), .ZN(_01908_ ) );
INV_X1 _09484_ ( .A(\IF_ID_pc [18] ), .ZN(_01909_ ) );
OAI21_X1 _09485_ ( .A(_01908_ ), .B1(_01909_ ), .B2(_01883_ ), .ZN(\io_master_araddr [18] ) );
OR2_X1 _09486_ ( .A1(\io_master_araddr [17] ), .A2(\io_master_araddr [18] ), .ZN(_01910_ ) );
OR3_X1 _09487_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(_01873_ ), .ZN(_01911_ ) );
OAI211_X1 _09488_ ( .A(_01878_ ), .B(_01911_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01881_ ), .ZN(_01912_ ) );
INV_X1 _09489_ ( .A(\IF_ID_pc [20] ), .ZN(_01913_ ) );
OAI21_X2 _09490_ ( .A(_01912_ ), .B1(_01913_ ), .B2(_01883_ ), .ZN(\io_master_araddr [20] ) );
OR4_X1 _09491_ ( .A1(\io_master_araddr [23] ), .A2(_01904_ ), .A3(_01910_ ), .A4(\io_master_araddr [20] ), .ZN(_01914_ ) );
CLKBUF_X2 _09492_ ( .A(_01869_ ), .Z(_01915_ ) );
CLKBUF_X2 _09493_ ( .A(_01915_ ), .Z(_01916_ ) );
CLKBUF_X2 _09494_ ( .A(_01916_ ), .Z(_01917_ ) );
CLKBUF_X2 _09495_ ( .A(_01917_ ), .Z(_01918_ ) );
OR2_X1 _09496_ ( .A1(\EX_LS_dest_csreg_mem [27] ), .A2(\EX_LS_dest_csreg_mem [26] ), .ZN(_01919_ ) );
NOR3_X1 _09497_ ( .A1(_01919_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(\EX_LS_dest_csreg_mem [25] ), .ZN(_01920_ ) );
NOR4_X1 _09498_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\EX_LS_dest_csreg_mem [29] ), .A4(\EX_LS_dest_csreg_mem [28] ), .ZN(_01921_ ) );
AND2_X1 _09499_ ( .A1(_01920_ ), .A2(_01921_ ), .ZN(_01922_ ) );
AND2_X1 _09500_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_01923_ ) );
INV_X1 _09501_ ( .A(\EX_LS_flag [2] ), .ZN(_01924_ ) );
AND2_X1 _09502_ ( .A1(_01923_ ), .A2(_01924_ ), .ZN(_01925_ ) );
AND2_X1 _09503_ ( .A1(_01922_ ), .A2(_01925_ ), .ZN(_01926_ ) );
INV_X1 _09504_ ( .A(_01926_ ), .ZN(_01927_ ) );
INV_X1 _09505_ ( .A(\EX_LS_typ [4] ), .ZN(_01928_ ) );
AND2_X1 _09506_ ( .A1(_01925_ ), .A2(_01928_ ), .ZN(_01929_ ) );
NOR2_X1 _09507_ ( .A1(fanout_net_3 ), .A2(fanout_net_4 ), .ZN(_01930_ ) );
INV_X1 _09508_ ( .A(_01930_ ), .ZN(_01931_ ) );
INV_X1 _09509_ ( .A(\EX_LS_typ [1] ), .ZN(_01932_ ) );
INV_X1 _09510_ ( .A(\EX_LS_typ [3] ), .ZN(_01933_ ) );
NAND4_X1 _09511_ ( .A1(_01931_ ), .A2(_01932_ ), .A3(_01933_ ), .A4(\EX_LS_typ [2] ), .ZN(_01934_ ) );
AND2_X1 _09512_ ( .A1(fanout_net_3 ), .A2(\EX_LS_typ [1] ), .ZN(_01935_ ) );
NOR2_X1 _09513_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_01936_ ) );
NAND2_X1 _09514_ ( .A1(_01935_ ), .A2(_01936_ ), .ZN(_01937_ ) );
AOI21_X1 _09515_ ( .A(\EX_LS_typ [0] ), .B1(_01934_ ), .B2(_01937_ ), .ZN(_01938_ ) );
AND3_X1 _09516_ ( .A1(_01935_ ), .A2(\EX_LS_typ [0] ), .A3(_01936_ ), .ZN(_01939_ ) );
OAI21_X1 _09517_ ( .A(_01929_ ), .B1(_01938_ ), .B2(_01939_ ), .ZN(_01940_ ) );
AND2_X2 _09518_ ( .A1(_01927_ ), .A2(_01940_ ), .ZN(_01941_ ) );
NOR2_X4 _09519_ ( .A1(_01870_ ), .A2(\EX_LS_flag [0] ), .ZN(_01942_ ) );
BUF_X2 _09520_ ( .A(_01942_ ), .Z(_01943_ ) );
AND2_X1 _09521_ ( .A1(_01943_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_01944_ ) );
AND2_X1 _09522_ ( .A1(_01922_ ), .A2(_01944_ ), .ZN(_01945_ ) );
NAND3_X1 _09523_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_01946_ ) );
OAI21_X1 _09524_ ( .A(_01937_ ), .B1(_01930_ ), .B2(_01946_ ), .ZN(_01947_ ) );
NAND3_X1 _09525_ ( .A1(_01924_ ), .A2(_01928_ ), .A3(\EX_LS_typ [0] ), .ZN(_01948_ ) );
NOR3_X1 _09526_ ( .A1(_01948_ ), .A2(_01870_ ), .A3(\EX_LS_flag [0] ), .ZN(_01949_ ) );
AND2_X1 _09527_ ( .A1(_01947_ ), .A2(_01949_ ), .ZN(_01950_ ) );
NOR2_X1 _09528_ ( .A1(_01945_ ), .A2(_01950_ ), .ZN(_01951_ ) );
AND2_X1 _09529_ ( .A1(_01941_ ), .A2(_01951_ ), .ZN(_01952_ ) );
AOI21_X1 _09530_ ( .A(_01918_ ), .B1(_01888_ ), .B2(_01952_ ), .ZN(_01953_ ) );
OR3_X1 _09531_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(_01886_ ), .ZN(_01954_ ) );
OAI211_X1 _09532_ ( .A(_01878_ ), .B(_01954_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01881_ ), .ZN(_01955_ ) );
OAI221_X1 _09533_ ( .A(\IF_ID_pc [28] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01890_ ), .C2(_01891_ ), .ZN(_01956_ ) );
AND2_X1 _09534_ ( .A1(_01955_ ), .A2(_01956_ ), .ZN(_01957_ ) );
OR3_X1 _09535_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(_01886_ ), .ZN(_01958_ ) );
OAI211_X1 _09536_ ( .A(_01878_ ), .B(_01958_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01881_ ), .ZN(_01959_ ) );
OAI221_X1 _09537_ ( .A(\IF_ID_pc [26] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01890_ ), .C2(_01891_ ), .ZN(_01960_ ) );
AND2_X1 _09538_ ( .A1(_01959_ ), .A2(_01960_ ), .ZN(_01961_ ) );
OR3_X1 _09539_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(_01873_ ), .ZN(_01962_ ) );
OAI211_X1 _09540_ ( .A(_01877_ ), .B(_01962_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01881_ ), .ZN(_01963_ ) );
OAI221_X1 _09541_ ( .A(\IF_ID_pc [21] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01865_ ), .C2(_01866_ ), .ZN(_01964_ ) );
AND2_X1 _09542_ ( .A1(_01963_ ), .A2(_01964_ ), .ZN(_01965_ ) );
OR3_X1 _09543_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(_01873_ ), .ZN(_01966_ ) );
OAI211_X1 _09544_ ( .A(_01877_ ), .B(_01966_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01874_ ), .ZN(_01967_ ) );
OAI221_X1 _09545_ ( .A(\IF_ID_pc [19] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01865_ ), .C2(_01866_ ), .ZN(_01968_ ) );
AND2_X1 _09546_ ( .A1(_01967_ ), .A2(_01968_ ), .ZN(_01969_ ) );
AND4_X1 _09547_ ( .A1(_01957_ ), .A2(_01961_ ), .A3(_01965_ ), .A4(_01969_ ), .ZN(_01970_ ) );
OR3_X1 _09548_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(_01886_ ), .ZN(_01971_ ) );
OAI211_X1 _09549_ ( .A(_01878_ ), .B(_01971_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01881_ ), .ZN(_01972_ ) );
OAI221_X1 _09550_ ( .A(\IF_ID_pc [29] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01890_ ), .C2(_01891_ ), .ZN(_01973_ ) );
AND2_X1 _09551_ ( .A1(_01972_ ), .A2(_01973_ ), .ZN(_01974_ ) );
OR3_X1 _09552_ ( .A1(_01879_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(_01886_ ), .ZN(_01975_ ) );
OAI211_X1 _09553_ ( .A(_01878_ ), .B(_01975_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01881_ ), .ZN(_01976_ ) );
OAI221_X1 _09554_ ( .A(\IF_ID_pc [27] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01865_ ), .C2(_01891_ ), .ZN(_01977_ ) );
AND2_X1 _09555_ ( .A1(_01976_ ), .A2(_01977_ ), .ZN(_01978_ ) );
OR3_X1 _09556_ ( .A1(_01872_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(_01873_ ), .ZN(_01979_ ) );
OAI211_X1 _09557_ ( .A(_01877_ ), .B(_01979_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01874_ ), .ZN(_01980_ ) );
OAI221_X1 _09558_ ( .A(\IF_ID_pc [22] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01865_ ), .C2(_01866_ ), .ZN(_01981_ ) );
AND2_X1 _09559_ ( .A1(_01980_ ), .A2(_01981_ ), .ZN(_01982_ ) );
OR3_X1 _09560_ ( .A1(_01872_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(_01873_ ), .ZN(_01983_ ) );
OAI211_X1 _09561_ ( .A(_01877_ ), .B(_01983_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01874_ ), .ZN(_01984_ ) );
OAI221_X1 _09562_ ( .A(\IF_ID_pc [16] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01865_ ), .C2(_01866_ ), .ZN(_01985_ ) );
AND2_X1 _09563_ ( .A1(_01984_ ), .A2(_01985_ ), .ZN(_01986_ ) );
AND4_X1 _09564_ ( .A1(_01974_ ), .A2(_01978_ ), .A3(_01982_ ), .A4(_01986_ ), .ZN(_01987_ ) );
NAND2_X1 _09565_ ( .A1(_01970_ ), .A2(_01987_ ), .ZN(_01988_ ) );
NOR2_X1 _09566_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_01989_ ) );
AOI211_X1 _09567_ ( .A(_01868_ ), .B(_01867_ ), .C1(\myifu.state [0] ), .C2(_01989_ ), .ZN(_01990_ ) );
NOR4_X1 _09568_ ( .A1(_01914_ ), .A2(_01953_ ), .A3(_01988_ ), .A4(_01990_ ), .ZN(_01991_ ) );
OAI21_X1 _09569_ ( .A(_01459_ ), .B1(_01991_ ), .B2(\myclint.rvalid ), .ZN(_01992_ ) );
BUF_X4 _09570_ ( .A(_01883_ ), .Z(_01993_ ) );
AOI211_X1 _09571_ ( .A(_01891_ ), .B(_01993_ ), .C1(_01890_ ), .C2(_01989_ ), .ZN(_01994_ ) );
AOI211_X1 _09572_ ( .A(_01875_ ), .B(_01918_ ), .C1(_01888_ ), .C2(_01952_ ), .ZN(_01995_ ) );
NOR2_X1 _09573_ ( .A1(_01994_ ), .A2(_01995_ ), .ZN(_01996_ ) );
NAND4_X1 _09574_ ( .A1(_01893_ ), .A2(_01974_ ), .A3(_01978_ ), .A4(\io_master_araddr [25] ), .ZN(_01997_ ) );
NOR4_X1 _09575_ ( .A1(_01997_ ), .A2(_01910_ ), .A3(\io_master_araddr [23] ), .A4(\io_master_araddr [20] ), .ZN(_01998_ ) );
NAND4_X1 _09576_ ( .A1(_01897_ ), .A2(_01901_ ), .A3(_01957_ ), .A4(_01961_ ), .ZN(_01999_ ) );
NAND4_X1 _09577_ ( .A1(_01965_ ), .A2(_01969_ ), .A3(_01982_ ), .A4(_01986_ ), .ZN(_02000_ ) );
NOR2_X1 _09578_ ( .A1(_01999_ ), .A2(_02000_ ), .ZN(_02001_ ) );
AND3_X1 _09579_ ( .A1(_01998_ ), .A2(\myclint.rvalid ), .A3(_02001_ ), .ZN(_02002_ ) );
AOI21_X1 _09580_ ( .A(_01992_ ), .B1(_01996_ ), .B2(_02002_ ), .ZN(_00064_ ) );
INV_X1 _09581_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02003_ ) );
CLKBUF_X2 _09582_ ( .A(_02003_ ), .Z(_02004_ ) );
AND2_X1 _09583_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00065_ ) );
AND2_X1 _09584_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00066_ ) );
AND2_X1 _09585_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00067_ ) );
AND2_X1 _09586_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [20] ), .ZN(_00068_ ) );
INV_X1 _09587_ ( .A(\LS_WB_wdata_csreg [19] ), .ZN(_02005_ ) );
NOR2_X1 _09588_ ( .A1(_02005_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00069_ ) );
AND2_X1 _09589_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [18] ), .ZN(_00070_ ) );
INV_X1 _09590_ ( .A(\LS_WB_wdata_csreg [17] ), .ZN(_02006_ ) );
NOR2_X1 _09591_ ( .A1(_02006_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00071_ ) );
AND2_X1 _09592_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00072_ ) );
AND2_X1 _09593_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00073_ ) );
AND2_X1 _09594_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00074_ ) );
INV_X1 _09595_ ( .A(\LS_WB_wdata_csreg [13] ), .ZN(_02007_ ) );
NOR2_X1 _09596_ ( .A1(_02007_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00075_ ) );
AND2_X1 _09597_ ( .A1(_02004_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00076_ ) );
CLKBUF_X2 _09598_ ( .A(_02003_ ), .Z(_02008_ ) );
AND2_X1 _09599_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00077_ ) );
AND2_X1 _09600_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00078_ ) );
AND2_X1 _09601_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00079_ ) );
AND2_X1 _09602_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00080_ ) );
AND2_X1 _09603_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00081_ ) );
AND2_X1 _09604_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00082_ ) );
AND2_X1 _09605_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [6] ), .ZN(_00083_ ) );
AND2_X1 _09606_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00084_ ) );
AND2_X1 _09607_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [4] ), .ZN(_00085_ ) );
AND2_X1 _09608_ ( .A1(_02008_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00086_ ) );
AND2_X1 _09609_ ( .A1(_02003_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00087_ ) );
AND2_X1 _09610_ ( .A1(_02003_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00088_ ) );
AND2_X1 _09611_ ( .A1(_02003_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00089_ ) );
AND2_X1 _09612_ ( .A1(_02003_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00090_ ) );
AND2_X1 _09613_ ( .A1(_02003_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00091_ ) );
AND2_X1 _09614_ ( .A1(_02003_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00092_ ) );
AOI21_X1 _09615_ ( .A(excp_written ), .B1(\LS_WB_wen_csreg [6] ), .B2(\LS_WB_wen_csreg [7] ), .ZN(_02009_ ) );
NOR2_X1 _09616_ ( .A1(_02009_ ), .A2(fanout_net_2 ), .ZN(_00093_ ) );
OR2_X1 _09617_ ( .A1(\myexu.pc_jump [25] ), .A2(\myexu.pc_jump [24] ), .ZN(_02010_ ) );
NOR3_X1 _09618_ ( .A1(_02010_ ), .A2(\myexu.pc_jump [27] ), .A3(\myexu.pc_jump [26] ), .ZN(_02011_ ) );
NOR4_X1 _09619_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02012_ ) );
AND2_X1 _09620_ ( .A1(_02011_ ), .A2(_02012_ ), .ZN(_02013_ ) );
NOR2_X1 _09621_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02014_ ) );
INV_X1 _09622_ ( .A(_02014_ ), .ZN(_02015_ ) );
OR3_X1 _09623_ ( .A1(_02013_ ), .A2(exception_quest_IDU ), .A3(_02015_ ), .ZN(_02016_ ) );
NOR2_X1 _09624_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02017_ ) );
AND2_X1 _09625_ ( .A1(_02017_ ), .A2(_01458_ ), .ZN(_02018_ ) );
AND4_X1 _09626_ ( .A1(_01951_ ), .A2(_01941_ ), .A3(_02016_ ), .A4(_02018_ ), .ZN(_00094_ ) );
INV_X1 _09627_ ( .A(_02018_ ), .ZN(_02019_ ) );
AOI21_X1 _09628_ ( .A(_02019_ ), .B1(_01952_ ), .B2(exception_quest_IDU ), .ZN(_00095_ ) );
INV_X32 _09629_ ( .A(\EX_LS_dest_reg [4] ), .ZN(_02020_ ) );
INV_X4 _09630_ ( .A(\ID_EX_rs1 [2] ), .ZN(_02021_ ) );
AOI22_X1 _09631_ ( .A1(\ID_EX_rs1 [4] ), .A2(_02020_ ), .B1(_02021_ ), .B2(\EX_LS_dest_reg [2] ), .ZN(_02022_ ) );
INV_X1 _09632_ ( .A(\ID_EX_rs1 [3] ), .ZN(_02023_ ) );
OAI221_X1 _09633_ ( .A(_02022_ ), .B1(\ID_EX_rs1 [4] ), .B2(_02020_ ), .C1(_02023_ ), .C2(\EX_LS_dest_reg [3] ), .ZN(_02024_ ) );
XOR2_X1 _09634_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .Z(_02025_ ) );
INV_X1 _09635_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .ZN(_02026_ ) );
NOR2_X1 _09636_ ( .A1(_02021_ ), .A2(\EX_LS_dest_reg [2] ), .ZN(_02027_ ) );
NOR4_X1 _09637_ ( .A1(_02024_ ), .A2(_02025_ ), .A3(_02026_ ), .A4(_02027_ ), .ZN(_02028_ ) );
NOR4_X1 _09638_ ( .A1(\EX_LS_dest_reg [3] ), .A2(\EX_LS_dest_reg [2] ), .A3(\EX_LS_dest_reg [1] ), .A4(\EX_LS_dest_reg [0] ), .ZN(_02029_ ) );
NAND2_X1 _09639_ ( .A1(_02029_ ), .A2(_02020_ ), .ZN(_02030_ ) );
INV_X1 _09640_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02031_ ) );
NAND2_X1 _09641_ ( .A1(_02031_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02032_ ) );
NOR2_X1 _09642_ ( .A1(_02031_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02033_ ) );
AOI21_X1 _09643_ ( .A(_02033_ ), .B1(_02023_ ), .B2(\EX_LS_dest_reg [3] ), .ZN(_02034_ ) );
NAND4_X1 _09644_ ( .A1(_02028_ ), .A2(_02030_ ), .A3(_02032_ ), .A4(_02034_ ), .ZN(_02035_ ) );
CLKBUF_X2 _09645_ ( .A(_02035_ ), .Z(_02036_ ) );
CLKBUF_X2 _09646_ ( .A(_02036_ ), .Z(_02037_ ) );
AND2_X2 _09647_ ( .A1(_01942_ ), .A2(\EX_LS_flag [2] ), .ZN(_02038_ ) );
BUF_X4 _09648_ ( .A(_02038_ ), .Z(_02039_ ) );
NOR2_X2 _09649_ ( .A1(_02039_ ), .A2(_01925_ ), .ZN(_02040_ ) );
OAI211_X1 _09650_ ( .A(_01870_ ), .B(\EX_LS_flag [0] ), .C1(\EX_LS_flag [2] ), .C2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02041_ ) );
AND2_X2 _09651_ ( .A1(_02040_ ), .A2(_02041_ ), .ZN(_02042_ ) );
BUF_X8 _09652_ ( .A(_02042_ ), .Z(_02043_ ) );
CLKBUF_X2 _09653_ ( .A(_02043_ ), .Z(_02044_ ) );
BUF_X2 _09654_ ( .A(_02044_ ), .Z(_02045_ ) );
OR3_X1 _09655_ ( .A1(_02037_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02045_ ), .ZN(_02046_ ) );
INV_X1 _09656_ ( .A(fanout_net_28 ), .ZN(_02047_ ) );
BUF_X4 _09657_ ( .A(_02047_ ), .Z(_02048_ ) );
BUF_X4 _09658_ ( .A(_02048_ ), .Z(_02049_ ) );
BUF_X4 _09659_ ( .A(_02049_ ), .Z(_02050_ ) );
INV_X1 _09660_ ( .A(fanout_net_27 ), .ZN(_02051_ ) );
BUF_X4 _09661_ ( .A(_02051_ ), .Z(_02052_ ) );
BUF_X4 _09662_ ( .A(_02052_ ), .Z(_02053_ ) );
BUF_X4 _09663_ ( .A(_02053_ ), .Z(_02054_ ) );
BUF_X4 _09664_ ( .A(_02054_ ), .Z(_02055_ ) );
INV_X1 _09665_ ( .A(fanout_net_16 ), .ZN(_02056_ ) );
CLKBUF_X2 _09666_ ( .A(_02056_ ), .Z(_02057_ ) );
BUF_X2 _09667_ ( .A(_02057_ ), .Z(_02058_ ) );
BUF_X4 _09668_ ( .A(_02058_ ), .Z(_02059_ ) );
BUF_X2 _09669_ ( .A(_02059_ ), .Z(_02060_ ) );
OAI21_X1 _09670_ ( .A(fanout_net_25 ), .B1(_02060_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02061_ ) );
NOR2_X1 _09671_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02062_ ) );
NOR2_X1 _09672_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02063_ ) );
INV_X2 _09673_ ( .A(fanout_net_25 ), .ZN(_02064_ ) );
BUF_X4 _09674_ ( .A(_02064_ ), .Z(_02065_ ) );
BUF_X4 _09675_ ( .A(_02065_ ), .Z(_02066_ ) );
BUF_X4 _09676_ ( .A(_02066_ ), .Z(_02067_ ) );
BUF_X4 _09677_ ( .A(_02067_ ), .Z(_02068_ ) );
OAI21_X1 _09678_ ( .A(_02068_ ), .B1(_02060_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02069_ ) );
OAI221_X1 _09679_ ( .A(_02055_ ), .B1(_02061_ ), .B2(_02062_ ), .C1(_02063_ ), .C2(_02069_ ), .ZN(_02070_ ) );
MUX2_X1 _09680_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02071_ ) );
MUX2_X1 _09681_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02072_ ) );
MUX2_X1 _09682_ ( .A(_02071_ ), .B(_02072_ ), .S(fanout_net_25 ), .Z(_02073_ ) );
BUF_X4 _09683_ ( .A(_02055_ ), .Z(_02074_ ) );
OAI211_X1 _09684_ ( .A(_02050_ ), .B(_02070_ ), .C1(_02073_ ), .C2(_02074_ ), .ZN(_02075_ ) );
NOR2_X1 _09685_ ( .A1(_02060_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02076_ ) );
OAI21_X1 _09686_ ( .A(fanout_net_25 ), .B1(fanout_net_16 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02077_ ) );
NOR2_X1 _09687_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02078_ ) );
OAI21_X1 _09688_ ( .A(_02068_ ), .B1(_02060_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02079_ ) );
OAI221_X1 _09689_ ( .A(fanout_net_27 ), .B1(_02076_ ), .B2(_02077_ ), .C1(_02078_ ), .C2(_02079_ ), .ZN(_02080_ ) );
MUX2_X1 _09690_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02081_ ) );
MUX2_X1 _09691_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02082_ ) );
MUX2_X1 _09692_ ( .A(_02081_ ), .B(_02082_ ), .S(_02068_ ), .Z(_02083_ ) );
OAI211_X1 _09693_ ( .A(fanout_net_28 ), .B(_02080_ ), .C1(_02083_ ), .C2(fanout_net_27 ), .ZN(_02084_ ) );
BUF_X2 _09694_ ( .A(_02035_ ), .Z(_02085_ ) );
BUF_X2 _09695_ ( .A(_02085_ ), .Z(_02086_ ) );
BUF_X2 _09696_ ( .A(_02086_ ), .Z(_02087_ ) );
BUF_X2 _09697_ ( .A(_02045_ ), .Z(_02088_ ) );
OAI211_X1 _09698_ ( .A(_02075_ ), .B(_02084_ ), .C1(_02087_ ), .C2(_02088_ ), .ZN(_02089_ ) );
AND2_X2 _09699_ ( .A1(_02046_ ), .A2(_02089_ ), .ZN(_02090_ ) );
XOR2_X1 _09700_ ( .A(_02090_ ), .B(\ID_EX_imm [30] ), .Z(_02091_ ) );
INV_X1 _09701_ ( .A(_02091_ ), .ZN(_02092_ ) );
BUF_X4 _09702_ ( .A(_02043_ ), .Z(_02093_ ) );
BUF_X2 _09703_ ( .A(_02093_ ), .Z(_02094_ ) );
CLKBUF_X3 _09704_ ( .A(_02094_ ), .Z(_02095_ ) );
OR3_X1 _09705_ ( .A1(_02037_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02095_ ), .ZN(_02096_ ) );
INV_X1 _09706_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02097_ ) );
NAND2_X1 _09707_ ( .A1(_02097_ ), .A2(fanout_net_16 ), .ZN(_02098_ ) );
BUF_X4 _09708_ ( .A(_02066_ ), .Z(_02099_ ) );
BUF_X4 _09709_ ( .A(_02099_ ), .Z(_02100_ ) );
OAI211_X1 _09710_ ( .A(_02098_ ), .B(_02100_ ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02101_ ) );
INV_X1 _09711_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02102_ ) );
NAND2_X1 _09712_ ( .A1(_02102_ ), .A2(fanout_net_16 ), .ZN(_02103_ ) );
OAI211_X1 _09713_ ( .A(_02103_ ), .B(fanout_net_25 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02104_ ) );
BUF_X4 _09714_ ( .A(_02052_ ), .Z(_02105_ ) );
BUF_X4 _09715_ ( .A(_02105_ ), .Z(_02106_ ) );
BUF_X4 _09716_ ( .A(_02106_ ), .Z(_02107_ ) );
NAND3_X1 _09717_ ( .A1(_02101_ ), .A2(_02104_ ), .A3(_02107_ ), .ZN(_02108_ ) );
MUX2_X1 _09718_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02109_ ) );
MUX2_X1 _09719_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02110_ ) );
MUX2_X1 _09720_ ( .A(_02109_ ), .B(_02110_ ), .S(_02068_ ), .Z(_02111_ ) );
OAI211_X1 _09721_ ( .A(fanout_net_28 ), .B(_02108_ ), .C1(_02111_ ), .C2(_02074_ ), .ZN(_02112_ ) );
INV_X1 _09722_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02113_ ) );
NAND2_X1 _09723_ ( .A1(_02113_ ), .A2(fanout_net_16 ), .ZN(_02114_ ) );
OAI211_X1 _09724_ ( .A(_02114_ ), .B(_02100_ ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02115_ ) );
INV_X1 _09725_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02116_ ) );
NAND2_X1 _09726_ ( .A1(_02116_ ), .A2(fanout_net_16 ), .ZN(_02117_ ) );
OAI211_X1 _09727_ ( .A(_02117_ ), .B(fanout_net_25 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02118_ ) );
NAND3_X1 _09728_ ( .A1(_02115_ ), .A2(_02118_ ), .A3(_02055_ ), .ZN(_02119_ ) );
MUX2_X1 _09729_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02120_ ) );
MUX2_X1 _09730_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02121_ ) );
MUX2_X1 _09731_ ( .A(_02120_ ), .B(_02121_ ), .S(_02068_ ), .Z(_02122_ ) );
OAI211_X1 _09732_ ( .A(_02050_ ), .B(_02119_ ), .C1(_02122_ ), .C2(_02074_ ), .ZN(_02123_ ) );
OAI211_X1 _09733_ ( .A(_02112_ ), .B(_02123_ ), .C1(_02087_ ), .C2(_02088_ ), .ZN(_02124_ ) );
NAND2_X1 _09734_ ( .A1(_02096_ ), .A2(_02124_ ), .ZN(_02125_ ) );
XNOR2_X1 _09735_ ( .A(_02125_ ), .B(\ID_EX_imm [28] ), .ZN(_02126_ ) );
BUF_X2 _09736_ ( .A(_02043_ ), .Z(_02127_ ) );
BUF_X2 _09737_ ( .A(_02127_ ), .Z(_02128_ ) );
OR3_X1 _09738_ ( .A1(_02086_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02128_ ), .ZN(_02129_ ) );
BUF_X2 _09739_ ( .A(_02056_ ), .Z(_02130_ ) );
BUF_X2 _09740_ ( .A(_02130_ ), .Z(_02131_ ) );
BUF_X2 _09741_ ( .A(_02131_ ), .Z(_02132_ ) );
OR2_X1 _09742_ ( .A1(_02132_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02133_ ) );
OAI211_X1 _09743_ ( .A(_02133_ ), .B(fanout_net_25 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02134_ ) );
OR2_X1 _09744_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02135_ ) );
BUF_X2 _09745_ ( .A(_02057_ ), .Z(_02136_ ) );
BUF_X2 _09746_ ( .A(_02136_ ), .Z(_02137_ ) );
OAI211_X1 _09747_ ( .A(_02135_ ), .B(_02099_ ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02138_ ) );
NAND3_X1 _09748_ ( .A1(_02134_ ), .A2(_02106_ ), .A3(_02138_ ), .ZN(_02139_ ) );
MUX2_X1 _09749_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02140_ ) );
MUX2_X1 _09750_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02141_ ) );
MUX2_X1 _09751_ ( .A(_02140_ ), .B(_02141_ ), .S(_02067_ ), .Z(_02142_ ) );
OAI211_X1 _09752_ ( .A(_02049_ ), .B(_02139_ ), .C1(_02142_ ), .C2(_02055_ ), .ZN(_02143_ ) );
OR2_X1 _09753_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02144_ ) );
BUF_X2 _09754_ ( .A(_02132_ ), .Z(_02145_ ) );
OAI211_X1 _09755_ ( .A(_02144_ ), .B(fanout_net_25 ), .C1(_02145_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02146_ ) );
OR2_X1 _09756_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02147_ ) );
OAI211_X1 _09757_ ( .A(_02147_ ), .B(_02099_ ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02148_ ) );
NAND3_X1 _09758_ ( .A1(_02146_ ), .A2(_02148_ ), .A3(fanout_net_27 ), .ZN(_02149_ ) );
MUX2_X1 _09759_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02150_ ) );
MUX2_X1 _09760_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02151_ ) );
MUX2_X1 _09761_ ( .A(_02150_ ), .B(_02151_ ), .S(fanout_net_25 ), .Z(_02152_ ) );
OAI211_X1 _09762_ ( .A(fanout_net_28 ), .B(_02149_ ), .C1(_02152_ ), .C2(fanout_net_27 ), .ZN(_02153_ ) );
OAI211_X1 _09763_ ( .A(_02143_ ), .B(_02153_ ), .C1(_02037_ ), .C2(_02045_ ), .ZN(_02154_ ) );
NAND2_X1 _09764_ ( .A1(_02129_ ), .A2(_02154_ ), .ZN(_02155_ ) );
XOR2_X1 _09765_ ( .A(_02155_ ), .B(\ID_EX_imm [22] ), .Z(_02156_ ) );
OR3_X1 _09766_ ( .A1(_02086_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02128_ ), .ZN(_02157_ ) );
OR2_X1 _09767_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02158_ ) );
OAI211_X1 _09768_ ( .A(_02158_ ), .B(_02099_ ), .C1(_02145_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02159_ ) );
OR2_X1 _09769_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02160_ ) );
OAI211_X1 _09770_ ( .A(_02160_ ), .B(fanout_net_25 ), .C1(_02145_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02161_ ) );
NAND3_X1 _09771_ ( .A1(_02159_ ), .A2(_02161_ ), .A3(_02106_ ), .ZN(_02162_ ) );
MUX2_X1 _09772_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02163_ ) );
MUX2_X1 _09773_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02164_ ) );
MUX2_X1 _09774_ ( .A(_02163_ ), .B(_02164_ ), .S(_02067_ ), .Z(_02165_ ) );
OAI211_X1 _09775_ ( .A(fanout_net_28 ), .B(_02162_ ), .C1(_02165_ ), .C2(_02055_ ), .ZN(_02166_ ) );
OR2_X1 _09776_ ( .A1(_02132_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02167_ ) );
OAI211_X1 _09777_ ( .A(_02167_ ), .B(_02099_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02168_ ) );
OR2_X1 _09778_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02169_ ) );
OAI211_X1 _09779_ ( .A(_02169_ ), .B(fanout_net_25 ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02170_ ) );
NAND3_X1 _09780_ ( .A1(_02168_ ), .A2(_02106_ ), .A3(_02170_ ), .ZN(_02171_ ) );
MUX2_X1 _09781_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02172_ ) );
MUX2_X1 _09782_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02173_ ) );
MUX2_X1 _09783_ ( .A(_02172_ ), .B(_02173_ ), .S(_02067_ ), .Z(_02174_ ) );
OAI211_X1 _09784_ ( .A(_02050_ ), .B(_02171_ ), .C1(_02174_ ), .C2(_02055_ ), .ZN(_02175_ ) );
OAI211_X1 _09785_ ( .A(_02166_ ), .B(_02175_ ), .C1(_02037_ ), .C2(_02045_ ), .ZN(_02176_ ) );
INV_X1 _09786_ ( .A(\ID_EX_imm [23] ), .ZN(_02177_ ) );
NAND3_X1 _09787_ ( .A1(_02157_ ), .A2(_02176_ ), .A3(_02177_ ), .ZN(_02178_ ) );
NAND2_X1 _09788_ ( .A1(_02157_ ), .A2(_02176_ ), .ZN(_02179_ ) );
NAND2_X1 _09789_ ( .A1(_02179_ ), .A2(\ID_EX_imm [23] ), .ZN(_02180_ ) );
AND3_X1 _09790_ ( .A1(_02156_ ), .A2(_02178_ ), .A3(_02180_ ), .ZN(_02181_ ) );
OR3_X1 _09791_ ( .A1(_02037_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02045_ ), .ZN(_02182_ ) );
OR2_X1 _09792_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02183_ ) );
OAI211_X1 _09793_ ( .A(_02183_ ), .B(_02100_ ), .C1(_02060_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02184_ ) );
OR2_X1 _09794_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02185_ ) );
OAI211_X1 _09795_ ( .A(_02185_ ), .B(fanout_net_25 ), .C1(_02060_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02186_ ) );
NAND3_X1 _09796_ ( .A1(_02184_ ), .A2(_02186_ ), .A3(_02055_ ), .ZN(_02187_ ) );
MUX2_X1 _09797_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02188_ ) );
MUX2_X1 _09798_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02189_ ) );
MUX2_X1 _09799_ ( .A(_02188_ ), .B(_02189_ ), .S(_02068_ ), .Z(_02190_ ) );
OAI211_X1 _09800_ ( .A(fanout_net_28 ), .B(_02187_ ), .C1(_02190_ ), .C2(_02107_ ), .ZN(_02191_ ) );
OR2_X1 _09801_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02192_ ) );
OAI211_X1 _09802_ ( .A(_02192_ ), .B(_02068_ ), .C1(_02060_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02193_ ) );
OR2_X1 _09803_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02194_ ) );
OAI211_X1 _09804_ ( .A(_02194_ ), .B(fanout_net_25 ), .C1(_02060_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02195_ ) );
NAND3_X1 _09805_ ( .A1(_02193_ ), .A2(_02195_ ), .A3(_02055_ ), .ZN(_02196_ ) );
MUX2_X1 _09806_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02197_ ) );
MUX2_X1 _09807_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02198_ ) );
MUX2_X1 _09808_ ( .A(_02197_ ), .B(_02198_ ), .S(_02068_ ), .Z(_02199_ ) );
OAI211_X1 _09809_ ( .A(_02050_ ), .B(_02196_ ), .C1(_02199_ ), .C2(_02107_ ), .ZN(_02200_ ) );
OAI211_X1 _09810_ ( .A(_02191_ ), .B(_02200_ ), .C1(_02087_ ), .C2(_02088_ ), .ZN(_02201_ ) );
NAND2_X1 _09811_ ( .A1(_02182_ ), .A2(_02201_ ), .ZN(_02202_ ) );
INV_X1 _09812_ ( .A(\ID_EX_imm [20] ), .ZN(_02203_ ) );
XNOR2_X1 _09813_ ( .A(_02202_ ), .B(_02203_ ), .ZN(_02204_ ) );
OR3_X1 _09814_ ( .A1(_02036_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02094_ ), .ZN(_02205_ ) );
INV_X1 _09815_ ( .A(\ID_EX_imm [21] ), .ZN(_02206_ ) );
OR2_X1 _09816_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02207_ ) );
OAI211_X1 _09817_ ( .A(_02207_ ), .B(_02067_ ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02208_ ) );
OR2_X1 _09818_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02209_ ) );
OAI211_X1 _09819_ ( .A(_02209_ ), .B(fanout_net_25 ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02210_ ) );
NAND3_X1 _09820_ ( .A1(_02208_ ), .A2(_02210_ ), .A3(_02054_ ), .ZN(_02211_ ) );
MUX2_X1 _09821_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02212_ ) );
MUX2_X1 _09822_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02213_ ) );
BUF_X4 _09823_ ( .A(_02065_ ), .Z(_02214_ ) );
BUF_X4 _09824_ ( .A(_02214_ ), .Z(_02215_ ) );
MUX2_X1 _09825_ ( .A(_02212_ ), .B(_02213_ ), .S(_02215_ ), .Z(_02216_ ) );
OAI211_X1 _09826_ ( .A(_02049_ ), .B(_02211_ ), .C1(_02216_ ), .C2(_02106_ ), .ZN(_02217_ ) );
OR2_X1 _09827_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02218_ ) );
OAI211_X1 _09828_ ( .A(_02218_ ), .B(fanout_net_25 ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02219_ ) );
OR2_X1 _09829_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02220_ ) );
OAI211_X1 _09830_ ( .A(_02220_ ), .B(_02067_ ), .C1(_02059_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02221_ ) );
NAND3_X1 _09831_ ( .A1(_02219_ ), .A2(_02221_ ), .A3(fanout_net_27 ), .ZN(_02222_ ) );
MUX2_X1 _09832_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02223_ ) );
MUX2_X1 _09833_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02224_ ) );
MUX2_X1 _09834_ ( .A(_02223_ ), .B(_02224_ ), .S(fanout_net_25 ), .Z(_02225_ ) );
OAI211_X1 _09835_ ( .A(fanout_net_28 ), .B(_02222_ ), .C1(_02225_ ), .C2(fanout_net_27 ), .ZN(_02226_ ) );
OAI211_X1 _09836_ ( .A(_02217_ ), .B(_02226_ ), .C1(_02086_ ), .C2(_02128_ ), .ZN(_02227_ ) );
AND3_X1 _09837_ ( .A1(_02205_ ), .A2(_02206_ ), .A3(_02227_ ), .ZN(_02228_ ) );
AOI21_X1 _09838_ ( .A(_02206_ ), .B1(_02205_ ), .B2(_02227_ ), .ZN(_02229_ ) );
NOR2_X1 _09839_ ( .A1(_02228_ ), .A2(_02229_ ), .ZN(_02230_ ) );
AND2_X1 _09840_ ( .A1(_02204_ ), .A2(_02230_ ), .ZN(_02231_ ) );
NAND2_X1 _09841_ ( .A1(_02181_ ), .A2(_02231_ ), .ZN(_02232_ ) );
OR2_X1 _09842_ ( .A1(_02132_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02233_ ) );
OAI211_X1 _09843_ ( .A(_02233_ ), .B(fanout_net_25 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02234_ ) );
OR2_X1 _09844_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02235_ ) );
OAI211_X1 _09845_ ( .A(_02235_ ), .B(_02099_ ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02236_ ) );
NAND3_X1 _09846_ ( .A1(_02234_ ), .A2(_02054_ ), .A3(_02236_ ), .ZN(_02237_ ) );
MUX2_X1 _09847_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02238_ ) );
MUX2_X1 _09848_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02239_ ) );
MUX2_X1 _09849_ ( .A(_02238_ ), .B(_02239_ ), .S(_02067_ ), .Z(_02240_ ) );
OAI211_X1 _09850_ ( .A(fanout_net_28 ), .B(_02237_ ), .C1(_02240_ ), .C2(_02106_ ), .ZN(_02241_ ) );
MUX2_X1 _09851_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02242_ ) );
AND2_X1 _09852_ ( .A1(_02242_ ), .A2(_02215_ ), .ZN(_02243_ ) );
MUX2_X1 _09853_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02244_ ) );
AOI211_X1 _09854_ ( .A(fanout_net_27 ), .B(_02243_ ), .C1(fanout_net_25 ), .C2(_02244_ ), .ZN(_02245_ ) );
MUX2_X1 _09855_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02246_ ) );
MUX2_X1 _09856_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02247_ ) );
MUX2_X1 _09857_ ( .A(_02246_ ), .B(_02247_ ), .S(_02215_ ), .Z(_02248_ ) );
OAI21_X1 _09858_ ( .A(_02049_ ), .B1(_02248_ ), .B2(_02106_ ), .ZN(_02249_ ) );
OAI221_X1 _09859_ ( .A(_02241_ ), .B1(_02245_ ), .B2(_02249_ ), .C1(_02086_ ), .C2(_02045_ ), .ZN(_02250_ ) );
OR3_X1 _09860_ ( .A1(_02086_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02128_ ), .ZN(_02251_ ) );
NAND2_X2 _09861_ ( .A1(_02250_ ), .A2(_02251_ ), .ZN(_02252_ ) );
INV_X1 _09862_ ( .A(\ID_EX_imm [19] ), .ZN(_02253_ ) );
XNOR2_X1 _09863_ ( .A(_02252_ ), .B(_02253_ ), .ZN(_02254_ ) );
OR3_X1 _09864_ ( .A1(_02086_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02128_ ), .ZN(_02255_ ) );
OR2_X1 _09865_ ( .A1(_02132_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02256_ ) );
OAI211_X1 _09866_ ( .A(_02256_ ), .B(_02099_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02257_ ) );
OR2_X1 _09867_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02258_ ) );
OAI211_X1 _09868_ ( .A(_02258_ ), .B(fanout_net_25 ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02259_ ) );
NAND3_X1 _09869_ ( .A1(_02257_ ), .A2(_02106_ ), .A3(_02259_ ), .ZN(_02260_ ) );
MUX2_X1 _09870_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02261_ ) );
MUX2_X1 _09871_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02262_ ) );
MUX2_X1 _09872_ ( .A(_02261_ ), .B(_02262_ ), .S(_02067_ ), .Z(_02263_ ) );
OAI211_X1 _09873_ ( .A(_02049_ ), .B(_02260_ ), .C1(_02263_ ), .C2(_02055_ ), .ZN(_02264_ ) );
OR2_X1 _09874_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02265_ ) );
OAI211_X1 _09875_ ( .A(_02265_ ), .B(fanout_net_25 ), .C1(_02145_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02266_ ) );
OR2_X1 _09876_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02267_ ) );
OAI211_X1 _09877_ ( .A(_02267_ ), .B(_02099_ ), .C1(_02137_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02268_ ) );
NAND3_X1 _09878_ ( .A1(_02266_ ), .A2(_02268_ ), .A3(fanout_net_27 ), .ZN(_02269_ ) );
MUX2_X1 _09879_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02270_ ) );
MUX2_X1 _09880_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02271_ ) );
MUX2_X1 _09881_ ( .A(_02270_ ), .B(_02271_ ), .S(fanout_net_25 ), .Z(_02272_ ) );
OAI211_X1 _09882_ ( .A(fanout_net_28 ), .B(_02269_ ), .C1(_02272_ ), .C2(fanout_net_27 ), .ZN(_02273_ ) );
OAI211_X1 _09883_ ( .A(_02264_ ), .B(_02273_ ), .C1(_02037_ ), .C2(_02045_ ), .ZN(_02274_ ) );
NAND2_X1 _09884_ ( .A1(_02255_ ), .A2(_02274_ ), .ZN(_02275_ ) );
INV_X1 _09885_ ( .A(\ID_EX_imm [18] ), .ZN(_02276_ ) );
XNOR2_X1 _09886_ ( .A(_02275_ ), .B(_02276_ ), .ZN(_02277_ ) );
AND2_X1 _09887_ ( .A1(_02254_ ), .A2(_02277_ ), .ZN(_02278_ ) );
OR3_X1 _09888_ ( .A1(_02036_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02044_ ), .ZN(_02279_ ) );
OR2_X1 _09889_ ( .A1(_02136_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02280_ ) );
OAI211_X1 _09890_ ( .A(_02280_ ), .B(_02215_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02281_ ) );
OR2_X1 _09891_ ( .A1(_02136_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02282_ ) );
OAI211_X1 _09892_ ( .A(_02282_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02283_ ) );
NAND3_X1 _09893_ ( .A1(_02281_ ), .A2(_02283_ ), .A3(fanout_net_27 ), .ZN(_02284_ ) );
MUX2_X1 _09894_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02285_ ) );
MUX2_X1 _09895_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02286_ ) );
MUX2_X1 _09896_ ( .A(_02285_ ), .B(_02286_ ), .S(_02215_ ), .Z(_02287_ ) );
OAI211_X1 _09897_ ( .A(_02049_ ), .B(_02284_ ), .C1(_02287_ ), .C2(fanout_net_27 ), .ZN(_02288_ ) );
NOR2_X1 _09898_ ( .A1(_02059_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02289_ ) );
OAI21_X1 _09899_ ( .A(fanout_net_25 ), .B1(fanout_net_18 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02290_ ) );
NOR2_X1 _09900_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02291_ ) );
OAI21_X1 _09901_ ( .A(_02215_ ), .B1(_02059_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02292_ ) );
OAI221_X1 _09902_ ( .A(_02105_ ), .B1(_02289_ ), .B2(_02290_ ), .C1(_02291_ ), .C2(_02292_ ), .ZN(_02293_ ) );
MUX2_X1 _09903_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02294_ ) );
MUX2_X1 _09904_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02295_ ) );
MUX2_X1 _09905_ ( .A(_02294_ ), .B(_02295_ ), .S(fanout_net_25 ), .Z(_02296_ ) );
OAI211_X1 _09906_ ( .A(fanout_net_28 ), .B(_02293_ ), .C1(_02296_ ), .C2(_02106_ ), .ZN(_02297_ ) );
OAI211_X1 _09907_ ( .A(_02288_ ), .B(_02297_ ), .C1(_02086_ ), .C2(_02128_ ), .ZN(_02298_ ) );
NAND2_X1 _09908_ ( .A1(_02279_ ), .A2(_02298_ ), .ZN(_02299_ ) );
INV_X1 _09909_ ( .A(\ID_EX_imm [17] ), .ZN(_02300_ ) );
XNOR2_X1 _09910_ ( .A(_02299_ ), .B(_02300_ ), .ZN(_02301_ ) );
OR3_X1 _09911_ ( .A1(_02036_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02094_ ), .ZN(_02302_ ) );
OR2_X1 _09912_ ( .A1(_02132_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02303_ ) );
OAI211_X1 _09913_ ( .A(_02303_ ), .B(_02099_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02304_ ) );
OR2_X1 _09914_ ( .A1(_02136_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02305_ ) );
OAI211_X1 _09915_ ( .A(_02305_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02306_ ) );
NAND3_X1 _09916_ ( .A1(_02304_ ), .A2(_02306_ ), .A3(fanout_net_27 ), .ZN(_02307_ ) );
MUX2_X1 _09917_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02308_ ) );
MUX2_X1 _09918_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02309_ ) );
MUX2_X1 _09919_ ( .A(_02308_ ), .B(_02309_ ), .S(_02067_ ), .Z(_02310_ ) );
OAI211_X1 _09920_ ( .A(_02049_ ), .B(_02307_ ), .C1(_02310_ ), .C2(fanout_net_27 ), .ZN(_02311_ ) );
NOR2_X1 _09921_ ( .A1(_02059_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02312_ ) );
OAI21_X1 _09922_ ( .A(fanout_net_25 ), .B1(fanout_net_18 ), .B2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02313_ ) );
NOR2_X1 _09923_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02314_ ) );
OAI21_X1 _09924_ ( .A(_02067_ ), .B1(_02059_ ), .B2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02315_ ) );
OAI221_X1 _09925_ ( .A(_02054_ ), .B1(_02312_ ), .B2(_02313_ ), .C1(_02314_ ), .C2(_02315_ ), .ZN(_02316_ ) );
MUX2_X1 _09926_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02317_ ) );
MUX2_X1 _09927_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02318_ ) );
MUX2_X1 _09928_ ( .A(_02317_ ), .B(_02318_ ), .S(fanout_net_25 ), .Z(_02319_ ) );
OAI211_X1 _09929_ ( .A(fanout_net_28 ), .B(_02316_ ), .C1(_02319_ ), .C2(_02106_ ), .ZN(_02320_ ) );
OAI211_X1 _09930_ ( .A(_02311_ ), .B(_02320_ ), .C1(_02086_ ), .C2(_02045_ ), .ZN(_02321_ ) );
NAND2_X1 _09931_ ( .A1(_02302_ ), .A2(_02321_ ), .ZN(_02322_ ) );
INV_X1 _09932_ ( .A(\ID_EX_imm [16] ), .ZN(_02323_ ) );
XNOR2_X1 _09933_ ( .A(_02322_ ), .B(_02323_ ), .ZN(_02324_ ) );
NAND3_X1 _09934_ ( .A1(_02278_ ), .A2(_02301_ ), .A3(_02324_ ), .ZN(_02325_ ) );
BUF_X2 _09935_ ( .A(_02035_ ), .Z(_02326_ ) );
CLKBUF_X2 _09936_ ( .A(_02042_ ), .Z(_02327_ ) );
OR3_X1 _09937_ ( .A1(_02326_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02328_ ) );
OR2_X1 _09938_ ( .A1(_02057_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02329_ ) );
BUF_X4 _09939_ ( .A(_02065_ ), .Z(_02330_ ) );
OAI211_X1 _09940_ ( .A(_02329_ ), .B(_02330_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02331_ ) );
BUF_X4 _09941_ ( .A(_02052_ ), .Z(_02332_ ) );
OR2_X1 _09942_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02333_ ) );
BUF_X2 _09943_ ( .A(_02130_ ), .Z(_02334_ ) );
OAI211_X1 _09944_ ( .A(_02333_ ), .B(fanout_net_25 ), .C1(_02334_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02335_ ) );
NAND3_X1 _09945_ ( .A1(_02331_ ), .A2(_02332_ ), .A3(_02335_ ), .ZN(_02336_ ) );
MUX2_X1 _09946_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02337_ ) );
MUX2_X1 _09947_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02338_ ) );
BUF_X4 _09948_ ( .A(_02065_ ), .Z(_02339_ ) );
MUX2_X1 _09949_ ( .A(_02337_ ), .B(_02338_ ), .S(_02339_ ), .Z(_02340_ ) );
OAI211_X1 _09950_ ( .A(fanout_net_28 ), .B(_02336_ ), .C1(_02340_ ), .C2(_02053_ ), .ZN(_02341_ ) );
OR2_X1 _09951_ ( .A1(_02057_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02342_ ) );
OAI211_X1 _09952_ ( .A(_02342_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02343_ ) );
OR2_X1 _09953_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02344_ ) );
OAI211_X1 _09954_ ( .A(_02344_ ), .B(_02339_ ), .C1(_02334_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02345_ ) );
NAND3_X1 _09955_ ( .A1(_02343_ ), .A2(_02332_ ), .A3(_02345_ ), .ZN(_02346_ ) );
MUX2_X1 _09956_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02347_ ) );
MUX2_X1 _09957_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02348_ ) );
MUX2_X1 _09958_ ( .A(_02347_ ), .B(_02348_ ), .S(_02339_ ), .Z(_02349_ ) );
OAI211_X1 _09959_ ( .A(_02048_ ), .B(_02346_ ), .C1(_02349_ ), .C2(_02053_ ), .ZN(_02350_ ) );
OAI211_X1 _09960_ ( .A(_02341_ ), .B(_02350_ ), .C1(_02326_ ), .C2(_02093_ ), .ZN(_02351_ ) );
NAND2_X1 _09961_ ( .A1(_02328_ ), .A2(_02351_ ), .ZN(_02352_ ) );
XNOR2_X1 _09962_ ( .A(_02352_ ), .B(\ID_EX_imm [3] ), .ZN(_02353_ ) );
BUF_X2 _09963_ ( .A(_02042_ ), .Z(_02354_ ) );
CLKBUF_X2 _09964_ ( .A(_02354_ ), .Z(_02355_ ) );
OR3_X1 _09965_ ( .A1(_02085_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02356_ ) );
OR2_X1 _09966_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02357_ ) );
OAI211_X1 _09967_ ( .A(_02357_ ), .B(_02214_ ), .C1(_02136_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02358_ ) );
OR2_X1 _09968_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02359_ ) );
OAI211_X1 _09969_ ( .A(_02359_ ), .B(fanout_net_25 ), .C1(_02136_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02360_ ) );
NAND3_X1 _09970_ ( .A1(_02358_ ), .A2(_02360_ ), .A3(_02053_ ), .ZN(_02361_ ) );
MUX2_X1 _09971_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02362_ ) );
MUX2_X1 _09972_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02363_ ) );
MUX2_X1 _09973_ ( .A(_02362_ ), .B(_02363_ ), .S(_02214_ ), .Z(_02364_ ) );
OAI211_X1 _09974_ ( .A(_02048_ ), .B(_02361_ ), .C1(_02364_ ), .C2(_02105_ ), .ZN(_02365_ ) );
OR2_X1 _09975_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02366_ ) );
OAI211_X1 _09976_ ( .A(_02366_ ), .B(fanout_net_26 ), .C1(_02136_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02367_ ) );
OR2_X1 _09977_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02368_ ) );
OAI211_X1 _09978_ ( .A(_02368_ ), .B(_02214_ ), .C1(_02136_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02369_ ) );
NAND3_X1 _09979_ ( .A1(_02367_ ), .A2(_02369_ ), .A3(fanout_net_27 ), .ZN(_02370_ ) );
MUX2_X1 _09980_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02371_ ) );
MUX2_X1 _09981_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02372_ ) );
MUX2_X1 _09982_ ( .A(_02371_ ), .B(_02372_ ), .S(fanout_net_26 ), .Z(_02373_ ) );
OAI211_X1 _09983_ ( .A(fanout_net_28 ), .B(_02370_ ), .C1(_02373_ ), .C2(fanout_net_27 ), .ZN(_02374_ ) );
OAI211_X1 _09984_ ( .A(_02365_ ), .B(_02374_ ), .C1(_02085_ ), .C2(_02044_ ), .ZN(_02375_ ) );
NAND2_X1 _09985_ ( .A1(_02356_ ), .A2(_02375_ ), .ZN(_02376_ ) );
INV_X1 _09986_ ( .A(\ID_EX_imm [2] ), .ZN(_02377_ ) );
XNOR2_X1 _09987_ ( .A(_02376_ ), .B(_02377_ ), .ZN(_02378_ ) );
OR3_X1 _09988_ ( .A1(_02035_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02354_ ), .ZN(_02379_ ) );
OR2_X1 _09989_ ( .A1(_02130_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02380_ ) );
OAI211_X1 _09990_ ( .A(_02380_ ), .B(fanout_net_26 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02381_ ) );
OR2_X1 _09991_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02382_ ) );
OAI211_X1 _09992_ ( .A(_02382_ ), .B(_02064_ ), .C1(_02130_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02383_ ) );
NAND3_X1 _09993_ ( .A1(_02381_ ), .A2(_02051_ ), .A3(_02383_ ), .ZN(_02384_ ) );
MUX2_X1 _09994_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02385_ ) );
MUX2_X1 _09995_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02386_ ) );
MUX2_X1 _09996_ ( .A(_02385_ ), .B(_02386_ ), .S(_02064_ ), .Z(_02387_ ) );
OAI211_X1 _09997_ ( .A(fanout_net_28 ), .B(_02384_ ), .C1(_02387_ ), .C2(_02052_ ), .ZN(_02388_ ) );
OR2_X1 _09998_ ( .A1(_02130_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02389_ ) );
OAI211_X1 _09999_ ( .A(_02389_ ), .B(_02064_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02390_ ) );
OR2_X1 _10000_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02391_ ) );
OAI211_X1 _10001_ ( .A(_02391_ ), .B(fanout_net_26 ), .C1(_02130_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02392_ ) );
NAND3_X1 _10002_ ( .A1(_02390_ ), .A2(_02051_ ), .A3(_02392_ ), .ZN(_02393_ ) );
MUX2_X1 _10003_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02394_ ) );
MUX2_X1 _10004_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02395_ ) );
MUX2_X1 _10005_ ( .A(_02394_ ), .B(_02395_ ), .S(_02064_ ), .Z(_02396_ ) );
OAI211_X1 _10006_ ( .A(_02047_ ), .B(_02393_ ), .C1(_02396_ ), .C2(_02052_ ), .ZN(_02397_ ) );
OAI211_X1 _10007_ ( .A(_02388_ ), .B(_02397_ ), .C1(_02035_ ), .C2(_02043_ ), .ZN(_02398_ ) );
NAND2_X2 _10008_ ( .A1(_02379_ ), .A2(_02398_ ), .ZN(_02399_ ) );
INV_X1 _10009_ ( .A(\ID_EX_imm [1] ), .ZN(_02400_ ) );
XNOR2_X1 _10010_ ( .A(_02399_ ), .B(_02400_ ), .ZN(_02401_ ) );
NOR2_X1 _10011_ ( .A1(_02035_ ), .A2(_02354_ ), .ZN(_02402_ ) );
NAND2_X1 _10012_ ( .A1(_02402_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_02403_ ) );
OR2_X1 _10013_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02404_ ) );
OAI211_X1 _10014_ ( .A(_02404_ ), .B(_02065_ ), .C1(_02130_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02405_ ) );
OR2_X1 _10015_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02406_ ) );
OAI211_X1 _10016_ ( .A(_02406_ ), .B(fanout_net_26 ), .C1(_02130_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02407_ ) );
NAND3_X1 _10017_ ( .A1(_02405_ ), .A2(_02407_ ), .A3(_02051_ ), .ZN(_02408_ ) );
MUX2_X1 _10018_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02409_ ) );
MUX2_X1 _10019_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02410_ ) );
MUX2_X1 _10020_ ( .A(_02409_ ), .B(_02410_ ), .S(_02064_ ), .Z(_02411_ ) );
OAI211_X1 _10021_ ( .A(fanout_net_28 ), .B(_02408_ ), .C1(_02411_ ), .C2(_02052_ ), .ZN(_02412_ ) );
OR2_X1 _10022_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(fanout_net_19 ), .ZN(_02413_ ) );
OAI211_X1 _10023_ ( .A(_02413_ ), .B(_02064_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_02130_ ), .ZN(_02414_ ) );
OR2_X1 _10024_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02415_ ) );
OAI211_X1 _10025_ ( .A(_02415_ ), .B(fanout_net_26 ), .C1(_02130_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02416_ ) );
NAND3_X1 _10026_ ( .A1(_02414_ ), .A2(_02416_ ), .A3(_02051_ ), .ZN(_02417_ ) );
MUX2_X1 _10027_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02418_ ) );
MUX2_X1 _10028_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02419_ ) );
MUX2_X1 _10029_ ( .A(_02418_ ), .B(_02419_ ), .S(_02064_ ), .Z(_02420_ ) );
OAI211_X1 _10030_ ( .A(_02047_ ), .B(_02417_ ), .C1(_02420_ ), .C2(_02052_ ), .ZN(_02421_ ) );
NAND2_X1 _10031_ ( .A1(_02412_ ), .A2(_02421_ ), .ZN(_02422_ ) );
OAI21_X1 _10032_ ( .A(_02422_ ), .B1(_02035_ ), .B2(_02043_ ), .ZN(_02423_ ) );
AND3_X1 _10033_ ( .A1(_02403_ ), .A2(\ID_EX_imm [0] ), .A3(_02423_ ), .ZN(_02424_ ) );
AND2_X1 _10034_ ( .A1(_02401_ ), .A2(_02424_ ), .ZN(_02425_ ) );
AOI21_X1 _10035_ ( .A(_02400_ ), .B1(_02379_ ), .B2(_02398_ ), .ZN(_02426_ ) );
OAI21_X4 _10036_ ( .A(_02378_ ), .B1(_02425_ ), .B2(_02426_ ), .ZN(_02427_ ) );
NAND2_X1 _10037_ ( .A1(_02376_ ), .A2(\ID_EX_imm [2] ), .ZN(_02428_ ) );
AOI21_X1 _10038_ ( .A(_02353_ ), .B1(_02427_ ), .B2(_02428_ ), .ZN(_02429_ ) );
AOI21_X1 _10039_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B1(_02328_ ), .B2(_02351_ ), .ZN(_02430_ ) );
NOR2_X2 _10040_ ( .A1(_02429_ ), .A2(_02430_ ), .ZN(_02431_ ) );
OR3_X1 _10041_ ( .A1(_02326_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02432_ ) );
OR2_X1 _10042_ ( .A1(_02057_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02433_ ) );
OAI211_X1 _10043_ ( .A(_02433_ ), .B(fanout_net_26 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02434_ ) );
OR2_X1 _10044_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02435_ ) );
OAI211_X1 _10045_ ( .A(_02435_ ), .B(_02330_ ), .C1(_02334_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02436_ ) );
NAND3_X1 _10046_ ( .A1(_02434_ ), .A2(_02332_ ), .A3(_02436_ ), .ZN(_02437_ ) );
MUX2_X1 _10047_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02438_ ) );
MUX2_X1 _10048_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02439_ ) );
MUX2_X1 _10049_ ( .A(_02438_ ), .B(_02439_ ), .S(_02339_ ), .Z(_02440_ ) );
OAI211_X1 _10050_ ( .A(fanout_net_28 ), .B(_02437_ ), .C1(_02440_ ), .C2(_02053_ ), .ZN(_02441_ ) );
OR2_X1 _10051_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02442_ ) );
OAI211_X1 _10052_ ( .A(_02442_ ), .B(_02330_ ), .C1(_02334_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02443_ ) );
OR2_X1 _10053_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02444_ ) );
OAI211_X1 _10054_ ( .A(_02444_ ), .B(fanout_net_26 ), .C1(_02334_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02445_ ) );
NAND3_X1 _10055_ ( .A1(_02443_ ), .A2(_02445_ ), .A3(_02332_ ), .ZN(_02446_ ) );
MUX2_X1 _10056_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02447_ ) );
MUX2_X1 _10057_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02448_ ) );
MUX2_X1 _10058_ ( .A(_02447_ ), .B(_02448_ ), .S(_02339_ ), .Z(_02449_ ) );
OAI211_X1 _10059_ ( .A(_02048_ ), .B(_02446_ ), .C1(_02449_ ), .C2(_02053_ ), .ZN(_02450_ ) );
OAI211_X1 _10060_ ( .A(_02441_ ), .B(_02450_ ), .C1(_02085_ ), .C2(_02093_ ), .ZN(_02451_ ) );
NAND2_X1 _10061_ ( .A1(_02432_ ), .A2(_02451_ ), .ZN(_02452_ ) );
INV_X1 _10062_ ( .A(\ID_EX_imm [4] ), .ZN(_02453_ ) );
XNOR2_X1 _10063_ ( .A(_02452_ ), .B(_02453_ ), .ZN(_02454_ ) );
INV_X1 _10064_ ( .A(_02454_ ), .ZN(_02455_ ) );
NOR2_X1 _10065_ ( .A1(_02431_ ), .A2(_02455_ ), .ZN(_02456_ ) );
OR3_X1 _10066_ ( .A1(_02326_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02457_ ) );
OR2_X1 _10067_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02458_ ) );
OAI211_X1 _10068_ ( .A(_02458_ ), .B(_02330_ ), .C1(_02058_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02459_ ) );
OR2_X1 _10069_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02460_ ) );
OAI211_X1 _10070_ ( .A(_02460_ ), .B(fanout_net_26 ), .C1(_02058_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02461_ ) );
NAND3_X1 _10071_ ( .A1(_02459_ ), .A2(_02461_ ), .A3(fanout_net_27 ), .ZN(_02462_ ) );
MUX2_X1 _10072_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02463_ ) );
MUX2_X1 _10073_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02464_ ) );
MUX2_X1 _10074_ ( .A(_02463_ ), .B(_02464_ ), .S(_02330_ ), .Z(_02465_ ) );
OAI211_X1 _10075_ ( .A(_02048_ ), .B(_02462_ ), .C1(_02465_ ), .C2(fanout_net_27 ), .ZN(_02466_ ) );
NOR2_X1 _10076_ ( .A1(_02131_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02467_ ) );
OAI21_X1 _10077_ ( .A(fanout_net_26 ), .B1(fanout_net_20 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02468_ ) );
NOR2_X1 _10078_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02469_ ) );
OAI21_X1 _10079_ ( .A(_02339_ ), .B1(_02131_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02470_ ) );
OAI221_X1 _10080_ ( .A(_02052_ ), .B1(_02467_ ), .B2(_02468_ ), .C1(_02469_ ), .C2(_02470_ ), .ZN(_02471_ ) );
MUX2_X1 _10081_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02472_ ) );
MUX2_X1 _10082_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02473_ ) );
MUX2_X1 _10083_ ( .A(_02472_ ), .B(_02473_ ), .S(fanout_net_26 ), .Z(_02474_ ) );
OAI211_X1 _10084_ ( .A(fanout_net_28 ), .B(_02471_ ), .C1(_02474_ ), .C2(_02053_ ), .ZN(_02475_ ) );
OAI211_X1 _10085_ ( .A(_02466_ ), .B(_02475_ ), .C1(_02085_ ), .C2(_02093_ ), .ZN(_02476_ ) );
NAND2_X2 _10086_ ( .A1(_02457_ ), .A2(_02476_ ), .ZN(_02477_ ) );
XOR2_X1 _10087_ ( .A(_02477_ ), .B(\ID_EX_imm [7] ), .Z(_02478_ ) );
OR3_X1 _10088_ ( .A1(_02326_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02479_ ) );
OR2_X1 _10089_ ( .A1(_02057_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02480_ ) );
OAI211_X1 _10090_ ( .A(_02480_ ), .B(_02214_ ), .C1(fanout_net_20 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02481_ ) );
OR2_X1 _10091_ ( .A1(fanout_net_20 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02482_ ) );
OAI211_X1 _10092_ ( .A(_02482_ ), .B(fanout_net_26 ), .C1(_02334_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02483_ ) );
NAND3_X1 _10093_ ( .A1(_02481_ ), .A2(fanout_net_27 ), .A3(_02483_ ), .ZN(_02484_ ) );
MUX2_X1 _10094_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02485_ ) );
MUX2_X1 _10095_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02486_ ) );
MUX2_X1 _10096_ ( .A(_02485_ ), .B(_02486_ ), .S(_02330_ ), .Z(_02487_ ) );
OAI211_X1 _10097_ ( .A(_02048_ ), .B(_02484_ ), .C1(_02487_ ), .C2(fanout_net_27 ), .ZN(_02488_ ) );
NOR2_X1 _10098_ ( .A1(_02131_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02489_ ) );
OAI21_X1 _10099_ ( .A(fanout_net_26 ), .B1(fanout_net_20 ), .B2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02490_ ) );
NOR2_X1 _10100_ ( .A1(fanout_net_20 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02491_ ) );
OAI21_X1 _10101_ ( .A(_02330_ ), .B1(_02334_ ), .B2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02492_ ) );
OAI221_X1 _10102_ ( .A(_02332_ ), .B1(_02489_ ), .B2(_02490_ ), .C1(_02491_ ), .C2(_02492_ ), .ZN(_02493_ ) );
MUX2_X1 _10103_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02494_ ) );
MUX2_X1 _10104_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02495_ ) );
MUX2_X1 _10105_ ( .A(_02494_ ), .B(_02495_ ), .S(fanout_net_26 ), .Z(_02496_ ) );
OAI211_X1 _10106_ ( .A(fanout_net_28 ), .B(_02493_ ), .C1(_02496_ ), .C2(_02105_ ), .ZN(_02497_ ) );
OAI211_X1 _10107_ ( .A(_02488_ ), .B(_02497_ ), .C1(_02085_ ), .C2(_02093_ ), .ZN(_02498_ ) );
NAND2_X1 _10108_ ( .A1(_02479_ ), .A2(_02498_ ), .ZN(_02499_ ) );
XOR2_X1 _10109_ ( .A(_02499_ ), .B(\ID_EX_imm [6] ), .Z(_02500_ ) );
AND2_X1 _10110_ ( .A1(_02478_ ), .A2(_02500_ ), .ZN(_02501_ ) );
NAND2_X1 _10111_ ( .A1(_02402_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02502_ ) );
OR2_X1 _10112_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02503_ ) );
OAI211_X1 _10113_ ( .A(_02503_ ), .B(fanout_net_26 ), .C1(_02057_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02504_ ) );
INV_X1 _10114_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02505_ ) );
NAND2_X1 _10115_ ( .A1(_02505_ ), .A2(fanout_net_20 ), .ZN(_02506_ ) );
OAI211_X1 _10116_ ( .A(_02506_ ), .B(_02065_ ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02507_ ) );
NAND3_X1 _10117_ ( .A1(_02504_ ), .A2(_02507_ ), .A3(_02052_ ), .ZN(_02508_ ) );
MUX2_X1 _10118_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02509_ ) );
MUX2_X1 _10119_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02510_ ) );
MUX2_X1 _10120_ ( .A(_02509_ ), .B(_02510_ ), .S(_02064_ ), .Z(_02511_ ) );
OAI211_X1 _10121_ ( .A(_02047_ ), .B(_02508_ ), .C1(_02511_ ), .C2(_02052_ ), .ZN(_02512_ ) );
OR2_X1 _10122_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02513_ ) );
OAI211_X1 _10123_ ( .A(_02513_ ), .B(_02065_ ), .C1(_02057_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02514_ ) );
INV_X1 _10124_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02515_ ) );
NAND2_X1 _10125_ ( .A1(_02515_ ), .A2(fanout_net_20 ), .ZN(_02516_ ) );
OAI211_X1 _10126_ ( .A(_02516_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02517_ ) );
NAND3_X1 _10127_ ( .A1(_02514_ ), .A2(_02517_ ), .A3(fanout_net_27 ), .ZN(_02518_ ) );
MUX2_X1 _10128_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02519_ ) );
MUX2_X1 _10129_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02520_ ) );
MUX2_X1 _10130_ ( .A(_02519_ ), .B(_02520_ ), .S(fanout_net_26 ), .Z(_02521_ ) );
OAI211_X1 _10131_ ( .A(fanout_net_28 ), .B(_02518_ ), .C1(_02521_ ), .C2(fanout_net_27 ), .ZN(_02522_ ) );
NAND2_X1 _10132_ ( .A1(_02512_ ), .A2(_02522_ ), .ZN(_02523_ ) );
OAI21_X1 _10133_ ( .A(_02523_ ), .B1(_02326_ ), .B2(_02355_ ), .ZN(_02524_ ) );
AND2_X2 _10134_ ( .A1(_02502_ ), .A2(_02524_ ), .ZN(_02525_ ) );
XNOR2_X1 _10135_ ( .A(_02525_ ), .B(\ID_EX_imm [5] ), .ZN(_02526_ ) );
INV_X1 _10136_ ( .A(_02526_ ), .ZN(_02527_ ) );
NAND3_X1 _10137_ ( .A1(_02456_ ), .A2(_02501_ ), .A3(_02527_ ), .ZN(_02528_ ) );
XNOR2_X1 _10138_ ( .A(_02477_ ), .B(\ID_EX_imm [7] ), .ZN(_02529_ ) );
BUF_X4 _10139_ ( .A(_02499_ ), .Z(_02530_ ) );
NAND2_X1 _10140_ ( .A1(_02530_ ), .A2(\ID_EX_imm [6] ), .ZN(_02531_ ) );
NOR2_X1 _10141_ ( .A1(_02529_ ), .A2(_02531_ ), .ZN(_02532_ ) );
INV_X1 _10142_ ( .A(_02452_ ), .ZN(_02533_ ) );
NOR3_X1 _10143_ ( .A1(_02526_ ), .A2(_02453_ ), .A3(_02533_ ), .ZN(_02534_ ) );
INV_X1 _10144_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02535_ ) );
AOI21_X1 _10145_ ( .A(_02534_ ), .B1(_02535_ ), .B2(_02525_ ), .ZN(_02536_ ) );
INV_X1 _10146_ ( .A(_02536_ ), .ZN(_02537_ ) );
AOI221_X4 _10147_ ( .A(_02532_ ), .B1(\ID_EX_imm [7] ), .B2(_02477_ ), .C1(_02537_ ), .C2(_02501_ ), .ZN(_02538_ ) );
NAND2_X2 _10148_ ( .A1(_02528_ ), .A2(_02538_ ), .ZN(_02539_ ) );
OR3_X1 _10149_ ( .A1(_02036_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02044_ ), .ZN(_02540_ ) );
OR2_X1 _10150_ ( .A1(_02058_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02541_ ) );
OAI211_X1 _10151_ ( .A(_02541_ ), .B(_02215_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02542_ ) );
OR2_X1 _10152_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02543_ ) );
OAI211_X1 _10153_ ( .A(_02543_ ), .B(fanout_net_26 ), .C1(_02059_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02544_ ) );
NAND3_X1 _10154_ ( .A1(_02542_ ), .A2(_02054_ ), .A3(_02544_ ), .ZN(_02545_ ) );
MUX2_X1 _10155_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02546_ ) );
MUX2_X1 _10156_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02547_ ) );
MUX2_X1 _10157_ ( .A(_02546_ ), .B(_02547_ ), .S(_02215_ ), .Z(_02548_ ) );
OAI211_X1 _10158_ ( .A(_02049_ ), .B(_02545_ ), .C1(_02548_ ), .C2(_02054_ ), .ZN(_02549_ ) );
OR2_X1 _10159_ ( .A1(_02058_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02550_ ) );
OAI211_X1 _10160_ ( .A(_02550_ ), .B(fanout_net_26 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02551_ ) );
OR2_X1 _10161_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02552_ ) );
OAI211_X1 _10162_ ( .A(_02552_ ), .B(_02215_ ), .C1(_02059_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02553_ ) );
NAND3_X1 _10163_ ( .A1(_02551_ ), .A2(fanout_net_27 ), .A3(_02553_ ), .ZN(_02554_ ) );
MUX2_X1 _10164_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02555_ ) );
MUX2_X1 _10165_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02556_ ) );
MUX2_X1 _10166_ ( .A(_02555_ ), .B(_02556_ ), .S(fanout_net_26 ), .Z(_02557_ ) );
OAI211_X1 _10167_ ( .A(fanout_net_28 ), .B(_02554_ ), .C1(_02557_ ), .C2(fanout_net_27 ), .ZN(_02558_ ) );
OAI211_X1 _10168_ ( .A(_02549_ ), .B(_02558_ ), .C1(_02086_ ), .C2(_02128_ ), .ZN(_02559_ ) );
NAND2_X1 _10169_ ( .A1(_02540_ ), .A2(_02559_ ), .ZN(_02560_ ) );
BUF_X4 _10170_ ( .A(_02560_ ), .Z(_02561_ ) );
INV_X1 _10171_ ( .A(\ID_EX_imm [12] ), .ZN(_02562_ ) );
XNOR2_X1 _10172_ ( .A(_02561_ ), .B(_02562_ ), .ZN(_02563_ ) );
OR3_X1 _10173_ ( .A1(_02326_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02564_ ) );
INV_X1 _10174_ ( .A(\ID_EX_imm [13] ), .ZN(_02565_ ) );
OR2_X1 _10175_ ( .A1(_02131_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02566_ ) );
OAI211_X1 _10176_ ( .A(_02566_ ), .B(fanout_net_26 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02567_ ) );
OR2_X1 _10177_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02568_ ) );
OAI211_X1 _10178_ ( .A(_02568_ ), .B(_02214_ ), .C1(_02058_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02569_ ) );
NAND3_X1 _10179_ ( .A1(_02567_ ), .A2(_02053_ ), .A3(_02569_ ), .ZN(_02570_ ) );
MUX2_X1 _10180_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02571_ ) );
MUX2_X1 _10181_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02572_ ) );
MUX2_X1 _10182_ ( .A(_02571_ ), .B(_02572_ ), .S(_02214_ ), .Z(_02573_ ) );
OAI211_X1 _10183_ ( .A(_02048_ ), .B(_02570_ ), .C1(_02573_ ), .C2(_02105_ ), .ZN(_02574_ ) );
OR2_X1 _10184_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02575_ ) );
OAI211_X1 _10185_ ( .A(_02575_ ), .B(fanout_net_26 ), .C1(_02136_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02576_ ) );
OR2_X1 _10186_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02577_ ) );
OAI211_X1 _10187_ ( .A(_02577_ ), .B(_02214_ ), .C1(_02058_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02578_ ) );
NAND3_X1 _10188_ ( .A1(_02576_ ), .A2(_02578_ ), .A3(fanout_net_27 ), .ZN(_02579_ ) );
MUX2_X1 _10189_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02580_ ) );
MUX2_X1 _10190_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02581_ ) );
MUX2_X1 _10191_ ( .A(_02580_ ), .B(_02581_ ), .S(fanout_net_26 ), .Z(_02582_ ) );
OAI211_X1 _10192_ ( .A(fanout_net_28 ), .B(_02579_ ), .C1(_02582_ ), .C2(fanout_net_27 ), .ZN(_02583_ ) );
OAI211_X1 _10193_ ( .A(_02574_ ), .B(_02583_ ), .C1(_02085_ ), .C2(_02127_ ), .ZN(_02584_ ) );
AND3_X1 _10194_ ( .A1(_02564_ ), .A2(_02565_ ), .A3(_02584_ ), .ZN(_02585_ ) );
AOI21_X1 _10195_ ( .A(_02565_ ), .B1(_02564_ ), .B2(_02584_ ), .ZN(_02586_ ) );
NOR2_X1 _10196_ ( .A1(_02585_ ), .A2(_02586_ ), .ZN(_02587_ ) );
AND2_X1 _10197_ ( .A1(_02563_ ), .A2(_02587_ ), .ZN(_02588_ ) );
OR3_X1 _10198_ ( .A1(_02085_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02127_ ), .ZN(_02589_ ) );
OR2_X1 _10199_ ( .A1(_02131_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02590_ ) );
OAI211_X1 _10200_ ( .A(_02590_ ), .B(_02066_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02591_ ) );
OR2_X1 _10201_ ( .A1(_02131_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02592_ ) );
OAI211_X1 _10202_ ( .A(_02592_ ), .B(fanout_net_26 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02593_ ) );
NAND3_X1 _10203_ ( .A1(_02591_ ), .A2(_02593_ ), .A3(_02105_ ), .ZN(_02594_ ) );
MUX2_X1 _10204_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02595_ ) );
MUX2_X1 _10205_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02596_ ) );
MUX2_X1 _10206_ ( .A(_02595_ ), .B(_02596_ ), .S(_02066_ ), .Z(_02597_ ) );
OAI211_X1 _10207_ ( .A(fanout_net_28 ), .B(_02594_ ), .C1(_02597_ ), .C2(_02054_ ), .ZN(_02598_ ) );
OR2_X1 _10208_ ( .A1(_02131_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02599_ ) );
OAI211_X1 _10209_ ( .A(_02599_ ), .B(_02066_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02600_ ) );
OR2_X1 _10210_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02601_ ) );
OAI211_X1 _10211_ ( .A(_02601_ ), .B(fanout_net_26 ), .C1(_02136_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02602_ ) );
NAND3_X1 _10212_ ( .A1(_02600_ ), .A2(_02105_ ), .A3(_02602_ ), .ZN(_02603_ ) );
MUX2_X1 _10213_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02604_ ) );
MUX2_X1 _10214_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02605_ ) );
MUX2_X1 _10215_ ( .A(_02604_ ), .B(_02605_ ), .S(_02214_ ), .Z(_02606_ ) );
OAI211_X1 _10216_ ( .A(_02048_ ), .B(_02603_ ), .C1(_02606_ ), .C2(_02054_ ), .ZN(_02607_ ) );
OAI211_X1 _10217_ ( .A(_02598_ ), .B(_02607_ ), .C1(_02036_ ), .C2(_02044_ ), .ZN(_02608_ ) );
NAND2_X1 _10218_ ( .A1(_02589_ ), .A2(_02608_ ), .ZN(_02609_ ) );
XOR2_X1 _10219_ ( .A(_02609_ ), .B(\ID_EX_imm [15] ), .Z(_02610_ ) );
OR3_X1 _10220_ ( .A1(_02036_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02044_ ), .ZN(_02611_ ) );
OR2_X1 _10221_ ( .A1(_02058_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02612_ ) );
OAI211_X1 _10222_ ( .A(_02612_ ), .B(_02215_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02613_ ) );
OR2_X1 _10223_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02614_ ) );
OAI211_X1 _10224_ ( .A(_02614_ ), .B(fanout_net_26 ), .C1(_02059_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02615_ ) );
NAND3_X1 _10225_ ( .A1(_02613_ ), .A2(_02105_ ), .A3(_02615_ ), .ZN(_02616_ ) );
MUX2_X1 _10226_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02617_ ) );
MUX2_X1 _10227_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02618_ ) );
MUX2_X1 _10228_ ( .A(_02617_ ), .B(_02618_ ), .S(_02066_ ), .Z(_02619_ ) );
OAI211_X1 _10229_ ( .A(_02049_ ), .B(_02616_ ), .C1(_02619_ ), .C2(_02054_ ), .ZN(_02620_ ) );
OR2_X1 _10230_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02621_ ) );
OAI211_X1 _10231_ ( .A(_02621_ ), .B(fanout_net_26 ), .C1(_02059_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02622_ ) );
OR2_X1 _10232_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02623_ ) );
OAI211_X1 _10233_ ( .A(_02623_ ), .B(_02066_ ), .C1(_02132_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02624_ ) );
NAND3_X1 _10234_ ( .A1(_02622_ ), .A2(_02624_ ), .A3(fanout_net_27 ), .ZN(_02625_ ) );
MUX2_X1 _10235_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02626_ ) );
MUX2_X1 _10236_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02627_ ) );
MUX2_X1 _10237_ ( .A(_02626_ ), .B(_02627_ ), .S(fanout_net_26 ), .Z(_02628_ ) );
OAI211_X1 _10238_ ( .A(fanout_net_28 ), .B(_02625_ ), .C1(_02628_ ), .C2(fanout_net_27 ), .ZN(_02629_ ) );
OAI211_X1 _10239_ ( .A(_02620_ ), .B(_02629_ ), .C1(_02036_ ), .C2(_02094_ ), .ZN(_02630_ ) );
NAND2_X2 _10240_ ( .A1(_02611_ ), .A2(_02630_ ), .ZN(_02631_ ) );
INV_X1 _10241_ ( .A(\ID_EX_imm [14] ), .ZN(_02632_ ) );
XNOR2_X1 _10242_ ( .A(_02631_ ), .B(_02632_ ), .ZN(_02633_ ) );
AND3_X1 _10243_ ( .A1(_02588_ ), .A2(_02610_ ), .A3(_02633_ ), .ZN(_02634_ ) );
OR3_X1 _10244_ ( .A1(_02036_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02127_ ), .ZN(_02635_ ) );
OR2_X1 _10245_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02636_ ) );
OAI211_X1 _10246_ ( .A(_02636_ ), .B(_02066_ ), .C1(_02132_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02637_ ) );
OR2_X1 _10247_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02638_ ) );
OAI211_X1 _10248_ ( .A(_02638_ ), .B(fanout_net_26 ), .C1(_02132_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02639_ ) );
NAND3_X1 _10249_ ( .A1(_02637_ ), .A2(_02639_ ), .A3(_02105_ ), .ZN(_02640_ ) );
MUX2_X1 _10250_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02641_ ) );
MUX2_X1 _10251_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02642_ ) );
MUX2_X1 _10252_ ( .A(_02641_ ), .B(_02642_ ), .S(_02066_ ), .Z(_02643_ ) );
OAI211_X1 _10253_ ( .A(_02049_ ), .B(_02640_ ), .C1(_02643_ ), .C2(_02054_ ), .ZN(_02644_ ) );
OR2_X1 _10254_ ( .A1(_02334_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02645_ ) );
OAI211_X1 _10255_ ( .A(_02645_ ), .B(fanout_net_26 ), .C1(fanout_net_22 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02646_ ) );
OR2_X1 _10256_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02647_ ) );
OAI211_X1 _10257_ ( .A(_02647_ ), .B(_02066_ ), .C1(_02132_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02648_ ) );
NAND3_X1 _10258_ ( .A1(_02646_ ), .A2(fanout_net_27 ), .A3(_02648_ ), .ZN(_02649_ ) );
MUX2_X1 _10259_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02650_ ) );
MUX2_X1 _10260_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02651_ ) );
MUX2_X1 _10261_ ( .A(_02650_ ), .B(_02651_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02652_ ) );
OAI211_X1 _10262_ ( .A(fanout_net_28 ), .B(_02649_ ), .C1(_02652_ ), .C2(fanout_net_27 ), .ZN(_02653_ ) );
OAI211_X1 _10263_ ( .A(_02644_ ), .B(_02653_ ), .C1(_02036_ ), .C2(_02094_ ), .ZN(_02654_ ) );
NAND2_X2 _10264_ ( .A1(_02635_ ), .A2(_02654_ ), .ZN(_02655_ ) );
XOR2_X1 _10265_ ( .A(_02655_ ), .B(\ID_EX_imm [8] ), .Z(_02656_ ) );
OR3_X1 _10266_ ( .A1(_02326_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02657_ ) );
OR2_X1 _10267_ ( .A1(_02057_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02658_ ) );
OAI211_X1 _10268_ ( .A(_02658_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_22 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02659_ ) );
OR2_X1 _10269_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02660_ ) );
OAI211_X1 _10270_ ( .A(_02660_ ), .B(_02330_ ), .C1(_02334_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02661_ ) );
NAND3_X1 _10271_ ( .A1(_02659_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02661_ ), .ZN(_02662_ ) );
MUX2_X1 _10272_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02663_ ) );
MUX2_X1 _10273_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02664_ ) );
MUX2_X1 _10274_ ( .A(_02663_ ), .B(_02664_ ), .S(_02330_ ), .Z(_02665_ ) );
OAI211_X1 _10275_ ( .A(_02048_ ), .B(_02662_ ), .C1(_02665_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02666_ ) );
NOR2_X1 _10276_ ( .A1(_02131_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02667_ ) );
OAI21_X1 _10277_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_22 ), .B2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02668_ ) );
NOR2_X1 _10278_ ( .A1(fanout_net_22 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02669_ ) );
OAI21_X1 _10279_ ( .A(_02339_ ), .B1(_02131_ ), .B2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02670_ ) );
OAI221_X1 _10280_ ( .A(_02332_ ), .B1(_02667_ ), .B2(_02668_ ), .C1(_02669_ ), .C2(_02670_ ), .ZN(_02671_ ) );
MUX2_X1 _10281_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02672_ ) );
MUX2_X1 _10282_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02673_ ) );
MUX2_X1 _10283_ ( .A(_02672_ ), .B(_02673_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02674_ ) );
OAI211_X1 _10284_ ( .A(fanout_net_28 ), .B(_02671_ ), .C1(_02674_ ), .C2(_02053_ ), .ZN(_02675_ ) );
OAI211_X1 _10285_ ( .A(_02666_ ), .B(_02675_ ), .C1(_02085_ ), .C2(_02127_ ), .ZN(_02676_ ) );
NAND2_X1 _10286_ ( .A1(_02657_ ), .A2(_02676_ ), .ZN(_02677_ ) );
BUF_X4 _10287_ ( .A(_02677_ ), .Z(_02678_ ) );
AND2_X1 _10288_ ( .A1(_02678_ ), .A2(\ID_EX_imm [9] ), .ZN(_02679_ ) );
INV_X1 _10289_ ( .A(_02679_ ), .ZN(_02680_ ) );
OR2_X1 _10290_ ( .A1(_02678_ ), .A2(\ID_EX_imm [9] ), .ZN(_02681_ ) );
AND3_X1 _10291_ ( .A1(_02656_ ), .A2(_02680_ ), .A3(_02681_ ), .ZN(_02682_ ) );
OR2_X1 _10292_ ( .A1(_02057_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02683_ ) );
OAI211_X1 _10293_ ( .A(_02683_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02684_ ) );
OR2_X1 _10294_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02685_ ) );
OAI211_X1 _10295_ ( .A(_02685_ ), .B(_02339_ ), .C1(_02334_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02686_ ) );
NAND3_X1 _10296_ ( .A1(_02684_ ), .A2(_02332_ ), .A3(_02686_ ), .ZN(_02687_ ) );
MUX2_X1 _10297_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02688_ ) );
MUX2_X1 _10298_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02689_ ) );
MUX2_X1 _10299_ ( .A(_02688_ ), .B(_02689_ ), .S(_02339_ ), .Z(_02690_ ) );
OAI211_X1 _10300_ ( .A(fanout_net_28 ), .B(_02687_ ), .C1(_02690_ ), .C2(_02053_ ), .ZN(_02691_ ) );
MUX2_X1 _10301_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02692_ ) );
AND2_X1 _10302_ ( .A1(_02692_ ), .A2(_02065_ ), .ZN(_02693_ ) );
MUX2_X1 _10303_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02694_ ) );
AOI211_X1 _10304_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_02693_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C2(_02694_ ), .ZN(_02695_ ) );
MUX2_X1 _10305_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02696_ ) );
MUX2_X1 _10306_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02697_ ) );
MUX2_X1 _10307_ ( .A(_02696_ ), .B(_02697_ ), .S(_02065_ ), .Z(_02698_ ) );
OAI21_X1 _10308_ ( .A(_02047_ ), .B1(_02698_ ), .B2(_02332_ ), .ZN(_02699_ ) );
OAI221_X1 _10309_ ( .A(_02691_ ), .B1(_02695_ ), .B2(_02699_ ), .C1(_02326_ ), .C2(_02093_ ), .ZN(_02700_ ) );
OR3_X1 _10310_ ( .A1(_02035_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02701_ ) );
NAND2_X2 _10311_ ( .A1(_02700_ ), .A2(_02701_ ), .ZN(_02702_ ) );
INV_X1 _10312_ ( .A(\ID_EX_imm [11] ), .ZN(_02703_ ) );
XNOR2_X1 _10313_ ( .A(_02702_ ), .B(_02703_ ), .ZN(_02704_ ) );
OR2_X1 _10314_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02705_ ) );
OAI211_X1 _10315_ ( .A(_02705_ ), .B(_02214_ ), .C1(_02058_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02706_ ) );
OR2_X1 _10316_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02707_ ) );
OAI211_X1 _10317_ ( .A(_02707_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02058_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02708_ ) );
NAND3_X1 _10318_ ( .A1(_02706_ ), .A2(_02708_ ), .A3(_02332_ ), .ZN(_02709_ ) );
MUX2_X1 _10319_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02710_ ) );
MUX2_X1 _10320_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02711_ ) );
MUX2_X1 _10321_ ( .A(_02710_ ), .B(_02711_ ), .S(_02330_ ), .Z(_02712_ ) );
OAI211_X1 _10322_ ( .A(fanout_net_28 ), .B(_02709_ ), .C1(_02712_ ), .C2(_02105_ ), .ZN(_02713_ ) );
MUX2_X1 _10323_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02714_ ) );
AND2_X1 _10324_ ( .A1(_02714_ ), .A2(_02339_ ), .ZN(_02715_ ) );
MUX2_X1 _10325_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02716_ ) );
AOI211_X1 _10326_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_02715_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C2(_02716_ ), .ZN(_02717_ ) );
MUX2_X1 _10327_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02718_ ) );
MUX2_X1 _10328_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02719_ ) );
MUX2_X1 _10329_ ( .A(_02718_ ), .B(_02719_ ), .S(_02065_ ), .Z(_02720_ ) );
OAI21_X1 _10330_ ( .A(_02048_ ), .B1(_02720_ ), .B2(_02332_ ), .ZN(_02721_ ) );
OAI221_X1 _10331_ ( .A(_02713_ ), .B1(_02717_ ), .B2(_02721_ ), .C1(_02085_ ), .C2(_02093_ ), .ZN(_02722_ ) );
OR3_X1 _10332_ ( .A1(_02326_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02723_ ) );
NAND2_X1 _10333_ ( .A1(_02722_ ), .A2(_02723_ ), .ZN(_02724_ ) );
INV_X1 _10334_ ( .A(\ID_EX_imm [10] ), .ZN(_02725_ ) );
XNOR2_X1 _10335_ ( .A(_02724_ ), .B(_02725_ ), .ZN(_02726_ ) );
AND3_X1 _10336_ ( .A1(_02682_ ), .A2(_02704_ ), .A3(_02726_ ), .ZN(_02727_ ) );
AND3_X1 _10337_ ( .A1(_02539_ ), .A2(_02634_ ), .A3(_02727_ ), .ZN(_02728_ ) );
INV_X2 _10338_ ( .A(_02728_ ), .ZN(_02729_ ) );
XNOR2_X1 _10339_ ( .A(_02678_ ), .B(\ID_EX_imm [9] ), .ZN(_02730_ ) );
NAND2_X1 _10340_ ( .A1(_02655_ ), .A2(\ID_EX_imm [8] ), .ZN(_02731_ ) );
OAI21_X1 _10341_ ( .A(_02680_ ), .B1(_02730_ ), .B2(_02731_ ), .ZN(_02732_ ) );
AND3_X1 _10342_ ( .A1(_02732_ ), .A2(_02704_ ), .A3(_02726_ ), .ZN(_02733_ ) );
AOI21_X1 _10343_ ( .A(_02703_ ), .B1(_02700_ ), .B2(_02701_ ), .ZN(_02734_ ) );
AND2_X1 _10344_ ( .A1(_02724_ ), .A2(\ID_EX_imm [10] ), .ZN(_02735_ ) );
AND2_X1 _10345_ ( .A1(_02704_ ), .A2(_02735_ ), .ZN(_02736_ ) );
NOR3_X1 _10346_ ( .A1(_02733_ ), .A2(_02734_ ), .A3(_02736_ ), .ZN(_02737_ ) );
INV_X1 _10347_ ( .A(_02737_ ), .ZN(_02738_ ) );
NAND2_X1 _10348_ ( .A1(_02738_ ), .A2(_02634_ ), .ZN(_02739_ ) );
OAI211_X1 _10349_ ( .A(\ID_EX_imm [14] ), .B(_02631_ ), .C1(_02609_ ), .C2(\ID_EX_imm [15] ), .ZN(_02740_ ) );
NAND2_X1 _10350_ ( .A1(_02561_ ), .A2(\ID_EX_imm [12] ), .ZN(_02741_ ) );
NOR3_X1 _10351_ ( .A1(_02741_ ), .A2(_02585_ ), .A3(_02586_ ), .ZN(_02742_ ) );
OR2_X1 _10352_ ( .A1(_02742_ ), .A2(_02586_ ), .ZN(_02743_ ) );
AND2_X1 _10353_ ( .A1(_02610_ ), .A2(_02633_ ), .ZN(_02744_ ) );
AOI22_X1 _10354_ ( .A1(_02743_ ), .A2(_02744_ ), .B1(\ID_EX_imm [15] ), .B2(_02609_ ), .ZN(_02745_ ) );
AND3_X1 _10355_ ( .A1(_02739_ ), .A2(_02740_ ), .A3(_02745_ ), .ZN(_02746_ ) );
AOI211_X1 _10356_ ( .A(_02232_ ), .B(_02325_ ), .C1(_02729_ ), .C2(_02746_ ), .ZN(_02747_ ) );
AND2_X1 _10357_ ( .A1(_02322_ ), .A2(\ID_EX_imm [16] ), .ZN(_02748_ ) );
AND2_X1 _10358_ ( .A1(_02301_ ), .A2(_02748_ ), .ZN(_02749_ ) );
AOI21_X1 _10359_ ( .A(_02749_ ), .B1(\ID_EX_imm [17] ), .B2(_02299_ ), .ZN(_02750_ ) );
INV_X1 _10360_ ( .A(_02750_ ), .ZN(_02751_ ) );
NAND2_X1 _10361_ ( .A1(_02751_ ), .A2(_02278_ ), .ZN(_02752_ ) );
AND2_X1 _10362_ ( .A1(_02275_ ), .A2(\ID_EX_imm [18] ), .ZN(_02753_ ) );
AND2_X1 _10363_ ( .A1(_02254_ ), .A2(_02753_ ), .ZN(_02754_ ) );
AOI21_X1 _10364_ ( .A(_02754_ ), .B1(\ID_EX_imm [19] ), .B2(_02252_ ), .ZN(_02755_ ) );
AND2_X1 _10365_ ( .A1(_02752_ ), .A2(_02755_ ), .ZN(_02756_ ) );
OR2_X1 _10366_ ( .A1(_02756_ ), .A2(_02232_ ), .ZN(_02757_ ) );
NAND2_X1 _10367_ ( .A1(_02202_ ), .A2(\ID_EX_imm [20] ), .ZN(_02758_ ) );
NOR3_X1 _10368_ ( .A1(_02758_ ), .A2(_02228_ ), .A3(_02229_ ), .ZN(_02759_ ) );
OR2_X1 _10369_ ( .A1(_02759_ ), .A2(_02229_ ), .ZN(_02760_ ) );
NAND2_X1 _10370_ ( .A1(_02181_ ), .A2(_02760_ ), .ZN(_02761_ ) );
NAND4_X1 _10371_ ( .A1(_02180_ ), .A2(\ID_EX_imm [22] ), .A3(_02178_ ), .A4(_02155_ ), .ZN(_02762_ ) );
NAND4_X1 _10372_ ( .A1(_02757_ ), .A2(_02180_ ), .A3(_02761_ ), .A4(_02762_ ), .ZN(_02763_ ) );
OR2_X1 _10373_ ( .A1(_02747_ ), .A2(_02763_ ), .ZN(_02764_ ) );
OR3_X1 _10374_ ( .A1(_02087_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02095_ ), .ZN(_02765_ ) );
OR2_X1 _10375_ ( .A1(_02060_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02766_ ) );
BUF_X4 _10376_ ( .A(_02099_ ), .Z(_02767_ ) );
OAI211_X1 _10377_ ( .A(_02766_ ), .B(_02767_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02768_ ) );
OR2_X1 _10378_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02769_ ) );
BUF_X4 _10379_ ( .A(_02145_ ), .Z(_02770_ ) );
OAI211_X1 _10380_ ( .A(_02769_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02771_ ) );
NAND3_X1 _10381_ ( .A1(_02768_ ), .A2(_02107_ ), .A3(_02771_ ), .ZN(_02772_ ) );
MUX2_X1 _10382_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02773_ ) );
MUX2_X1 _10383_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02774_ ) );
MUX2_X1 _10384_ ( .A(_02773_ ), .B(_02774_ ), .S(_02100_ ), .Z(_02775_ ) );
OAI211_X1 _10385_ ( .A(_02050_ ), .B(_02772_ ), .C1(_02775_ ), .C2(_02074_ ), .ZN(_02776_ ) );
OR2_X1 _10386_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02777_ ) );
OAI211_X1 _10387_ ( .A(_02777_ ), .B(_02767_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02778_ ) );
NOR2_X1 _10388_ ( .A1(_02770_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02779_ ) );
OAI21_X1 _10389_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_23 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02780_ ) );
OAI211_X1 _10390_ ( .A(_02778_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_02779_ ), .C2(_02780_ ), .ZN(_02781_ ) );
MUX2_X1 _10391_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02782_ ) );
MUX2_X1 _10392_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02783_ ) );
MUX2_X1 _10393_ ( .A(_02782_ ), .B(_02783_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02784_ ) );
OAI211_X1 _10394_ ( .A(_02781_ ), .B(fanout_net_28 ), .C1(_02784_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02785_ ) );
OAI211_X1 _10395_ ( .A(_02776_ ), .B(_02785_ ), .C1(_02087_ ), .C2(_02088_ ), .ZN(_02786_ ) );
NAND2_X1 _10396_ ( .A1(_02765_ ), .A2(_02786_ ), .ZN(_02787_ ) );
INV_X1 _10397_ ( .A(\ID_EX_imm [24] ), .ZN(_02788_ ) );
XNOR2_X1 _10398_ ( .A(_02787_ ), .B(_02788_ ), .ZN(_02789_ ) );
AND2_X1 _10399_ ( .A1(_02764_ ), .A2(_02789_ ), .ZN(_02790_ ) );
AOI21_X1 _10400_ ( .A(_02788_ ), .B1(_02765_ ), .B2(_02786_ ), .ZN(_02791_ ) );
NOR2_X2 _10401_ ( .A1(_02790_ ), .A2(_02791_ ), .ZN(_02792_ ) );
OR3_X1 _10402_ ( .A1(_02037_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02095_ ), .ZN(_02793_ ) );
OR2_X1 _10403_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02794_ ) );
OAI211_X1 _10404_ ( .A(_02794_ ), .B(_02767_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02795_ ) );
INV_X1 _10405_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02796_ ) );
NAND2_X1 _10406_ ( .A1(_02796_ ), .A2(fanout_net_23 ), .ZN(_02797_ ) );
OAI211_X1 _10407_ ( .A(_02797_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02798_ ) );
NAND3_X1 _10408_ ( .A1(_02795_ ), .A2(_02798_ ), .A3(_02107_ ), .ZN(_02799_ ) );
MUX2_X1 _10409_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02800_ ) );
MUX2_X1 _10410_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02801_ ) );
MUX2_X1 _10411_ ( .A(_02800_ ), .B(_02801_ ), .S(_02100_ ), .Z(_02802_ ) );
OAI211_X1 _10412_ ( .A(_02050_ ), .B(_02799_ ), .C1(_02802_ ), .C2(_02074_ ), .ZN(_02803_ ) );
OR2_X1 _10413_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02804_ ) );
OAI211_X1 _10414_ ( .A(_02804_ ), .B(_02767_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02805_ ) );
OR2_X1 _10415_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02806_ ) );
OAI211_X1 _10416_ ( .A(_02806_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02807_ ) );
NAND3_X1 _10417_ ( .A1(_02805_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02807_ ), .ZN(_02808_ ) );
MUX2_X1 _10418_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02809_ ) );
MUX2_X1 _10419_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02810_ ) );
MUX2_X1 _10420_ ( .A(_02809_ ), .B(_02810_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02811_ ) );
OAI211_X1 _10421_ ( .A(fanout_net_28 ), .B(_02808_ ), .C1(_02811_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02812_ ) );
OAI211_X1 _10422_ ( .A(_02803_ ), .B(_02812_ ), .C1(_02087_ ), .C2(_02088_ ), .ZN(_02813_ ) );
NAND2_X1 _10423_ ( .A1(_02793_ ), .A2(_02813_ ), .ZN(_02814_ ) );
BUF_X2 _10424_ ( .A(_02814_ ), .Z(_02815_ ) );
NAND2_X1 _10425_ ( .A1(_02815_ ), .A2(\ID_EX_imm [25] ), .ZN(_02816_ ) );
NAND2_X1 _10426_ ( .A1(_02792_ ), .A2(_02816_ ), .ZN(_02817_ ) );
OR3_X1 _10427_ ( .A1(_02037_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02095_ ), .ZN(_02818_ ) );
INV_X1 _10428_ ( .A(\ID_EX_imm [27] ), .ZN(_02819_ ) );
OR2_X1 _10429_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02820_ ) );
OAI211_X1 _10430_ ( .A(_02820_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02821_ ) );
INV_X1 _10431_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02822_ ) );
NAND2_X1 _10432_ ( .A1(_02822_ ), .A2(fanout_net_23 ), .ZN(_02823_ ) );
OAI211_X1 _10433_ ( .A(_02823_ ), .B(_02100_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02824_ ) );
NAND3_X1 _10434_ ( .A1(_02821_ ), .A2(_02107_ ), .A3(_02824_ ), .ZN(_02825_ ) );
MUX2_X1 _10435_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02826_ ) );
MUX2_X1 _10436_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02827_ ) );
MUX2_X1 _10437_ ( .A(_02826_ ), .B(_02827_ ), .S(_02100_ ), .Z(_02828_ ) );
OAI211_X1 _10438_ ( .A(fanout_net_28 ), .B(_02825_ ), .C1(_02828_ ), .C2(_02074_ ), .ZN(_02829_ ) );
OR2_X1 _10439_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02830_ ) );
OAI211_X1 _10440_ ( .A(_02830_ ), .B(_02767_ ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02831_ ) );
OR2_X1 _10441_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02832_ ) );
OAI211_X1 _10442_ ( .A(_02832_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02833_ ) );
NAND3_X1 _10443_ ( .A1(_02831_ ), .A2(_02833_ ), .A3(_02107_ ), .ZN(_02834_ ) );
MUX2_X1 _10444_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02835_ ) );
MUX2_X1 _10445_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02836_ ) );
MUX2_X1 _10446_ ( .A(_02835_ ), .B(_02836_ ), .S(_02100_ ), .Z(_02837_ ) );
OAI211_X1 _10447_ ( .A(_02050_ ), .B(_02834_ ), .C1(_02837_ ), .C2(_02074_ ), .ZN(_02838_ ) );
OAI211_X1 _10448_ ( .A(_02829_ ), .B(_02838_ ), .C1(_02087_ ), .C2(_02088_ ), .ZN(_02839_ ) );
AND3_X1 _10449_ ( .A1(_02818_ ), .A2(_02819_ ), .A3(_02839_ ), .ZN(_02840_ ) );
AOI21_X1 _10450_ ( .A(_02819_ ), .B1(_02818_ ), .B2(_02839_ ), .ZN(_02841_ ) );
NOR2_X1 _10451_ ( .A1(_02840_ ), .A2(_02841_ ), .ZN(_02842_ ) );
OR2_X1 _10452_ ( .A1(_02060_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02843_ ) );
OAI211_X1 _10453_ ( .A(_02843_ ), .B(_02767_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02844_ ) );
OR2_X1 _10454_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02845_ ) );
OAI211_X1 _10455_ ( .A(_02845_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02846_ ) );
NAND3_X1 _10456_ ( .A1(_02844_ ), .A2(_02846_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02847_ ) );
MUX2_X1 _10457_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02848_ ) );
MUX2_X1 _10458_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02849_ ) );
MUX2_X1 _10459_ ( .A(_02848_ ), .B(_02849_ ), .S(_02767_ ), .Z(_02850_ ) );
OAI211_X1 _10460_ ( .A(_02050_ ), .B(_02847_ ), .C1(_02850_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02851_ ) );
INV_X1 _10461_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02852_ ) );
AOI21_X1 _10462_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(_02852_ ), .B2(fanout_net_24 ), .ZN(_02853_ ) );
OR2_X1 _10463_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02854_ ) );
MUX2_X1 _10464_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02855_ ) );
AOI221_X4 _10465_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B1(_02853_ ), .B2(_02854_ ), .C1(_02855_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_02856_ ) );
MUX2_X1 _10466_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02857_ ) );
MUX2_X1 _10467_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02858_ ) );
MUX2_X1 _10468_ ( .A(_02857_ ), .B(_02858_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02859_ ) );
OAI21_X1 _10469_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B1(_02859_ ), .B2(_02074_ ), .ZN(_02860_ ) );
BUF_X4 _10470_ ( .A(_02095_ ), .Z(_02861_ ) );
OAI221_X1 _10471_ ( .A(_02851_ ), .B1(_02856_ ), .B2(_02860_ ), .C1(_02087_ ), .C2(_02861_ ), .ZN(_02862_ ) );
OR3_X1 _10472_ ( .A1(_02037_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02095_ ), .ZN(_02863_ ) );
NAND2_X1 _10473_ ( .A1(_02862_ ), .A2(_02863_ ), .ZN(_02864_ ) );
INV_X1 _10474_ ( .A(\ID_EX_imm [26] ), .ZN(_02865_ ) );
XNOR2_X1 _10475_ ( .A(_02864_ ), .B(_02865_ ), .ZN(_02866_ ) );
INV_X1 _10476_ ( .A(\ID_EX_imm [25] ), .ZN(_02867_ ) );
NAND3_X1 _10477_ ( .A1(_02793_ ), .A2(_02867_ ), .A3(_02813_ ), .ZN(_02868_ ) );
NAND4_X1 _10478_ ( .A1(_02817_ ), .A2(_02842_ ), .A3(_02866_ ), .A4(_02868_ ), .ZN(_02869_ ) );
NAND2_X1 _10479_ ( .A1(_02864_ ), .A2(\ID_EX_imm [26] ), .ZN(_02870_ ) );
NOR3_X1 _10480_ ( .A1(_02870_ ), .A2(_02840_ ), .A3(_02841_ ), .ZN(_02871_ ) );
NOR2_X1 _10481_ ( .A1(_02871_ ), .A2(_02841_ ), .ZN(_02872_ ) );
AOI21_X2 _10482_ ( .A(_02126_ ), .B1(_02869_ ), .B2(_02872_ ), .ZN(_02873_ ) );
OR3_X1 _10483_ ( .A1(_02037_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02045_ ), .ZN(_02874_ ) );
OR2_X1 _10484_ ( .A1(_02137_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02875_ ) );
OAI211_X1 _10485_ ( .A(_02875_ ), .B(_02100_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02876_ ) );
OR2_X1 _10486_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02877_ ) );
OAI211_X1 _10487_ ( .A(_02877_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02878_ ) );
NAND3_X1 _10488_ ( .A1(_02876_ ), .A2(_02878_ ), .A3(_02107_ ), .ZN(_02879_ ) );
MUX2_X1 _10489_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02880_ ) );
MUX2_X1 _10490_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02881_ ) );
MUX2_X1 _10491_ ( .A(_02880_ ), .B(_02881_ ), .S(_02068_ ), .Z(_02882_ ) );
OAI211_X1 _10492_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02879_ ), .C1(_02882_ ), .C2(_02074_ ), .ZN(_02883_ ) );
OR2_X1 _10493_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02884_ ) );
OAI211_X1 _10494_ ( .A(_02884_ ), .B(_02100_ ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02885_ ) );
OR2_X1 _10495_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02886_ ) );
OAI211_X1 _10496_ ( .A(_02886_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02887_ ) );
NAND3_X1 _10497_ ( .A1(_02885_ ), .A2(_02887_ ), .A3(_02055_ ), .ZN(_02888_ ) );
MUX2_X1 _10498_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02889_ ) );
MUX2_X1 _10499_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02890_ ) );
MUX2_X1 _10500_ ( .A(_02889_ ), .B(_02890_ ), .S(_02068_ ), .Z(_02891_ ) );
OAI211_X1 _10501_ ( .A(_02050_ ), .B(_02888_ ), .C1(_02891_ ), .C2(_02107_ ), .ZN(_02892_ ) );
OAI211_X1 _10502_ ( .A(_02883_ ), .B(_02892_ ), .C1(_02087_ ), .C2(_02088_ ), .ZN(_02893_ ) );
NAND2_X1 _10503_ ( .A1(_02874_ ), .A2(_02893_ ), .ZN(_02894_ ) );
INV_X1 _10504_ ( .A(\ID_EX_imm [29] ), .ZN(_02895_ ) );
XNOR2_X1 _10505_ ( .A(_02894_ ), .B(_02895_ ), .ZN(_02896_ ) );
AND2_X1 _10506_ ( .A1(_02873_ ), .A2(_02896_ ), .ZN(_02897_ ) );
AOI21_X1 _10507_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02096_ ), .B2(_02124_ ), .ZN(_02898_ ) );
NAND2_X1 _10508_ ( .A1(_02896_ ), .A2(_02898_ ), .ZN(_02899_ ) );
INV_X1 _10509_ ( .A(_02894_ ), .ZN(_02900_ ) );
OAI21_X1 _10510_ ( .A(_02899_ ), .B1(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_02900_ ), .ZN(_02901_ ) );
OAI21_X2 _10511_ ( .A(_02092_ ), .B1(_02897_ ), .B2(_02901_ ), .ZN(_02902_ ) );
OR2_X1 _10512_ ( .A1(_02090_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02903_ ) );
AND2_X1 _10513_ ( .A1(_02902_ ), .A2(_02903_ ), .ZN(_02904_ ) );
NAND2_X1 _10514_ ( .A1(_02402_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02905_ ) );
OR2_X1 _10515_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02906_ ) );
OAI211_X1 _10516_ ( .A(_02906_ ), .B(_02767_ ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02907_ ) );
INV_X1 _10517_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02908_ ) );
NAND2_X1 _10518_ ( .A1(_02908_ ), .A2(fanout_net_24 ), .ZN(_02909_ ) );
OAI211_X1 _10519_ ( .A(_02909_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02910_ ) );
NAND3_X1 _10520_ ( .A1(_02907_ ), .A2(_02910_ ), .A3(_02107_ ), .ZN(_02911_ ) );
MUX2_X1 _10521_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02912_ ) );
MUX2_X1 _10522_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02913_ ) );
MUX2_X1 _10523_ ( .A(_02912_ ), .B(_02913_ ), .S(_02767_ ), .Z(_02914_ ) );
OAI211_X1 _10524_ ( .A(_02050_ ), .B(_02911_ ), .C1(_02914_ ), .C2(_02074_ ), .ZN(_02915_ ) );
OR2_X1 _10525_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02916_ ) );
OAI211_X1 _10526_ ( .A(_02916_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02770_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02917_ ) );
INV_X1 _10527_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02918_ ) );
NAND2_X1 _10528_ ( .A1(_02918_ ), .A2(fanout_net_24 ), .ZN(_02919_ ) );
OAI211_X1 _10529_ ( .A(_02919_ ), .B(_02767_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02920_ ) );
NAND3_X1 _10530_ ( .A1(_02917_ ), .A2(_02920_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02921_ ) );
MUX2_X1 _10531_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02922_ ) );
MUX2_X1 _10532_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02923_ ) );
MUX2_X1 _10533_ ( .A(_02922_ ), .B(_02923_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02924_ ) );
OAI211_X1 _10534_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02921_ ), .C1(_02924_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02925_ ) );
NAND2_X1 _10535_ ( .A1(_02915_ ), .A2(_02925_ ), .ZN(_02926_ ) );
OAI21_X1 _10536_ ( .A(_02926_ ), .B1(_02087_ ), .B2(_02861_ ), .ZN(_02927_ ) );
AND2_X2 _10537_ ( .A1(_02905_ ), .A2(_02927_ ), .ZN(_02928_ ) );
XNOR2_X1 _10538_ ( .A(_02928_ ), .B(\ID_EX_imm [31] ), .ZN(_02929_ ) );
XNOR2_X1 _10539_ ( .A(_02904_ ), .B(_02929_ ), .ZN(_02930_ ) );
AND2_X2 _10540_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_02931_ ) );
BUF_X4 _10541_ ( .A(_02931_ ), .Z(_02932_ ) );
NOR2_X1 _10542_ ( .A1(_02930_ ), .A2(_02932_ ), .ZN(_00097_ ) );
OR3_X1 _10543_ ( .A1(_02897_ ), .A2(_02901_ ), .A3(_02092_ ), .ZN(_02933_ ) );
INV_X1 _10544_ ( .A(_02931_ ), .ZN(_02934_ ) );
CLKBUF_X2 _10545_ ( .A(_02934_ ), .Z(_02935_ ) );
AND3_X1 _10546_ ( .A1(_02933_ ), .A2(_02935_ ), .A3(_02902_ ), .ZN(_00098_ ) );
AOI21_X1 _10547_ ( .A(_02325_ ), .B1(_02729_ ), .B2(_02746_ ), .ZN(_02936_ ) );
INV_X1 _10548_ ( .A(_02756_ ), .ZN(_02937_ ) );
OAI21_X1 _10549_ ( .A(_02204_ ), .B1(_02936_ ), .B2(_02937_ ), .ZN(_02938_ ) );
NAND2_X1 _10550_ ( .A1(_02938_ ), .A2(_02758_ ), .ZN(_02939_ ) );
XNOR2_X1 _10551_ ( .A(_02939_ ), .B(_02230_ ), .ZN(_02940_ ) );
NOR2_X1 _10552_ ( .A1(_02940_ ), .A2(_02932_ ), .ZN(_00099_ ) );
OR3_X1 _10553_ ( .A1(_02936_ ), .A2(_02204_ ), .A3(_02937_ ), .ZN(_02941_ ) );
AND3_X1 _10554_ ( .A1(_02941_ ), .A2(_02935_ ), .A3(_02938_ ), .ZN(_00100_ ) );
INV_X1 _10555_ ( .A(_02324_ ), .ZN(_02942_ ) );
AOI21_X1 _10556_ ( .A(_02942_ ), .B1(_02729_ ), .B2(_02746_ ), .ZN(_02943_ ) );
AND2_X1 _10557_ ( .A1(_02943_ ), .A2(_02301_ ), .ZN(_02944_ ) );
NOR2_X1 _10558_ ( .A1(_02944_ ), .A2(_02751_ ), .ZN(_02945_ ) );
AND3_X1 _10559_ ( .A1(_02255_ ), .A2(_02276_ ), .A3(_02274_ ), .ZN(_02946_ ) );
NOR3_X1 _10560_ ( .A1(_02945_ ), .A2(_02753_ ), .A3(_02946_ ), .ZN(_02947_ ) );
OR2_X1 _10561_ ( .A1(_02947_ ), .A2(_02753_ ), .ZN(_02948_ ) );
XNOR2_X1 _10562_ ( .A(_02948_ ), .B(_02254_ ), .ZN(_02949_ ) );
NOR2_X1 _10563_ ( .A1(_02949_ ), .A2(_02932_ ), .ZN(_00101_ ) );
XNOR2_X1 _10564_ ( .A(_02945_ ), .B(_02277_ ), .ZN(_02950_ ) );
AND2_X1 _10565_ ( .A1(_02950_ ), .A2(_02935_ ), .ZN(_00102_ ) );
OR2_X1 _10566_ ( .A1(_02943_ ), .A2(_02748_ ), .ZN(_02951_ ) );
XNOR2_X1 _10567_ ( .A(_02951_ ), .B(_02301_ ), .ZN(_02952_ ) );
NOR2_X1 _10568_ ( .A1(_02952_ ), .A2(_02932_ ), .ZN(_00103_ ) );
AND3_X1 _10569_ ( .A1(_02729_ ), .A2(_02746_ ), .A3(_02942_ ), .ZN(_02953_ ) );
NOR3_X1 _10570_ ( .A1(_02953_ ), .A2(_02943_ ), .A3(_02931_ ), .ZN(_00104_ ) );
INV_X1 _10571_ ( .A(_02588_ ), .ZN(_02954_ ) );
INV_X1 _10572_ ( .A(_02727_ ), .ZN(_02955_ ) );
AOI21_X1 _10573_ ( .A(_02955_ ), .B1(_02528_ ), .B2(_02538_ ), .ZN(_02956_ ) );
INV_X1 _10574_ ( .A(_02956_ ), .ZN(_02957_ ) );
AOI21_X1 _10575_ ( .A(_02954_ ), .B1(_02957_ ), .B2(_02737_ ), .ZN(_02958_ ) );
OR2_X1 _10576_ ( .A1(_02958_ ), .A2(_02743_ ), .ZN(_02959_ ) );
AND2_X1 _10577_ ( .A1(_02959_ ), .A2(_02633_ ), .ZN(_02960_ ) );
AND2_X1 _10578_ ( .A1(_02631_ ), .A2(\ID_EX_imm [14] ), .ZN(_02961_ ) );
OR2_X1 _10579_ ( .A1(_02960_ ), .A2(_02961_ ), .ZN(_02962_ ) );
XNOR2_X1 _10580_ ( .A(_02962_ ), .B(_02610_ ), .ZN(_02963_ ) );
NOR2_X1 _10581_ ( .A1(_02963_ ), .A2(_02932_ ), .ZN(_00105_ ) );
XOR2_X1 _10582_ ( .A(_02959_ ), .B(_02633_ ), .Z(_02964_ ) );
AND2_X1 _10583_ ( .A1(_02964_ ), .A2(_02935_ ), .ZN(_00106_ ) );
OAI21_X1 _10584_ ( .A(_02563_ ), .B1(_02956_ ), .B2(_02738_ ), .ZN(_02965_ ) );
NAND2_X1 _10585_ ( .A1(_02965_ ), .A2(_02741_ ), .ZN(_02966_ ) );
XNOR2_X1 _10586_ ( .A(_02966_ ), .B(_02587_ ), .ZN(_02967_ ) );
NOR2_X1 _10587_ ( .A1(_02967_ ), .A2(_02932_ ), .ZN(_00107_ ) );
OR3_X1 _10588_ ( .A1(_02956_ ), .A2(_02563_ ), .A3(_02738_ ), .ZN(_02968_ ) );
AND3_X1 _10589_ ( .A1(_02968_ ), .A2(_02935_ ), .A3(_02965_ ), .ZN(_00108_ ) );
OR2_X1 _10590_ ( .A1(_02873_ ), .A2(_02898_ ), .ZN(_02969_ ) );
XNOR2_X1 _10591_ ( .A(_02969_ ), .B(_02896_ ), .ZN(_02970_ ) );
NOR2_X1 _10592_ ( .A1(_02970_ ), .A2(_02932_ ), .ZN(_00109_ ) );
AND3_X1 _10593_ ( .A1(_02869_ ), .A2(_02872_ ), .A3(_02126_ ), .ZN(_02971_ ) );
NOR3_X1 _10594_ ( .A1(_02971_ ), .A2(_02873_ ), .A3(_02931_ ), .ZN(_00110_ ) );
NAND3_X1 _10595_ ( .A1(_02817_ ), .A2(_02866_ ), .A3(_02868_ ), .ZN(_02972_ ) );
NAND2_X1 _10596_ ( .A1(_02972_ ), .A2(_02870_ ), .ZN(_02973_ ) );
XNOR2_X1 _10597_ ( .A(_02973_ ), .B(_02842_ ), .ZN(_02974_ ) );
NOR2_X1 _10598_ ( .A1(_02974_ ), .A2(_02932_ ), .ZN(_00111_ ) );
NAND2_X1 _10599_ ( .A1(_02817_ ), .A2(_02868_ ), .ZN(_02975_ ) );
XNOR2_X1 _10600_ ( .A(_02975_ ), .B(_02866_ ), .ZN(_02976_ ) );
AND2_X1 _10601_ ( .A1(_02976_ ), .A2(_02935_ ), .ZN(_00112_ ) );
NAND2_X1 _10602_ ( .A1(_02816_ ), .A2(_02868_ ), .ZN(_02977_ ) );
XNOR2_X1 _10603_ ( .A(_02792_ ), .B(_02977_ ), .ZN(_02978_ ) );
NOR2_X1 _10604_ ( .A1(_02978_ ), .A2(_02932_ ), .ZN(_00113_ ) );
XOR2_X1 _10605_ ( .A(_02764_ ), .B(_02789_ ), .Z(_02979_ ) );
AND2_X1 _10606_ ( .A1(_02979_ ), .A2(_02935_ ), .ZN(_00114_ ) );
OAI21_X1 _10607_ ( .A(_02231_ ), .B1(_02936_ ), .B2(_02937_ ), .ZN(_02980_ ) );
INV_X1 _10608_ ( .A(_02980_ ), .ZN(_02981_ ) );
OAI21_X1 _10609_ ( .A(_02156_ ), .B1(_02981_ ), .B2(_02760_ ), .ZN(_02982_ ) );
NAND2_X1 _10610_ ( .A1(_02155_ ), .A2(\ID_EX_imm [22] ), .ZN(_02983_ ) );
AND4_X1 _10611_ ( .A1(_02178_ ), .A2(_02982_ ), .A3(_02180_ ), .A4(_02983_ ), .ZN(_02984_ ) );
AOI22_X1 _10612_ ( .A1(_02982_ ), .A2(_02983_ ), .B1(_02178_ ), .B2(_02180_ ), .ZN(_02985_ ) );
NOR2_X1 _10613_ ( .A1(_02984_ ), .A2(_02985_ ), .ZN(_02986_ ) );
NOR2_X1 _10614_ ( .A1(_02986_ ), .A2(_02932_ ), .ZN(_00115_ ) );
OR3_X1 _10615_ ( .A1(_02981_ ), .A2(_02156_ ), .A3(_02760_ ), .ZN(_02987_ ) );
AND3_X1 _10616_ ( .A1(_02987_ ), .A2(_02935_ ), .A3(_02982_ ), .ZN(_00116_ ) );
INV_X1 _10617_ ( .A(\IF_ID_inst [31] ), .ZN(_02988_ ) );
AND2_X1 _10618_ ( .A1(_02018_ ), .A2(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02989_ ) );
INV_X1 _10619_ ( .A(_02989_ ), .ZN(_02990_ ) );
BUF_X4 _10620_ ( .A(_02990_ ), .Z(_02991_ ) );
AND2_X1 _10621_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_02992_ ) );
AND2_X1 _10622_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_02993_ ) );
NOR2_X1 _10623_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_02994_ ) );
AND3_X1 _10624_ ( .A1(_02992_ ), .A2(_02993_ ), .A3(_02994_ ), .ZN(_02995_ ) );
AND2_X2 _10625_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_02996_ ) );
AND2_X1 _10626_ ( .A1(_02995_ ), .A2(_02996_ ), .ZN(_02997_ ) );
INV_X1 _10627_ ( .A(_02997_ ), .ZN(_02998_ ) );
INV_X1 _10628_ ( .A(\IF_ID_inst [6] ), .ZN(_02999_ ) );
NOR2_X1 _10629_ ( .A1(_02999_ ), .A2(\IF_ID_inst [12] ), .ZN(_03000_ ) );
AND3_X1 _10630_ ( .A1(_03000_ ), .A2(\IF_ID_inst [13] ), .A3(_02996_ ), .ZN(_03001_ ) );
AND2_X1 _10631_ ( .A1(_02992_ ), .A2(_02994_ ), .ZN(_03002_ ) );
BUF_X2 _10632_ ( .A(_03002_ ), .Z(_03003_ ) );
NAND2_X2 _10633_ ( .A1(_03001_ ), .A2(_03003_ ), .ZN(_03004_ ) );
AOI211_X1 _10634_ ( .A(_02988_ ), .B(_02991_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00195_ ) );
INV_X1 _10635_ ( .A(\IF_ID_inst [30] ), .ZN(_03005_ ) );
AOI211_X1 _10636_ ( .A(_03005_ ), .B(_02991_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00196_ ) );
INV_X1 _10637_ ( .A(\IF_ID_inst [21] ), .ZN(_03006_ ) );
AOI211_X1 _10638_ ( .A(_03006_ ), .B(_02991_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00197_ ) );
BUF_X4 _10639_ ( .A(_02990_ ), .Z(_03007_ ) );
BUF_X4 _10640_ ( .A(_03007_ ), .Z(_03008_ ) );
AND2_X1 _10641_ ( .A1(_02998_ ), .A2(_03004_ ), .ZN(_03009_ ) );
INV_X1 _10642_ ( .A(_03009_ ), .ZN(_03010_ ) );
INV_X1 _10643_ ( .A(\IF_ID_inst [20] ), .ZN(_03011_ ) );
AOI21_X1 _10644_ ( .A(_03008_ ), .B1(_03010_ ), .B2(_03011_ ), .ZN(_00198_ ) );
INV_X1 _10645_ ( .A(\IF_ID_inst [29] ), .ZN(_03012_ ) );
AOI21_X1 _10646_ ( .A(_03008_ ), .B1(_03010_ ), .B2(_03012_ ), .ZN(_00199_ ) );
INV_X1 _10647_ ( .A(\IF_ID_inst [28] ), .ZN(_03013_ ) );
AOI21_X1 _10648_ ( .A(_03008_ ), .B1(_03010_ ), .B2(_03013_ ), .ZN(_00200_ ) );
INV_X1 _10649_ ( .A(\IF_ID_inst [27] ), .ZN(_03014_ ) );
AOI211_X1 _10650_ ( .A(_03014_ ), .B(_02991_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00201_ ) );
INV_X1 _10651_ ( .A(\IF_ID_inst [26] ), .ZN(_03015_ ) );
AOI21_X1 _10652_ ( .A(_03008_ ), .B1(_03010_ ), .B2(_03015_ ), .ZN(_00202_ ) );
INV_X1 _10653_ ( .A(\IF_ID_inst [25] ), .ZN(_03016_ ) );
AOI211_X1 _10654_ ( .A(_03016_ ), .B(_03007_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00203_ ) );
INV_X1 _10655_ ( .A(\IF_ID_inst [24] ), .ZN(_03017_ ) );
AOI211_X1 _10656_ ( .A(_03017_ ), .B(_03007_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00204_ ) );
INV_X1 _10657_ ( .A(\IF_ID_inst [23] ), .ZN(_03018_ ) );
AOI211_X1 _10658_ ( .A(_03018_ ), .B(_03007_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00205_ ) );
INV_X1 _10659_ ( .A(\IF_ID_inst [22] ), .ZN(_03019_ ) );
AOI211_X1 _10660_ ( .A(_03019_ ), .B(_03007_ ), .C1(_02998_ ), .C2(_03004_ ), .ZN(_00206_ ) );
AND4_X1 _10661_ ( .A1(_01516_ ), .A2(_02017_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .A4(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00207_ ) );
AND4_X1 _10662_ ( .A1(_01459_ ), .A2(_02017_ ), .A3(\myidu.state [2] ), .A4(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_00208_ ) );
NOR4_X1 _10663_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .A4(\IF_ID_inst [31] ), .ZN(_03020_ ) );
NOR2_X1 _10664_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_03021_ ) );
NOR2_X1 _10665_ ( .A1(\IF_ID_inst [27] ), .A2(\IF_ID_inst [24] ), .ZN(_03022_ ) );
AND2_X1 _10666_ ( .A1(_03021_ ), .A2(_03022_ ), .ZN(_03023_ ) );
AND2_X1 _10667_ ( .A1(_03020_ ), .A2(_03023_ ), .ZN(_03024_ ) );
NOR2_X1 _10668_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_03025_ ) );
NOR2_X1 _10669_ ( .A1(\IF_ID_inst [7] ), .A2(\IF_ID_inst [15] ), .ZN(_03026_ ) );
AND4_X1 _10670_ ( .A1(_02996_ ), .A2(_03000_ ), .A3(_03025_ ), .A4(_03026_ ), .ZN(_03027_ ) );
INV_X1 _10671_ ( .A(\IF_ID_inst [8] ), .ZN(_03028_ ) );
NOR3_X1 _10672_ ( .A1(\IF_ID_inst [11] ), .A2(\IF_ID_inst [10] ), .A3(\IF_ID_inst [9] ), .ZN(_03029_ ) );
AND4_X1 _10673_ ( .A1(_03028_ ), .A2(_03029_ ), .A3(_02992_ ), .A4(_02994_ ), .ZN(_03030_ ) );
AND3_X1 _10674_ ( .A1(_03024_ ), .A2(_03027_ ), .A3(_03030_ ), .ZN(_03031_ ) );
NOR2_X1 _10675_ ( .A1(\IF_ID_inst [18] ), .A2(\IF_ID_inst [17] ), .ZN(_03032_ ) );
NOR2_X1 _10676_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [16] ), .ZN(_03033_ ) );
NOR2_X1 _10677_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_03034_ ) );
AND3_X1 _10678_ ( .A1(_03032_ ), .A2(_03033_ ), .A3(_03034_ ), .ZN(_03035_ ) );
AND3_X1 _10679_ ( .A1(_03035_ ), .A2(_03006_ ), .A3(\IF_ID_inst [20] ), .ZN(_03036_ ) );
AND2_X1 _10680_ ( .A1(_03031_ ), .A2(_03036_ ), .ZN(_03037_ ) );
INV_X1 _10681_ ( .A(\IF_ID_inst [5] ), .ZN(_03038_ ) );
NOR2_X4 _10682_ ( .A1(_03038_ ), .A2(\IF_ID_inst [4] ), .ZN(_03039_ ) );
AND3_X1 _10683_ ( .A1(_03000_ ), .A2(_03039_ ), .A3(_03025_ ), .ZN(_03040_ ) );
AND2_X1 _10684_ ( .A1(_03040_ ), .A2(_03003_ ), .ZN(_03041_ ) );
INV_X1 _10685_ ( .A(_03041_ ), .ZN(_03042_ ) );
NOR2_X1 _10686_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03043_ ) );
AND4_X1 _10687_ ( .A1(\IF_ID_inst [12] ), .A2(_03025_ ), .A3(_03043_ ), .A4(_02999_ ), .ZN(_03044_ ) );
AND3_X1 _10688_ ( .A1(_02992_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_03045_ ) );
AND2_X1 _10689_ ( .A1(_03044_ ), .A2(_03045_ ), .ZN(_03046_ ) );
INV_X1 _10690_ ( .A(_03046_ ), .ZN(_03047_ ) );
AND2_X1 _10691_ ( .A1(_03030_ ), .A2(_03027_ ), .ZN(_03048_ ) );
INV_X1 _10692_ ( .A(_03048_ ), .ZN(_03049_ ) );
NAND4_X1 _10693_ ( .A1(_03011_ ), .A2(_03018_ ), .A3(_03019_ ), .A4(\IF_ID_inst [29] ), .ZN(_03050_ ) );
NAND4_X1 _10694_ ( .A1(_03005_ ), .A2(_02988_ ), .A3(\IF_ID_inst [21] ), .A4(\IF_ID_inst [28] ), .ZN(_03051_ ) );
NOR2_X1 _10695_ ( .A1(_03050_ ), .A2(_03051_ ), .ZN(_03052_ ) );
AND2_X1 _10696_ ( .A1(_03032_ ), .A2(_03033_ ), .ZN(_03053_ ) );
AND3_X1 _10697_ ( .A1(_03052_ ), .A2(_03053_ ), .A3(_03023_ ), .ZN(_03054_ ) );
INV_X1 _10698_ ( .A(_03054_ ), .ZN(_03055_ ) );
OAI211_X1 _10699_ ( .A(_03042_ ), .B(_03047_ ), .C1(_03049_ ), .C2(_03055_ ), .ZN(_03056_ ) );
AND2_X1 _10700_ ( .A1(_02995_ ), .A2(_03039_ ), .ZN(_03057_ ) );
AND2_X1 _10701_ ( .A1(_03057_ ), .A2(\IF_ID_inst [14] ), .ZN(_03058_ ) );
AOI211_X1 _10702_ ( .A(_03037_ ), .B(_03056_ ), .C1(\IF_ID_inst [13] ), .C2(_03058_ ), .ZN(_03059_ ) );
CLKBUF_X2 _10703_ ( .A(_02989_ ), .Z(_03060_ ) );
NOR2_X1 _10704_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03061_ ) );
AND3_X1 _10705_ ( .A1(_03003_ ), .A2(_03039_ ), .A3(_03061_ ), .ZN(_03062_ ) );
INV_X1 _10706_ ( .A(\IF_ID_inst [13] ), .ZN(_03063_ ) );
NOR2_X1 _10707_ ( .A1(_03063_ ), .A2(\IF_ID_inst [14] ), .ZN(_03064_ ) );
AND2_X1 _10708_ ( .A1(_03062_ ), .A2(_03064_ ), .ZN(_03065_ ) );
INV_X1 _10709_ ( .A(_03065_ ), .ZN(_03066_ ) );
INV_X1 _10710_ ( .A(\IF_ID_inst [12] ), .ZN(_03067_ ) );
NOR2_X1 _10711_ ( .A1(_03067_ ), .A2(\IF_ID_inst [6] ), .ZN(_03068_ ) );
AND3_X1 _10712_ ( .A1(_03003_ ), .A2(_03039_ ), .A3(_03068_ ), .ZN(_03069_ ) );
OAI21_X1 _10713_ ( .A(_03025_ ), .B1(_03062_ ), .B2(_03069_ ), .ZN(_03070_ ) );
AND2_X1 _10714_ ( .A1(_03066_ ), .A2(_03070_ ), .ZN(_03071_ ) );
INV_X1 _10715_ ( .A(_03071_ ), .ZN(_03072_ ) );
AND2_X1 _10716_ ( .A1(_03000_ ), .A2(_03039_ ), .ZN(_03073_ ) );
AND2_X1 _10717_ ( .A1(_03073_ ), .A2(_03003_ ), .ZN(_03074_ ) );
AND2_X1 _10718_ ( .A1(_03074_ ), .A2(\IF_ID_inst [14] ), .ZN(_03075_ ) );
AND3_X1 _10719_ ( .A1(_02995_ ), .A2(_03063_ ), .A3(_03039_ ), .ZN(_03076_ ) );
OR2_X1 _10720_ ( .A1(_03075_ ), .A2(_03076_ ), .ZN(_03077_ ) );
NOR2_X1 _10721_ ( .A1(_03072_ ), .A2(_03077_ ), .ZN(_03078_ ) );
AND4_X1 _10722_ ( .A1(\IF_ID_inst [11] ), .A2(_03059_ ), .A3(_03060_ ), .A4(_03078_ ), .ZN(_00209_ ) );
AND4_X1 _10723_ ( .A1(\IF_ID_inst [10] ), .A2(_03059_ ), .A3(_03060_ ), .A4(_03078_ ), .ZN(_00210_ ) );
AND4_X1 _10724_ ( .A1(\IF_ID_inst [9] ), .A2(_03059_ ), .A3(_03060_ ), .A4(_03078_ ), .ZN(_00211_ ) );
AND4_X1 _10725_ ( .A1(\IF_ID_inst [8] ), .A2(_03059_ ), .A3(_03060_ ), .A4(_03078_ ), .ZN(_00212_ ) );
AND4_X1 _10726_ ( .A1(\IF_ID_inst [7] ), .A2(_03059_ ), .A3(_03060_ ), .A4(_03078_ ), .ZN(_00213_ ) );
AND3_X1 _10727_ ( .A1(_03052_ ), .A2(_03053_ ), .A3(_03023_ ), .ZN(_03079_ ) );
INV_X1 _10728_ ( .A(_03003_ ), .ZN(_03080_ ) );
NAND4_X1 _10729_ ( .A1(_03000_ ), .A2(_02996_ ), .A3(_03025_ ), .A4(_03026_ ), .ZN(_03081_ ) );
NAND2_X1 _10730_ ( .A1(_03029_ ), .A2(_03028_ ), .ZN(_03082_ ) );
NOR3_X1 _10731_ ( .A1(_03080_ ), .A2(_03081_ ), .A3(_03082_ ), .ZN(_03083_ ) );
AND2_X1 _10732_ ( .A1(_03079_ ), .A2(_03083_ ), .ZN(_03084_ ) );
INV_X1 _10733_ ( .A(_03039_ ), .ZN(_03085_ ) );
NOR2_X2 _10734_ ( .A1(_03085_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03086_ ) );
AND2_X1 _10735_ ( .A1(_03086_ ), .A2(_03045_ ), .ZN(_03087_ ) );
CLKBUF_X2 _10736_ ( .A(_03087_ ), .Z(_03088_ ) );
BUF_X2 _10737_ ( .A(_03088_ ), .Z(_03089_ ) );
NAND3_X1 _10738_ ( .A1(\IF_ID_inst [2] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [1] ), .ZN(_03090_ ) );
NOR2_X1 _10739_ ( .A1(_03090_ ), .A2(\IF_ID_inst [3] ), .ZN(_03091_ ) );
INV_X1 _10740_ ( .A(\IF_ID_inst [4] ), .ZN(_03092_ ) );
NOR2_X1 _10741_ ( .A1(_03092_ ), .A2(\IF_ID_inst [6] ), .ZN(_03093_ ) );
AND2_X1 _10742_ ( .A1(_03091_ ), .A2(_03093_ ), .ZN(_03094_ ) );
NOR3_X1 _10743_ ( .A1(_03084_ ), .A2(_03089_ ), .A3(_03094_ ), .ZN(_03095_ ) );
CLKBUF_X2 _10744_ ( .A(_02989_ ), .Z(_03096_ ) );
NAND3_X1 _10745_ ( .A1(_03083_ ), .A2(_03036_ ), .A3(_03024_ ), .ZN(_03097_ ) );
AND2_X1 _10746_ ( .A1(_03097_ ), .A2(_03047_ ), .ZN(_03098_ ) );
AND4_X1 _10747_ ( .A1(\IF_ID_inst [19] ), .A2(_03095_ ), .A3(_03096_ ), .A4(_03098_ ), .ZN(_00214_ ) );
AND4_X1 _10748_ ( .A1(\IF_ID_inst [18] ), .A2(_03095_ ), .A3(_03096_ ), .A4(_03098_ ), .ZN(_00215_ ) );
AND4_X1 _10749_ ( .A1(\IF_ID_inst [17] ), .A2(_03095_ ), .A3(_03096_ ), .A4(_03098_ ), .ZN(_00216_ ) );
XNOR2_X1 _10750_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_03099_ ) );
XNOR2_X1 _10751_ ( .A(\myexu.pc_jump [2] ), .B(\IF_ID_pc [2] ), .ZN(_03100_ ) );
XNOR2_X1 _10752_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_03101_ ) );
XNOR2_X1 _10753_ ( .A(fanout_net_8 ), .B(\myexu.pc_jump [3] ), .ZN(_03102_ ) );
AND4_X1 _10754_ ( .A1(_03099_ ), .A2(_03100_ ), .A3(_03101_ ), .A4(_03102_ ), .ZN(_03103_ ) );
XNOR2_X1 _10755_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_03104_ ) );
XNOR2_X1 _10756_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_03105_ ) );
XNOR2_X1 _10757_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_03106_ ) );
XNOR2_X1 _10758_ ( .A(fanout_net_12 ), .B(\myexu.pc_jump [4] ), .ZN(_03107_ ) );
AND4_X1 _10759_ ( .A1(_03104_ ), .A2(_03105_ ), .A3(_03106_ ), .A4(_03107_ ), .ZN(_03108_ ) );
XNOR2_X1 _10760_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_03109_ ) );
XNOR2_X1 _10761_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_03110_ ) );
XNOR2_X1 _10762_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_03111_ ) );
XNOR2_X1 _10763_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_03112_ ) );
AND4_X1 _10764_ ( .A1(_03109_ ), .A2(_03110_ ), .A3(_03111_ ), .A4(_03112_ ), .ZN(_03113_ ) );
XNOR2_X1 _10765_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_03114_ ) );
XNOR2_X1 _10766_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_03115_ ) );
XNOR2_X1 _10767_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_03116_ ) );
XNOR2_X1 _10768_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_03117_ ) );
AND4_X1 _10769_ ( .A1(_03114_ ), .A2(_03115_ ), .A3(_03116_ ), .A4(_03117_ ), .ZN(_03118_ ) );
AND4_X1 _10770_ ( .A1(_03103_ ), .A2(_03108_ ), .A3(_03113_ ), .A4(_03118_ ), .ZN(_03119_ ) );
XNOR2_X1 _10771_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_03120_ ) );
XNOR2_X1 _10772_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_03121_ ) );
XNOR2_X1 _10773_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_03122_ ) );
XNOR2_X1 _10774_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_03123_ ) );
AND4_X1 _10775_ ( .A1(_03120_ ), .A2(_03121_ ), .A3(_03122_ ), .A4(_03123_ ), .ZN(_03124_ ) );
XNOR2_X1 _10776_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_03125_ ) );
XNOR2_X1 _10777_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_03126_ ) );
XNOR2_X1 _10778_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_03127_ ) );
XNOR2_X1 _10779_ ( .A(\IF_ID_pc [25] ), .B(\myexu.pc_jump [25] ), .ZN(_03128_ ) );
AND4_X1 _10780_ ( .A1(_03125_ ), .A2(_03126_ ), .A3(_03127_ ), .A4(_03128_ ), .ZN(_03129_ ) );
XNOR2_X1 _10781_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_03130_ ) );
XNOR2_X1 _10782_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_03131_ ) );
XNOR2_X1 _10783_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_03132_ ) );
XNOR2_X1 _10784_ ( .A(\IF_ID_pc [21] ), .B(\myexu.pc_jump [21] ), .ZN(_03133_ ) );
AND4_X1 _10785_ ( .A1(_03130_ ), .A2(_03131_ ), .A3(_03132_ ), .A4(_03133_ ), .ZN(_03134_ ) );
XNOR2_X1 _10786_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_03135_ ) );
XNOR2_X1 _10787_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_03136_ ) );
XNOR2_X1 _10788_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_03137_ ) );
XNOR2_X1 _10789_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_03138_ ) );
AND4_X1 _10790_ ( .A1(_03135_ ), .A2(_03136_ ), .A3(_03137_ ), .A4(_03138_ ), .ZN(_03139_ ) );
AND4_X1 _10791_ ( .A1(_03124_ ), .A2(_03129_ ), .A3(_03134_ ), .A4(_03139_ ), .ZN(_03140_ ) );
AND2_X1 _10792_ ( .A1(_03119_ ), .A2(_03140_ ), .ZN(_03141_ ) );
INV_X1 _10793_ ( .A(check_quest ), .ZN(_03142_ ) );
NOR2_X1 _10794_ ( .A1(_03141_ ), .A2(_03142_ ), .ZN(_03143_ ) );
INV_X1 _10795_ ( .A(\myifu.state [1] ), .ZN(_03144_ ) );
NOR2_X1 _10796_ ( .A1(_03144_ ), .A2(fanout_net_43 ), .ZN(_03145_ ) );
INV_X1 _10797_ ( .A(_03145_ ), .ZN(_03146_ ) );
NOR2_X1 _10798_ ( .A1(_03143_ ), .A2(_03146_ ), .ZN(_03147_ ) );
AND2_X1 _10799_ ( .A1(_03147_ ), .A2(IDU_ready_IFU ), .ZN(_03148_ ) );
INV_X1 _10800_ ( .A(_03148_ ), .ZN(_03149_ ) );
BUF_X4 _10801_ ( .A(_03149_ ), .Z(_03150_ ) );
AND2_X1 _10802_ ( .A1(_03095_ ), .A2(_03098_ ), .ZN(_03151_ ) );
NOR3_X1 _10803_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_03152_ ) );
AND2_X1 _10804_ ( .A1(_03152_ ), .A2(_03014_ ), .ZN(_03153_ ) );
AND2_X2 _10805_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_03154_ ) );
AND3_X1 _10806_ ( .A1(_03153_ ), .A2(_03154_ ), .A3(_03021_ ), .ZN(_03155_ ) );
AND2_X1 _10807_ ( .A1(_03155_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03156_ ) );
AND4_X1 _10808_ ( .A1(\IF_ID_inst [4] ), .A2(_02999_ ), .A3(\IF_ID_inst [5] ), .A4(\IF_ID_inst [12] ), .ZN(_03157_ ) );
AND2_X2 _10809_ ( .A1(_03003_ ), .A2(_03157_ ), .ZN(_03158_ ) );
NAND2_X1 _10810_ ( .A1(_03156_ ), .A2(_03158_ ), .ZN(_03159_ ) );
AND2_X1 _10811_ ( .A1(_03002_ ), .A2(_03061_ ), .ZN(_03160_ ) );
BUF_X2 _10812_ ( .A(_03160_ ), .Z(_03161_ ) );
AND2_X1 _10813_ ( .A1(_03161_ ), .A2(_02996_ ), .ZN(_03162_ ) );
NAND2_X1 _10814_ ( .A1(_03156_ ), .A2(_03162_ ), .ZN(_03163_ ) );
NOR2_X1 _10815_ ( .A1(_03005_ ), .A2(\IF_ID_inst [29] ), .ZN(_03164_ ) );
NOR2_X1 _10816_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_03165_ ) );
AND3_X1 _10817_ ( .A1(_03164_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03165_ ), .ZN(_03166_ ) );
INV_X1 _10818_ ( .A(\IF_ID_inst [14] ), .ZN(_03167_ ) );
NOR2_X1 _10819_ ( .A1(_03167_ ), .A2(\IF_ID_inst [13] ), .ZN(_03168_ ) );
AND2_X1 _10820_ ( .A1(_03168_ ), .A2(_03021_ ), .ZN(_03169_ ) );
AND2_X1 _10821_ ( .A1(_03166_ ), .A2(_03169_ ), .ZN(_03170_ ) );
AND2_X1 _10822_ ( .A1(_03170_ ), .A2(_03158_ ), .ZN(_03171_ ) );
INV_X1 _10823_ ( .A(_03171_ ), .ZN(_03172_ ) );
AND3_X1 _10824_ ( .A1(_03152_ ), .A2(_03014_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03173_ ) );
AND2_X1 _10825_ ( .A1(_03025_ ), .A2(_03021_ ), .ZN(_03174_ ) );
AND2_X1 _10826_ ( .A1(_03173_ ), .A2(_03174_ ), .ZN(_03175_ ) );
AND2_X1 _10827_ ( .A1(_03173_ ), .A2(_03169_ ), .ZN(_03176_ ) );
OAI211_X1 _10828_ ( .A(_02996_ ), .B(_03161_ ), .C1(_03175_ ), .C2(_03176_ ), .ZN(_03177_ ) );
NAND4_X1 _10829_ ( .A1(_03159_ ), .A2(_03163_ ), .A3(_03172_ ), .A4(_03177_ ), .ZN(_03178_ ) );
AND4_X1 _10830_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A2(_03021_ ), .A3(\IF_ID_inst [13] ), .A4(_03167_ ), .ZN(_03179_ ) );
AND2_X1 _10831_ ( .A1(_03153_ ), .A2(_03179_ ), .ZN(_03180_ ) );
OR3_X1 _10832_ ( .A1(_03175_ ), .A2(_03176_ ), .A3(_03180_ ), .ZN(_03181_ ) );
AND2_X1 _10833_ ( .A1(_03181_ ), .A2(_03158_ ), .ZN(_03182_ ) );
NOR2_X1 _10834_ ( .A1(_03178_ ), .A2(_03182_ ), .ZN(_03183_ ) );
INV_X1 _10835_ ( .A(_03183_ ), .ZN(_03184_ ) );
AND2_X1 _10836_ ( .A1(_03160_ ), .A2(_03043_ ), .ZN(_03185_ ) );
AOI21_X1 _10837_ ( .A(_03041_ ), .B1(_03185_ ), .B2(_03064_ ), .ZN(_03186_ ) );
BUF_X2 _10838_ ( .A(_03009_ ), .Z(_03187_ ) );
NAND2_X1 _10839_ ( .A1(_03186_ ), .A2(_03187_ ), .ZN(_03188_ ) );
NOR4_X1 _10840_ ( .A1(_03184_ ), .A2(_03077_ ), .A3(_03072_ ), .A4(_03188_ ), .ZN(_03189_ ) );
AND3_X1 _10841_ ( .A1(_03180_ ), .A2(_02996_ ), .A3(_03161_ ), .ZN(_03190_ ) );
INV_X1 _10842_ ( .A(_03190_ ), .ZN(_03191_ ) );
AND4_X1 _10843_ ( .A1(_02996_ ), .A2(_03161_ ), .A3(_03174_ ), .A4(_03166_ ), .ZN(_03192_ ) );
INV_X1 _10844_ ( .A(_03192_ ), .ZN(_03193_ ) );
NAND4_X1 _10845_ ( .A1(_03038_ ), .A2(_02999_ ), .A3(\IF_ID_inst [4] ), .A4(\IF_ID_inst [12] ), .ZN(_03194_ ) );
NOR2_X1 _10846_ ( .A1(_03080_ ), .A2(_03194_ ), .ZN(_03195_ ) );
BUF_X2 _10847_ ( .A(_03195_ ), .Z(_03196_ ) );
AND2_X1 _10848_ ( .A1(_03196_ ), .A2(_03154_ ), .ZN(_03197_ ) );
INV_X1 _10849_ ( .A(_03197_ ), .ZN(_03198_ ) );
INV_X1 _10850_ ( .A(_03064_ ), .ZN(_03199_ ) );
NOR2_X1 _10851_ ( .A1(_03092_ ), .A2(\IF_ID_inst [5] ), .ZN(_03200_ ) );
NAND3_X1 _10852_ ( .A1(_03161_ ), .A2(_03199_ ), .A3(_03200_ ), .ZN(_03201_ ) );
AND4_X1 _10853_ ( .A1(_03191_ ), .A2(_03193_ ), .A3(_03198_ ), .A4(_03201_ ), .ZN(_03202_ ) );
AND3_X1 _10854_ ( .A1(_03003_ ), .A2(_03068_ ), .A3(_03043_ ), .ZN(_03203_ ) );
NAND2_X1 _10855_ ( .A1(_03203_ ), .A2(_03063_ ), .ZN(_03204_ ) );
NAND3_X1 _10856_ ( .A1(_03196_ ), .A2(\IF_ID_inst [13] ), .A3(_03167_ ), .ZN(_03205_ ) );
NAND3_X1 _10857_ ( .A1(_03161_ ), .A2(_03063_ ), .A3(_03043_ ), .ZN(_03206_ ) );
NAND3_X1 _10858_ ( .A1(_03161_ ), .A2(_03064_ ), .A3(_03200_ ), .ZN(_03207_ ) );
AND4_X1 _10859_ ( .A1(_03204_ ), .A2(_03205_ ), .A3(_03206_ ), .A4(_03207_ ), .ZN(_03208_ ) );
NAND3_X1 _10860_ ( .A1(_02995_ ), .A2(_03154_ ), .A3(_03039_ ), .ZN(_03209_ ) );
OAI211_X1 _10861_ ( .A(_03196_ ), .B(_03169_ ), .C1(_03166_ ), .C2(_03173_ ), .ZN(_03210_ ) );
AND2_X1 _10862_ ( .A1(_03040_ ), .A2(_03091_ ), .ZN(_03211_ ) );
INV_X1 _10863_ ( .A(_03211_ ), .ZN(_03212_ ) );
NAND2_X1 _10864_ ( .A1(_03175_ ), .A2(_03195_ ), .ZN(_03213_ ) );
AND4_X1 _10865_ ( .A1(_03209_ ), .A2(_03210_ ), .A3(_03212_ ), .A4(_03213_ ), .ZN(_03214_ ) );
AND4_X1 _10866_ ( .A1(_03151_ ), .A2(_03202_ ), .A3(_03208_ ), .A4(_03214_ ), .ZN(_03215_ ) );
AOI221_X4 _10867_ ( .A(_03150_ ), .B1(\IF_ID_inst [18] ), .B2(_03151_ ), .C1(_03189_ ), .C2(_03215_ ), .ZN(_03216_ ) );
AND2_X2 _10868_ ( .A1(_03189_ ), .A2(_03215_ ), .ZN(_03217_ ) );
NOR2_X1 _10869_ ( .A1(_03217_ ), .A2(_03150_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _10870_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_03218_ ) );
AOI211_X1 _10871_ ( .A(_03007_ ), .B(_03216_ ), .C1(_03218_ ), .C2(_02023_ ), .ZN(_00217_ ) );
AND4_X1 _10872_ ( .A1(\IF_ID_inst [16] ), .A2(_03095_ ), .A3(_03096_ ), .A4(_03098_ ), .ZN(_00218_ ) );
AOI221_X4 _10873_ ( .A(_03150_ ), .B1(\IF_ID_inst [17] ), .B2(_03151_ ), .C1(_03189_ ), .C2(_03215_ ), .ZN(_03219_ ) );
AOI211_X1 _10874_ ( .A(_03007_ ), .B(_03219_ ), .C1(_03218_ ), .C2(_02021_ ), .ZN(_00219_ ) );
AND4_X1 _10875_ ( .A1(\IF_ID_inst [15] ), .A2(_03095_ ), .A3(_03096_ ), .A4(_03098_ ), .ZN(_00220_ ) );
INV_X1 _10876_ ( .A(_03217_ ), .ZN(_03220_ ) );
NAND4_X1 _10877_ ( .A1(_03220_ ), .A2(\IF_ID_inst [16] ), .A3(_03151_ ), .A4(_03148_ ), .ZN(_03221_ ) );
OAI21_X1 _10878_ ( .A(\ID_EX_rs1 [1] ), .B1(_03217_ ), .B2(_03150_ ), .ZN(_03222_ ) );
AOI21_X1 _10879_ ( .A(_03008_ ), .B1(_03221_ ), .B2(_03222_ ), .ZN(_00221_ ) );
AND2_X1 _10880_ ( .A1(_03048_ ), .A2(_03054_ ), .ZN(_03223_ ) );
NOR2_X1 _10881_ ( .A1(_03223_ ), .A2(_03046_ ), .ZN(_03224_ ) );
INV_X1 _10882_ ( .A(_03224_ ), .ZN(_03225_ ) );
NAND2_X1 _10883_ ( .A1(_03196_ ), .A2(\IF_ID_inst [13] ), .ZN(_03226_ ) );
NAND2_X1 _10884_ ( .A1(_03226_ ), .A2(_03201_ ), .ZN(_03227_ ) );
NOR4_X1 _10885_ ( .A1(_03225_ ), .A2(_03010_ ), .A3(_03037_ ), .A4(_03227_ ), .ZN(_03228_ ) );
AND2_X1 _10886_ ( .A1(_03185_ ), .A2(_03064_ ), .ZN(_03229_ ) );
NOR3_X1 _10887_ ( .A1(_03229_ ), .A2(_03089_ ), .A3(_03211_ ), .ZN(_03230_ ) );
AND2_X1 _10888_ ( .A1(_03206_ ), .A2(_03204_ ), .ZN(_03231_ ) );
NAND4_X1 _10889_ ( .A1(_03195_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03153_ ), .A4(_03169_ ), .ZN(_03232_ ) );
NAND2_X1 _10890_ ( .A1(_03170_ ), .A2(_03196_ ), .ZN(_03233_ ) );
NAND3_X1 _10891_ ( .A1(_03232_ ), .A2(_03213_ ), .A3(_03233_ ), .ZN(_03234_ ) );
INV_X1 _10892_ ( .A(_03094_ ), .ZN(_03235_ ) );
NAND2_X1 _10893_ ( .A1(_03207_ ), .A2(_03235_ ), .ZN(_03236_ ) );
NOR2_X1 _10894_ ( .A1(_03234_ ), .A2(_03236_ ), .ZN(_03237_ ) );
AND3_X1 _10895_ ( .A1(_03230_ ), .A2(_03231_ ), .A3(_03237_ ), .ZN(_03238_ ) );
AND4_X1 _10896_ ( .A1(\IF_ID_inst [24] ), .A2(_03228_ ), .A3(_03096_ ), .A4(_03238_ ), .ZN(_00222_ ) );
NAND4_X1 _10897_ ( .A1(_03220_ ), .A2(\IF_ID_inst [15] ), .A3(_03151_ ), .A4(_03148_ ), .ZN(_03239_ ) );
OAI21_X1 _10898_ ( .A(\ID_EX_rs1 [0] ), .B1(_03217_ ), .B2(_03150_ ), .ZN(_03240_ ) );
AOI21_X1 _10899_ ( .A(_03008_ ), .B1(_03239_ ), .B2(_03240_ ), .ZN(_00223_ ) );
AND4_X1 _10900_ ( .A1(\IF_ID_inst [23] ), .A2(_03228_ ), .A3(_03096_ ), .A4(_03238_ ), .ZN(_00224_ ) );
AND4_X1 _10901_ ( .A1(\IF_ID_inst [22] ), .A2(_03228_ ), .A3(_03096_ ), .A4(_03238_ ), .ZN(_00225_ ) );
AND2_X1 _10902_ ( .A1(_03228_ ), .A2(_03238_ ), .ZN(_03241_ ) );
NAND4_X1 _10903_ ( .A1(_03220_ ), .A2(\IF_ID_inst [23] ), .A3(_03148_ ), .A4(_03241_ ), .ZN(_03242_ ) );
OAI21_X1 _10904_ ( .A(\ID_EX_rs2 [3] ), .B1(_03217_ ), .B2(_03150_ ), .ZN(_03243_ ) );
AOI21_X1 _10905_ ( .A(_03008_ ), .B1(_03242_ ), .B2(_03243_ ), .ZN(_00226_ ) );
AND4_X1 _10906_ ( .A1(\IF_ID_inst [21] ), .A2(_03228_ ), .A3(_03096_ ), .A4(_03238_ ), .ZN(_00227_ ) );
NAND4_X1 _10907_ ( .A1(_03220_ ), .A2(\IF_ID_inst [22] ), .A3(_03148_ ), .A4(_03241_ ), .ZN(_03244_ ) );
OAI21_X1 _10908_ ( .A(\ID_EX_rs2 [2] ), .B1(_03217_ ), .B2(_03150_ ), .ZN(_03245_ ) );
AOI21_X1 _10909_ ( .A(_03008_ ), .B1(_03244_ ), .B2(_03245_ ), .ZN(_00228_ ) );
AND4_X1 _10910_ ( .A1(\IF_ID_inst [20] ), .A2(_03228_ ), .A3(_03096_ ), .A4(_03238_ ), .ZN(_00229_ ) );
AOI221_X4 _10911_ ( .A(_03149_ ), .B1(_03241_ ), .B2(\IF_ID_inst [21] ), .C1(_03189_ ), .C2(_03215_ ), .ZN(_03246_ ) );
INV_X1 _10912_ ( .A(\ID_EX_rs2 [1] ), .ZN(_03247_ ) );
AOI211_X1 _10913_ ( .A(_03007_ ), .B(_03246_ ), .C1(_03218_ ), .C2(_03247_ ), .ZN(_00230_ ) );
INV_X1 _10914_ ( .A(IDU_valid_EXU ), .ZN(_03248_ ) );
AND4_X1 _10915_ ( .A1(_03248_ ), .A2(_03060_ ), .A3(_03045_ ), .A4(_03044_ ), .ZN(_00231_ ) );
AOI221_X4 _10916_ ( .A(_03149_ ), .B1(_03241_ ), .B2(\IF_ID_inst [20] ), .C1(_03189_ ), .C2(_03215_ ), .ZN(_03249_ ) );
INV_X16 _10917_ ( .A(\ID_EX_rs2 [0] ), .ZN(_03250_ ) );
AOI211_X1 _10918_ ( .A(_03007_ ), .B(_03249_ ), .C1(_03218_ ), .C2(_03250_ ), .ZN(_00232_ ) );
XNOR2_X1 _10919_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_03251_ ) );
XNOR2_X1 _10920_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_03252_ ) );
XNOR2_X1 _10921_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_03253_ ) );
XNOR2_X1 _10922_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_03254_ ) );
AND4_X1 _10923_ ( .A1(_03251_ ), .A2(_03252_ ), .A3(_03253_ ), .A4(_03254_ ), .ZN(_03255_ ) );
XNOR2_X1 _10924_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_03256_ ) );
AND2_X1 _10925_ ( .A1(_03255_ ), .A2(_03256_ ), .ZN(_03257_ ) );
AND2_X1 _10926_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03258_ ) );
INV_X1 _10927_ ( .A(\ID_EX_typ [7] ), .ZN(_03259_ ) );
AND2_X1 _10928_ ( .A1(_03258_ ), .A2(_03259_ ), .ZN(_03260_ ) );
AND2_X1 _10929_ ( .A1(_03257_ ), .A2(_03260_ ), .ZN(_03261_ ) );
XNOR2_X1 _10930_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_03262_ ) );
XNOR2_X1 _10931_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_03263_ ) );
XNOR2_X1 _10932_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_03264_ ) );
NAND4_X1 _10933_ ( .A1(_03260_ ), .A2(_03262_ ), .A3(_03263_ ), .A4(_03264_ ), .ZN(_03265_ ) );
XOR2_X1 _10934_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .Z(_03266_ ) );
XOR2_X1 _10935_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .Z(_03267_ ) );
NOR3_X1 _10936_ ( .A1(_03265_ ), .A2(_03266_ ), .A3(_03267_ ), .ZN(_03268_ ) );
NOR2_X1 _10937_ ( .A1(_03261_ ), .A2(_03268_ ), .ZN(_03269_ ) );
INV_X1 _10938_ ( .A(_03269_ ), .ZN(_03270_ ) );
AND2_X1 _10939_ ( .A1(_03151_ ), .A2(_03270_ ), .ZN(_03271_ ) );
INV_X1 _10940_ ( .A(_03154_ ), .ZN(_03272_ ) );
NAND3_X1 _10941_ ( .A1(_03161_ ), .A2(_03272_ ), .A3(_03043_ ), .ZN(_03273_ ) );
AND3_X1 _10942_ ( .A1(_03212_ ), .A2(_03204_ ), .A3(_03273_ ), .ZN(_03274_ ) );
NAND3_X1 _10943_ ( .A1(_03274_ ), .A2(_03198_ ), .A3(_03201_ ), .ZN(_03275_ ) );
NAND2_X1 _10944_ ( .A1(_03196_ ), .A2(_03064_ ), .ZN(_03276_ ) );
NAND2_X1 _10945_ ( .A1(_03276_ ), .A2(_03207_ ), .ZN(_03277_ ) );
NOR2_X2 _10946_ ( .A1(_03275_ ), .A2(_03277_ ), .ZN(_03278_ ) );
INV_X1 _10947_ ( .A(_03278_ ), .ZN(_03279_ ) );
NOR3_X1 _10948_ ( .A1(_03271_ ), .A2(_03010_ ), .A3(_03279_ ), .ZN(_03280_ ) );
AOI21_X1 _10949_ ( .A(_03261_ ), .B1(_03278_ ), .B2(_03187_ ), .ZN(_03281_ ) );
INV_X1 _10950_ ( .A(IDU_ready_IFU ), .ZN(_03282_ ) );
NOR4_X1 _10951_ ( .A1(_03280_ ), .A2(_03281_ ), .A3(_03282_ ), .A4(_03007_ ), .ZN(_00233_ ) );
AND3_X1 _10952_ ( .A1(_03035_ ), .A2(_03006_ ), .A3(_03011_ ), .ZN(_03283_ ) );
AND3_X1 _10953_ ( .A1(_03048_ ), .A2(_03024_ ), .A3(_03283_ ), .ZN(_03284_ ) );
NOR2_X1 _10954_ ( .A1(_03010_ ), .A2(_03284_ ), .ZN(_03285_ ) );
INV_X1 _10955_ ( .A(_03089_ ), .ZN(_03286_ ) );
AND4_X1 _10956_ ( .A1(_03224_ ), .A2(_03285_ ), .A3(_03286_ ), .A4(_03212_ ), .ZN(_03287_ ) );
OAI21_X1 _10957_ ( .A(\IF_ID_inst [14] ), .B1(_03074_ ), .B2(_03057_ ), .ZN(_03288_ ) );
AND3_X1 _10958_ ( .A1(_02995_ ), .A2(_03025_ ), .A3(_03039_ ), .ZN(_03289_ ) );
NOR2_X1 _10959_ ( .A1(_03041_ ), .A2(_03289_ ), .ZN(_03290_ ) );
AND2_X1 _10960_ ( .A1(_03288_ ), .A2(_03290_ ), .ZN(_03291_ ) );
AOI21_X1 _10961_ ( .A(_03008_ ), .B1(_03287_ ), .B2(_03291_ ), .ZN(_00234_ ) );
NAND2_X1 _10962_ ( .A1(_03203_ ), .A2(_03168_ ), .ZN(_03292_ ) );
AOI22_X1 _10963_ ( .A1(_03185_ ), .A2(_03272_ ), .B1(_03025_ ), .B2(_03203_ ), .ZN(_03293_ ) );
AND3_X1 _10964_ ( .A1(_03071_ ), .A2(_03292_ ), .A3(_03293_ ), .ZN(_03294_ ) );
AOI21_X1 _10965_ ( .A(_03008_ ), .B1(_03294_ ), .B2(_03285_ ), .ZN(_00235_ ) );
NOR2_X1 _10966_ ( .A1(_03190_ ), .A2(_03192_ ), .ZN(_03295_ ) );
INV_X1 _10967_ ( .A(_03295_ ), .ZN(_03296_ ) );
NOR4_X1 _10968_ ( .A1(_03184_ ), .A2(_03296_ ), .A3(_03227_ ), .A4(_03284_ ), .ZN(_03297_ ) );
AOI21_X1 _10969_ ( .A(_02991_ ), .B1(_03297_ ), .B2(_03238_ ), .ZN(_00236_ ) );
AND3_X1 _10970_ ( .A1(_03226_ ), .A2(_03047_ ), .A3(_03201_ ), .ZN(_03298_ ) );
AOI21_X1 _10971_ ( .A(_02991_ ), .B1(_03237_ ), .B2(_03298_ ), .ZN(_00237_ ) );
NOR4_X1 _10972_ ( .A1(_03190_ ), .A2(_03236_ ), .A3(_03192_ ), .A4(_03065_ ), .ZN(_03299_ ) );
INV_X1 _10973_ ( .A(_03084_ ), .ZN(_03300_ ) );
AOI21_X1 _10974_ ( .A(_02991_ ), .B1(_03299_ ), .B2(_03300_ ), .ZN(_00238_ ) );
AOI211_X1 _10975_ ( .A(_03058_ ), .B(_03234_ ), .C1(\IF_ID_inst [13] ), .C2(_02997_ ), .ZN(_03301_ ) );
OAI21_X1 _10976_ ( .A(_03064_ ), .B1(_03185_ ), .B2(_03196_ ), .ZN(_03302_ ) );
AOI21_X1 _10977_ ( .A(_03171_ ), .B1(_03181_ ), .B2(_03158_ ), .ZN(_03303_ ) );
AND4_X1 _10978_ ( .A1(_03235_ ), .A2(_03301_ ), .A3(_03302_ ), .A4(_03303_ ), .ZN(_03304_ ) );
AOI21_X1 _10979_ ( .A(_02991_ ), .B1(_03304_ ), .B2(_03066_ ), .ZN(_00239_ ) );
AND2_X1 _10980_ ( .A1(_03069_ ), .A2(_03025_ ), .ZN(_03305_ ) );
AND3_X1 _10981_ ( .A1(_02999_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_03306_ ) );
AOI221_X4 _10982_ ( .A(_03305_ ), .B1(_03025_ ), .B2(_03203_ ), .C1(_03091_ ), .C2(_03306_ ), .ZN(_03307_ ) );
NAND3_X1 _10983_ ( .A1(_03176_ ), .A2(_02996_ ), .A3(_03161_ ), .ZN(_03308_ ) );
AND4_X1 _10984_ ( .A1(_03066_ ), .A2(_03307_ ), .A3(_03292_ ), .A4(_03308_ ), .ZN(_03309_ ) );
AND2_X1 _10985_ ( .A1(_03161_ ), .A2(_03200_ ), .ZN(_03310_ ) );
NAND2_X1 _10986_ ( .A1(_03310_ ), .A2(\IF_ID_inst [14] ), .ZN(_03311_ ) );
OAI22_X1 _10987_ ( .A1(_03176_ ), .A2(_03170_ ), .B1(_03196_ ), .B2(_03158_ ), .ZN(_03312_ ) );
AOI22_X1 _10988_ ( .A1(_03074_ ), .A2(\IF_ID_inst [14] ), .B1(_03003_ ), .B2(_03001_ ), .ZN(_03313_ ) );
AND4_X1 _10989_ ( .A1(_03163_ ), .A2(_03311_ ), .A3(_03312_ ), .A4(_03313_ ), .ZN(_03314_ ) );
AOI21_X1 _10990_ ( .A(_02991_ ), .B1(_03309_ ), .B2(_03314_ ), .ZN(_00240_ ) );
INV_X1 _10991_ ( .A(_03037_ ), .ZN(_03315_ ) );
AOI22_X1 _10992_ ( .A1(_03162_ ), .A2(_03180_ ), .B1(_03154_ ), .B2(_03196_ ), .ZN(_03316_ ) );
NAND4_X1 _10993_ ( .A1(_03315_ ), .A2(_03070_ ), .A3(_03308_ ), .A4(_03316_ ), .ZN(_03317_ ) );
OAI21_X1 _10994_ ( .A(_03158_ ), .B1(_03156_ ), .B2(_03170_ ), .ZN(_03318_ ) );
NAND2_X1 _10995_ ( .A1(_03076_ ), .A2(_03167_ ), .ZN(_03319_ ) );
OAI211_X1 _10996_ ( .A(_03318_ ), .B(_03319_ ), .C1(_03167_ ), .C2(_03004_ ), .ZN(_03320_ ) );
AND3_X1 _10997_ ( .A1(_03003_ ), .A2(_02993_ ), .A3(_03039_ ), .ZN(_03321_ ) );
AND2_X1 _10998_ ( .A1(_03321_ ), .A2(_03154_ ), .ZN(_03322_ ) );
OR2_X1 _10999_ ( .A1(_03322_ ), .A2(_03211_ ), .ZN(_03323_ ) );
NAND3_X1 _11000_ ( .A1(_03310_ ), .A2(_03063_ ), .A3(\IF_ID_inst [14] ), .ZN(_03324_ ) );
NAND3_X1 _11001_ ( .A1(_03158_ ), .A2(_03174_ ), .A3(_03173_ ), .ZN(_03325_ ) );
NAND4_X1 _11002_ ( .A1(_03324_ ), .A2(_03066_ ), .A3(_03292_ ), .A4(_03325_ ), .ZN(_03326_ ) );
NOR4_X1 _11003_ ( .A1(_03317_ ), .A2(_03320_ ), .A3(_03323_ ), .A4(_03326_ ), .ZN(_03327_ ) );
OAI21_X1 _11004_ ( .A(_03168_ ), .B1(_03185_ ), .B2(_02997_ ), .ZN(_03328_ ) );
OAI21_X1 _11005_ ( .A(_03154_ ), .B1(_03074_ ), .B2(_02997_ ), .ZN(_03329_ ) );
OAI21_X1 _11006_ ( .A(_03196_ ), .B1(_03175_ ), .B2(_03170_ ), .ZN(_03330_ ) );
AND3_X1 _11007_ ( .A1(_03328_ ), .A2(_03329_ ), .A3(_03330_ ), .ZN(_03331_ ) );
AOI21_X1 _11008_ ( .A(_02991_ ), .B1(_03327_ ), .B2(_03331_ ), .ZN(_00241_ ) );
INV_X1 _11009_ ( .A(_03141_ ), .ZN(_03332_ ) );
INV_X1 _11010_ ( .A(fanout_net_43 ), .ZN(_03333_ ) );
BUF_X4 _11011_ ( .A(_03333_ ), .Z(_03334_ ) );
NAND4_X1 _11012_ ( .A1(_03332_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_03334_ ), .ZN(_03335_ ) );
NAND2_X1 _11013_ ( .A1(\mtvec [0] ), .A2(fanout_net_43 ), .ZN(_03336_ ) );
AOI21_X1 _11014_ ( .A(fanout_net_2 ), .B1(_03335_ ), .B2(_03336_ ), .ZN(_00245_ ) );
NOR4_X1 _11015_ ( .A1(_02988_ ), .A2(_03038_ ), .A3(\IF_ID_inst [4] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03337_ ) );
AND2_X1 _11016_ ( .A1(_03337_ ), .A2(_03002_ ), .ZN(_03338_ ) );
AND2_X1 _11017_ ( .A1(_03338_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03339_ ) );
OAI211_X1 _11018_ ( .A(_03086_ ), .B(\IF_ID_inst [31] ), .C1(_03002_ ), .C2(_03045_ ), .ZN(_03340_ ) );
NOR2_X1 _11019_ ( .A1(_03339_ ), .A2(_03340_ ), .ZN(_03341_ ) );
BUF_X4 _11020_ ( .A(_03341_ ), .Z(_03342_ ) );
XNOR2_X1 _11021_ ( .A(_03342_ ), .B(\IF_ID_pc [29] ), .ZN(_03343_ ) );
NAND2_X1 _11022_ ( .A1(_03086_ ), .A2(_03002_ ), .ZN(_03344_ ) );
NOR2_X4 _11023_ ( .A1(_03344_ ), .A2(_02988_ ), .ZN(_03345_ ) );
AND2_X1 _11024_ ( .A1(_03345_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03346_ ) );
INV_X1 _11025_ ( .A(_03346_ ), .ZN(_03347_ ) );
AND2_X1 _11026_ ( .A1(_03089_ ), .A2(\IF_ID_inst [16] ), .ZN(_03348_ ) );
OAI21_X1 _11027_ ( .A(_03347_ ), .B1(_03345_ ), .B2(_03348_ ), .ZN(_03349_ ) );
INV_X1 _11028_ ( .A(\IF_ID_pc [16] ), .ZN(_03350_ ) );
XNOR2_X1 _11029_ ( .A(_03349_ ), .B(_03350_ ), .ZN(_03351_ ) );
AND3_X1 _11030_ ( .A1(_02992_ ), .A2(\IF_ID_inst [31] ), .A3(_02994_ ), .ZN(_03352_ ) );
AND2_X1 _11031_ ( .A1(_03086_ ), .A2(_03352_ ), .ZN(_03353_ ) );
NAND2_X1 _11032_ ( .A1(_03353_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03354_ ) );
AND2_X1 _11033_ ( .A1(_03088_ ), .A2(\IF_ID_inst [15] ), .ZN(_03355_ ) );
OAI21_X1 _11034_ ( .A(_03354_ ), .B1(_03355_ ), .B2(_03345_ ), .ZN(_03356_ ) );
XNOR2_X1 _11035_ ( .A(_03356_ ), .B(\IF_ID_pc [15] ), .ZN(_03357_ ) );
INV_X1 _11036_ ( .A(_03357_ ), .ZN(_03358_ ) );
NOR2_X1 _11037_ ( .A1(_03351_ ), .A2(_03358_ ), .ZN(_03359_ ) );
AND2_X1 _11038_ ( .A1(_03087_ ), .A2(\IF_ID_inst [24] ), .ZN(_03360_ ) );
INV_X1 _11039_ ( .A(_03360_ ), .ZN(_03361_ ) );
INV_X1 _11040_ ( .A(_03338_ ), .ZN(_03362_ ) );
OAI21_X1 _11041_ ( .A(_03361_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_03362_ ), .ZN(_03363_ ) );
OR2_X1 _11042_ ( .A1(_03363_ ), .A2(fanout_net_12 ), .ZN(_03364_ ) );
AND4_X1 _11043_ ( .A1(\IF_ID_inst [31] ), .A2(_03086_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .A4(_03002_ ), .ZN(_03365_ ) );
AND3_X1 _11044_ ( .A1(_03086_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .A3(_03045_ ), .ZN(_03366_ ) );
NOR2_X1 _11045_ ( .A1(_03365_ ), .A2(_03366_ ), .ZN(_03367_ ) );
INV_X1 _11046_ ( .A(\IF_ID_pc [2] ), .ZN(_03368_ ) );
XNOR2_X1 _11047_ ( .A(_03367_ ), .B(_03368_ ), .ZN(_03369_ ) );
AND2_X1 _11048_ ( .A1(_03087_ ), .A2(\IF_ID_inst [21] ), .ZN(_03370_ ) );
NOR2_X1 _11049_ ( .A1(_03362_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03371_ ) );
OR2_X1 _11050_ ( .A1(_03370_ ), .A2(_03371_ ), .ZN(_03372_ ) );
AND3_X1 _11051_ ( .A1(_03369_ ), .A2(\IF_ID_pc [1] ), .A3(_03372_ ), .ZN(_03373_ ) );
NOR3_X1 _11052_ ( .A1(_03365_ ), .A2(_03366_ ), .A3(_03368_ ), .ZN(_03374_ ) );
NOR2_X1 _11053_ ( .A1(_03373_ ), .A2(_03374_ ), .ZN(_03375_ ) );
AND2_X1 _11054_ ( .A1(_03087_ ), .A2(\IF_ID_inst [23] ), .ZN(_03376_ ) );
INV_X1 _11055_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03377_ ) );
MUX2_X1 _11056_ ( .A(_03376_ ), .B(_03377_ ), .S(_03345_ ), .Z(_03378_ ) );
XNOR2_X1 _11057_ ( .A(_03378_ ), .B(fanout_net_8 ), .ZN(_03379_ ) );
NOR2_X2 _11058_ ( .A1(_03375_ ), .A2(_03379_ ), .ZN(_03380_ ) );
INV_X1 _11059_ ( .A(_03378_ ), .ZN(_03381_ ) );
NOR2_X1 _11060_ ( .A1(_03381_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03382_ ) );
OAI21_X1 _11061_ ( .A(_03364_ ), .B1(_03380_ ), .B2(_03382_ ), .ZN(_03383_ ) );
NAND2_X1 _11062_ ( .A1(_03363_ ), .A2(fanout_net_12 ), .ZN(_03384_ ) );
AND2_X1 _11063_ ( .A1(_03383_ ), .A2(_03384_ ), .ZN(_03385_ ) );
AND2_X1 _11064_ ( .A1(_03087_ ), .A2(\IF_ID_inst [25] ), .ZN(_03386_ ) );
INV_X1 _11065_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03387_ ) );
AOI21_X1 _11066_ ( .A(_03386_ ), .B1(_03353_ ), .B2(_03387_ ), .ZN(_03388_ ) );
INV_X1 _11067_ ( .A(\IF_ID_pc [5] ), .ZN(_03389_ ) );
XNOR2_X1 _11068_ ( .A(_03388_ ), .B(_03389_ ), .ZN(_03390_ ) );
NOR2_X1 _11069_ ( .A1(_03385_ ), .A2(_03390_ ), .ZN(_03391_ ) );
NOR2_X1 _11070_ ( .A1(_03388_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03392_ ) );
NOR2_X1 _11071_ ( .A1(_03391_ ), .A2(_03392_ ), .ZN(_03393_ ) );
AND2_X1 _11072_ ( .A1(_03088_ ), .A2(\IF_ID_inst [26] ), .ZN(_03394_ ) );
INV_X1 _11073_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03395_ ) );
AOI21_X1 _11074_ ( .A(_03394_ ), .B1(_03395_ ), .B2(_03338_ ), .ZN(_03396_ ) );
OAI21_X1 _11075_ ( .A(_03393_ ), .B1(_01808_ ), .B2(_03396_ ), .ZN(_03397_ ) );
AND2_X1 _11076_ ( .A1(_03087_ ), .A2(\IF_ID_inst [27] ), .ZN(_03398_ ) );
INV_X1 _11077_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03399_ ) );
AOI21_X1 _11078_ ( .A(_03398_ ), .B1(_03399_ ), .B2(_03338_ ), .ZN(_03400_ ) );
XNOR2_X1 _11079_ ( .A(_03400_ ), .B(\IF_ID_pc [7] ), .ZN(_03401_ ) );
NAND2_X1 _11080_ ( .A1(_03396_ ), .A2(_01808_ ), .ZN(_03402_ ) );
AND3_X2 _11081_ ( .A1(_03397_ ), .A2(_03401_ ), .A3(_03402_ ), .ZN(_03403_ ) );
INV_X1 _11082_ ( .A(\IF_ID_pc [7] ), .ZN(_03404_ ) );
NOR2_X1 _11083_ ( .A1(_03400_ ), .A2(_03404_ ), .ZN(_03405_ ) );
NOR2_X1 _11084_ ( .A1(_03403_ ), .A2(_03405_ ), .ZN(_03406_ ) );
INV_X1 _11085_ ( .A(\IF_ID_pc [8] ), .ZN(_03407_ ) );
AND2_X1 _11086_ ( .A1(_03088_ ), .A2(\IF_ID_inst [28] ), .ZN(_03408_ ) );
INV_X1 _11087_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03409_ ) );
AOI21_X1 _11088_ ( .A(_03408_ ), .B1(_03409_ ), .B2(_03338_ ), .ZN(_03410_ ) );
AOI21_X1 _11089_ ( .A(_03406_ ), .B1(_03407_ ), .B2(_03410_ ), .ZN(_03411_ ) );
NOR2_X1 _11090_ ( .A1(_03410_ ), .A2(_03407_ ), .ZN(_03412_ ) );
OR2_X2 _11091_ ( .A1(_03411_ ), .A2(_03412_ ), .ZN(_03413_ ) );
AND2_X1 _11092_ ( .A1(_03088_ ), .A2(\IF_ID_inst [13] ), .ZN(_03414_ ) );
INV_X1 _11093_ ( .A(_03414_ ), .ZN(_03415_ ) );
AOI21_X1 _11094_ ( .A(_03339_ ), .B1(_03415_ ), .B2(_03362_ ), .ZN(_03416_ ) );
XNOR2_X1 _11095_ ( .A(_03416_ ), .B(_01838_ ), .ZN(_03417_ ) );
AND2_X1 _11096_ ( .A1(_03088_ ), .A2(\IF_ID_inst [14] ), .ZN(_03418_ ) );
INV_X1 _11097_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03419_ ) );
MUX2_X1 _11098_ ( .A(_03418_ ), .B(_03419_ ), .S(_03345_ ), .Z(_03420_ ) );
NOR2_X1 _11099_ ( .A1(_03420_ ), .A2(\IF_ID_pc [14] ), .ZN(_03421_ ) );
INV_X1 _11100_ ( .A(_03421_ ), .ZN(_03422_ ) );
NAND2_X1 _11101_ ( .A1(_03420_ ), .A2(\IF_ID_pc [14] ), .ZN(_03423_ ) );
AND3_X1 _11102_ ( .A1(_03417_ ), .A2(_03422_ ), .A3(_03423_ ), .ZN(_03424_ ) );
AND2_X1 _11103_ ( .A1(_03088_ ), .A2(\IF_ID_inst [12] ), .ZN(_03425_ ) );
MUX2_X1 _11104_ ( .A(_03425_ ), .B(_03419_ ), .S(_03345_ ), .Z(_03426_ ) );
XNOR2_X1 _11105_ ( .A(_03426_ ), .B(\IF_ID_pc [12] ), .ZN(_03427_ ) );
NAND2_X1 _11106_ ( .A1(_03088_ ), .A2(\IF_ID_inst [20] ), .ZN(_03428_ ) );
OAI21_X1 _11107_ ( .A(_03428_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03362_ ), .ZN(_03429_ ) );
XNOR2_X1 _11108_ ( .A(_03429_ ), .B(_01741_ ), .ZN(_03430_ ) );
INV_X1 _11109_ ( .A(_03430_ ), .ZN(_03431_ ) );
NOR2_X1 _11110_ ( .A1(_03427_ ), .A2(_03431_ ), .ZN(_03432_ ) );
AND2_X1 _11111_ ( .A1(_03088_ ), .A2(\IF_ID_inst [29] ), .ZN(_03433_ ) );
INV_X1 _11112_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03434_ ) );
AOI21_X1 _11113_ ( .A(_03433_ ), .B1(_03353_ ), .B2(_03434_ ), .ZN(_03435_ ) );
XNOR2_X1 _11114_ ( .A(_03435_ ), .B(\IF_ID_pc [9] ), .ZN(_03436_ ) );
AND2_X1 _11115_ ( .A1(_03088_ ), .A2(\IF_ID_inst [30] ), .ZN(_03437_ ) );
INV_X1 _11116_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03438_ ) );
AOI21_X1 _11117_ ( .A(_03437_ ), .B1(_03353_ ), .B2(_03438_ ), .ZN(_03439_ ) );
XNOR2_X1 _11118_ ( .A(_03439_ ), .B(\IF_ID_pc [10] ), .ZN(_03440_ ) );
AND2_X1 _11119_ ( .A1(_03436_ ), .A2(_03440_ ), .ZN(_03441_ ) );
AND2_X1 _11120_ ( .A1(_03432_ ), .A2(_03441_ ), .ZN(_03442_ ) );
AND4_X1 _11121_ ( .A1(_03359_ ), .A2(_03413_ ), .A3(_03424_ ), .A4(_03442_ ), .ZN(_03443_ ) );
MUX2_X1 _11122_ ( .A(_03433_ ), .B(_03434_ ), .S(_03345_ ), .Z(_03444_ ) );
NAND3_X1 _11123_ ( .A1(_03440_ ), .A2(\IF_ID_pc [9] ), .A3(_03444_ ), .ZN(_03445_ ) );
INV_X1 _11124_ ( .A(\IF_ID_pc [10] ), .ZN(_03446_ ) );
OAI21_X1 _11125_ ( .A(_03445_ ), .B1(_03446_ ), .B2(_03439_ ), .ZN(_03447_ ) );
AND2_X1 _11126_ ( .A1(_03447_ ), .A2(_03432_ ), .ZN(_03448_ ) );
NAND2_X1 _11127_ ( .A1(_03426_ ), .A2(\IF_ID_pc [12] ), .ZN(_03449_ ) );
NAND2_X1 _11128_ ( .A1(_03429_ ), .A2(\IF_ID_pc [11] ), .ZN(_03450_ ) );
OAI21_X1 _11129_ ( .A(_03449_ ), .B1(_03427_ ), .B2(_03450_ ), .ZN(_03451_ ) );
OAI211_X1 _11130_ ( .A(_03359_ ), .B(_03424_ ), .C1(_03448_ ), .C2(_03451_ ), .ZN(_03452_ ) );
OR2_X1 _11131_ ( .A1(_03349_ ), .A2(_03350_ ), .ZN(_03453_ ) );
INV_X1 _11132_ ( .A(_03345_ ), .ZN(_03454_ ) );
AOI21_X1 _11133_ ( .A(_03346_ ), .B1(_03454_ ), .B2(_03415_ ), .ZN(_03455_ ) );
NAND4_X1 _11134_ ( .A1(_03422_ ), .A2(\IF_ID_pc [13] ), .A3(_03455_ ), .A4(_03423_ ), .ZN(_03456_ ) );
NAND2_X1 _11135_ ( .A1(_03456_ ), .A2(_03423_ ), .ZN(_03457_ ) );
NAND2_X1 _11136_ ( .A1(_03457_ ), .A2(_03359_ ), .ZN(_03458_ ) );
INV_X1 _11137_ ( .A(\IF_ID_pc [15] ), .ZN(_03459_ ) );
OR3_X1 _11138_ ( .A1(_03351_ ), .A2(_03459_ ), .A3(_03356_ ), .ZN(_03460_ ) );
NAND4_X1 _11139_ ( .A1(_03452_ ), .A2(_03453_ ), .A3(_03458_ ), .A4(_03460_ ), .ZN(_03461_ ) );
NOR2_X2 _11140_ ( .A1(_03443_ ), .A2(_03461_ ), .ZN(_03462_ ) );
INV_X1 _11141_ ( .A(_03462_ ), .ZN(_03463_ ) );
AND2_X1 _11142_ ( .A1(_03089_ ), .A2(\IF_ID_inst [18] ), .ZN(_03464_ ) );
MUX2_X1 _11143_ ( .A(_03419_ ), .B(_03464_ ), .S(_03362_ ), .Z(_03465_ ) );
XNOR2_X1 _11144_ ( .A(_03465_ ), .B(_01909_ ), .ZN(_03466_ ) );
AND2_X1 _11145_ ( .A1(_03089_ ), .A2(\IF_ID_inst [17] ), .ZN(_03467_ ) );
INV_X1 _11146_ ( .A(_03467_ ), .ZN(_03468_ ) );
AOI21_X1 _11147_ ( .A(_03339_ ), .B1(_03468_ ), .B2(_03362_ ), .ZN(_03469_ ) );
XNOR2_X1 _11148_ ( .A(_03469_ ), .B(_01699_ ), .ZN(_03470_ ) );
AND2_X1 _11149_ ( .A1(_03089_ ), .A2(\IF_ID_inst [19] ), .ZN(_03471_ ) );
MUX2_X1 _11150_ ( .A(_03419_ ), .B(_03471_ ), .S(_03362_ ), .Z(_03472_ ) );
XOR2_X1 _11151_ ( .A(_03472_ ), .B(\IF_ID_pc [19] ), .Z(_03473_ ) );
XNOR2_X1 _11152_ ( .A(_03341_ ), .B(_01913_ ), .ZN(_03474_ ) );
AND2_X1 _11153_ ( .A1(_03473_ ), .A2(_03474_ ), .ZN(_03475_ ) );
NAND4_X1 _11154_ ( .A1(_03463_ ), .A2(_03466_ ), .A3(_03470_ ), .A4(_03475_ ), .ZN(_03476_ ) );
AOI21_X1 _11155_ ( .A(_03346_ ), .B1(_03454_ ), .B2(_03468_ ), .ZN(_03477_ ) );
AND3_X1 _11156_ ( .A1(_03466_ ), .A2(\IF_ID_pc [17] ), .A3(_03477_ ), .ZN(_03478_ ) );
AND2_X1 _11157_ ( .A1(_03465_ ), .A2(\IF_ID_pc [18] ), .ZN(_03479_ ) );
OR2_X1 _11158_ ( .A1(_03478_ ), .A2(_03479_ ), .ZN(_03480_ ) );
AND2_X1 _11159_ ( .A1(_03480_ ), .A2(_03475_ ), .ZN(_03481_ ) );
AOI21_X1 _11160_ ( .A(_02988_ ), .B1(_03286_ ), .B2(_03344_ ), .ZN(_03482_ ) );
AND2_X1 _11161_ ( .A1(_03482_ ), .A2(_03354_ ), .ZN(_03483_ ) );
AND2_X1 _11162_ ( .A1(_03483_ ), .A2(\IF_ID_pc [20] ), .ZN(_03484_ ) );
AND3_X1 _11163_ ( .A1(_03474_ ), .A2(\IF_ID_pc [19] ), .A3(_03472_ ), .ZN(_03485_ ) );
NOR3_X1 _11164_ ( .A1(_03481_ ), .A2(_03484_ ), .A3(_03485_ ), .ZN(_03486_ ) );
NAND2_X1 _11165_ ( .A1(_03476_ ), .A2(_03486_ ), .ZN(_03487_ ) );
XNOR2_X1 _11166_ ( .A(_03341_ ), .B(_01861_ ), .ZN(_03488_ ) );
XNOR2_X1 _11167_ ( .A(_03341_ ), .B(_01790_ ), .ZN(_03489_ ) );
AND2_X1 _11168_ ( .A1(_03488_ ), .A2(_03489_ ), .ZN(_03490_ ) );
XNOR2_X1 _11169_ ( .A(_03342_ ), .B(_01847_ ), .ZN(_03491_ ) );
XNOR2_X1 _11170_ ( .A(_03342_ ), .B(_01728_ ), .ZN(_03492_ ) );
AND2_X1 _11171_ ( .A1(_03491_ ), .A2(_03492_ ), .ZN(_03493_ ) );
AND3_X2 _11172_ ( .A1(_03487_ ), .A2(_03490_ ), .A3(_03493_ ), .ZN(_03494_ ) );
OAI211_X1 _11173_ ( .A(_03490_ ), .B(_03483_ ), .C1(\IF_ID_pc [22] ), .C2(\IF_ID_pc [21] ), .ZN(_03495_ ) );
AND2_X1 _11174_ ( .A1(_03089_ ), .A2(\IF_ID_inst [31] ), .ZN(_03496_ ) );
OAI221_X1 _11175_ ( .A(_03354_ ), .B1(\IF_ID_pc [24] ), .B2(\IF_ID_pc [23] ), .C1(_03496_ ), .C2(_03345_ ), .ZN(_03497_ ) );
NAND2_X1 _11176_ ( .A1(_03495_ ), .A2(_03497_ ), .ZN(_03498_ ) );
NOR2_X1 _11177_ ( .A1(_03494_ ), .A2(_03498_ ), .ZN(_03499_ ) );
INV_X1 _11178_ ( .A(_03499_ ), .ZN(_03500_ ) );
XNOR2_X1 _11179_ ( .A(_03342_ ), .B(_01775_ ), .ZN(_03501_ ) );
XNOR2_X1 _11180_ ( .A(_03342_ ), .B(_01788_ ), .ZN(_03502_ ) );
AND3_X4 _11181_ ( .A1(_03500_ ), .A2(_03501_ ), .A3(_03502_ ), .ZN(_03503_ ) );
XOR2_X1 _11182_ ( .A(_03342_ ), .B(\IF_ID_pc [28] ), .Z(_03504_ ) );
XNOR2_X1 _11183_ ( .A(_03342_ ), .B(_01850_ ), .ZN(_03505_ ) );
NAND3_X1 _11184_ ( .A1(_03503_ ), .A2(_03504_ ), .A3(_03505_ ), .ZN(_03506_ ) );
INV_X1 _11185_ ( .A(_03483_ ), .ZN(_03507_ ) );
AOI21_X1 _11186_ ( .A(_03507_ ), .B1(_01775_ ), .B2(_01788_ ), .ZN(_03508_ ) );
NAND3_X1 _11187_ ( .A1(_03508_ ), .A2(_03504_ ), .A3(_03505_ ), .ZN(_03509_ ) );
NAND3_X1 _11188_ ( .A1(_03482_ ), .A2(\IF_ID_pc [28] ), .A3(_03354_ ), .ZN(_03510_ ) );
AND2_X1 _11189_ ( .A1(_03483_ ), .A2(\IF_ID_pc [27] ), .ZN(_03511_ ) );
INV_X1 _11190_ ( .A(_03511_ ), .ZN(_03512_ ) );
AND3_X1 _11191_ ( .A1(_03509_ ), .A2(_03510_ ), .A3(_03512_ ), .ZN(_03513_ ) );
AOI21_X2 _11192_ ( .A(_03343_ ), .B1(_03506_ ), .B2(_03513_ ), .ZN(_03514_ ) );
AND3_X1 _11193_ ( .A1(_03482_ ), .A2(\IF_ID_pc [29] ), .A3(_03354_ ), .ZN(_03515_ ) );
NOR2_X1 _11194_ ( .A1(_03514_ ), .A2(_03515_ ), .ZN(_03516_ ) );
XNOR2_X1 _11195_ ( .A(_03342_ ), .B(\IF_ID_pc [30] ), .ZN(_03517_ ) );
OR2_X1 _11196_ ( .A1(_03516_ ), .A2(_03517_ ), .ZN(_03518_ ) );
AOI21_X1 _11197_ ( .A(_03143_ ), .B1(_03516_ ), .B2(_03517_ ), .ZN(_03519_ ) );
AOI221_X1 _11198_ ( .A(fanout_net_43 ), .B1(\myexu.pc_jump [30] ), .B2(_03143_ ), .C1(_03518_ ), .C2(_03519_ ), .ZN(_03520_ ) );
BUF_X4 _11199_ ( .A(_03334_ ), .Z(_03521_ ) );
NOR2_X1 _11200_ ( .A1(_03521_ ), .A2(\mtvec [30] ), .ZN(_03522_ ) );
NOR3_X1 _11201_ ( .A1(_03520_ ), .A2(fanout_net_2 ), .A3(_03522_ ), .ZN(_00246_ ) );
OR2_X1 _11202_ ( .A1(_03487_ ), .A2(_03492_ ), .ZN(_03523_ ) );
INV_X2 _11203_ ( .A(_03143_ ), .ZN(_03524_ ) );
NAND2_X1 _11204_ ( .A1(_03487_ ), .A2(_03492_ ), .ZN(_03525_ ) );
AND3_X1 _11205_ ( .A1(_03523_ ), .A2(_03524_ ), .A3(_03525_ ), .ZN(_03526_ ) );
BUF_X4 _11206_ ( .A(_03143_ ), .Z(_03527_ ) );
AOI211_X1 _11207_ ( .A(fanout_net_43 ), .B(_03526_ ), .C1(\myexu.pc_jump [21] ), .C2(_03527_ ), .ZN(_03528_ ) );
NOR2_X1 _11208_ ( .A1(_03521_ ), .A2(\mtvec [21] ), .ZN(_03529_ ) );
NOR3_X1 _11209_ ( .A1(_03528_ ), .A2(fanout_net_2 ), .A3(_03529_ ), .ZN(_00247_ ) );
INV_X1 _11210_ ( .A(_03466_ ), .ZN(_03530_ ) );
INV_X1 _11211_ ( .A(_03470_ ), .ZN(_03531_ ) );
NOR3_X1 _11212_ ( .A1(_03462_ ), .A2(_03530_ ), .A3(_03531_ ), .ZN(_03532_ ) );
OAI21_X1 _11213_ ( .A(_03473_ ), .B1(_03532_ ), .B2(_03480_ ), .ZN(_03533_ ) );
AND2_X1 _11214_ ( .A1(_03472_ ), .A2(\IF_ID_pc [19] ), .ZN(_03534_ ) );
INV_X1 _11215_ ( .A(_03534_ ), .ZN(_03535_ ) );
AND2_X1 _11216_ ( .A1(_03533_ ), .A2(_03535_ ), .ZN(_03536_ ) );
XNOR2_X1 _11217_ ( .A(_03536_ ), .B(_03474_ ), .ZN(_03537_ ) );
BUF_X4 _11218_ ( .A(_03524_ ), .Z(_03538_ ) );
AND2_X1 _11219_ ( .A1(_03537_ ), .A2(_03538_ ), .ZN(_03539_ ) );
AOI211_X1 _11220_ ( .A(fanout_net_43 ), .B(_03539_ ), .C1(\myexu.pc_jump [20] ), .C2(_03527_ ), .ZN(_03540_ ) );
NOR2_X1 _11221_ ( .A1(_03521_ ), .A2(\mtvec [20] ), .ZN(_03541_ ) );
NOR3_X1 _11222_ ( .A1(_03540_ ), .A2(fanout_net_2 ), .A3(_03541_ ), .ZN(_00248_ ) );
NOR2_X1 _11223_ ( .A1(_03532_ ), .A2(_03480_ ), .ZN(_03542_ ) );
XOR2_X1 _11224_ ( .A(_03542_ ), .B(_03473_ ), .Z(_03543_ ) );
BUF_X4 _11225_ ( .A(_03538_ ), .Z(_03544_ ) );
NAND2_X1 _11226_ ( .A1(_03543_ ), .A2(_03544_ ), .ZN(_03545_ ) );
BUF_X4 _11227_ ( .A(_03538_ ), .Z(_03546_ ) );
OAI211_X1 _11228_ ( .A(_03545_ ), .B(_03521_ ), .C1(\myexu.pc_jump [19] ), .C2(_03546_ ), .ZN(_03547_ ) );
NAND2_X1 _11229_ ( .A1(\mtvec [19] ), .A2(fanout_net_43 ), .ZN(_03548_ ) );
AOI21_X1 _11230_ ( .A(fanout_net_2 ), .B1(_03547_ ), .B2(_03548_ ), .ZN(_00249_ ) );
OR3_X1 _11231_ ( .A1(_03141_ ), .A2(_03142_ ), .A3(\myexu.pc_jump [18] ), .ZN(_03549_ ) );
NAND2_X1 _11232_ ( .A1(_03477_ ), .A2(\IF_ID_pc [17] ), .ZN(_03550_ ) );
OAI21_X1 _11233_ ( .A(_03550_ ), .B1(_03462_ ), .B2(_03531_ ), .ZN(_03551_ ) );
XNOR2_X1 _11234_ ( .A(_03551_ ), .B(_03530_ ), .ZN(_03552_ ) );
OAI211_X1 _11235_ ( .A(_03521_ ), .B(_03549_ ), .C1(_03552_ ), .C2(_03527_ ), .ZN(_03553_ ) );
NAND2_X1 _11236_ ( .A1(\mtvec [18] ), .A2(fanout_net_43 ), .ZN(_03554_ ) );
AOI21_X1 _11237_ ( .A(fanout_net_2 ), .B1(_03553_ ), .B2(_03554_ ), .ZN(_00250_ ) );
XNOR2_X1 _11238_ ( .A(_03462_ ), .B(_03531_ ), .ZN(_03555_ ) );
NAND2_X1 _11239_ ( .A1(_03555_ ), .A2(_03544_ ), .ZN(_03556_ ) );
BUF_X4 _11240_ ( .A(_03334_ ), .Z(_03557_ ) );
OAI211_X1 _11241_ ( .A(_03556_ ), .B(_03557_ ), .C1(\myexu.pc_jump [17] ), .C2(_03546_ ), .ZN(_03558_ ) );
NAND2_X1 _11242_ ( .A1(\mtvec [17] ), .A2(fanout_net_43 ), .ZN(_03559_ ) );
AOI21_X1 _11243_ ( .A(fanout_net_2 ), .B1(_03558_ ), .B2(_03559_ ), .ZN(_00251_ ) );
OAI21_X1 _11244_ ( .A(_03442_ ), .B1(_03411_ ), .B2(_03412_ ), .ZN(_03560_ ) );
NAND2_X1 _11245_ ( .A1(_03447_ ), .A2(_03432_ ), .ZN(_03561_ ) );
OR2_X1 _11246_ ( .A1(_03427_ ), .A2(_03450_ ), .ZN(_03562_ ) );
AND3_X1 _11247_ ( .A1(_03561_ ), .A2(_03449_ ), .A3(_03562_ ), .ZN(_03563_ ) );
NAND2_X1 _11248_ ( .A1(_03560_ ), .A2(_03563_ ), .ZN(_03564_ ) );
AOI21_X1 _11249_ ( .A(_03457_ ), .B1(_03564_ ), .B2(_03424_ ), .ZN(_03565_ ) );
NOR2_X1 _11250_ ( .A1(_03565_ ), .A2(_03358_ ), .ZN(_03566_ ) );
NOR2_X1 _11251_ ( .A1(_03356_ ), .A2(_03459_ ), .ZN(_03567_ ) );
OR3_X1 _11252_ ( .A1(_03566_ ), .A2(_03351_ ), .A3(_03567_ ), .ZN(_03568_ ) );
BUF_X4 _11253_ ( .A(_03524_ ), .Z(_03569_ ) );
OAI21_X1 _11254_ ( .A(_03351_ ), .B1(_03566_ ), .B2(_03567_ ), .ZN(_03570_ ) );
NAND3_X1 _11255_ ( .A1(_03568_ ), .A2(_03569_ ), .A3(_03570_ ), .ZN(_03571_ ) );
OAI211_X1 _11256_ ( .A(_03571_ ), .B(_03557_ ), .C1(\myexu.pc_jump [16] ), .C2(_03546_ ), .ZN(_03572_ ) );
NAND2_X1 _11257_ ( .A1(\mtvec [16] ), .A2(fanout_net_43 ), .ZN(_03573_ ) );
AOI21_X1 _11258_ ( .A(fanout_net_2 ), .B1(_03572_ ), .B2(_03573_ ), .ZN(_00252_ ) );
XNOR2_X1 _11259_ ( .A(_03565_ ), .B(_03357_ ), .ZN(_03574_ ) );
MUX2_X1 _11260_ ( .A(\myexu.pc_jump [15] ), .B(_03574_ ), .S(_03524_ ), .Z(_03575_ ) );
MUX2_X1 _11261_ ( .A(\mtvec [15] ), .B(_03575_ ), .S(_03334_ ), .Z(_03576_ ) );
AND2_X1 _11262_ ( .A1(_03576_ ), .A2(_01545_ ), .ZN(_00253_ ) );
AND2_X1 _11263_ ( .A1(_03416_ ), .A2(\IF_ID_pc [13] ), .ZN(_03577_ ) );
AND2_X1 _11264_ ( .A1(_03564_ ), .A2(_03417_ ), .ZN(_03578_ ) );
AND2_X1 _11265_ ( .A1(_03420_ ), .A2(\IF_ID_pc [14] ), .ZN(_03579_ ) );
OR4_X1 _11266_ ( .A1(_03577_ ), .A2(_03578_ ), .A3(_03421_ ), .A4(_03579_ ), .ZN(_03580_ ) );
OAI22_X1 _11267_ ( .A1(_03578_ ), .A2(_03577_ ), .B1(_03421_ ), .B2(_03579_ ), .ZN(_03581_ ) );
NAND3_X1 _11268_ ( .A1(_03580_ ), .A2(_03569_ ), .A3(_03581_ ), .ZN(_03582_ ) );
OAI211_X1 _11269_ ( .A(_03582_ ), .B(_03557_ ), .C1(\myexu.pc_jump [14] ), .C2(_03546_ ), .ZN(_03583_ ) );
NAND2_X1 _11270_ ( .A1(\mtvec [14] ), .A2(fanout_net_43 ), .ZN(_03584_ ) );
AOI21_X1 _11271_ ( .A(fanout_net_2 ), .B1(_03583_ ), .B2(_03584_ ), .ZN(_00254_ ) );
NOR2_X1 _11272_ ( .A1(_03564_ ), .A2(_03417_ ), .ZN(_03585_ ) );
OAI21_X1 _11273_ ( .A(_03569_ ), .B1(_03578_ ), .B2(_03585_ ), .ZN(_03586_ ) );
OAI211_X1 _11274_ ( .A(_03586_ ), .B(_03557_ ), .C1(\myexu.pc_jump [13] ), .C2(_03546_ ), .ZN(_03587_ ) );
NAND2_X1 _11275_ ( .A1(\mtvec [13] ), .A2(fanout_net_43 ), .ZN(_03588_ ) );
AOI21_X1 _11276_ ( .A(fanout_net_2 ), .B1(_03587_ ), .B2(_03588_ ), .ZN(_00255_ ) );
AOI21_X1 _11277_ ( .A(_03447_ ), .B1(_03413_ ), .B2(_03441_ ), .ZN(_03589_ ) );
OR2_X1 _11278_ ( .A1(_03589_ ), .A2(_03431_ ), .ZN(_03590_ ) );
AND3_X1 _11279_ ( .A1(_03590_ ), .A2(_03450_ ), .A3(_03427_ ), .ZN(_03591_ ) );
AOI21_X1 _11280_ ( .A(_03427_ ), .B1(_03590_ ), .B2(_03450_ ), .ZN(_03592_ ) );
OAI21_X1 _11281_ ( .A(_03569_ ), .B1(_03591_ ), .B2(_03592_ ), .ZN(_03593_ ) );
OAI211_X1 _11282_ ( .A(_03593_ ), .B(_03557_ ), .C1(\myexu.pc_jump [12] ), .C2(_03546_ ), .ZN(_03594_ ) );
NAND2_X1 _11283_ ( .A1(\mtvec [12] ), .A2(fanout_net_43 ), .ZN(_03595_ ) );
AOI21_X1 _11284_ ( .A(fanout_net_2 ), .B1(_03594_ ), .B2(_03595_ ), .ZN(_00256_ ) );
AND3_X1 _11285_ ( .A1(_03506_ ), .A2(_03513_ ), .A3(_03343_ ), .ZN(_03596_ ) );
OAI21_X1 _11286_ ( .A(_03569_ ), .B1(_03596_ ), .B2(_03514_ ), .ZN(_03597_ ) );
OAI211_X1 _11287_ ( .A(_03597_ ), .B(_03557_ ), .C1(\myexu.pc_jump [29] ), .C2(_03546_ ), .ZN(_03598_ ) );
NAND2_X1 _11288_ ( .A1(\mtvec [29] ), .A2(fanout_net_43 ), .ZN(_03599_ ) );
AOI21_X1 _11289_ ( .A(fanout_net_2 ), .B1(_03598_ ), .B2(_03599_ ), .ZN(_00257_ ) );
XNOR2_X1 _11290_ ( .A(_03589_ ), .B(_03431_ ), .ZN(_03600_ ) );
NAND2_X1 _11291_ ( .A1(_03600_ ), .A2(_03569_ ), .ZN(_03601_ ) );
OAI211_X1 _11292_ ( .A(_03601_ ), .B(_03557_ ), .C1(\myexu.pc_jump [11] ), .C2(_03546_ ), .ZN(_03602_ ) );
NAND2_X1 _11293_ ( .A1(\mtvec [11] ), .A2(fanout_net_43 ), .ZN(_03603_ ) );
AOI21_X1 _11294_ ( .A(fanout_net_2 ), .B1(_03602_ ), .B2(_03603_ ), .ZN(_00258_ ) );
AND2_X1 _11295_ ( .A1(_03413_ ), .A2(_03436_ ), .ZN(_03604_ ) );
NOR2_X1 _11296_ ( .A1(_03435_ ), .A2(_01686_ ), .ZN(_03605_ ) );
OR2_X1 _11297_ ( .A1(_03604_ ), .A2(_03605_ ), .ZN(_03606_ ) );
OAI21_X1 _11298_ ( .A(_03524_ ), .B1(_03606_ ), .B2(_03440_ ), .ZN(_03607_ ) );
AOI21_X1 _11299_ ( .A(_03607_ ), .B1(_03606_ ), .B2(_03440_ ), .ZN(_03608_ ) );
AOI211_X1 _11300_ ( .A(fanout_net_43 ), .B(_03608_ ), .C1(\myexu.pc_jump [10] ), .C2(_03527_ ), .ZN(_03609_ ) );
NOR2_X1 _11301_ ( .A1(_03521_ ), .A2(\mtvec [10] ), .ZN(_03610_ ) );
NOR3_X1 _11302_ ( .A1(_03609_ ), .A2(fanout_net_2 ), .A3(_03610_ ), .ZN(_00259_ ) );
NOR3_X1 _11303_ ( .A1(_03411_ ), .A2(_03412_ ), .A3(_03436_ ), .ZN(_03611_ ) );
OAI21_X1 _11304_ ( .A(_03538_ ), .B1(_03604_ ), .B2(_03611_ ), .ZN(_03612_ ) );
OAI211_X1 _11305_ ( .A(_03612_ ), .B(_03557_ ), .C1(\myexu.pc_jump [9] ), .C2(_03544_ ), .ZN(_03613_ ) );
NAND2_X1 _11306_ ( .A1(\mtvec [9] ), .A2(fanout_net_43 ), .ZN(_03614_ ) );
AOI21_X1 _11307_ ( .A(fanout_net_2 ), .B1(_03613_ ), .B2(_03614_ ), .ZN(_00260_ ) );
INV_X1 _11308_ ( .A(_03406_ ), .ZN(_03615_ ) );
XNOR2_X1 _11309_ ( .A(_03410_ ), .B(\IF_ID_pc [8] ), .ZN(_03616_ ) );
OAI21_X1 _11310_ ( .A(_03524_ ), .B1(_03615_ ), .B2(_03616_ ), .ZN(_03617_ ) );
AOI21_X1 _11311_ ( .A(_03617_ ), .B1(_03615_ ), .B2(_03616_ ), .ZN(_03618_ ) );
AOI211_X1 _11312_ ( .A(fanout_net_43 ), .B(_03618_ ), .C1(\myexu.pc_jump [8] ), .C2(_03527_ ), .ZN(_03619_ ) );
NOR2_X1 _11313_ ( .A1(_03521_ ), .A2(\mtvec [8] ), .ZN(_03620_ ) );
NOR3_X1 _11314_ ( .A1(_03619_ ), .A2(fanout_net_2 ), .A3(_03620_ ), .ZN(_00261_ ) );
AOI21_X1 _11315_ ( .A(_03401_ ), .B1(_03397_ ), .B2(_03402_ ), .ZN(_03621_ ) );
OAI21_X1 _11316_ ( .A(_03538_ ), .B1(_03403_ ), .B2(_03621_ ), .ZN(_03622_ ) );
OAI211_X1 _11317_ ( .A(_03622_ ), .B(_03557_ ), .C1(\myexu.pc_jump [7] ), .C2(_03544_ ), .ZN(_03623_ ) );
NAND2_X1 _11318_ ( .A1(\mtvec [7] ), .A2(fanout_net_43 ), .ZN(_03624_ ) );
AOI21_X1 _11319_ ( .A(fanout_net_2 ), .B1(_03623_ ), .B2(_03624_ ), .ZN(_00262_ ) );
XNOR2_X1 _11320_ ( .A(_03396_ ), .B(_01808_ ), .ZN(_03625_ ) );
XNOR2_X1 _11321_ ( .A(_03393_ ), .B(_03625_ ), .ZN(_03626_ ) );
NAND2_X1 _11322_ ( .A1(_03626_ ), .A2(_03569_ ), .ZN(_03627_ ) );
OAI211_X1 _11323_ ( .A(_03627_ ), .B(_03557_ ), .C1(\myexu.pc_jump [6] ), .C2(_03544_ ), .ZN(_03628_ ) );
NAND2_X1 _11324_ ( .A1(\mtvec [6] ), .A2(fanout_net_43 ), .ZN(_03629_ ) );
AOI21_X1 _11325_ ( .A(fanout_net_2 ), .B1(_03628_ ), .B2(_03629_ ), .ZN(_00263_ ) );
AND3_X1 _11326_ ( .A1(_03383_ ), .A2(_03384_ ), .A3(_03390_ ), .ZN(_03630_ ) );
OAI21_X1 _11327_ ( .A(_03538_ ), .B1(_03391_ ), .B2(_03630_ ), .ZN(_03631_ ) );
OAI211_X1 _11328_ ( .A(_03631_ ), .B(_03334_ ), .C1(\myexu.pc_jump [5] ), .C2(_03544_ ), .ZN(_03632_ ) );
NAND2_X1 _11329_ ( .A1(\mtvec [5] ), .A2(fanout_net_43 ), .ZN(_03633_ ) );
AOI21_X1 _11330_ ( .A(fanout_net_2 ), .B1(_03632_ ), .B2(_03633_ ), .ZN(_00264_ ) );
NOR2_X1 _11331_ ( .A1(_03380_ ), .A2(_03382_ ), .ZN(_03634_ ) );
INV_X1 _11332_ ( .A(fanout_net_12 ), .ZN(_03635_ ) );
BUF_X2 _11333_ ( .A(_03635_ ), .Z(_03636_ ) );
XNOR2_X1 _11334_ ( .A(_03363_ ), .B(_03636_ ), .ZN(_03637_ ) );
XNOR2_X1 _11335_ ( .A(_03634_ ), .B(_03637_ ), .ZN(_03638_ ) );
NAND2_X1 _11336_ ( .A1(_03638_ ), .A2(_03538_ ), .ZN(_03639_ ) );
NAND3_X1 _11337_ ( .A1(_03332_ ), .A2(check_quest ), .A3(\myexu.pc_jump [4] ), .ZN(_03640_ ) );
AOI21_X1 _11338_ ( .A(fanout_net_43 ), .B1(_03639_ ), .B2(_03640_ ), .ZN(_03641_ ) );
AOI21_X1 _11339_ ( .A(_03641_ ), .B1(\mtvec [4] ), .B2(fanout_net_43 ), .ZN(_03642_ ) );
NOR2_X1 _11340_ ( .A1(_03642_ ), .A2(fanout_net_2 ), .ZN(_00265_ ) );
AND2_X1 _11341_ ( .A1(_03375_ ), .A2(_03379_ ), .ZN(_03643_ ) );
OAI21_X1 _11342_ ( .A(_03524_ ), .B1(_03643_ ), .B2(_03380_ ), .ZN(_03644_ ) );
OAI211_X1 _11343_ ( .A(_03644_ ), .B(_03333_ ), .C1(\myexu.pc_jump [3] ), .C2(_03524_ ), .ZN(_03645_ ) );
NAND2_X1 _11344_ ( .A1(\mtvec [3] ), .A2(fanout_net_43 ), .ZN(_03646_ ) );
AOI21_X1 _11345_ ( .A(fanout_net_2 ), .B1(_03645_ ), .B2(_03646_ ), .ZN(_00266_ ) );
AOI21_X1 _11346_ ( .A(fanout_net_12 ), .B1(IDU_ready_IFU ), .B2(\myifu.state [1] ), .ZN(_03647_ ) );
AND2_X1 _11347_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
AOI211_X1 _11348_ ( .A(fanout_net_2 ), .B(_03647_ ), .C1(_03642_ ), .C2(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_00267_ ) );
AOI21_X1 _11349_ ( .A(_03369_ ), .B1(\IF_ID_pc [1] ), .B2(_03372_ ), .ZN(_03648_ ) );
OAI21_X1 _11350_ ( .A(_03538_ ), .B1(_03373_ ), .B2(_03648_ ), .ZN(_03649_ ) );
OAI211_X1 _11351_ ( .A(_03649_ ), .B(_03334_ ), .C1(\myexu.pc_jump [2] ), .C2(_03544_ ), .ZN(_03650_ ) );
NAND2_X1 _11352_ ( .A1(\mtvec [2] ), .A2(fanout_net_43 ), .ZN(_03651_ ) );
AOI21_X1 _11353_ ( .A(reset ), .B1(_03650_ ), .B2(_03651_ ), .ZN(_00268_ ) );
AND3_X1 _11354_ ( .A1(_03645_ ), .A2(_03646_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_03652_ ) );
INV_X1 _11355_ ( .A(fanout_net_8 ), .ZN(_03653_ ) );
BUF_X4 _11356_ ( .A(_03653_ ), .Z(_03654_ ) );
BUF_X2 _11357_ ( .A(_03654_ ), .Z(_03655_ ) );
INV_X1 _11358_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_03656_ ) );
AOI211_X1 _11359_ ( .A(reset ), .B(_03652_ ), .C1(_03655_ ), .C2(_03656_ ), .ZN(_00269_ ) );
OAI21_X1 _11360_ ( .A(_03505_ ), .B1(_03503_ ), .B2(_03508_ ), .ZN(_03657_ ) );
AND2_X1 _11361_ ( .A1(_03657_ ), .A2(_03512_ ), .ZN(_03658_ ) );
XNOR2_X1 _11362_ ( .A(_03658_ ), .B(_03504_ ), .ZN(_03659_ ) );
MUX2_X1 _11363_ ( .A(\myexu.pc_jump [28] ), .B(_03659_ ), .S(_03524_ ), .Z(_03660_ ) );
MUX2_X1 _11364_ ( .A(\mtvec [28] ), .B(_03660_ ), .S(_03333_ ), .Z(_03661_ ) );
AND2_X1 _11365_ ( .A1(_03661_ ), .A2(_01545_ ), .ZN(_00270_ ) );
XNOR2_X1 _11366_ ( .A(_03372_ ), .B(\IF_ID_pc [1] ), .ZN(_03662_ ) );
NAND2_X1 _11367_ ( .A1(_03662_ ), .A2(_03569_ ), .ZN(_03663_ ) );
OAI211_X1 _11368_ ( .A(_03663_ ), .B(_03334_ ), .C1(\myexu.pc_jump [1] ), .C2(_03544_ ), .ZN(_03664_ ) );
NAND2_X1 _11369_ ( .A1(\mtvec [1] ), .A2(fanout_net_43 ), .ZN(_03665_ ) );
AOI21_X1 _11370_ ( .A(reset ), .B1(_03664_ ), .B2(_03665_ ), .ZN(_00271_ ) );
NOR2_X1 _11371_ ( .A1(_03503_ ), .A2(_03508_ ), .ZN(_03666_ ) );
XOR2_X1 _11372_ ( .A(_03666_ ), .B(_03505_ ), .Z(_03667_ ) );
NAND2_X1 _11373_ ( .A1(_03667_ ), .A2(_03569_ ), .ZN(_03668_ ) );
OAI211_X1 _11374_ ( .A(_03668_ ), .B(_03334_ ), .C1(\myexu.pc_jump [27] ), .C2(_03544_ ), .ZN(_03669_ ) );
NAND2_X1 _11375_ ( .A1(\mtvec [27] ), .A2(fanout_net_43 ), .ZN(_03670_ ) );
AOI21_X1 _11376_ ( .A(reset ), .B1(_03669_ ), .B2(_03670_ ), .ZN(_00272_ ) );
OAI21_X1 _11377_ ( .A(_03502_ ), .B1(_03494_ ), .B2(_03498_ ), .ZN(_03671_ ) );
OAI21_X1 _11378_ ( .A(_03671_ ), .B1(_01788_ ), .B2(_03507_ ), .ZN(_03672_ ) );
XOR2_X1 _11379_ ( .A(_03672_ ), .B(_03501_ ), .Z(_03673_ ) );
MUX2_X1 _11380_ ( .A(\myexu.pc_jump [26] ), .B(_03673_ ), .S(_03524_ ), .Z(_03674_ ) );
MUX2_X1 _11381_ ( .A(\mtvec [26] ), .B(_03674_ ), .S(_03333_ ), .Z(_03675_ ) );
AND2_X1 _11382_ ( .A1(_03675_ ), .A2(_01545_ ), .ZN(_00273_ ) );
XOR2_X1 _11383_ ( .A(_03499_ ), .B(_03502_ ), .Z(_03676_ ) );
NAND2_X1 _11384_ ( .A1(_03676_ ), .A2(_03569_ ), .ZN(_03677_ ) );
OAI211_X1 _11385_ ( .A(_03677_ ), .B(_03334_ ), .C1(\myexu.pc_jump [25] ), .C2(_03544_ ), .ZN(_03678_ ) );
NAND2_X1 _11386_ ( .A1(\mtvec [25] ), .A2(fanout_net_43 ), .ZN(_03679_ ) );
AOI21_X1 _11387_ ( .A(reset ), .B1(_03678_ ), .B2(_03679_ ), .ZN(_00274_ ) );
NAND2_X1 _11388_ ( .A1(_03487_ ), .A2(_03493_ ), .ZN(_03680_ ) );
OAI21_X1 _11389_ ( .A(_03483_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_03681_ ) );
NAND2_X1 _11390_ ( .A1(_03680_ ), .A2(_03681_ ), .ZN(_03682_ ) );
AND2_X1 _11391_ ( .A1(_03682_ ), .A2(_03489_ ), .ZN(_03683_ ) );
AND2_X1 _11392_ ( .A1(_03483_ ), .A2(\IF_ID_pc [23] ), .ZN(_03684_ ) );
NOR2_X1 _11393_ ( .A1(_03683_ ), .A2(_03684_ ), .ZN(_03685_ ) );
XNOR2_X1 _11394_ ( .A(_03685_ ), .B(_03488_ ), .ZN(_03686_ ) );
AND2_X1 _11395_ ( .A1(_03686_ ), .A2(_03538_ ), .ZN(_03687_ ) );
AOI211_X1 _11396_ ( .A(fanout_net_43 ), .B(_03687_ ), .C1(\myexu.pc_jump [24] ), .C2(_03527_ ), .ZN(_03688_ ) );
NOR2_X1 _11397_ ( .A1(_03521_ ), .A2(\mtvec [24] ), .ZN(_03689_ ) );
NOR3_X1 _11398_ ( .A1(_03688_ ), .A2(reset ), .A3(_03689_ ), .ZN(_00275_ ) );
NOR2_X1 _11399_ ( .A1(_03682_ ), .A2(_03489_ ), .ZN(_03690_ ) );
NOR3_X1 _11400_ ( .A1(_03683_ ), .A2(_03690_ ), .A3(_03143_ ), .ZN(_03691_ ) );
AOI211_X1 _11401_ ( .A(fanout_net_43 ), .B(_03691_ ), .C1(\myexu.pc_jump [23] ), .C2(_03527_ ), .ZN(_03692_ ) );
NOR2_X1 _11402_ ( .A1(_03521_ ), .A2(\mtvec [23] ), .ZN(_03693_ ) );
NOR3_X1 _11403_ ( .A1(_03692_ ), .A2(reset ), .A3(_03693_ ), .ZN(_00276_ ) );
OAI21_X1 _11404_ ( .A(_03525_ ), .B1(_01728_ ), .B2(_03507_ ), .ZN(_03694_ ) );
XNOR2_X1 _11405_ ( .A(_03694_ ), .B(_03491_ ), .ZN(_03695_ ) );
NOR2_X1 _11406_ ( .A1(_03695_ ), .A2(_03143_ ), .ZN(_03696_ ) );
AOI211_X1 _11407_ ( .A(\myifu.to_reset ), .B(_03696_ ), .C1(\myexu.pc_jump [22] ), .C2(_03527_ ), .ZN(_03697_ ) );
NOR2_X1 _11408_ ( .A1(_03521_ ), .A2(\mtvec [22] ), .ZN(_03698_ ) );
NOR3_X1 _11409_ ( .A1(_03697_ ), .A2(reset ), .A3(_03698_ ), .ZN(_00277_ ) );
NAND2_X1 _11410_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_03699_ ) );
OAI22_X1 _11411_ ( .A1(_03514_ ), .A2(_03515_ ), .B1(\IF_ID_pc [30] ), .B2(_03342_ ), .ZN(_03700_ ) );
NAND3_X1 _11412_ ( .A1(_03482_ ), .A2(\IF_ID_pc [30] ), .A3(_03354_ ), .ZN(_03701_ ) );
NAND2_X1 _11413_ ( .A1(_03700_ ), .A2(_03701_ ), .ZN(_03702_ ) );
XNOR2_X1 _11414_ ( .A(_03342_ ), .B(\IF_ID_pc [31] ), .ZN(_03703_ ) );
OAI21_X1 _11415_ ( .A(_03538_ ), .B1(_03702_ ), .B2(_03703_ ), .ZN(_03704_ ) );
AOI21_X1 _11416_ ( .A(_03704_ ), .B1(_03702_ ), .B2(_03703_ ), .ZN(_03705_ ) );
OAI21_X1 _11417_ ( .A(_03334_ ), .B1(_03546_ ), .B2(\myexu.pc_jump [31] ), .ZN(_03706_ ) );
OAI211_X1 _11418_ ( .A(_01545_ ), .B(_03699_ ), .C1(_03705_ ), .C2(_03706_ ), .ZN(_00278_ ) );
NOR2_X2 _11419_ ( .A1(_01914_ ), .A2(_01988_ ), .ZN(_03707_ ) );
INV_X1 _11420_ ( .A(_03707_ ), .ZN(_03708_ ) );
NOR2_X1 _11421_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_03709_ ) );
NOR2_X1 _11422_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_03710_ ) );
INV_X1 _11423_ ( .A(\io_master_rid [1] ), .ZN(_03711_ ) );
NAND4_X1 _11424_ ( .A1(_03709_ ), .A2(_03710_ ), .A3(_03711_ ), .A4(\io_master_rid [0] ), .ZN(_03712_ ) );
AOI21_X1 _11425_ ( .A(_01883_ ), .B1(_03708_ ), .B2(_03712_ ), .ZN(_03713_ ) );
AND2_X1 _11426_ ( .A1(_01998_ ), .A2(_02001_ ), .ZN(_03714_ ) );
NOR2_X1 _11427_ ( .A1(_03714_ ), .A2(io_master_rlast ), .ZN(_03715_ ) );
INV_X1 _11428_ ( .A(_03715_ ), .ZN(_03716_ ) );
INV_X1 _11429_ ( .A(_01965_ ), .ZN(\io_master_araddr [21] ) );
INV_X1 _11430_ ( .A(_01982_ ), .ZN(\io_master_araddr [22] ) );
NOR4_X1 _11431_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [22] ), .A3(\io_master_araddr [23] ), .A4(\io_master_araddr [20] ), .ZN(_03717_ ) );
INV_X1 _11432_ ( .A(_01969_ ), .ZN(\io_master_araddr [19] ) );
INV_X1 _11433_ ( .A(_01986_ ), .ZN(\io_master_araddr [16] ) );
NOR4_X1 _11434_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [16] ), .A3(\io_master_araddr [17] ), .A4(\io_master_araddr [18] ), .ZN(_03718_ ) );
AND2_X2 _11435_ ( .A1(_03717_ ), .A2(_03718_ ), .ZN(_03719_ ) );
NAND4_X1 _11436_ ( .A1(_01893_ ), .A2(_01897_ ), .A3(_01957_ ), .A4(_01974_ ), .ZN(_03720_ ) );
NAND4_X4 _11437_ ( .A1(_01901_ ), .A2(_01961_ ), .A3(_01978_ ), .A4(\io_master_araddr [25] ), .ZN(_03721_ ) );
NOR2_X2 _11438_ ( .A1(_03720_ ), .A2(_03721_ ), .ZN(_03722_ ) );
AOI21_X1 _11439_ ( .A(io_master_rvalid ), .B1(_03719_ ), .B2(_03722_ ), .ZN(_03723_ ) );
AND4_X1 _11440_ ( .A1(\myclint.state_r_$_NOT__A_Y ), .A2(_03717_ ), .A3(_03718_ ), .A4(_03722_ ), .ZN(_03724_ ) );
NOR2_X1 _11441_ ( .A1(_03723_ ), .A2(_03724_ ), .ZN(_03725_ ) );
NAND3_X1 _11442_ ( .A1(_03713_ ), .A2(_03716_ ), .A3(_03725_ ), .ZN(_03726_ ) );
INV_X1 _11443_ ( .A(\myifu.tmp_offset [2] ), .ZN(_03727_ ) );
AND3_X1 _11444_ ( .A1(_03726_ ), .A2(_01460_ ), .A3(_03727_ ), .ZN(_00279_ ) );
NOR3_X1 _11445_ ( .A1(reset ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00280_ ) );
AND3_X1 _11446_ ( .A1(_02017_ ), .A2(_03144_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_03728_ ) );
INV_X1 _11447_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_03729_ ) );
MUX2_X1 _11448_ ( .A(_02017_ ), .B(_03729_ ), .S(\myifu.to_reset ), .Z(_03730_ ) );
AOI211_X1 _11449_ ( .A(reset ), .B(_03728_ ), .C1(_03730_ ), .C2(\myifu.state [1] ), .ZN(_00281_ ) );
INV_X1 _11450_ ( .A(_01944_ ), .ZN(_03731_ ) );
NOR2_X1 _11451_ ( .A1(_01951_ ), .A2(_03731_ ), .ZN(_03732_ ) );
INV_X1 _11452_ ( .A(_03732_ ), .ZN(_03733_ ) );
BUF_X2 _11453_ ( .A(_03733_ ), .Z(_03734_ ) );
BUF_X4 _11454_ ( .A(_02039_ ), .Z(_03735_ ) );
MUX2_X1 _11455_ ( .A(\LS_WB_waddr_csreg [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_03735_ ), .Z(_03736_ ) );
NOR2_X1 _11456_ ( .A1(_01924_ ), .A2(\EX_LS_flag [1] ), .ZN(_03737_ ) );
OR2_X1 _11457_ ( .A1(_03737_ ), .A2(_01923_ ), .ZN(_03738_ ) );
NOR2_X1 _11458_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_03739_ ) );
AND2_X2 _11459_ ( .A1(_03739_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_03740_ ) );
NOR2_X2 _11460_ ( .A1(_03738_ ), .A2(_03740_ ), .ZN(_03741_ ) );
BUF_X4 _11461_ ( .A(_03741_ ), .Z(_03742_ ) );
BUF_X2 _11462_ ( .A(_03742_ ), .Z(_03743_ ) );
AND3_X1 _11463_ ( .A1(_03734_ ), .A2(_03736_ ), .A3(_03743_ ), .ZN(_00284_ ) );
BUF_X4 _11464_ ( .A(_01925_ ), .Z(_03744_ ) );
NOR2_X1 _11465_ ( .A1(_03732_ ), .A2(_03740_ ), .ZN(_03745_ ) );
INV_X1 _11466_ ( .A(_03745_ ), .ZN(_03746_ ) );
NAND3_X1 _11467_ ( .A1(_01943_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_03747_ ) );
BUF_X4 _11468_ ( .A(_01924_ ), .Z(_03748_ ) );
BUF_X4 _11469_ ( .A(_03748_ ), .Z(_03749_ ) );
NAND2_X1 _11470_ ( .A1(_03749_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03750_ ) );
AOI211_X1 _11471_ ( .A(_03744_ ), .B(_03746_ ), .C1(_03747_ ), .C2(_03750_ ), .ZN(_00285_ ) );
NAND3_X1 _11472_ ( .A1(_01943_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_03751_ ) );
NAND2_X1 _11473_ ( .A1(_03749_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_03752_ ) );
AOI211_X1 _11474_ ( .A(_03744_ ), .B(_03746_ ), .C1(_03751_ ), .C2(_03752_ ), .ZN(_00286_ ) );
NAND3_X1 _11475_ ( .A1(_01943_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_03753_ ) );
NAND2_X1 _11476_ ( .A1(_03749_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_03754_ ) );
AOI211_X1 _11477_ ( .A(_03744_ ), .B(_03746_ ), .C1(_03753_ ), .C2(_03754_ ), .ZN(_00287_ ) );
NAND3_X1 _11478_ ( .A1(_01943_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_03755_ ) );
NAND2_X1 _11479_ ( .A1(_03749_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03756_ ) );
AOI211_X1 _11480_ ( .A(_03744_ ), .B(_03746_ ), .C1(_03755_ ), .C2(_03756_ ), .ZN(_00288_ ) );
NAND3_X1 _11481_ ( .A1(_01943_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_03757_ ) );
NAND2_X1 _11482_ ( .A1(_03749_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_03758_ ) );
AOI211_X1 _11483_ ( .A(_03744_ ), .B(_03746_ ), .C1(_03757_ ), .C2(_03758_ ), .ZN(_00289_ ) );
NAND3_X1 _11484_ ( .A1(_01943_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_03759_ ) );
NAND2_X1 _11485_ ( .A1(_03749_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_03760_ ) );
AOI211_X1 _11486_ ( .A(_03744_ ), .B(_03746_ ), .C1(_03759_ ), .C2(_03760_ ), .ZN(_00290_ ) );
NAND3_X1 _11487_ ( .A1(_01943_ ), .A2(fanout_net_4 ), .A3(\EX_LS_flag [2] ), .ZN(_03761_ ) );
NAND2_X1 _11488_ ( .A1(_03749_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_03762_ ) );
AOI211_X1 _11489_ ( .A(_03744_ ), .B(_03746_ ), .C1(_03761_ ), .C2(_03762_ ), .ZN(_00291_ ) );
INV_X1 _11490_ ( .A(_03744_ ), .ZN(_03763_ ) );
INV_X1 _11491_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_03764_ ) );
AND4_X1 _11492_ ( .A1(_03764_ ), .A2(_01871_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03765_ ) );
NOR2_X1 _11493_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_03766_ ) );
OAI211_X1 _11494_ ( .A(_03745_ ), .B(_03763_ ), .C1(_03765_ ), .C2(_03766_ ), .ZN(_00292_ ) );
NOR4_X1 _11495_ ( .A1(_03749_ ), .A2(_01870_ ), .A3(\EX_LS_dest_csreg_mem [8] ), .A4(\EX_LS_flag [0] ), .ZN(_03767_ ) );
NOR2_X1 _11496_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_03768_ ) );
OAI211_X1 _11497_ ( .A(_03745_ ), .B(_03763_ ), .C1(_03767_ ), .C2(_03768_ ), .ZN(_00293_ ) );
NOR4_X1 _11498_ ( .A1(_03749_ ), .A2(_01870_ ), .A3(\EX_LS_dest_csreg_mem [6] ), .A4(\EX_LS_flag [0] ), .ZN(_03769_ ) );
NOR2_X1 _11499_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_03770_ ) );
OAI211_X1 _11500_ ( .A(_03745_ ), .B(_03763_ ), .C1(_03769_ ), .C2(_03770_ ), .ZN(_00294_ ) );
INV_X1 _11501_ ( .A(fanout_net_3 ), .ZN(_03771_ ) );
AND4_X1 _11502_ ( .A1(_03771_ ), .A2(_01871_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03772_ ) );
NOR2_X1 _11503_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_03773_ ) );
OAI211_X1 _11504_ ( .A(_03745_ ), .B(_03763_ ), .C1(_03772_ ), .C2(_03773_ ), .ZN(_00295_ ) );
INV_X1 _11505_ ( .A(\mysc.state [2] ), .ZN(_03774_ ) );
NOR2_X1 _11506_ ( .A1(_03774_ ), .A2(reset ), .ZN(_00303_ ) );
NOR2_X1 _11507_ ( .A1(_03248_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _11508_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_03775_ ) );
NOR2_X1 _11509_ ( .A1(_03259_ ), .A2(\ID_EX_typ [6] ), .ZN(_03776_ ) );
AND2_X1 _11510_ ( .A1(_03776_ ), .A2(\ID_EX_typ [5] ), .ZN(_03777_ ) );
BUF_X2 _11511_ ( .A(_03777_ ), .Z(_03778_ ) );
INV_X2 _11512_ ( .A(fanout_net_5 ), .ZN(_03779_ ) );
AND2_X2 _11513_ ( .A1(_03778_ ), .A2(_03779_ ), .ZN(_03780_ ) );
INV_X1 _11514_ ( .A(_03780_ ), .ZN(_03781_ ) );
INV_X1 _11515_ ( .A(\ID_EX_typ [5] ), .ZN(_03782_ ) );
INV_X1 _11516_ ( .A(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03783_ ) );
NAND3_X1 _11517_ ( .A1(_03776_ ), .A2(_03782_ ), .A3(_03783_ ), .ZN(_03784_ ) );
AOI21_X1 _11518_ ( .A(_03775_ ), .B1(_03781_ ), .B2(_03784_ ), .ZN(_03785_ ) );
INV_X1 _11519_ ( .A(\myec.state [1] ), .ZN(_03786_ ) );
NAND2_X1 _11520_ ( .A1(_03786_ ), .A2(\myec.state [0] ), .ZN(_03787_ ) );
NOR2_X1 _11521_ ( .A1(reset ), .A2(excp_written ), .ZN(_03788_ ) );
AND2_X1 _11522_ ( .A1(_03787_ ), .A2(_03788_ ), .ZN(_03789_ ) );
BUF_X2 _11523_ ( .A(_03789_ ), .Z(_03790_ ) );
INV_X1 _11524_ ( .A(\ID_EX_typ [6] ), .ZN(_03791_ ) );
CLKBUF_X2 _11525_ ( .A(_01886_ ), .Z(_03792_ ) );
CLKBUF_X2 _11526_ ( .A(_03792_ ), .Z(_03793_ ) );
AND4_X1 _11527_ ( .A1(\ID_EX_typ [7] ), .A2(_03791_ ), .A3(_03793_ ), .A4(IDU_valid_EXU ), .ZN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _11528_ ( .A1(_03142_ ), .A2(check_assert ), .ZN(_03794_ ) );
OAI21_X1 _11529_ ( .A(_03790_ ), .B1(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(_03794_ ), .ZN(_03795_ ) );
NOR2_X1 _11530_ ( .A1(_03785_ ), .A2(_03795_ ), .ZN(_00096_ ) );
CLKBUF_X2 _11531_ ( .A(_03787_ ), .Z(_03796_ ) );
CLKBUF_X2 _11532_ ( .A(_03796_ ), .Z(_03797_ ) );
CLKBUF_X2 _11533_ ( .A(_03788_ ), .Z(_03798_ ) );
CLKBUF_X2 _11534_ ( .A(_03798_ ), .Z(_03799_ ) );
AND3_X1 _11535_ ( .A1(_03797_ ), .A2(\ID_EX_rd [4] ), .A3(_03799_ ), .ZN(_00117_ ) );
AND3_X1 _11536_ ( .A1(_03797_ ), .A2(\ID_EX_rd [3] ), .A3(_03799_ ), .ZN(_00118_ ) );
AND3_X1 _11537_ ( .A1(_03797_ ), .A2(\ID_EX_rd [2] ), .A3(_03799_ ), .ZN(_00119_ ) );
AND3_X1 _11538_ ( .A1(_03797_ ), .A2(\ID_EX_rd [1] ), .A3(_03799_ ), .ZN(_00120_ ) );
AND3_X1 _11539_ ( .A1(_03797_ ), .A2(\ID_EX_rd [0] ), .A3(_03799_ ), .ZN(_00121_ ) );
INV_X2 _11540_ ( .A(_03789_ ), .ZN(_03800_ ) );
BUF_X4 _11541_ ( .A(_03800_ ), .Z(_03801_ ) );
INV_X1 _11542_ ( .A(\EX_LS_dest_csreg_mem [7] ), .ZN(_03802_ ) );
AOI22_X1 _11543_ ( .A1(_03764_ ), .A2(\ID_EX_csr [9] ), .B1(_03802_ ), .B2(\ID_EX_csr [7] ), .ZN(_03803_ ) );
XNOR2_X1 _11544_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_03804_ ) );
INV_X1 _11545_ ( .A(\ID_EX_csr [0] ), .ZN(_03805_ ) );
INV_X1 _11546_ ( .A(\ID_EX_csr [7] ), .ZN(_03806_ ) );
AOI22_X1 _11547_ ( .A1(fanout_net_3 ), .A2(_03805_ ), .B1(_03806_ ), .B2(\EX_LS_dest_csreg_mem [7] ), .ZN(_03807_ ) );
NAND4_X1 _11548_ ( .A1(_02039_ ), .A2(_03803_ ), .A3(_03804_ ), .A4(_03807_ ), .ZN(_03808_ ) );
XOR2_X1 _11549_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .Z(_03809_ ) );
XNOR2_X1 _11550_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_03810_ ) );
XNOR2_X1 _11551_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_03811_ ) );
NAND2_X1 _11552_ ( .A1(_03810_ ), .A2(_03811_ ), .ZN(_03812_ ) );
NOR3_X1 _11553_ ( .A1(_03808_ ), .A2(_03809_ ), .A3(_03812_ ), .ZN(_03813_ ) );
BUF_X2 _11554_ ( .A(_03813_ ), .Z(_03814_ ) );
BUF_X2 _11555_ ( .A(_03814_ ), .Z(_03815_ ) );
INV_X1 _11556_ ( .A(\ID_EX_csr [5] ), .ZN(_03816_ ) );
AOI22_X1 _11557_ ( .A1(_03771_ ), .A2(\ID_EX_csr [0] ), .B1(_03816_ ), .B2(\EX_LS_dest_csreg_mem [5] ), .ZN(_03817_ ) );
INV_X1 _11558_ ( .A(fanout_net_4 ), .ZN(_03818_ ) );
OAI221_X1 _11559_ ( .A(_03817_ ), .B1(_03818_ ), .B2(\ID_EX_csr [1] ), .C1(\EX_LS_dest_csreg_mem [5] ), .C2(_03816_ ), .ZN(_03819_ ) );
XNOR2_X1 _11560_ ( .A(\EX_LS_dest_csreg_mem [8] ), .B(\ID_EX_csr [8] ), .ZN(_03820_ ) );
INV_X1 _11561_ ( .A(\ID_EX_csr [3] ), .ZN(_03821_ ) );
OR2_X1 _11562_ ( .A1(_03821_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .ZN(_03822_ ) );
OAI211_X1 _11563_ ( .A(_03820_ ), .B(_03822_ ), .C1(_03764_ ), .C2(\ID_EX_csr [9] ), .ZN(_03823_ ) );
INV_X1 _11564_ ( .A(\ID_EX_csr [4] ), .ZN(_03824_ ) );
AOI22_X1 _11565_ ( .A1(_03818_ ), .A2(\ID_EX_csr [1] ), .B1(_03824_ ), .B2(\EX_LS_dest_csreg_mem [4] ), .ZN(_03825_ ) );
NAND2_X1 _11566_ ( .A1(_03821_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .ZN(_03826_ ) );
OAI211_X1 _11567_ ( .A(_03825_ ), .B(_03826_ ), .C1(\EX_LS_dest_csreg_mem [4] ), .C2(_03824_ ), .ZN(_03827_ ) );
NOR3_X1 _11568_ ( .A1(_03819_ ), .A2(_03823_ ), .A3(_03827_ ), .ZN(_03828_ ) );
BUF_X2 _11569_ ( .A(_03828_ ), .Z(_03829_ ) );
BUF_X2 _11570_ ( .A(_03829_ ), .Z(_03830_ ) );
NAND3_X1 _11571_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(\EX_LS_result_csreg_mem [30] ), .ZN(_03831_ ) );
NOR2_X1 _11572_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_03832_ ) );
NAND3_X1 _11573_ ( .A1(_03832_ ), .A2(_03816_ ), .A3(_03824_ ), .ZN(_03833_ ) );
INV_X1 _11574_ ( .A(\ID_EX_csr [11] ), .ZN(_03834_ ) );
NAND3_X1 _11575_ ( .A1(_03834_ ), .A2(\ID_EX_csr [9] ), .A3(\ID_EX_csr [8] ), .ZN(_03835_ ) );
NOR3_X1 _11576_ ( .A1(_03833_ ), .A2(\ID_EX_csr [10] ), .A3(_03835_ ), .ZN(_03836_ ) );
CLKBUF_X2 _11577_ ( .A(_03836_ ), .Z(_03837_ ) );
BUF_X2 _11578_ ( .A(_03837_ ), .Z(_03838_ ) );
NOR2_X1 _11579_ ( .A1(_03805_ ), .A2(\ID_EX_csr [1] ), .ZN(_03839_ ) );
AND3_X1 _11580_ ( .A1(_03839_ ), .A2(_03821_ ), .A3(\ID_EX_csr [2] ), .ZN(_03840_ ) );
BUF_X2 _11581_ ( .A(_03840_ ), .Z(_03841_ ) );
BUF_X2 _11582_ ( .A(_03841_ ), .Z(_03842_ ) );
NAND3_X1 _11583_ ( .A1(_03838_ ), .A2(\mtvec [30] ), .A3(_03842_ ), .ZN(_03843_ ) );
INV_X1 _11584_ ( .A(\ID_EX_csr [6] ), .ZN(_03844_ ) );
NOR3_X1 _11585_ ( .A1(_03844_ ), .A2(\ID_EX_csr [5] ), .A3(\ID_EX_csr [4] ), .ZN(_03845_ ) );
NAND2_X1 _11586_ ( .A1(_03845_ ), .A2(_03806_ ), .ZN(_03846_ ) );
NOR3_X1 _11587_ ( .A1(_03846_ ), .A2(\ID_EX_csr [10] ), .A3(_03835_ ), .ZN(_03847_ ) );
CLKBUF_X2 _11588_ ( .A(_03847_ ), .Z(_03848_ ) );
NOR2_X1 _11589_ ( .A1(\ID_EX_csr [3] ), .A2(\ID_EX_csr [2] ), .ZN(_03849_ ) );
AND2_X1 _11590_ ( .A1(_03839_ ), .A2(_03849_ ), .ZN(_03850_ ) );
BUF_X2 _11591_ ( .A(_03850_ ), .Z(_03851_ ) );
NAND3_X1 _11592_ ( .A1(_03848_ ), .A2(\mepc [30] ), .A3(_03851_ ), .ZN(_03852_ ) );
INV_X1 _11593_ ( .A(\ID_EX_csr [2] ), .ZN(_03853_ ) );
NAND3_X1 _11594_ ( .A1(_03821_ ), .A2(_03853_ ), .A3(\ID_EX_csr [1] ), .ZN(_03854_ ) );
NOR2_X1 _11595_ ( .A1(_03854_ ), .A2(\ID_EX_csr [0] ), .ZN(_03855_ ) );
CLKBUF_X3 _11596_ ( .A(_03855_ ), .Z(_03856_ ) );
NAND3_X1 _11597_ ( .A1(_03848_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_03856_ ), .ZN(_03857_ ) );
AND2_X1 _11598_ ( .A1(_03852_ ), .A2(_03857_ ), .ZN(_03858_ ) );
AND4_X1 _11599_ ( .A1(\ID_EX_csr [10] ), .A2(_03816_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_03859_ ) );
AND2_X1 _11600_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_03860_ ) );
AND3_X2 _11601_ ( .A1(_03859_ ), .A2(_03860_ ), .A3(_03832_ ), .ZN(_03861_ ) );
AND2_X1 _11602_ ( .A1(_03861_ ), .A2(_03850_ ), .ZN(_03862_ ) );
INV_X1 _11603_ ( .A(_03862_ ), .ZN(_03863_ ) );
BUF_X2 _11604_ ( .A(_03837_ ), .Z(_03864_ ) );
INV_X1 _11605_ ( .A(\ID_EX_csr [1] ), .ZN(_03865_ ) );
AND3_X2 _11606_ ( .A1(_03849_ ), .A2(_03865_ ), .A3(_03805_ ), .ZN(_03866_ ) );
BUF_X2 _11607_ ( .A(_03866_ ), .Z(_03867_ ) );
NAND3_X1 _11608_ ( .A1(_03864_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_03867_ ), .ZN(_03868_ ) );
AND4_X1 _11609_ ( .A1(_03843_ ), .A2(_03858_ ), .A3(_03863_ ), .A4(_03868_ ), .ZN(_03869_ ) );
AND2_X1 _11610_ ( .A1(_03813_ ), .A2(_03828_ ), .ZN(_03870_ ) );
BUF_X4 _11611_ ( .A(_03870_ ), .Z(_03871_ ) );
OAI21_X1 _11612_ ( .A(_03831_ ), .B1(_03869_ ), .B2(_03871_ ), .ZN(_03872_ ) );
AND2_X1 _11613_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_03873_ ) );
AND2_X1 _11614_ ( .A1(_03873_ ), .A2(\ID_EX_pc [4] ), .ZN(_03874_ ) );
AND2_X1 _11615_ ( .A1(_03874_ ), .A2(\ID_EX_pc [5] ), .ZN(_03875_ ) );
AND2_X1 _11616_ ( .A1(_03875_ ), .A2(\ID_EX_pc [6] ), .ZN(_03876_ ) );
AND2_X1 _11617_ ( .A1(_03876_ ), .A2(\ID_EX_pc [7] ), .ZN(_03877_ ) );
AND2_X1 _11618_ ( .A1(_03877_ ), .A2(\ID_EX_pc [8] ), .ZN(_03878_ ) );
AND2_X2 _11619_ ( .A1(_03878_ ), .A2(\ID_EX_pc [9] ), .ZN(_03879_ ) );
AND2_X1 _11620_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_03880_ ) );
AND2_X1 _11621_ ( .A1(_03879_ ), .A2(_03880_ ), .ZN(_03881_ ) );
AND3_X1 _11622_ ( .A1(_03881_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_03882_ ) );
AND3_X1 _11623_ ( .A1(_03882_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_03883_ ) );
AND3_X1 _11624_ ( .A1(_03883_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_03884_ ) );
AND3_X1 _11625_ ( .A1(_03884_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_03885_ ) );
AND3_X1 _11626_ ( .A1(_03885_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_03886_ ) );
AND3_X1 _11627_ ( .A1(_03886_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_03887_ ) );
AND3_X1 _11628_ ( .A1(_03887_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_03888_ ) );
AND3_X1 _11629_ ( .A1(_03888_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_03889_ ) );
NAND3_X1 _11630_ ( .A1(_03889_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_03890_ ) );
XNOR2_X1 _11631_ ( .A(_03890_ ), .B(\ID_EX_pc [30] ), .ZN(_03891_ ) );
NOR2_X1 _11632_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_03892_ ) );
XOR2_X1 _11633_ ( .A(\ID_EX_pc [25] ), .B(\ID_EX_imm [25] ), .Z(_03893_ ) );
XOR2_X1 _11634_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_03894_ ) );
XOR2_X1 _11635_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_03895_ ) );
XOR2_X1 _11636_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_03896_ ) );
AND2_X1 _11637_ ( .A1(_03895_ ), .A2(_03896_ ), .ZN(_03897_ ) );
XOR2_X1 _11638_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_03898_ ) );
NOR2_X1 _11639_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03899_ ) );
XOR2_X1 _11640_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_03900_ ) );
XOR2_X1 _11641_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_03901_ ) );
AND2_X1 _11642_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_03902_ ) );
AND2_X1 _11643_ ( .A1(_03901_ ), .A2(_03902_ ), .ZN(_03903_ ) );
AND2_X1 _11644_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_03904_ ) );
OAI21_X1 _11645_ ( .A(_03900_ ), .B1(_03903_ ), .B2(_03904_ ), .ZN(_03905_ ) );
NAND2_X1 _11646_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_03906_ ) );
AOI21_X1 _11647_ ( .A(_03899_ ), .B1(_03905_ ), .B2(_03906_ ), .ZN(_03907_ ) );
AND2_X1 _11648_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03908_ ) );
OAI21_X1 _11649_ ( .A(_03898_ ), .B1(_03907_ ), .B2(_03908_ ), .ZN(_03909_ ) );
NAND2_X1 _11650_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03910_ ) );
NAND2_X1 _11651_ ( .A1(_03909_ ), .A2(_03910_ ), .ZN(_03911_ ) );
OAI21_X1 _11652_ ( .A(_03911_ ), .B1(\ID_EX_pc [5] ), .B2(\ID_EX_imm [5] ), .ZN(_03912_ ) );
AND2_X1 _11653_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03913_ ) );
INV_X1 _11654_ ( .A(_03913_ ), .ZN(_03914_ ) );
NAND2_X1 _11655_ ( .A1(_03912_ ), .A2(_03914_ ), .ZN(_03915_ ) );
XOR2_X1 _11656_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_03916_ ) );
NAND2_X1 _11657_ ( .A1(_03915_ ), .A2(_03916_ ), .ZN(_03917_ ) );
NAND2_X1 _11658_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03918_ ) );
NAND2_X1 _11659_ ( .A1(_03917_ ), .A2(_03918_ ), .ZN(_03919_ ) );
OAI21_X1 _11660_ ( .A(_03919_ ), .B1(\ID_EX_pc [7] ), .B2(\ID_EX_imm [7] ), .ZN(_03920_ ) );
AND2_X1 _11661_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03921_ ) );
INV_X1 _11662_ ( .A(_03921_ ), .ZN(_03922_ ) );
NAND2_X1 _11663_ ( .A1(_03920_ ), .A2(_03922_ ), .ZN(_03923_ ) );
XOR2_X1 _11664_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_03924_ ) );
XOR2_X1 _11665_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_03925_ ) );
AND2_X1 _11666_ ( .A1(_03924_ ), .A2(_03925_ ), .ZN(_03926_ ) );
XOR2_X1 _11667_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_03927_ ) );
XOR2_X1 _11668_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_03928_ ) );
AND2_X1 _11669_ ( .A1(_03927_ ), .A2(_03928_ ), .ZN(_03929_ ) );
AND3_X1 _11670_ ( .A1(_03923_ ), .A2(_03926_ ), .A3(_03929_ ), .ZN(_03930_ ) );
AND2_X1 _11671_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_03931_ ) );
AND2_X1 _11672_ ( .A1(_03924_ ), .A2(_03931_ ), .ZN(_03932_ ) );
AOI21_X1 _11673_ ( .A(_03932_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_03933_ ) );
AND2_X1 _11674_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_03934_ ) );
AND2_X1 _11675_ ( .A1(_03928_ ), .A2(_03934_ ), .ZN(_03935_ ) );
AOI21_X1 _11676_ ( .A(_03935_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_03936_ ) );
INV_X1 _11677_ ( .A(_03926_ ), .ZN(_03937_ ) );
OAI21_X1 _11678_ ( .A(_03933_ ), .B1(_03936_ ), .B2(_03937_ ), .ZN(_03938_ ) );
OR2_X1 _11679_ ( .A1(_03930_ ), .A2(_03938_ ), .ZN(_03939_ ) );
XOR2_X1 _11680_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_03940_ ) );
XOR2_X1 _11681_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_03941_ ) );
XOR2_X1 _11682_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_03942_ ) );
XOR2_X1 _11683_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .Z(_03943_ ) );
AND2_X1 _11684_ ( .A1(_03942_ ), .A2(_03943_ ), .ZN(_03944_ ) );
NAND4_X1 _11685_ ( .A1(_03939_ ), .A2(_03940_ ), .A3(_03941_ ), .A4(_03944_ ), .ZN(_03945_ ) );
AND2_X1 _11686_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_03946_ ) );
AND2_X1 _11687_ ( .A1(_03943_ ), .A2(_03946_ ), .ZN(_03947_ ) );
AOI21_X1 _11688_ ( .A(_03947_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_03948_ ) );
NAND2_X1 _11689_ ( .A1(_03940_ ), .A2(_03941_ ), .ZN(_03949_ ) );
NOR2_X1 _11690_ ( .A1(_03948_ ), .A2(_03949_ ), .ZN(_03950_ ) );
AND2_X1 _11691_ ( .A1(\ID_EX_pc [15] ), .A2(\ID_EX_imm [15] ), .ZN(_03951_ ) );
AND2_X1 _11692_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_03952_ ) );
AND2_X1 _11693_ ( .A1(_03940_ ), .A2(_03952_ ), .ZN(_03953_ ) );
NOR3_X1 _11694_ ( .A1(_03950_ ), .A2(_03951_ ), .A3(_03953_ ), .ZN(_03954_ ) );
NAND2_X1 _11695_ ( .A1(_03945_ ), .A2(_03954_ ), .ZN(_03955_ ) );
XOR2_X1 _11696_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_03956_ ) );
XOR2_X1 _11697_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_03957_ ) );
AND4_X1 _11698_ ( .A1(_03897_ ), .A2(_03955_ ), .A3(_03956_ ), .A4(_03957_ ), .ZN(_03958_ ) );
AND2_X1 _11699_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_03959_ ) );
AND2_X1 _11700_ ( .A1(_03895_ ), .A2(_03959_ ), .ZN(_03960_ ) );
AOI21_X1 _11701_ ( .A(_03960_ ), .B1(\ID_EX_pc [19] ), .B2(\ID_EX_imm [19] ), .ZN(_03961_ ) );
AND2_X1 _11702_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_imm [17] ), .ZN(_03962_ ) );
AND2_X1 _11703_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_03963_ ) );
AOI21_X1 _11704_ ( .A(_03962_ ), .B1(_03957_ ), .B2(_03963_ ), .ZN(_03964_ ) );
INV_X1 _11705_ ( .A(_03897_ ), .ZN(_03965_ ) );
OAI21_X1 _11706_ ( .A(_03961_ ), .B1(_03964_ ), .B2(_03965_ ), .ZN(_03966_ ) );
OR2_X1 _11707_ ( .A1(_03958_ ), .A2(_03966_ ), .ZN(_03967_ ) );
XOR2_X1 _11708_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_03968_ ) );
XOR2_X1 _11709_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_03969_ ) );
AND2_X1 _11710_ ( .A1(_03968_ ), .A2(_03969_ ), .ZN(_03970_ ) );
XOR2_X1 _11711_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_03971_ ) );
XOR2_X1 _11712_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_03972_ ) );
AND2_X1 _11713_ ( .A1(_03971_ ), .A2(_03972_ ), .ZN(_03973_ ) );
AND3_X1 _11714_ ( .A1(_03967_ ), .A2(_03970_ ), .A3(_03973_ ), .ZN(_03974_ ) );
AND2_X1 _11715_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_03975_ ) );
AND2_X1 _11716_ ( .A1(_03968_ ), .A2(_03975_ ), .ZN(_03976_ ) );
AOI21_X1 _11717_ ( .A(_03976_ ), .B1(\ID_EX_pc [23] ), .B2(\ID_EX_imm [23] ), .ZN(_03977_ ) );
AND3_X1 _11718_ ( .A1(_03971_ ), .A2(\ID_EX_pc [20] ), .A3(\ID_EX_imm [20] ), .ZN(_03978_ ) );
AOI21_X1 _11719_ ( .A(_03978_ ), .B1(\ID_EX_pc [21] ), .B2(\ID_EX_imm [21] ), .ZN(_03979_ ) );
INV_X1 _11720_ ( .A(_03970_ ), .ZN(_03980_ ) );
OAI21_X1 _11721_ ( .A(_03977_ ), .B1(_03979_ ), .B2(_03980_ ), .ZN(_03981_ ) );
OAI211_X1 _11722_ ( .A(_03893_ ), .B(_03894_ ), .C1(_03974_ ), .C2(_03981_ ), .ZN(_03982_ ) );
AND2_X1 _11723_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_03983_ ) );
AND2_X1 _11724_ ( .A1(_03893_ ), .A2(_03983_ ), .ZN(_03984_ ) );
AOI21_X1 _11725_ ( .A(_03984_ ), .B1(\ID_EX_pc [25] ), .B2(\ID_EX_imm [25] ), .ZN(_03985_ ) );
NAND2_X1 _11726_ ( .A1(_03982_ ), .A2(_03985_ ), .ZN(_03986_ ) );
XOR2_X1 _11727_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_03987_ ) );
XOR2_X1 _11728_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_03988_ ) );
NAND3_X1 _11729_ ( .A1(_03986_ ), .A2(_03987_ ), .A3(_03988_ ), .ZN(_03989_ ) );
AND3_X1 _11730_ ( .A1(_03987_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_03990_ ) );
AOI21_X1 _11731_ ( .A(_03990_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_03991_ ) );
NAND2_X1 _11732_ ( .A1(_03989_ ), .A2(_03991_ ), .ZN(_03992_ ) );
XOR2_X1 _11733_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_03993_ ) );
NAND2_X1 _11734_ ( .A1(_03992_ ), .A2(_03993_ ), .ZN(_03994_ ) );
NAND2_X1 _11735_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_03995_ ) );
AOI21_X1 _11736_ ( .A(_03892_ ), .B1(_03994_ ), .B2(_03995_ ), .ZN(_03996_ ) );
AND2_X1 _11737_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_03997_ ) );
OR2_X1 _11738_ ( .A1(_03996_ ), .A2(_03997_ ), .ZN(_03998_ ) );
XOR2_X1 _11739_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_03999_ ) );
XOR2_X1 _11740_ ( .A(_03998_ ), .B(_03999_ ), .Z(_04000_ ) );
NOR2_X1 _11741_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_5 ), .ZN(_04001_ ) );
AND2_X1 _11742_ ( .A1(_04001_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04002_ ) );
AND2_X1 _11743_ ( .A1(_02029_ ), .A2(_02020_ ), .ZN(_04003_ ) );
AOI22_X4 _11744_ ( .A1(_02020_ ), .A2(\ID_EX_rs2 [4] ), .B1(_03250_ ), .B2(\EX_LS_dest_reg [0] ), .ZN(_04004_ ) );
INV_X2 _11745_ ( .A(\EX_LS_dest_reg [2] ), .ZN(_04005_ ) );
NAND2_X1 _11746_ ( .A1(_04005_ ), .A2(\ID_EX_rs2 [2] ), .ZN(_04006_ ) );
OAI211_X1 _11747_ ( .A(_04004_ ), .B(_04006_ ), .C1(_02020_ ), .C2(\ID_EX_rs2 [4] ), .ZN(_04007_ ) );
XOR2_X2 _11748_ ( .A(\EX_LS_dest_reg [3] ), .B(\ID_EX_rs2 [3] ), .Z(_04008_ ) );
NOR2_X1 _11749_ ( .A1(_04005_ ), .A2(\ID_EX_rs2 [2] ), .ZN(_04009_ ) );
OR4_X2 _11750_ ( .A1(_02026_ ), .A2(_04007_ ), .A3(_04008_ ), .A4(_04009_ ), .ZN(_04010_ ) );
NOR2_X1 _11751_ ( .A1(_02031_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_04011_ ) );
OAI22_X1 _11752_ ( .A1(\EX_LS_dest_reg [1] ), .A2(_03247_ ), .B1(_03250_ ), .B2(\EX_LS_dest_reg [0] ), .ZN(_04012_ ) );
OR4_X4 _11753_ ( .A1(_04003_ ), .A2(_04010_ ), .A3(_04011_ ), .A4(_04012_ ), .ZN(_04013_ ) );
BUF_X8 _11754_ ( .A(_04013_ ), .Z(_04014_ ) );
INV_X1 _11755_ ( .A(\EX_LS_result_reg [23] ), .ZN(_04015_ ) );
OR3_X1 _11756_ ( .A1(_04014_ ), .A2(_04015_ ), .A3(_02327_ ), .ZN(_04016_ ) );
INV_X1 _11757_ ( .A(fanout_net_41 ), .ZN(_04017_ ) );
BUF_X4 _11758_ ( .A(_04017_ ), .Z(_04018_ ) );
OR2_X1 _11759_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][23] ), .ZN(_04019_ ) );
INV_X1 _11760_ ( .A(fanout_net_38 ), .ZN(_04020_ ) );
BUF_X4 _11761_ ( .A(_04020_ ), .Z(_04021_ ) );
BUF_X4 _11762_ ( .A(_04021_ ), .Z(_04022_ ) );
INV_X1 _11763_ ( .A(fanout_net_29 ), .ZN(_04023_ ) );
BUF_X2 _11764_ ( .A(_04023_ ), .Z(_04024_ ) );
BUF_X4 _11765_ ( .A(_04024_ ), .Z(_04025_ ) );
OAI211_X1 _11766_ ( .A(_04019_ ), .B(_04022_ ), .C1(_04025_ ), .C2(\myreg.Reg[1][23] ), .ZN(_04026_ ) );
OR2_X1 _11767_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[2][23] ), .ZN(_04027_ ) );
OAI211_X1 _11768_ ( .A(_04027_ ), .B(fanout_net_38 ), .C1(_04025_ ), .C2(\myreg.Reg[3][23] ), .ZN(_04028_ ) );
INV_X2 _11769_ ( .A(fanout_net_40 ), .ZN(_04029_ ) );
BUF_X4 _11770_ ( .A(_04029_ ), .Z(_04030_ ) );
NAND3_X1 _11771_ ( .A1(_04026_ ), .A2(_04028_ ), .A3(_04030_ ), .ZN(_04031_ ) );
MUX2_X1 _11772_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_29 ), .Z(_04032_ ) );
MUX2_X1 _11773_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_29 ), .Z(_04033_ ) );
MUX2_X1 _11774_ ( .A(_04032_ ), .B(_04033_ ), .S(_04022_ ), .Z(_04034_ ) );
BUF_X4 _11775_ ( .A(_04029_ ), .Z(_04035_ ) );
OAI211_X1 _11776_ ( .A(_04018_ ), .B(_04031_ ), .C1(_04034_ ), .C2(_04035_ ), .ZN(_04036_ ) );
OR2_X1 _11777_ ( .A1(_04024_ ), .A2(\myreg.Reg[15][23] ), .ZN(_04037_ ) );
OAI211_X1 _11778_ ( .A(_04037_ ), .B(fanout_net_38 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[14][23] ), .ZN(_04038_ ) );
OR2_X1 _11779_ ( .A1(_04024_ ), .A2(\myreg.Reg[13][23] ), .ZN(_04039_ ) );
OAI211_X1 _11780_ ( .A(_04039_ ), .B(_04022_ ), .C1(fanout_net_29 ), .C2(\myreg.Reg[12][23] ), .ZN(_04040_ ) );
NAND3_X1 _11781_ ( .A1(_04038_ ), .A2(_04040_ ), .A3(fanout_net_40 ), .ZN(_04041_ ) );
MUX2_X1 _11782_ ( .A(\myreg.Reg[8][23] ), .B(\myreg.Reg[9][23] ), .S(fanout_net_29 ), .Z(_04042_ ) );
MUX2_X1 _11783_ ( .A(\myreg.Reg[10][23] ), .B(\myreg.Reg[11][23] ), .S(fanout_net_29 ), .Z(_04043_ ) );
MUX2_X1 _11784_ ( .A(_04042_ ), .B(_04043_ ), .S(fanout_net_38 ), .Z(_04044_ ) );
OAI211_X1 _11785_ ( .A(fanout_net_41 ), .B(_04041_ ), .C1(_04044_ ), .C2(fanout_net_40 ), .ZN(_04045_ ) );
NAND2_X1 _11786_ ( .A1(_04036_ ), .A2(_04045_ ), .ZN(_04046_ ) );
BUF_X8 _11787_ ( .A(_04013_ ), .Z(_04047_ ) );
BUF_X16 _11788_ ( .A(_04047_ ), .Z(_04048_ ) );
OAI21_X4 _11789_ ( .A(_04046_ ), .B1(_04048_ ), .B2(_02127_ ), .ZN(_04049_ ) );
AND2_X2 _11790_ ( .A1(_04016_ ), .A2(_04049_ ), .ZN(_04050_ ) );
INV_X1 _11791_ ( .A(_02179_ ), .ZN(_04051_ ) );
XNOR2_X1 _11792_ ( .A(_04050_ ), .B(_04051_ ), .ZN(_04052_ ) );
BUF_X8 _11793_ ( .A(_04014_ ), .Z(_04053_ ) );
OR3_X4 _11794_ ( .A1(_04053_ ), .A2(\EX_LS_result_reg [22] ), .A3(_02094_ ), .ZN(_04054_ ) );
OR2_X1 _11795_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][22] ), .ZN(_04055_ ) );
BUF_X4 _11796_ ( .A(_04020_ ), .Z(_04056_ ) );
BUF_X4 _11797_ ( .A(_04056_ ), .Z(_04057_ ) );
BUF_X4 _11798_ ( .A(_04057_ ), .Z(_04058_ ) );
BUF_X2 _11799_ ( .A(_04023_ ), .Z(_04059_ ) );
CLKBUF_X2 _11800_ ( .A(_04059_ ), .Z(_04060_ ) );
BUF_X2 _11801_ ( .A(_04060_ ), .Z(_04061_ ) );
BUF_X2 _11802_ ( .A(_04061_ ), .Z(_04062_ ) );
OAI211_X1 _11803_ ( .A(_04055_ ), .B(_04058_ ), .C1(_04062_ ), .C2(\myreg.Reg[9][22] ), .ZN(_04063_ ) );
OR2_X1 _11804_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[10][22] ), .ZN(_04064_ ) );
OAI211_X1 _11805_ ( .A(_04064_ ), .B(fanout_net_38 ), .C1(_04062_ ), .C2(\myreg.Reg[11][22] ), .ZN(_04065_ ) );
BUF_X4 _11806_ ( .A(_04030_ ), .Z(_04066_ ) );
BUF_X4 _11807_ ( .A(_04066_ ), .Z(_04067_ ) );
NAND3_X1 _11808_ ( .A1(_04063_ ), .A2(_04065_ ), .A3(_04067_ ), .ZN(_04068_ ) );
MUX2_X1 _11809_ ( .A(\myreg.Reg[14][22] ), .B(\myreg.Reg[15][22] ), .S(fanout_net_29 ), .Z(_04069_ ) );
MUX2_X1 _11810_ ( .A(\myreg.Reg[12][22] ), .B(\myreg.Reg[13][22] ), .S(fanout_net_29 ), .Z(_04070_ ) );
BUF_X4 _11811_ ( .A(_04057_ ), .Z(_04071_ ) );
MUX2_X1 _11812_ ( .A(_04069_ ), .B(_04070_ ), .S(_04071_ ), .Z(_04072_ ) );
OAI211_X1 _11813_ ( .A(fanout_net_41 ), .B(_04068_ ), .C1(_04072_ ), .C2(_04067_ ), .ZN(_04073_ ) );
BUF_X4 _11814_ ( .A(_04018_ ), .Z(_04074_ ) );
BUF_X4 _11815_ ( .A(_04035_ ), .Z(_04075_ ) );
NOR2_X1 _11816_ ( .A1(_04062_ ), .A2(\myreg.Reg[3][22] ), .ZN(_04076_ ) );
OAI21_X1 _11817_ ( .A(fanout_net_38 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[2][22] ), .ZN(_04077_ ) );
NOR2_X1 _11818_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][22] ), .ZN(_04078_ ) );
OAI21_X1 _11819_ ( .A(_04071_ ), .B1(_04062_ ), .B2(\myreg.Reg[1][22] ), .ZN(_04079_ ) );
OAI221_X1 _11820_ ( .A(_04075_ ), .B1(_04076_ ), .B2(_04077_ ), .C1(_04078_ ), .C2(_04079_ ), .ZN(_04080_ ) );
MUX2_X1 _11821_ ( .A(\myreg.Reg[6][22] ), .B(\myreg.Reg[7][22] ), .S(fanout_net_29 ), .Z(_04081_ ) );
MUX2_X1 _11822_ ( .A(\myreg.Reg[4][22] ), .B(\myreg.Reg[5][22] ), .S(fanout_net_29 ), .Z(_04082_ ) );
MUX2_X1 _11823_ ( .A(_04081_ ), .B(_04082_ ), .S(_04071_ ), .Z(_04083_ ) );
OAI211_X1 _11824_ ( .A(_04074_ ), .B(_04080_ ), .C1(_04083_ ), .C2(_04067_ ), .ZN(_04084_ ) );
BUF_X8 _11825_ ( .A(_04048_ ), .Z(_04085_ ) );
OAI211_X1 _11826_ ( .A(_04073_ ), .B(_04084_ ), .C1(_04085_ ), .C2(_02128_ ), .ZN(_04086_ ) );
NAND2_X1 _11827_ ( .A1(_04054_ ), .A2(_04086_ ), .ZN(_04087_ ) );
INV_X1 _11828_ ( .A(_02155_ ), .ZN(_04088_ ) );
XNOR2_X1 _11829_ ( .A(_04087_ ), .B(_04088_ ), .ZN(_04089_ ) );
AND2_X1 _11830_ ( .A1(_04052_ ), .A2(_04089_ ), .ZN(_04090_ ) );
OR3_X4 _11831_ ( .A1(_04053_ ), .A2(\EX_LS_result_reg [21] ), .A3(_02044_ ), .ZN(_04091_ ) );
OR2_X1 _11832_ ( .A1(_04061_ ), .A2(\myreg.Reg[5][21] ), .ZN(_04092_ ) );
OAI211_X1 _11833_ ( .A(_04092_ ), .B(_04071_ ), .C1(fanout_net_29 ), .C2(\myreg.Reg[4][21] ), .ZN(_04093_ ) );
OR2_X1 _11834_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[6][21] ), .ZN(_04094_ ) );
OAI211_X1 _11835_ ( .A(_04094_ ), .B(fanout_net_38 ), .C1(_04062_ ), .C2(\myreg.Reg[7][21] ), .ZN(_04095_ ) );
NAND3_X1 _11836_ ( .A1(_04093_ ), .A2(fanout_net_40 ), .A3(_04095_ ), .ZN(_04096_ ) );
MUX2_X1 _11837_ ( .A(\myreg.Reg[2][21] ), .B(\myreg.Reg[3][21] ), .S(fanout_net_29 ), .Z(_04097_ ) );
MUX2_X1 _11838_ ( .A(\myreg.Reg[0][21] ), .B(\myreg.Reg[1][21] ), .S(fanout_net_29 ), .Z(_04098_ ) );
MUX2_X1 _11839_ ( .A(_04097_ ), .B(_04098_ ), .S(_04071_ ), .Z(_04099_ ) );
OAI211_X1 _11840_ ( .A(_04074_ ), .B(_04096_ ), .C1(_04099_ ), .C2(fanout_net_40 ), .ZN(_04100_ ) );
BUF_X4 _11841_ ( .A(_04025_ ), .Z(_04101_ ) );
NOR2_X1 _11842_ ( .A1(_04101_ ), .A2(\myreg.Reg[11][21] ), .ZN(_04102_ ) );
OAI21_X1 _11843_ ( .A(fanout_net_38 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[10][21] ), .ZN(_04103_ ) );
NOR2_X1 _11844_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][21] ), .ZN(_04104_ ) );
OAI21_X1 _11845_ ( .A(_04071_ ), .B1(_04062_ ), .B2(\myreg.Reg[9][21] ), .ZN(_04105_ ) );
OAI221_X1 _11846_ ( .A(_04075_ ), .B1(_04102_ ), .B2(_04103_ ), .C1(_04104_ ), .C2(_04105_ ), .ZN(_04106_ ) );
MUX2_X1 _11847_ ( .A(\myreg.Reg[12][21] ), .B(\myreg.Reg[13][21] ), .S(fanout_net_29 ), .Z(_04107_ ) );
MUX2_X1 _11848_ ( .A(\myreg.Reg[14][21] ), .B(\myreg.Reg[15][21] ), .S(fanout_net_29 ), .Z(_04108_ ) );
MUX2_X1 _11849_ ( .A(_04107_ ), .B(_04108_ ), .S(fanout_net_38 ), .Z(_04109_ ) );
OAI211_X1 _11850_ ( .A(fanout_net_41 ), .B(_04106_ ), .C1(_04109_ ), .C2(_04067_ ), .ZN(_04110_ ) );
OAI211_X1 _11851_ ( .A(_04100_ ), .B(_04110_ ), .C1(_04085_ ), .C2(_02128_ ), .ZN(_04111_ ) );
NAND2_X1 _11852_ ( .A1(_04091_ ), .A2(_04111_ ), .ZN(_04112_ ) );
NAND2_X1 _11853_ ( .A1(_02205_ ), .A2(_02227_ ), .ZN(_04113_ ) );
INV_X1 _11854_ ( .A(_04113_ ), .ZN(_04114_ ) );
XNOR2_X1 _11855_ ( .A(_04112_ ), .B(_04114_ ), .ZN(_04115_ ) );
OR3_X4 _11856_ ( .A1(_04085_ ), .A2(\EX_LS_result_reg [20] ), .A3(_02045_ ), .ZN(_04116_ ) );
BUF_X4 _11857_ ( .A(_04074_ ), .Z(_04117_ ) );
OR2_X1 _11858_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[4][20] ), .ZN(_04118_ ) );
BUF_X4 _11859_ ( .A(_04101_ ), .Z(_04119_ ) );
OAI211_X1 _11860_ ( .A(_04118_ ), .B(_04058_ ), .C1(_04119_ ), .C2(\myreg.Reg[5][20] ), .ZN(_04120_ ) );
OR2_X1 _11861_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[6][20] ), .ZN(_04121_ ) );
OAI211_X1 _11862_ ( .A(_04121_ ), .B(fanout_net_38 ), .C1(_04119_ ), .C2(\myreg.Reg[7][20] ), .ZN(_04122_ ) );
NAND3_X1 _11863_ ( .A1(_04120_ ), .A2(_04122_ ), .A3(fanout_net_40 ), .ZN(_04123_ ) );
MUX2_X1 _11864_ ( .A(\myreg.Reg[2][20] ), .B(\myreg.Reg[3][20] ), .S(fanout_net_29 ), .Z(_04124_ ) );
MUX2_X1 _11865_ ( .A(\myreg.Reg[0][20] ), .B(\myreg.Reg[1][20] ), .S(fanout_net_29 ), .Z(_04125_ ) );
MUX2_X1 _11866_ ( .A(_04124_ ), .B(_04125_ ), .S(_04058_ ), .Z(_04126_ ) );
OAI211_X1 _11867_ ( .A(_04117_ ), .B(_04123_ ), .C1(_04126_ ), .C2(fanout_net_40 ), .ZN(_04127_ ) );
NOR2_X1 _11868_ ( .A1(_04119_ ), .A2(\myreg.Reg[11][20] ), .ZN(_04128_ ) );
OAI21_X1 _11869_ ( .A(fanout_net_38 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[10][20] ), .ZN(_04129_ ) );
NOR2_X1 _11870_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][20] ), .ZN(_04130_ ) );
OAI21_X1 _11871_ ( .A(_04058_ ), .B1(_04119_ ), .B2(\myreg.Reg[9][20] ), .ZN(_04131_ ) );
OAI221_X1 _11872_ ( .A(_04067_ ), .B1(_04128_ ), .B2(_04129_ ), .C1(_04130_ ), .C2(_04131_ ), .ZN(_04132_ ) );
MUX2_X1 _11873_ ( .A(\myreg.Reg[12][20] ), .B(\myreg.Reg[13][20] ), .S(fanout_net_30 ), .Z(_04133_ ) );
MUX2_X1 _11874_ ( .A(\myreg.Reg[14][20] ), .B(\myreg.Reg[15][20] ), .S(fanout_net_30 ), .Z(_04134_ ) );
MUX2_X1 _11875_ ( .A(_04133_ ), .B(_04134_ ), .S(fanout_net_38 ), .Z(_04135_ ) );
BUF_X4 _11876_ ( .A(_04067_ ), .Z(_04136_ ) );
OAI211_X1 _11877_ ( .A(fanout_net_41 ), .B(_04132_ ), .C1(_04135_ ), .C2(_04136_ ), .ZN(_04137_ ) );
OAI211_X1 _11878_ ( .A(_04127_ ), .B(_04137_ ), .C1(_04085_ ), .C2(_02095_ ), .ZN(_04138_ ) );
NAND2_X1 _11879_ ( .A1(_04116_ ), .A2(_04138_ ), .ZN(_04139_ ) );
INV_X1 _11880_ ( .A(_02202_ ), .ZN(_04140_ ) );
XNOR2_X1 _11881_ ( .A(_04139_ ), .B(_04140_ ), .ZN(_04141_ ) );
AND3_X1 _11882_ ( .A1(_04090_ ), .A2(_04115_ ), .A3(_04141_ ), .ZN(_04142_ ) );
OR3_X4 _11883_ ( .A1(_04053_ ), .A2(\EX_LS_result_reg [19] ), .A3(_02044_ ), .ZN(_04143_ ) );
CLKBUF_X2 _11884_ ( .A(_04024_ ), .Z(_04144_ ) );
OR2_X1 _11885_ ( .A1(_04144_ ), .A2(\myreg.Reg[5][19] ), .ZN(_04145_ ) );
BUF_X4 _11886_ ( .A(_04021_ ), .Z(_04146_ ) );
BUF_X4 _11887_ ( .A(_04146_ ), .Z(_04147_ ) );
OAI211_X1 _11888_ ( .A(_04145_ ), .B(_04147_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[4][19] ), .ZN(_04148_ ) );
OR2_X1 _11889_ ( .A1(_04144_ ), .A2(\myreg.Reg[7][19] ), .ZN(_04149_ ) );
OAI211_X1 _11890_ ( .A(_04149_ ), .B(fanout_net_38 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[6][19] ), .ZN(_04150_ ) );
NAND3_X1 _11891_ ( .A1(_04148_ ), .A2(_04150_ ), .A3(fanout_net_40 ), .ZN(_04151_ ) );
MUX2_X1 _11892_ ( .A(\myreg.Reg[2][19] ), .B(\myreg.Reg[3][19] ), .S(fanout_net_30 ), .Z(_04152_ ) );
MUX2_X1 _11893_ ( .A(\myreg.Reg[0][19] ), .B(\myreg.Reg[1][19] ), .S(fanout_net_30 ), .Z(_04153_ ) );
MUX2_X1 _11894_ ( .A(_04152_ ), .B(_04153_ ), .S(_04147_ ), .Z(_04154_ ) );
OAI211_X1 _11895_ ( .A(_04074_ ), .B(_04151_ ), .C1(_04154_ ), .C2(fanout_net_40 ), .ZN(_04155_ ) );
NOR2_X1 _11896_ ( .A1(_04101_ ), .A2(\myreg.Reg[11][19] ), .ZN(_04156_ ) );
OAI21_X1 _11897_ ( .A(fanout_net_38 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][19] ), .ZN(_04157_ ) );
NOR2_X1 _11898_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][19] ), .ZN(_04158_ ) );
OAI21_X1 _11899_ ( .A(_04147_ ), .B1(_04101_ ), .B2(\myreg.Reg[9][19] ), .ZN(_04159_ ) );
OAI221_X1 _11900_ ( .A(_04066_ ), .B1(_04156_ ), .B2(_04157_ ), .C1(_04158_ ), .C2(_04159_ ), .ZN(_04160_ ) );
MUX2_X1 _11901_ ( .A(\myreg.Reg[12][19] ), .B(\myreg.Reg[13][19] ), .S(fanout_net_30 ), .Z(_04161_ ) );
MUX2_X1 _11902_ ( .A(\myreg.Reg[14][19] ), .B(\myreg.Reg[15][19] ), .S(fanout_net_30 ), .Z(_04162_ ) );
MUX2_X1 _11903_ ( .A(_04161_ ), .B(_04162_ ), .S(fanout_net_38 ), .Z(_04163_ ) );
OAI211_X1 _11904_ ( .A(fanout_net_41 ), .B(_04160_ ), .C1(_04163_ ), .C2(_04075_ ), .ZN(_04164_ ) );
OAI211_X1 _11905_ ( .A(_04155_ ), .B(_04164_ ), .C1(_04053_ ), .C2(_02094_ ), .ZN(_04165_ ) );
NAND2_X1 _11906_ ( .A1(_04143_ ), .A2(_04165_ ), .ZN(_04166_ ) );
INV_X1 _11907_ ( .A(_02252_ ), .ZN(_04167_ ) );
XNOR2_X2 _11908_ ( .A(_04166_ ), .B(_04167_ ), .ZN(_04168_ ) );
OR3_X4 _11909_ ( .A1(_04053_ ), .A2(\EX_LS_result_reg [18] ), .A3(_02094_ ), .ZN(_04169_ ) );
OR2_X1 _11910_ ( .A1(_04061_ ), .A2(\myreg.Reg[11][18] ), .ZN(_04170_ ) );
OAI211_X1 _11911_ ( .A(_04170_ ), .B(fanout_net_38 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[10][18] ), .ZN(_04171_ ) );
OR2_X1 _11912_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][18] ), .ZN(_04172_ ) );
OAI211_X1 _11913_ ( .A(_04172_ ), .B(_04058_ ), .C1(_04062_ ), .C2(\myreg.Reg[9][18] ), .ZN(_04173_ ) );
NAND3_X1 _11914_ ( .A1(_04171_ ), .A2(_04067_ ), .A3(_04173_ ), .ZN(_04174_ ) );
MUX2_X1 _11915_ ( .A(\myreg.Reg[14][18] ), .B(\myreg.Reg[15][18] ), .S(fanout_net_30 ), .Z(_04175_ ) );
MUX2_X1 _11916_ ( .A(\myreg.Reg[12][18] ), .B(\myreg.Reg[13][18] ), .S(fanout_net_30 ), .Z(_04176_ ) );
MUX2_X1 _11917_ ( .A(_04175_ ), .B(_04176_ ), .S(_04071_ ), .Z(_04177_ ) );
OAI211_X1 _11918_ ( .A(fanout_net_41 ), .B(_04174_ ), .C1(_04177_ ), .C2(_04067_ ), .ZN(_04178_ ) );
OR2_X1 _11919_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[0][18] ), .ZN(_04179_ ) );
OAI211_X1 _11920_ ( .A(_04179_ ), .B(_04071_ ), .C1(_04062_ ), .C2(\myreg.Reg[1][18] ), .ZN(_04180_ ) );
NOR2_X1 _11921_ ( .A1(_04062_ ), .A2(\myreg.Reg[3][18] ), .ZN(_04181_ ) );
OAI21_X1 _11922_ ( .A(fanout_net_38 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[2][18] ), .ZN(_04182_ ) );
OAI211_X1 _11923_ ( .A(_04180_ ), .B(_04075_ ), .C1(_04181_ ), .C2(_04182_ ), .ZN(_04183_ ) );
MUX2_X1 _11924_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_30 ), .Z(_04184_ ) );
MUX2_X1 _11925_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_30 ), .Z(_04185_ ) );
MUX2_X1 _11926_ ( .A(_04184_ ), .B(_04185_ ), .S(_04071_ ), .Z(_04186_ ) );
OAI211_X1 _11927_ ( .A(_04074_ ), .B(_04183_ ), .C1(_04186_ ), .C2(_04067_ ), .ZN(_04187_ ) );
OAI211_X1 _11928_ ( .A(_04178_ ), .B(_04187_ ), .C1(_04085_ ), .C2(_02128_ ), .ZN(_04188_ ) );
NAND2_X1 _11929_ ( .A1(_04169_ ), .A2(_04188_ ), .ZN(_04189_ ) );
INV_X1 _11930_ ( .A(_02275_ ), .ZN(_04190_ ) );
XNOR2_X1 _11931_ ( .A(_04189_ ), .B(_04190_ ), .ZN(_04191_ ) );
AND2_X1 _11932_ ( .A1(_04168_ ), .A2(_04191_ ), .ZN(_04192_ ) );
OR3_X1 _11933_ ( .A1(_04085_ ), .A2(\EX_LS_result_reg [16] ), .A3(_02095_ ), .ZN(_04193_ ) );
OR2_X1 _11934_ ( .A1(_04119_ ), .A2(\myreg.Reg[3][16] ), .ZN(_04194_ ) );
OAI211_X1 _11935_ ( .A(_04194_ ), .B(fanout_net_38 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[2][16] ), .ZN(_04195_ ) );
OR2_X1 _11936_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[0][16] ), .ZN(_04196_ ) );
BUF_X4 _11937_ ( .A(_04058_ ), .Z(_04197_ ) );
BUF_X4 _11938_ ( .A(_04119_ ), .Z(_04198_ ) );
OAI211_X1 _11939_ ( .A(_04196_ ), .B(_04197_ ), .C1(_04198_ ), .C2(\myreg.Reg[1][16] ), .ZN(_04199_ ) );
NAND3_X1 _11940_ ( .A1(_04195_ ), .A2(_04136_ ), .A3(_04199_ ), .ZN(_04200_ ) );
MUX2_X1 _11941_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_30 ), .Z(_04201_ ) );
MUX2_X1 _11942_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_30 ), .Z(_04202_ ) );
MUX2_X1 _11943_ ( .A(_04201_ ), .B(_04202_ ), .S(_04058_ ), .Z(_04203_ ) );
BUF_X4 _11944_ ( .A(_04136_ ), .Z(_04204_ ) );
OAI211_X1 _11945_ ( .A(_04117_ ), .B(_04200_ ), .C1(_04203_ ), .C2(_04204_ ), .ZN(_04205_ ) );
OR2_X1 _11946_ ( .A1(_04062_ ), .A2(\myreg.Reg[13][16] ), .ZN(_04206_ ) );
OAI211_X1 _11947_ ( .A(_04206_ ), .B(_04197_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[12][16] ), .ZN(_04207_ ) );
OR2_X1 _11948_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[14][16] ), .ZN(_04208_ ) );
OAI211_X1 _11949_ ( .A(_04208_ ), .B(fanout_net_38 ), .C1(_04119_ ), .C2(\myreg.Reg[15][16] ), .ZN(_04209_ ) );
NAND3_X1 _11950_ ( .A1(_04207_ ), .A2(fanout_net_40 ), .A3(_04209_ ), .ZN(_04210_ ) );
MUX2_X1 _11951_ ( .A(\myreg.Reg[8][16] ), .B(\myreg.Reg[9][16] ), .S(fanout_net_30 ), .Z(_04211_ ) );
MUX2_X1 _11952_ ( .A(\myreg.Reg[10][16] ), .B(\myreg.Reg[11][16] ), .S(fanout_net_30 ), .Z(_04212_ ) );
MUX2_X1 _11953_ ( .A(_04211_ ), .B(_04212_ ), .S(fanout_net_38 ), .Z(_04213_ ) );
OAI211_X1 _11954_ ( .A(fanout_net_41 ), .B(_04210_ ), .C1(_04213_ ), .C2(fanout_net_40 ), .ZN(_04214_ ) );
BUF_X2 _11955_ ( .A(_04085_ ), .Z(_04215_ ) );
OAI211_X4 _11956_ ( .A(_04205_ ), .B(_04214_ ), .C1(_04215_ ), .C2(_02088_ ), .ZN(_04216_ ) );
NAND2_X1 _11957_ ( .A1(_04193_ ), .A2(_04216_ ), .ZN(_04217_ ) );
INV_X1 _11958_ ( .A(_02322_ ), .ZN(_04218_ ) );
XNOR2_X1 _11959_ ( .A(_04217_ ), .B(_04218_ ), .ZN(_04219_ ) );
OR3_X2 _11960_ ( .A1(_04053_ ), .A2(\EX_LS_result_reg [17] ), .A3(_02127_ ), .ZN(_04220_ ) );
OR2_X1 _11961_ ( .A1(_04144_ ), .A2(\myreg.Reg[7][17] ), .ZN(_04221_ ) );
OAI211_X1 _11962_ ( .A(_04221_ ), .B(fanout_net_38 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[6][17] ), .ZN(_04222_ ) );
OR2_X1 _11963_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[4][17] ), .ZN(_04223_ ) );
OAI211_X1 _11964_ ( .A(_04223_ ), .B(_04147_ ), .C1(_04101_ ), .C2(\myreg.Reg[5][17] ), .ZN(_04224_ ) );
NAND3_X1 _11965_ ( .A1(_04222_ ), .A2(fanout_net_40 ), .A3(_04224_ ), .ZN(_04225_ ) );
MUX2_X1 _11966_ ( .A(\myreg.Reg[2][17] ), .B(\myreg.Reg[3][17] ), .S(fanout_net_30 ), .Z(_04226_ ) );
MUX2_X1 _11967_ ( .A(\myreg.Reg[0][17] ), .B(\myreg.Reg[1][17] ), .S(fanout_net_31 ), .Z(_04227_ ) );
MUX2_X1 _11968_ ( .A(_04226_ ), .B(_04227_ ), .S(_04147_ ), .Z(_04228_ ) );
OAI211_X1 _11969_ ( .A(_04074_ ), .B(_04225_ ), .C1(_04228_ ), .C2(fanout_net_40 ), .ZN(_04229_ ) );
NOR2_X1 _11970_ ( .A1(_04061_ ), .A2(\myreg.Reg[11][17] ), .ZN(_04230_ ) );
OAI21_X1 _11971_ ( .A(fanout_net_38 ), .B1(fanout_net_31 ), .B2(\myreg.Reg[10][17] ), .ZN(_04231_ ) );
NOR2_X1 _11972_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][17] ), .ZN(_04232_ ) );
OAI21_X1 _11973_ ( .A(_04057_ ), .B1(_04101_ ), .B2(\myreg.Reg[9][17] ), .ZN(_04233_ ) );
OAI221_X1 _11974_ ( .A(_04066_ ), .B1(_04230_ ), .B2(_04231_ ), .C1(_04232_ ), .C2(_04233_ ), .ZN(_04234_ ) );
MUX2_X1 _11975_ ( .A(\myreg.Reg[12][17] ), .B(\myreg.Reg[13][17] ), .S(fanout_net_31 ), .Z(_04235_ ) );
MUX2_X1 _11976_ ( .A(\myreg.Reg[14][17] ), .B(\myreg.Reg[15][17] ), .S(fanout_net_31 ), .Z(_04236_ ) );
MUX2_X1 _11977_ ( .A(_04235_ ), .B(_04236_ ), .S(fanout_net_38 ), .Z(_04237_ ) );
OAI211_X1 _11978_ ( .A(fanout_net_41 ), .B(_04234_ ), .C1(_04237_ ), .C2(_04075_ ), .ZN(_04238_ ) );
OAI211_X1 _11979_ ( .A(_04229_ ), .B(_04238_ ), .C1(_04053_ ), .C2(_02044_ ), .ZN(_04239_ ) );
NAND2_X1 _11980_ ( .A1(_04220_ ), .A2(_04239_ ), .ZN(_04240_ ) );
INV_X1 _11981_ ( .A(_02299_ ), .ZN(_04241_ ) );
XNOR2_X1 _11982_ ( .A(_04240_ ), .B(_04241_ ), .ZN(_04242_ ) );
AND3_X1 _11983_ ( .A1(_04192_ ), .A2(_04219_ ), .A3(_04242_ ), .ZN(_04243_ ) );
AND2_X1 _11984_ ( .A1(_04142_ ), .A2(_04243_ ), .ZN(_04244_ ) );
OR3_X1 _11985_ ( .A1(_04085_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02095_ ), .ZN(_04245_ ) );
NAND2_X1 _11986_ ( .A1(_02097_ ), .A2(fanout_net_31 ), .ZN(_04246_ ) );
BUF_X4 _11987_ ( .A(_04058_ ), .Z(_04247_ ) );
OAI211_X1 _11988_ ( .A(_04246_ ), .B(_04247_ ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04248_ ) );
NAND2_X1 _11989_ ( .A1(_02102_ ), .A2(fanout_net_31 ), .ZN(_04249_ ) );
OAI211_X1 _11990_ ( .A(_04249_ ), .B(fanout_net_38 ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04250_ ) );
NAND3_X1 _11991_ ( .A1(_04248_ ), .A2(_04250_ ), .A3(_04136_ ), .ZN(_04251_ ) );
MUX2_X1 _11992_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04252_ ) );
MUX2_X1 _11993_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04253_ ) );
MUX2_X1 _11994_ ( .A(_04252_ ), .B(_04253_ ), .S(_04197_ ), .Z(_04254_ ) );
BUF_X4 _11995_ ( .A(_04136_ ), .Z(_04255_ ) );
OAI211_X1 _11996_ ( .A(fanout_net_41 ), .B(_04251_ ), .C1(_04254_ ), .C2(_04255_ ), .ZN(_04256_ ) );
NAND2_X1 _11997_ ( .A1(_02113_ ), .A2(fanout_net_31 ), .ZN(_04257_ ) );
BUF_X4 _11998_ ( .A(_04058_ ), .Z(_04258_ ) );
OAI211_X1 _11999_ ( .A(_04257_ ), .B(_04258_ ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04259_ ) );
NAND2_X1 _12000_ ( .A1(_02116_ ), .A2(fanout_net_31 ), .ZN(_04260_ ) );
OAI211_X1 _12001_ ( .A(_04260_ ), .B(fanout_net_38 ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04261_ ) );
NAND3_X1 _12002_ ( .A1(_04259_ ), .A2(_04261_ ), .A3(_04136_ ), .ZN(_04262_ ) );
MUX2_X1 _12003_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04263_ ) );
MUX2_X1 _12004_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04264_ ) );
MUX2_X1 _12005_ ( .A(_04263_ ), .B(_04264_ ), .S(_04197_ ), .Z(_04265_ ) );
OAI211_X1 _12006_ ( .A(_04117_ ), .B(_04262_ ), .C1(_04265_ ), .C2(_04255_ ), .ZN(_04266_ ) );
OAI211_X1 _12007_ ( .A(_04256_ ), .B(_04266_ ), .C1(_04215_ ), .C2(_02861_ ), .ZN(_04267_ ) );
NAND2_X1 _12008_ ( .A1(_04245_ ), .A2(_04267_ ), .ZN(_04268_ ) );
XNOR2_X1 _12009_ ( .A(_04268_ ), .B(_02125_ ), .ZN(_04269_ ) );
OR3_X1 _12010_ ( .A1(_04085_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02095_ ), .ZN(_04270_ ) );
OR2_X1 _12011_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04271_ ) );
OAI211_X1 _12012_ ( .A(_04271_ ), .B(_04258_ ), .C1(_04198_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04272_ ) );
OR2_X1 _12013_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04273_ ) );
OAI211_X1 _12014_ ( .A(_04273_ ), .B(fanout_net_38 ), .C1(_04198_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04274_ ) );
NAND3_X1 _12015_ ( .A1(_04272_ ), .A2(_04274_ ), .A3(_04136_ ), .ZN(_04275_ ) );
MUX2_X1 _12016_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04276_ ) );
MUX2_X1 _12017_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04277_ ) );
MUX2_X1 _12018_ ( .A(_04276_ ), .B(_04277_ ), .S(_04197_ ), .Z(_04278_ ) );
OAI211_X1 _12019_ ( .A(fanout_net_41 ), .B(_04275_ ), .C1(_04278_ ), .C2(_04204_ ), .ZN(_04279_ ) );
OR2_X1 _12020_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04280_ ) );
OAI211_X1 _12021_ ( .A(_04280_ ), .B(_04258_ ), .C1(_04198_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04281_ ) );
OR2_X1 _12022_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04282_ ) );
OAI211_X1 _12023_ ( .A(_04282_ ), .B(fanout_net_38 ), .C1(_04198_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04283_ ) );
NAND3_X1 _12024_ ( .A1(_04281_ ), .A2(_04283_ ), .A3(_04136_ ), .ZN(_04284_ ) );
MUX2_X1 _12025_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04285_ ) );
MUX2_X1 _12026_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04286_ ) );
MUX2_X1 _12027_ ( .A(_04285_ ), .B(_04286_ ), .S(_04197_ ), .Z(_04287_ ) );
OAI211_X1 _12028_ ( .A(_04117_ ), .B(_04284_ ), .C1(_04287_ ), .C2(_04204_ ), .ZN(_04288_ ) );
OAI211_X1 _12029_ ( .A(_04279_ ), .B(_04288_ ), .C1(_04215_ ), .C2(_02861_ ), .ZN(_04289_ ) );
NAND2_X1 _12030_ ( .A1(_04270_ ), .A2(_04289_ ), .ZN(_04290_ ) );
XNOR2_X1 _12031_ ( .A(_04290_ ), .B(_02894_ ), .ZN(_04291_ ) );
AND2_X1 _12032_ ( .A1(_04269_ ), .A2(_04291_ ), .ZN(_04292_ ) );
NOR2_X4 _12033_ ( .A1(_04047_ ), .A2(_02354_ ), .ZN(_04293_ ) );
NAND2_X1 _12034_ ( .A1(_04293_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04294_ ) );
OR2_X1 _12035_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04295_ ) );
BUF_X4 _12036_ ( .A(_04119_ ), .Z(_04296_ ) );
OAI211_X1 _12037_ ( .A(_04295_ ), .B(_04247_ ), .C1(_04296_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04297_ ) );
NAND2_X1 _12038_ ( .A1(_02908_ ), .A2(fanout_net_31 ), .ZN(_04298_ ) );
OAI211_X1 _12039_ ( .A(_04298_ ), .B(fanout_net_38 ), .C1(fanout_net_31 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04299_ ) );
NAND3_X1 _12040_ ( .A1(_04297_ ), .A2(_04299_ ), .A3(_04204_ ), .ZN(_04300_ ) );
MUX2_X1 _12041_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04301_ ) );
MUX2_X1 _12042_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04302_ ) );
MUX2_X1 _12043_ ( .A(_04301_ ), .B(_04302_ ), .S(_04258_ ), .Z(_04303_ ) );
OAI211_X1 _12044_ ( .A(_04117_ ), .B(_04300_ ), .C1(_04303_ ), .C2(_04255_ ), .ZN(_04304_ ) );
OR2_X1 _12045_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04305_ ) );
OAI211_X1 _12046_ ( .A(_04305_ ), .B(fanout_net_38 ), .C1(_04296_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04306_ ) );
NAND2_X1 _12047_ ( .A1(_02918_ ), .A2(fanout_net_32 ), .ZN(_04307_ ) );
OAI211_X1 _12048_ ( .A(_04307_ ), .B(_04247_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04308_ ) );
NAND3_X1 _12049_ ( .A1(_04306_ ), .A2(_04308_ ), .A3(fanout_net_40 ), .ZN(_04309_ ) );
MUX2_X1 _12050_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04310_ ) );
MUX2_X1 _12051_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04311_ ) );
MUX2_X1 _12052_ ( .A(_04310_ ), .B(_04311_ ), .S(fanout_net_38 ), .Z(_04312_ ) );
OAI211_X1 _12053_ ( .A(fanout_net_41 ), .B(_04309_ ), .C1(_04312_ ), .C2(fanout_net_40 ), .ZN(_04313_ ) );
NAND2_X1 _12054_ ( .A1(_04304_ ), .A2(_04313_ ), .ZN(_04314_ ) );
OAI21_X1 _12055_ ( .A(_04314_ ), .B1(_04215_ ), .B2(_02861_ ), .ZN(_04315_ ) );
AND2_X1 _12056_ ( .A1(_04294_ ), .A2(_04315_ ), .ZN(_04316_ ) );
XNOR2_X1 _12057_ ( .A(_04316_ ), .B(_02928_ ), .ZN(_04317_ ) );
NAND2_X1 _12058_ ( .A1(_04293_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_04318_ ) );
OR2_X1 _12059_ ( .A1(_04119_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04319_ ) );
OAI211_X1 _12060_ ( .A(_04319_ ), .B(_04247_ ), .C1(fanout_net_32 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04320_ ) );
OR2_X1 _12061_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04321_ ) );
OAI211_X1 _12062_ ( .A(_04321_ ), .B(fanout_net_39 ), .C1(_04296_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04322_ ) );
NAND3_X1 _12063_ ( .A1(_04320_ ), .A2(_04204_ ), .A3(_04322_ ), .ZN(_04323_ ) );
MUX2_X1 _12064_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04324_ ) );
MUX2_X1 _12065_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04325_ ) );
MUX2_X1 _12066_ ( .A(_04324_ ), .B(_04325_ ), .S(_04258_ ), .Z(_04326_ ) );
OAI211_X1 _12067_ ( .A(_04117_ ), .B(_04323_ ), .C1(_04326_ ), .C2(_04255_ ), .ZN(_04327_ ) );
OR2_X1 _12068_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04328_ ) );
OAI211_X1 _12069_ ( .A(_04328_ ), .B(fanout_net_39 ), .C1(_04296_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04329_ ) );
OR2_X1 _12070_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04330_ ) );
OAI211_X1 _12071_ ( .A(_04330_ ), .B(_04247_ ), .C1(_04198_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04331_ ) );
NAND3_X1 _12072_ ( .A1(_04329_ ), .A2(_04331_ ), .A3(fanout_net_40 ), .ZN(_04332_ ) );
MUX2_X1 _12073_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04333_ ) );
MUX2_X1 _12074_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04334_ ) );
MUX2_X1 _12075_ ( .A(_04333_ ), .B(_04334_ ), .S(fanout_net_39 ), .Z(_04335_ ) );
OAI211_X1 _12076_ ( .A(fanout_net_41 ), .B(_04332_ ), .C1(_04335_ ), .C2(fanout_net_40 ), .ZN(_04336_ ) );
NAND2_X1 _12077_ ( .A1(_04327_ ), .A2(_04336_ ), .ZN(_04337_ ) );
OAI21_X1 _12078_ ( .A(_04337_ ), .B1(_04215_ ), .B2(_02861_ ), .ZN(_04338_ ) );
AND2_X1 _12079_ ( .A1(_04318_ ), .A2(_04338_ ), .ZN(_04339_ ) );
INV_X1 _12080_ ( .A(_02090_ ), .ZN(_04340_ ) );
XNOR2_X1 _12081_ ( .A(_04339_ ), .B(_04340_ ), .ZN(_04341_ ) );
AND3_X1 _12082_ ( .A1(_04292_ ), .A2(_04317_ ), .A3(_04341_ ), .ZN(_04342_ ) );
OR2_X1 _12083_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04343_ ) );
OAI211_X1 _12084_ ( .A(_04343_ ), .B(fanout_net_39 ), .C1(_04296_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04344_ ) );
NAND2_X1 _12085_ ( .A1(_02822_ ), .A2(fanout_net_32 ), .ZN(_04345_ ) );
OAI211_X1 _12086_ ( .A(_04345_ ), .B(_04247_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04346_ ) );
NAND3_X1 _12087_ ( .A1(_04344_ ), .A2(_04346_ ), .A3(_04204_ ), .ZN(_04347_ ) );
MUX2_X1 _12088_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04348_ ) );
MUX2_X1 _12089_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04349_ ) );
MUX2_X1 _12090_ ( .A(_04348_ ), .B(_04349_ ), .S(_04197_ ), .Z(_04350_ ) );
OAI211_X1 _12091_ ( .A(fanout_net_41 ), .B(_04347_ ), .C1(_04350_ ), .C2(_04255_ ), .ZN(_04351_ ) );
MUX2_X1 _12092_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04352_ ) );
AND2_X1 _12093_ ( .A1(_04352_ ), .A2(_04197_ ), .ZN(_04353_ ) );
MUX2_X1 _12094_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04354_ ) );
AOI211_X1 _12095_ ( .A(fanout_net_40 ), .B(_04353_ ), .C1(fanout_net_39 ), .C2(_04354_ ), .ZN(_04355_ ) );
MUX2_X1 _12096_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04356_ ) );
MUX2_X1 _12097_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04357_ ) );
MUX2_X1 _12098_ ( .A(_04356_ ), .B(_04357_ ), .S(_04058_ ), .Z(_04358_ ) );
OAI21_X1 _12099_ ( .A(_04117_ ), .B1(_04358_ ), .B2(_04204_ ), .ZN(_04359_ ) );
OAI221_X1 _12100_ ( .A(_04351_ ), .B1(_04355_ ), .B2(_04359_ ), .C1(_04215_ ), .C2(_02861_ ), .ZN(_04360_ ) );
INV_X1 _12101_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04361_ ) );
OR3_X4 _12102_ ( .A1(_04215_ ), .A2(_04361_ ), .A3(_02088_ ), .ZN(_04362_ ) );
NAND2_X1 _12103_ ( .A1(_04360_ ), .A2(_04362_ ), .ZN(_04363_ ) );
NAND2_X1 _12104_ ( .A1(_02818_ ), .A2(_02839_ ), .ZN(_04364_ ) );
XNOR2_X2 _12105_ ( .A(_04363_ ), .B(_04364_ ), .ZN(_04365_ ) );
NAND2_X1 _12106_ ( .A1(_04293_ ), .A2(\EX_LS_result_reg [26] ), .ZN(_04366_ ) );
OR2_X1 _12107_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04367_ ) );
OAI211_X1 _12108_ ( .A(_04367_ ), .B(fanout_net_39 ), .C1(_04296_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04368_ ) );
NAND2_X1 _12109_ ( .A1(_02852_ ), .A2(fanout_net_32 ), .ZN(_04369_ ) );
OAI211_X1 _12110_ ( .A(_04369_ ), .B(_04247_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04370_ ) );
NAND3_X1 _12111_ ( .A1(_04368_ ), .A2(_04370_ ), .A3(_04204_ ), .ZN(_04371_ ) );
MUX2_X1 _12112_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04372_ ) );
MUX2_X1 _12113_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04373_ ) );
MUX2_X1 _12114_ ( .A(_04372_ ), .B(_04373_ ), .S(_04258_ ), .Z(_04374_ ) );
OAI211_X1 _12115_ ( .A(fanout_net_41 ), .B(_04371_ ), .C1(_04374_ ), .C2(_04255_ ), .ZN(_04375_ ) );
OR2_X1 _12116_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04376_ ) );
OAI211_X1 _12117_ ( .A(_04376_ ), .B(_04258_ ), .C1(_04198_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04377_ ) );
NOR2_X1 _12118_ ( .A1(_04296_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04378_ ) );
OAI21_X1 _12119_ ( .A(fanout_net_39 ), .B1(fanout_net_32 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04379_ ) );
OAI211_X1 _12120_ ( .A(_04377_ ), .B(_04136_ ), .C1(_04378_ ), .C2(_04379_ ), .ZN(_04380_ ) );
MUX2_X1 _12121_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04381_ ) );
MUX2_X1 _12122_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04382_ ) );
MUX2_X1 _12123_ ( .A(_04381_ ), .B(_04382_ ), .S(_04258_ ), .Z(_04383_ ) );
OAI211_X1 _12124_ ( .A(_04117_ ), .B(_04380_ ), .C1(_04383_ ), .C2(_04255_ ), .ZN(_04384_ ) );
OAI211_X1 _12125_ ( .A(_04375_ ), .B(_04384_ ), .C1(_04215_ ), .C2(_02861_ ), .ZN(_04385_ ) );
NAND2_X1 _12126_ ( .A1(_04366_ ), .A2(_04385_ ), .ZN(_04386_ ) );
XNOR2_X1 _12127_ ( .A(_04386_ ), .B(_02864_ ), .ZN(_04387_ ) );
AND2_X1 _12128_ ( .A1(_04365_ ), .A2(_04387_ ), .ZN(_04388_ ) );
NAND2_X1 _12129_ ( .A1(_04293_ ), .A2(\EX_LS_result_reg [24] ), .ZN(_04389_ ) );
OR2_X1 _12130_ ( .A1(_04119_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04390_ ) );
OAI211_X1 _12131_ ( .A(_04390_ ), .B(_04247_ ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04391_ ) );
OR2_X1 _12132_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04392_ ) );
OAI211_X1 _12133_ ( .A(_04392_ ), .B(fanout_net_39 ), .C1(_04296_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04393_ ) );
NAND3_X1 _12134_ ( .A1(_04391_ ), .A2(fanout_net_40 ), .A3(_04393_ ), .ZN(_04394_ ) );
MUX2_X1 _12135_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04395_ ) );
MUX2_X1 _12136_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04396_ ) );
MUX2_X1 _12137_ ( .A(_04395_ ), .B(_04396_ ), .S(_04258_ ), .Z(_04397_ ) );
OAI211_X1 _12138_ ( .A(_04117_ ), .B(_04394_ ), .C1(_04397_ ), .C2(fanout_net_40 ), .ZN(_04398_ ) );
NOR2_X1 _12139_ ( .A1(_04198_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04399_ ) );
OAI21_X1 _12140_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04400_ ) );
NOR2_X1 _12141_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04401_ ) );
OAI21_X1 _12142_ ( .A(_04258_ ), .B1(_04198_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04402_ ) );
OAI221_X1 _12143_ ( .A(_04136_ ), .B1(_04399_ ), .B2(_04400_ ), .C1(_04401_ ), .C2(_04402_ ), .ZN(_04403_ ) );
MUX2_X1 _12144_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04404_ ) );
MUX2_X1 _12145_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04405_ ) );
MUX2_X1 _12146_ ( .A(_04404_ ), .B(_04405_ ), .S(fanout_net_39 ), .Z(_04406_ ) );
OAI211_X1 _12147_ ( .A(fanout_net_41 ), .B(_04403_ ), .C1(_04406_ ), .C2(_04255_ ), .ZN(_04407_ ) );
OAI211_X1 _12148_ ( .A(_04398_ ), .B(_04407_ ), .C1(_04215_ ), .C2(_02861_ ), .ZN(_04408_ ) );
NAND2_X1 _12149_ ( .A1(_04389_ ), .A2(_04408_ ), .ZN(_04409_ ) );
XNOR2_X1 _12150_ ( .A(_04409_ ), .B(_02787_ ), .ZN(_04410_ ) );
INV_X1 _12151_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04411_ ) );
OR3_X1 _12152_ ( .A1(_04085_ ), .A2(_04411_ ), .A3(_02088_ ), .ZN(_04412_ ) );
OR2_X1 _12153_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04413_ ) );
OAI211_X1 _12154_ ( .A(_04413_ ), .B(_04247_ ), .C1(_04296_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04414_ ) );
OR2_X1 _12155_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04415_ ) );
OAI211_X1 _12156_ ( .A(_04415_ ), .B(fanout_net_39 ), .C1(_04198_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04416_ ) );
NAND3_X1 _12157_ ( .A1(_04414_ ), .A2(_04416_ ), .A3(_04204_ ), .ZN(_04417_ ) );
MUX2_X1 _12158_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04418_ ) );
MUX2_X1 _12159_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04419_ ) );
MUX2_X1 _12160_ ( .A(_04418_ ), .B(_04419_ ), .S(_04197_ ), .Z(_04420_ ) );
OAI211_X1 _12161_ ( .A(fanout_net_41 ), .B(_04417_ ), .C1(_04420_ ), .C2(_04255_ ), .ZN(_04421_ ) );
OR2_X1 _12162_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04422_ ) );
OAI211_X1 _12163_ ( .A(_04422_ ), .B(_04247_ ), .C1(_04296_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04423_ ) );
NAND2_X1 _12164_ ( .A1(_02796_ ), .A2(fanout_net_33 ), .ZN(_04424_ ) );
OAI211_X1 _12165_ ( .A(_04424_ ), .B(fanout_net_39 ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04425_ ) );
NAND3_X1 _12166_ ( .A1(_04423_ ), .A2(_04425_ ), .A3(_04204_ ), .ZN(_04426_ ) );
MUX2_X1 _12167_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04427_ ) );
MUX2_X1 _12168_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04428_ ) );
MUX2_X1 _12169_ ( .A(_04427_ ), .B(_04428_ ), .S(_04197_ ), .Z(_04429_ ) );
OAI211_X1 _12170_ ( .A(_04117_ ), .B(_04426_ ), .C1(_04429_ ), .C2(_04255_ ), .ZN(_04430_ ) );
OAI211_X1 _12171_ ( .A(_04421_ ), .B(_04430_ ), .C1(_04215_ ), .C2(_02861_ ), .ZN(_04431_ ) );
NAND2_X1 _12172_ ( .A1(_04412_ ), .A2(_04431_ ), .ZN(_04432_ ) );
XNOR2_X1 _12173_ ( .A(_04432_ ), .B(_02814_ ), .ZN(_04433_ ) );
AND2_X1 _12174_ ( .A1(_04410_ ), .A2(_04433_ ), .ZN(_04434_ ) );
AND2_X1 _12175_ ( .A1(_04388_ ), .A2(_04434_ ), .ZN(_04435_ ) );
AND2_X2 _12176_ ( .A1(_04342_ ), .A2(_04435_ ), .ZN(_04436_ ) );
AND2_X1 _12177_ ( .A1(_04244_ ), .A2(_04436_ ), .ZN(_04437_ ) );
OR3_X2 _12178_ ( .A1(_04013_ ), .A2(\EX_LS_result_reg [1] ), .A3(_02354_ ), .ZN(_04438_ ) );
OR2_X1 _12179_ ( .A1(_04059_ ), .A2(\myreg.Reg[1][1] ), .ZN(_04439_ ) );
OAI211_X1 _12180_ ( .A(_04439_ ), .B(_04021_ ), .C1(fanout_net_33 ), .C2(\myreg.Reg[0][1] ), .ZN(_04440_ ) );
OR2_X1 _12181_ ( .A1(_04023_ ), .A2(\myreg.Reg[3][1] ), .ZN(_04441_ ) );
OAI211_X1 _12182_ ( .A(_04441_ ), .B(fanout_net_39 ), .C1(fanout_net_33 ), .C2(\myreg.Reg[2][1] ), .ZN(_04442_ ) );
NAND3_X1 _12183_ ( .A1(_04440_ ), .A2(_04442_ ), .A3(_04029_ ), .ZN(_04443_ ) );
MUX2_X1 _12184_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(fanout_net_33 ), .Z(_04444_ ) );
MUX2_X1 _12185_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(fanout_net_33 ), .Z(_04445_ ) );
MUX2_X1 _12186_ ( .A(_04444_ ), .B(_04445_ ), .S(_04021_ ), .Z(_04446_ ) );
OAI211_X1 _12187_ ( .A(_04017_ ), .B(_04443_ ), .C1(_04446_ ), .C2(_04030_ ), .ZN(_04447_ ) );
OR2_X1 _12188_ ( .A1(_04059_ ), .A2(\myreg.Reg[15][1] ), .ZN(_04448_ ) );
OAI211_X1 _12189_ ( .A(_04448_ ), .B(fanout_net_39 ), .C1(fanout_net_33 ), .C2(\myreg.Reg[14][1] ), .ZN(_04449_ ) );
OR2_X1 _12190_ ( .A1(_04023_ ), .A2(\myreg.Reg[13][1] ), .ZN(_04450_ ) );
OAI211_X1 _12191_ ( .A(_04450_ ), .B(_04021_ ), .C1(fanout_net_33 ), .C2(\myreg.Reg[12][1] ), .ZN(_04451_ ) );
NAND3_X1 _12192_ ( .A1(_04449_ ), .A2(_04451_ ), .A3(fanout_net_40 ), .ZN(_04452_ ) );
MUX2_X1 _12193_ ( .A(\myreg.Reg[8][1] ), .B(\myreg.Reg[9][1] ), .S(fanout_net_33 ), .Z(_04453_ ) );
MUX2_X1 _12194_ ( .A(\myreg.Reg[10][1] ), .B(\myreg.Reg[11][1] ), .S(fanout_net_33 ), .Z(_04454_ ) );
MUX2_X1 _12195_ ( .A(_04453_ ), .B(_04454_ ), .S(fanout_net_39 ), .Z(_04455_ ) );
OAI211_X1 _12196_ ( .A(fanout_net_41 ), .B(_04452_ ), .C1(_04455_ ), .C2(fanout_net_40 ), .ZN(_04456_ ) );
OAI211_X2 _12197_ ( .A(_04447_ ), .B(_04456_ ), .C1(_04047_ ), .C2(_02354_ ), .ZN(_04457_ ) );
NAND2_X2 _12198_ ( .A1(_04438_ ), .A2(_04457_ ), .ZN(_04458_ ) );
NAND2_X1 _12199_ ( .A1(_04458_ ), .A2(_02399_ ), .ZN(_04459_ ) );
NAND4_X1 _12200_ ( .A1(_04438_ ), .A2(_02379_ ), .A3(_02398_ ), .A4(_04457_ ), .ZN(_04460_ ) );
AND2_X1 _12201_ ( .A1(_04459_ ), .A2(_04460_ ), .ZN(_04461_ ) );
INV_X1 _12202_ ( .A(_04461_ ), .ZN(_04462_ ) );
INV_X1 _12203_ ( .A(\EX_LS_result_reg [0] ), .ZN(_04463_ ) );
OR3_X4 _12204_ ( .A1(_04047_ ), .A2(_04463_ ), .A3(_02354_ ), .ZN(_04464_ ) );
OR2_X1 _12205_ ( .A1(_04023_ ), .A2(\myreg.Reg[3][0] ), .ZN(_04465_ ) );
OAI211_X1 _12206_ ( .A(_04465_ ), .B(fanout_net_39 ), .C1(fanout_net_33 ), .C2(\myreg.Reg[2][0] ), .ZN(_04466_ ) );
OR2_X1 _12207_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[0][0] ), .ZN(_04467_ ) );
OAI211_X1 _12208_ ( .A(_04467_ ), .B(_04021_ ), .C1(_04024_ ), .C2(\myreg.Reg[1][0] ), .ZN(_04468_ ) );
NAND3_X1 _12209_ ( .A1(_04466_ ), .A2(_04029_ ), .A3(_04468_ ), .ZN(_04469_ ) );
MUX2_X1 _12210_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_33 ), .Z(_04470_ ) );
MUX2_X1 _12211_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_33 ), .Z(_04471_ ) );
MUX2_X1 _12212_ ( .A(_04470_ ), .B(_04471_ ), .S(_04020_ ), .Z(_04472_ ) );
OAI211_X1 _12213_ ( .A(_04017_ ), .B(_04469_ ), .C1(_04472_ ), .C2(_04030_ ), .ZN(_04473_ ) );
OR2_X1 _12214_ ( .A1(_04023_ ), .A2(\myreg.Reg[13][0] ), .ZN(_04474_ ) );
OAI211_X1 _12215_ ( .A(_04474_ ), .B(_04021_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[12][0] ), .ZN(_04475_ ) );
OR2_X1 _12216_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[14][0] ), .ZN(_04476_ ) );
OAI211_X1 _12217_ ( .A(_04476_ ), .B(fanout_net_39 ), .C1(_04024_ ), .C2(\myreg.Reg[15][0] ), .ZN(_04477_ ) );
NAND3_X1 _12218_ ( .A1(_04475_ ), .A2(fanout_net_40 ), .A3(_04477_ ), .ZN(_04478_ ) );
MUX2_X1 _12219_ ( .A(\myreg.Reg[8][0] ), .B(\myreg.Reg[9][0] ), .S(fanout_net_34 ), .Z(_04479_ ) );
MUX2_X1 _12220_ ( .A(\myreg.Reg[10][0] ), .B(\myreg.Reg[11][0] ), .S(fanout_net_34 ), .Z(_04480_ ) );
MUX2_X1 _12221_ ( .A(_04479_ ), .B(_04480_ ), .S(fanout_net_39 ), .Z(_04481_ ) );
OAI211_X1 _12222_ ( .A(fanout_net_41 ), .B(_04478_ ), .C1(_04481_ ), .C2(fanout_net_40 ), .ZN(_04482_ ) );
NAND2_X1 _12223_ ( .A1(_04473_ ), .A2(_04482_ ), .ZN(_04483_ ) );
OAI21_X4 _12224_ ( .A(_04483_ ), .B1(_04047_ ), .B2(_02043_ ), .ZN(_04484_ ) );
AND2_X1 _12225_ ( .A1(_04464_ ), .A2(_04484_ ), .ZN(_04485_ ) );
AND2_X2 _12226_ ( .A1(_02403_ ), .A2(_02423_ ), .ZN(_04486_ ) );
XNOR2_X1 _12227_ ( .A(_04485_ ), .B(_04486_ ), .ZN(_04487_ ) );
NOR2_X1 _12228_ ( .A1(_04462_ ), .A2(_04487_ ), .ZN(_04488_ ) );
OR3_X4 _12229_ ( .A1(_04047_ ), .A2(\EX_LS_result_reg [2] ), .A3(_02043_ ), .ZN(_04489_ ) );
OR2_X1 _12230_ ( .A1(_04024_ ), .A2(\myreg.Reg[1][2] ), .ZN(_04490_ ) );
OAI211_X1 _12231_ ( .A(_04490_ ), .B(_04022_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[0][2] ), .ZN(_04491_ ) );
OR2_X1 _12232_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[2][2] ), .ZN(_04492_ ) );
BUF_X4 _12233_ ( .A(_04059_ ), .Z(_04493_ ) );
OAI211_X1 _12234_ ( .A(_04492_ ), .B(fanout_net_39 ), .C1(_04493_ ), .C2(\myreg.Reg[3][2] ), .ZN(_04494_ ) );
NAND3_X1 _12235_ ( .A1(_04491_ ), .A2(_04030_ ), .A3(_04494_ ), .ZN(_04495_ ) );
MUX2_X1 _12236_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_34 ), .Z(_04496_ ) );
MUX2_X1 _12237_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_34 ), .Z(_04497_ ) );
MUX2_X1 _12238_ ( .A(_04496_ ), .B(_04497_ ), .S(_04056_ ), .Z(_04498_ ) );
OAI211_X1 _12239_ ( .A(_04018_ ), .B(_04495_ ), .C1(_04498_ ), .C2(_04035_ ), .ZN(_04499_ ) );
OR2_X1 _12240_ ( .A1(_04024_ ), .A2(\myreg.Reg[15][2] ), .ZN(_04500_ ) );
OAI211_X1 _12241_ ( .A(_04500_ ), .B(fanout_net_39 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[14][2] ), .ZN(_04501_ ) );
OR2_X1 _12242_ ( .A1(_04059_ ), .A2(\myreg.Reg[13][2] ), .ZN(_04502_ ) );
OAI211_X1 _12243_ ( .A(_04502_ ), .B(_04056_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[12][2] ), .ZN(_04503_ ) );
NAND3_X1 _12244_ ( .A1(_04501_ ), .A2(_04503_ ), .A3(fanout_net_40 ), .ZN(_04504_ ) );
MUX2_X1 _12245_ ( .A(\myreg.Reg[8][2] ), .B(\myreg.Reg[9][2] ), .S(fanout_net_34 ), .Z(_04505_ ) );
MUX2_X1 _12246_ ( .A(\myreg.Reg[10][2] ), .B(\myreg.Reg[11][2] ), .S(fanout_net_34 ), .Z(_04506_ ) );
MUX2_X1 _12247_ ( .A(_04505_ ), .B(_04506_ ), .S(fanout_net_39 ), .Z(_04507_ ) );
OAI211_X1 _12248_ ( .A(fanout_net_41 ), .B(_04504_ ), .C1(_04507_ ), .C2(fanout_net_40 ), .ZN(_04508_ ) );
OAI211_X4 _12249_ ( .A(_04499_ ), .B(_04508_ ), .C1(_04014_ ), .C2(_02327_ ), .ZN(_04509_ ) );
NAND2_X1 _12250_ ( .A1(_04489_ ), .A2(_04509_ ), .ZN(_04510_ ) );
INV_X1 _12251_ ( .A(_02376_ ), .ZN(_04511_ ) );
XNOR2_X1 _12252_ ( .A(_04510_ ), .B(_04511_ ), .ZN(_04512_ ) );
OR2_X1 _12253_ ( .A1(_04060_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04513_ ) );
OAI211_X1 _12254_ ( .A(_04513_ ), .B(_04146_ ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04514_ ) );
OR2_X1 _12255_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04515_ ) );
OAI211_X1 _12256_ ( .A(_04515_ ), .B(fanout_net_39 ), .C1(_04144_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04516_ ) );
NAND3_X1 _12257_ ( .A1(_04514_ ), .A2(_04035_ ), .A3(_04516_ ), .ZN(_04517_ ) );
MUX2_X1 _12258_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04518_ ) );
MUX2_X1 _12259_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04519_ ) );
MUX2_X1 _12260_ ( .A(_04518_ ), .B(_04519_ ), .S(_04146_ ), .Z(_04520_ ) );
OAI211_X1 _12261_ ( .A(_04018_ ), .B(_04517_ ), .C1(_04520_ ), .C2(_04066_ ), .ZN(_04521_ ) );
OR2_X1 _12262_ ( .A1(_04024_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04522_ ) );
OAI211_X1 _12263_ ( .A(_04522_ ), .B(_04146_ ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04523_ ) );
OR2_X1 _12264_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04524_ ) );
OAI211_X1 _12265_ ( .A(_04524_ ), .B(fanout_net_39 ), .C1(_04025_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04525_ ) );
NAND3_X1 _12266_ ( .A1(_04523_ ), .A2(fanout_net_40 ), .A3(_04525_ ), .ZN(_04526_ ) );
MUX2_X1 _12267_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04527_ ) );
MUX2_X1 _12268_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04528_ ) );
MUX2_X1 _12269_ ( .A(_04527_ ), .B(_04528_ ), .S(fanout_net_39 ), .Z(_04529_ ) );
OAI211_X1 _12270_ ( .A(fanout_net_41 ), .B(_04526_ ), .C1(_04529_ ), .C2(fanout_net_40 ), .ZN(_04530_ ) );
AOI21_X2 _12271_ ( .A(_04293_ ), .B1(_04521_ ), .B2(_04530_ ), .ZN(_04531_ ) );
AND2_X1 _12272_ ( .A1(_04293_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04532_ ) );
NOR2_X1 _12273_ ( .A1(_04531_ ), .A2(_04532_ ), .ZN(_04533_ ) );
XNOR2_X1 _12274_ ( .A(_04533_ ), .B(_02352_ ), .ZN(_04534_ ) );
AND3_X1 _12275_ ( .A1(_04488_ ), .A2(_04512_ ), .A3(_04534_ ), .ZN(_04535_ ) );
OR3_X4 _12276_ ( .A1(_04048_ ), .A2(\EX_LS_result_reg [12] ), .A3(_02127_ ), .ZN(_04536_ ) );
OR2_X1 _12277_ ( .A1(_04144_ ), .A2(\myreg.Reg[1][12] ), .ZN(_04537_ ) );
OAI211_X1 _12278_ ( .A(_04537_ ), .B(_04147_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[0][12] ), .ZN(_04538_ ) );
OR2_X1 _12279_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[2][12] ), .ZN(_04539_ ) );
OAI211_X1 _12280_ ( .A(_04539_ ), .B(fanout_net_39 ), .C1(_04101_ ), .C2(\myreg.Reg[3][12] ), .ZN(_04540_ ) );
NAND3_X1 _12281_ ( .A1(_04538_ ), .A2(_04075_ ), .A3(_04540_ ), .ZN(_04541_ ) );
MUX2_X1 _12282_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_34 ), .Z(_04542_ ) );
MUX2_X1 _12283_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_34 ), .Z(_04543_ ) );
MUX2_X1 _12284_ ( .A(_04542_ ), .B(_04543_ ), .S(_04147_ ), .Z(_04544_ ) );
OAI211_X1 _12285_ ( .A(_04074_ ), .B(_04541_ ), .C1(_04544_ ), .C2(_04075_ ), .ZN(_04545_ ) );
OR2_X1 _12286_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[14][12] ), .ZN(_04546_ ) );
OAI211_X1 _12287_ ( .A(_04546_ ), .B(fanout_net_39 ), .C1(_04101_ ), .C2(\myreg.Reg[15][12] ), .ZN(_04547_ ) );
OR2_X1 _12288_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[12][12] ), .ZN(_04548_ ) );
OAI211_X1 _12289_ ( .A(_04548_ ), .B(_04147_ ), .C1(_04101_ ), .C2(\myreg.Reg[13][12] ), .ZN(_04549_ ) );
NAND3_X1 _12290_ ( .A1(_04547_ ), .A2(_04549_ ), .A3(fanout_net_40 ), .ZN(_04550_ ) );
MUX2_X1 _12291_ ( .A(\myreg.Reg[8][12] ), .B(\myreg.Reg[9][12] ), .S(fanout_net_34 ), .Z(_04551_ ) );
MUX2_X1 _12292_ ( .A(\myreg.Reg[10][12] ), .B(\myreg.Reg[11][12] ), .S(fanout_net_34 ), .Z(_04552_ ) );
MUX2_X1 _12293_ ( .A(_04551_ ), .B(_04552_ ), .S(fanout_net_39 ), .Z(_04553_ ) );
OAI211_X1 _12294_ ( .A(fanout_net_41 ), .B(_04550_ ), .C1(_04553_ ), .C2(fanout_net_40 ), .ZN(_04554_ ) );
OAI211_X1 _12295_ ( .A(_04545_ ), .B(_04554_ ), .C1(_04053_ ), .C2(_02094_ ), .ZN(_04555_ ) );
NAND2_X1 _12296_ ( .A1(_04536_ ), .A2(_04555_ ), .ZN(_04556_ ) );
XNOR2_X1 _12297_ ( .A(_04556_ ), .B(_02561_ ), .ZN(_04557_ ) );
OR3_X4 _12298_ ( .A1(_04048_ ), .A2(\EX_LS_result_reg [13] ), .A3(_02355_ ), .ZN(_04558_ ) );
OR2_X1 _12299_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[8][13] ), .ZN(_04559_ ) );
OAI211_X1 _12300_ ( .A(_04559_ ), .B(_04057_ ), .C1(_04061_ ), .C2(\myreg.Reg[9][13] ), .ZN(_04560_ ) );
OR2_X1 _12301_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[10][13] ), .ZN(_04561_ ) );
OAI211_X1 _12302_ ( .A(_04561_ ), .B(fanout_net_39 ), .C1(_04061_ ), .C2(\myreg.Reg[11][13] ), .ZN(_04562_ ) );
NAND3_X1 _12303_ ( .A1(_04560_ ), .A2(_04562_ ), .A3(_04035_ ), .ZN(_04563_ ) );
MUX2_X1 _12304_ ( .A(\myreg.Reg[14][13] ), .B(\myreg.Reg[15][13] ), .S(fanout_net_35 ), .Z(_04564_ ) );
MUX2_X1 _12305_ ( .A(\myreg.Reg[12][13] ), .B(\myreg.Reg[13][13] ), .S(fanout_net_35 ), .Z(_04565_ ) );
MUX2_X1 _12306_ ( .A(_04564_ ), .B(_04565_ ), .S(_04057_ ), .Z(_04566_ ) );
OAI211_X1 _12307_ ( .A(fanout_net_41 ), .B(_04563_ ), .C1(_04566_ ), .C2(_04075_ ), .ZN(_04567_ ) );
NOR2_X1 _12308_ ( .A1(_04144_ ), .A2(\myreg.Reg[3][13] ), .ZN(_04568_ ) );
OAI21_X1 _12309_ ( .A(fanout_net_39 ), .B1(fanout_net_35 ), .B2(\myreg.Reg[2][13] ), .ZN(_04569_ ) );
NOR2_X1 _12310_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][13] ), .ZN(_04570_ ) );
OAI21_X1 _12311_ ( .A(_04057_ ), .B1(_04061_ ), .B2(\myreg.Reg[1][13] ), .ZN(_04571_ ) );
OAI221_X1 _12312_ ( .A(_04035_ ), .B1(_04568_ ), .B2(_04569_ ), .C1(_04570_ ), .C2(_04571_ ), .ZN(_04572_ ) );
MUX2_X1 _12313_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_35 ), .Z(_04573_ ) );
MUX2_X1 _12314_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_35 ), .Z(_04574_ ) );
MUX2_X1 _12315_ ( .A(_04573_ ), .B(_04574_ ), .S(_04057_ ), .Z(_04575_ ) );
OAI211_X1 _12316_ ( .A(_04074_ ), .B(_04572_ ), .C1(_04575_ ), .C2(_04075_ ), .ZN(_04576_ ) );
OAI211_X1 _12317_ ( .A(_04567_ ), .B(_04576_ ), .C1(_04048_ ), .C2(_02127_ ), .ZN(_04577_ ) );
NAND2_X1 _12318_ ( .A1(_04558_ ), .A2(_04577_ ), .ZN(_04578_ ) );
NAND2_X1 _12319_ ( .A1(_02564_ ), .A2(_02584_ ), .ZN(_04579_ ) );
AND2_X1 _12320_ ( .A1(_04578_ ), .A2(_04579_ ), .ZN(_04580_ ) );
NOR2_X1 _12321_ ( .A1(_04578_ ), .A2(_04579_ ), .ZN(_04581_ ) );
NOR3_X1 _12322_ ( .A1(_04557_ ), .A2(_04580_ ), .A3(_04581_ ), .ZN(_04582_ ) );
INV_X1 _12323_ ( .A(\EX_LS_result_reg [15] ), .ZN(_04583_ ) );
OR3_X4 _12324_ ( .A1(_04047_ ), .A2(_04583_ ), .A3(_02354_ ), .ZN(_04584_ ) );
OR2_X1 _12325_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][15] ), .ZN(_04585_ ) );
OAI211_X1 _12326_ ( .A(_04585_ ), .B(_04056_ ), .C1(_04060_ ), .C2(\myreg.Reg[1][15] ), .ZN(_04586_ ) );
OR2_X1 _12327_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][15] ), .ZN(_04587_ ) );
OAI211_X1 _12328_ ( .A(_04587_ ), .B(fanout_net_39 ), .C1(_04060_ ), .C2(\myreg.Reg[3][15] ), .ZN(_04588_ ) );
NAND3_X1 _12329_ ( .A1(_04586_ ), .A2(_04588_ ), .A3(_04029_ ), .ZN(_04589_ ) );
MUX2_X1 _12330_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_35 ), .Z(_04590_ ) );
MUX2_X1 _12331_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_35 ), .Z(_04591_ ) );
MUX2_X1 _12332_ ( .A(_04590_ ), .B(_04591_ ), .S(_04021_ ), .Z(_04592_ ) );
OAI211_X1 _12333_ ( .A(_04017_ ), .B(_04589_ ), .C1(_04592_ ), .C2(_04030_ ), .ZN(_04593_ ) );
OR2_X1 _12334_ ( .A1(_04059_ ), .A2(\myreg.Reg[15][15] ), .ZN(_04594_ ) );
OAI211_X1 _12335_ ( .A(_04594_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_35 ), .C2(\myreg.Reg[14][15] ), .ZN(_04595_ ) );
OR2_X1 _12336_ ( .A1(_04059_ ), .A2(\myreg.Reg[13][15] ), .ZN(_04596_ ) );
OAI211_X1 _12337_ ( .A(_04596_ ), .B(_04021_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[12][15] ), .ZN(_04597_ ) );
NAND3_X1 _12338_ ( .A1(_04595_ ), .A2(_04597_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04598_ ) );
MUX2_X1 _12339_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_35 ), .Z(_04599_ ) );
MUX2_X1 _12340_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_35 ), .Z(_04600_ ) );
MUX2_X1 _12341_ ( .A(_04599_ ), .B(_04600_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04601_ ) );
OAI211_X1 _12342_ ( .A(fanout_net_41 ), .B(_04598_ ), .C1(_04601_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04602_ ) );
NAND2_X1 _12343_ ( .A1(_04593_ ), .A2(_04602_ ), .ZN(_04603_ ) );
OAI21_X1 _12344_ ( .A(_04603_ ), .B1(_04014_ ), .B2(_02327_ ), .ZN(_04604_ ) );
AND2_X2 _12345_ ( .A1(_04584_ ), .A2(_04604_ ), .ZN(_04605_ ) );
INV_X1 _12346_ ( .A(_02609_ ), .ZN(_04606_ ) );
XNOR2_X1 _12347_ ( .A(_04605_ ), .B(_04606_ ), .ZN(_04607_ ) );
OR3_X4 _12348_ ( .A1(_04014_ ), .A2(\EX_LS_result_reg [14] ), .A3(_02327_ ), .ZN(_04608_ ) );
OR2_X1 _12349_ ( .A1(_04060_ ), .A2(\myreg.Reg[1][14] ), .ZN(_04609_ ) );
OAI211_X1 _12350_ ( .A(_04609_ ), .B(_04057_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[0][14] ), .ZN(_04610_ ) );
OR2_X1 _12351_ ( .A1(_04060_ ), .A2(\myreg.Reg[3][14] ), .ZN(_04611_ ) );
OAI211_X1 _12352_ ( .A(_04611_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_35 ), .C2(\myreg.Reg[2][14] ), .ZN(_04612_ ) );
NAND3_X1 _12353_ ( .A1(_04610_ ), .A2(_04612_ ), .A3(_04035_ ), .ZN(_04613_ ) );
MUX2_X1 _12354_ ( .A(\myreg.Reg[6][14] ), .B(\myreg.Reg[7][14] ), .S(fanout_net_35 ), .Z(_04614_ ) );
MUX2_X1 _12355_ ( .A(\myreg.Reg[4][14] ), .B(\myreg.Reg[5][14] ), .S(fanout_net_35 ), .Z(_04615_ ) );
MUX2_X1 _12356_ ( .A(_04614_ ), .B(_04615_ ), .S(_04146_ ), .Z(_04616_ ) );
OAI211_X1 _12357_ ( .A(_04018_ ), .B(_04613_ ), .C1(_04616_ ), .C2(_04066_ ), .ZN(_04617_ ) );
OR2_X1 _12358_ ( .A1(_04060_ ), .A2(\myreg.Reg[13][14] ), .ZN(_04618_ ) );
OAI211_X1 _12359_ ( .A(_04618_ ), .B(_04057_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[12][14] ), .ZN(_04619_ ) );
OR2_X1 _12360_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[14][14] ), .ZN(_04620_ ) );
OAI211_X1 _12361_ ( .A(_04620_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04144_ ), .C2(\myreg.Reg[15][14] ), .ZN(_04621_ ) );
NAND3_X1 _12362_ ( .A1(_04619_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04621_ ), .ZN(_04622_ ) );
MUX2_X1 _12363_ ( .A(\myreg.Reg[8][14] ), .B(\myreg.Reg[9][14] ), .S(fanout_net_35 ), .Z(_04623_ ) );
MUX2_X1 _12364_ ( .A(\myreg.Reg[10][14] ), .B(\myreg.Reg[11][14] ), .S(fanout_net_35 ), .Z(_04624_ ) );
MUX2_X1 _12365_ ( .A(_04623_ ), .B(_04624_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04625_ ) );
OAI211_X1 _12366_ ( .A(fanout_net_41 ), .B(_04622_ ), .C1(_04625_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04626_ ) );
OAI211_X1 _12367_ ( .A(_04617_ ), .B(_04626_ ), .C1(_04048_ ), .C2(_02093_ ), .ZN(_04627_ ) );
NAND2_X2 _12368_ ( .A1(_04608_ ), .A2(_04627_ ), .ZN(_04628_ ) );
INV_X1 _12369_ ( .A(_02631_ ), .ZN(_04629_ ) );
XNOR2_X1 _12370_ ( .A(_04628_ ), .B(_04629_ ), .ZN(_04630_ ) );
AND3_X1 _12371_ ( .A1(_04582_ ), .A2(_04607_ ), .A3(_04630_ ), .ZN(_04631_ ) );
OR3_X4 _12372_ ( .A1(_04047_ ), .A2(\EX_LS_result_reg [11] ), .A3(_02043_ ), .ZN(_04632_ ) );
OR2_X1 _12373_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[4][11] ), .ZN(_04633_ ) );
OAI211_X1 _12374_ ( .A(_04633_ ), .B(_04056_ ), .C1(_04493_ ), .C2(\myreg.Reg[5][11] ), .ZN(_04634_ ) );
OR2_X1 _12375_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[6][11] ), .ZN(_04635_ ) );
OAI211_X1 _12376_ ( .A(_04635_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04493_ ), .C2(\myreg.Reg[7][11] ), .ZN(_04636_ ) );
NAND3_X1 _12377_ ( .A1(_04634_ ), .A2(_04636_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04637_ ) );
MUX2_X1 _12378_ ( .A(\myreg.Reg[2][11] ), .B(\myreg.Reg[3][11] ), .S(fanout_net_35 ), .Z(_04638_ ) );
MUX2_X1 _12379_ ( .A(\myreg.Reg[0][11] ), .B(\myreg.Reg[1][11] ), .S(fanout_net_35 ), .Z(_04639_ ) );
MUX2_X1 _12380_ ( .A(_04638_ ), .B(_04639_ ), .S(_04056_ ), .Z(_04640_ ) );
OAI211_X1 _12381_ ( .A(_04018_ ), .B(_04637_ ), .C1(_04640_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04641_ ) );
NOR2_X1 _12382_ ( .A1(_04060_ ), .A2(\myreg.Reg[11][11] ), .ZN(_04642_ ) );
OAI21_X1 _12383_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_35 ), .B2(\myreg.Reg[10][11] ), .ZN(_04643_ ) );
NOR2_X1 _12384_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[8][11] ), .ZN(_04644_ ) );
OAI21_X1 _12385_ ( .A(_04056_ ), .B1(_04493_ ), .B2(\myreg.Reg[9][11] ), .ZN(_04645_ ) );
OAI221_X1 _12386_ ( .A(_04029_ ), .B1(_04642_ ), .B2(_04643_ ), .C1(_04644_ ), .C2(_04645_ ), .ZN(_04646_ ) );
MUX2_X1 _12387_ ( .A(\myreg.Reg[12][11] ), .B(\myreg.Reg[13][11] ), .S(fanout_net_35 ), .Z(_04647_ ) );
MUX2_X1 _12388_ ( .A(\myreg.Reg[14][11] ), .B(\myreg.Reg[15][11] ), .S(fanout_net_35 ), .Z(_04648_ ) );
MUX2_X1 _12389_ ( .A(_04647_ ), .B(_04648_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04649_ ) );
OAI211_X1 _12390_ ( .A(fanout_net_41 ), .B(_04646_ ), .C1(_04649_ ), .C2(_04035_ ), .ZN(_04650_ ) );
OAI211_X1 _12391_ ( .A(_04641_ ), .B(_04650_ ), .C1(_04014_ ), .C2(_02327_ ), .ZN(_04651_ ) );
NAND2_X1 _12392_ ( .A1(_04632_ ), .A2(_04651_ ), .ZN(_04652_ ) );
INV_X1 _12393_ ( .A(_02702_ ), .ZN(_04653_ ) );
XNOR2_X2 _12394_ ( .A(_04652_ ), .B(_04653_ ), .ZN(_04654_ ) );
OR3_X4 _12395_ ( .A1(_04014_ ), .A2(\EX_LS_result_reg [10] ), .A3(_02355_ ), .ZN(_04655_ ) );
OR2_X1 _12396_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[4][10] ), .ZN(_04656_ ) );
OAI211_X1 _12397_ ( .A(_04656_ ), .B(_04057_ ), .C1(_04061_ ), .C2(\myreg.Reg[5][10] ), .ZN(_04657_ ) );
OR2_X1 _12398_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[6][10] ), .ZN(_04658_ ) );
OAI211_X1 _12399_ ( .A(_04658_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04061_ ), .C2(\myreg.Reg[7][10] ), .ZN(_04659_ ) );
NAND3_X1 _12400_ ( .A1(_04657_ ), .A2(_04659_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04660_ ) );
MUX2_X1 _12401_ ( .A(\myreg.Reg[2][10] ), .B(\myreg.Reg[3][10] ), .S(fanout_net_36 ), .Z(_04661_ ) );
MUX2_X1 _12402_ ( .A(\myreg.Reg[0][10] ), .B(\myreg.Reg[1][10] ), .S(fanout_net_36 ), .Z(_04662_ ) );
MUX2_X1 _12403_ ( .A(_04661_ ), .B(_04662_ ), .S(_04146_ ), .Z(_04663_ ) );
OAI211_X1 _12404_ ( .A(_04074_ ), .B(_04660_ ), .C1(_04663_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04664_ ) );
NOR2_X1 _12405_ ( .A1(_04025_ ), .A2(\myreg.Reg[11][10] ), .ZN(_04665_ ) );
OAI21_X1 _12406_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_36 ), .B2(\myreg.Reg[10][10] ), .ZN(_04666_ ) );
NOR2_X1 _12407_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[8][10] ), .ZN(_04667_ ) );
OAI21_X1 _12408_ ( .A(_04146_ ), .B1(_04025_ ), .B2(\myreg.Reg[9][10] ), .ZN(_04668_ ) );
OAI221_X1 _12409_ ( .A(_04035_ ), .B1(_04665_ ), .B2(_04666_ ), .C1(_04667_ ), .C2(_04668_ ), .ZN(_04669_ ) );
MUX2_X1 _12410_ ( .A(\myreg.Reg[12][10] ), .B(\myreg.Reg[13][10] ), .S(fanout_net_36 ), .Z(_04670_ ) );
MUX2_X1 _12411_ ( .A(\myreg.Reg[14][10] ), .B(\myreg.Reg[15][10] ), .S(fanout_net_36 ), .Z(_04671_ ) );
MUX2_X1 _12412_ ( .A(_04670_ ), .B(_04671_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04672_ ) );
OAI211_X1 _12413_ ( .A(fanout_net_41 ), .B(_04669_ ), .C1(_04672_ ), .C2(_04066_ ), .ZN(_04673_ ) );
OAI211_X1 _12414_ ( .A(_04664_ ), .B(_04673_ ), .C1(_04048_ ), .C2(_02127_ ), .ZN(_04674_ ) );
NAND2_X1 _12415_ ( .A1(_04655_ ), .A2(_04674_ ), .ZN(_04675_ ) );
INV_X1 _12416_ ( .A(_02724_ ), .ZN(_04676_ ) );
XNOR2_X1 _12417_ ( .A(_04675_ ), .B(_04676_ ), .ZN(_04677_ ) );
AND2_X1 _12418_ ( .A1(_04654_ ), .A2(_04677_ ), .ZN(_04678_ ) );
OR3_X2 _12419_ ( .A1(_04053_ ), .A2(\EX_LS_result_reg [8] ), .A3(_02044_ ), .ZN(_04679_ ) );
OR2_X1 _12420_ ( .A1(_04061_ ), .A2(\myreg.Reg[1][8] ), .ZN(_04680_ ) );
OAI211_X1 _12421_ ( .A(_04680_ ), .B(_04071_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[0][8] ), .ZN(_04681_ ) );
OR2_X1 _12422_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[2][8] ), .ZN(_04682_ ) );
OAI211_X1 _12423_ ( .A(_04682_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04101_ ), .C2(\myreg.Reg[3][8] ), .ZN(_04683_ ) );
NAND3_X1 _12424_ ( .A1(_04681_ ), .A2(_04075_ ), .A3(_04683_ ), .ZN(_04684_ ) );
MUX2_X1 _12425_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_36 ), .Z(_04685_ ) );
MUX2_X1 _12426_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_36 ), .Z(_04686_ ) );
MUX2_X1 _12427_ ( .A(_04685_ ), .B(_04686_ ), .S(_04147_ ), .Z(_04687_ ) );
OAI211_X1 _12428_ ( .A(_04074_ ), .B(_04684_ ), .C1(_04687_ ), .C2(_04067_ ), .ZN(_04688_ ) );
OR2_X1 _12429_ ( .A1(_04144_ ), .A2(\myreg.Reg[15][8] ), .ZN(_04689_ ) );
OAI211_X1 _12430_ ( .A(_04689_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_36 ), .C2(\myreg.Reg[14][8] ), .ZN(_04690_ ) );
OR2_X1 _12431_ ( .A1(_04144_ ), .A2(\myreg.Reg[13][8] ), .ZN(_04691_ ) );
OAI211_X1 _12432_ ( .A(_04691_ ), .B(_04147_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[12][8] ), .ZN(_04692_ ) );
NAND3_X1 _12433_ ( .A1(_04690_ ), .A2(_04692_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04693_ ) );
MUX2_X1 _12434_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_36 ), .Z(_04694_ ) );
MUX2_X1 _12435_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_36 ), .Z(_04695_ ) );
MUX2_X1 _12436_ ( .A(_04694_ ), .B(_04695_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04696_ ) );
OAI211_X1 _12437_ ( .A(fanout_net_41 ), .B(_04693_ ), .C1(_04696_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04697_ ) );
OAI211_X1 _12438_ ( .A(_04688_ ), .B(_04697_ ), .C1(_04053_ ), .C2(_02094_ ), .ZN(_04698_ ) );
NAND2_X1 _12439_ ( .A1(_04679_ ), .A2(_04698_ ), .ZN(_04699_ ) );
INV_X1 _12440_ ( .A(_02655_ ), .ZN(_04700_ ) );
XNOR2_X1 _12441_ ( .A(_04699_ ), .B(_04700_ ), .ZN(_04701_ ) );
OR3_X4 _12442_ ( .A1(_04014_ ), .A2(\EX_LS_result_reg [9] ), .A3(_02043_ ), .ZN(_04702_ ) );
OR2_X1 _12443_ ( .A1(_04024_ ), .A2(\myreg.Reg[9][9] ), .ZN(_04703_ ) );
OAI211_X1 _12444_ ( .A(_04703_ ), .B(_04146_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[8][9] ), .ZN(_04704_ ) );
OR2_X1 _12445_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[10][9] ), .ZN(_04705_ ) );
OAI211_X1 _12446_ ( .A(_04705_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04025_ ), .C2(\myreg.Reg[11][9] ), .ZN(_04706_ ) );
NAND3_X1 _12447_ ( .A1(_04704_ ), .A2(_04035_ ), .A3(_04706_ ), .ZN(_04707_ ) );
MUX2_X1 _12448_ ( .A(\myreg.Reg[14][9] ), .B(\myreg.Reg[15][9] ), .S(fanout_net_36 ), .Z(_04708_ ) );
MUX2_X1 _12449_ ( .A(\myreg.Reg[12][9] ), .B(\myreg.Reg[13][9] ), .S(fanout_net_36 ), .Z(_04709_ ) );
MUX2_X1 _12450_ ( .A(_04708_ ), .B(_04709_ ), .S(_04022_ ), .Z(_04710_ ) );
OAI211_X1 _12451_ ( .A(fanout_net_41 ), .B(_04707_ ), .C1(_04710_ ), .C2(_04066_ ), .ZN(_04711_ ) );
OAI21_X1 _12452_ ( .A(_04056_ ), .B1(_04493_ ), .B2(\myreg.Reg[1][9] ), .ZN(_04712_ ) );
NOR2_X1 _12453_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[0][9] ), .ZN(_04713_ ) );
NOR2_X1 _12454_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[2][9] ), .ZN(_04714_ ) );
OAI21_X1 _12455_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(_04493_ ), .B2(\myreg.Reg[3][9] ), .ZN(_04715_ ) );
OAI221_X1 _12456_ ( .A(_04030_ ), .B1(_04712_ ), .B2(_04713_ ), .C1(_04714_ ), .C2(_04715_ ), .ZN(_04716_ ) );
MUX2_X1 _12457_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_36 ), .Z(_04717_ ) );
MUX2_X1 _12458_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_36 ), .Z(_04718_ ) );
MUX2_X1 _12459_ ( .A(_04717_ ), .B(_04718_ ), .S(_04022_ ), .Z(_04719_ ) );
OAI211_X1 _12460_ ( .A(_04018_ ), .B(_04716_ ), .C1(_04719_ ), .C2(_04066_ ), .ZN(_04720_ ) );
OAI211_X4 _12461_ ( .A(_04711_ ), .B(_04720_ ), .C1(_04048_ ), .C2(_02355_ ), .ZN(_04721_ ) );
NAND2_X1 _12462_ ( .A1(_04702_ ), .A2(_04721_ ), .ZN(_04722_ ) );
INV_X1 _12463_ ( .A(_02677_ ), .ZN(_04723_ ) );
XNOR2_X1 _12464_ ( .A(_04722_ ), .B(_04723_ ), .ZN(_04724_ ) );
AND3_X1 _12465_ ( .A1(_04678_ ), .A2(_04701_ ), .A3(_04724_ ), .ZN(_04725_ ) );
INV_X1 _12466_ ( .A(\EX_LS_result_reg [7] ), .ZN(_04726_ ) );
OR3_X4 _12467_ ( .A1(_04013_ ), .A2(_04726_ ), .A3(_02042_ ), .ZN(_04727_ ) );
OR2_X1 _12468_ ( .A1(_04023_ ), .A2(\myreg.Reg[1][7] ), .ZN(_04728_ ) );
OAI211_X1 _12469_ ( .A(_04728_ ), .B(_04020_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[0][7] ), .ZN(_04729_ ) );
OR2_X1 _12470_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[2][7] ), .ZN(_04730_ ) );
OAI211_X1 _12471_ ( .A(_04730_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04059_ ), .C2(\myreg.Reg[3][7] ), .ZN(_04731_ ) );
NAND3_X1 _12472_ ( .A1(_04729_ ), .A2(_04029_ ), .A3(_04731_ ), .ZN(_04732_ ) );
MUX2_X1 _12473_ ( .A(\myreg.Reg[6][7] ), .B(\myreg.Reg[7][7] ), .S(fanout_net_36 ), .Z(_04733_ ) );
MUX2_X1 _12474_ ( .A(\myreg.Reg[4][7] ), .B(\myreg.Reg[5][7] ), .S(fanout_net_36 ), .Z(_04734_ ) );
MUX2_X1 _12475_ ( .A(_04733_ ), .B(_04734_ ), .S(_04020_ ), .Z(_04735_ ) );
OAI211_X1 _12476_ ( .A(_04017_ ), .B(_04732_ ), .C1(_04735_ ), .C2(_04029_ ), .ZN(_04736_ ) );
OR2_X1 _12477_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][7] ), .ZN(_04737_ ) );
OAI211_X1 _12478_ ( .A(_04737_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04059_ ), .C2(\myreg.Reg[15][7] ), .ZN(_04738_ ) );
OR2_X1 _12479_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[12][7] ), .ZN(_04739_ ) );
OAI211_X1 _12480_ ( .A(_04739_ ), .B(_04020_ ), .C1(_04059_ ), .C2(\myreg.Reg[13][7] ), .ZN(_04740_ ) );
NAND3_X1 _12481_ ( .A1(_04738_ ), .A2(_04740_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04741_ ) );
MUX2_X1 _12482_ ( .A(\myreg.Reg[8][7] ), .B(\myreg.Reg[9][7] ), .S(fanout_net_37 ), .Z(_04742_ ) );
MUX2_X1 _12483_ ( .A(\myreg.Reg[10][7] ), .B(\myreg.Reg[11][7] ), .S(fanout_net_37 ), .Z(_04743_ ) );
MUX2_X1 _12484_ ( .A(_04742_ ), .B(_04743_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04744_ ) );
OAI211_X1 _12485_ ( .A(fanout_net_41 ), .B(_04741_ ), .C1(_04744_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04745_ ) );
NAND2_X1 _12486_ ( .A1(_04736_ ), .A2(_04745_ ), .ZN(_04746_ ) );
OAI21_X1 _12487_ ( .A(_04746_ ), .B1(_04013_ ), .B2(_02354_ ), .ZN(_04747_ ) );
AND2_X2 _12488_ ( .A1(_04727_ ), .A2(_04747_ ), .ZN(_04748_ ) );
INV_X1 _12489_ ( .A(_02477_ ), .ZN(_04749_ ) );
XNOR2_X1 _12490_ ( .A(_04748_ ), .B(_04749_ ), .ZN(_04750_ ) );
INV_X1 _12491_ ( .A(_04750_ ), .ZN(_04751_ ) );
OR3_X2 _12492_ ( .A1(_04014_ ), .A2(\EX_LS_result_reg [6] ), .A3(_02327_ ), .ZN(_04752_ ) );
OR2_X1 _12493_ ( .A1(_04060_ ), .A2(\myreg.Reg[7][6] ), .ZN(_04753_ ) );
OAI211_X1 _12494_ ( .A(_04753_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[6][6] ), .ZN(_04754_ ) );
OR2_X1 _12495_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[4][6] ), .ZN(_04755_ ) );
OAI211_X1 _12496_ ( .A(_04755_ ), .B(_04146_ ), .C1(_04144_ ), .C2(\myreg.Reg[5][6] ), .ZN(_04756_ ) );
NAND3_X1 _12497_ ( .A1(_04754_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04756_ ), .ZN(_04757_ ) );
MUX2_X1 _12498_ ( .A(\myreg.Reg[2][6] ), .B(\myreg.Reg[3][6] ), .S(fanout_net_37 ), .Z(_04758_ ) );
MUX2_X1 _12499_ ( .A(\myreg.Reg[0][6] ), .B(\myreg.Reg[1][6] ), .S(fanout_net_37 ), .Z(_04759_ ) );
MUX2_X1 _12500_ ( .A(_04758_ ), .B(_04759_ ), .S(_04022_ ), .Z(_04760_ ) );
OAI211_X1 _12501_ ( .A(_04018_ ), .B(_04757_ ), .C1(_04760_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04761_ ) );
NOR2_X1 _12502_ ( .A1(_04493_ ), .A2(\myreg.Reg[11][6] ), .ZN(_04762_ ) );
OAI21_X1 _12503_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_37 ), .B2(\myreg.Reg[10][6] ), .ZN(_04763_ ) );
NOR2_X1 _12504_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][6] ), .ZN(_04764_ ) );
OAI21_X1 _12505_ ( .A(_04022_ ), .B1(_04025_ ), .B2(\myreg.Reg[9][6] ), .ZN(_04765_ ) );
OAI221_X1 _12506_ ( .A(_04030_ ), .B1(_04762_ ), .B2(_04763_ ), .C1(_04764_ ), .C2(_04765_ ), .ZN(_04766_ ) );
MUX2_X1 _12507_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(fanout_net_37 ), .Z(_04767_ ) );
MUX2_X1 _12508_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(fanout_net_37 ), .Z(_04768_ ) );
MUX2_X1 _12509_ ( .A(_04767_ ), .B(_04768_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04769_ ) );
OAI211_X1 _12510_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04766_ ), .C1(_04769_ ), .C2(_04066_ ), .ZN(_04770_ ) );
OAI211_X4 _12511_ ( .A(_04761_ ), .B(_04770_ ), .C1(_04048_ ), .C2(_02093_ ), .ZN(_04771_ ) );
NAND2_X1 _12512_ ( .A1(_04752_ ), .A2(_04771_ ), .ZN(_04772_ ) );
XNOR2_X1 _12513_ ( .A(_04772_ ), .B(_02530_ ), .ZN(_04773_ ) );
NOR2_X1 _12514_ ( .A1(_04751_ ), .A2(_04773_ ), .ZN(_04774_ ) );
OR3_X2 _12515_ ( .A1(_04047_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02354_ ), .ZN(_04775_ ) );
OR2_X1 _12516_ ( .A1(fanout_net_37 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04776_ ) );
OAI211_X1 _12517_ ( .A(_04776_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04493_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04777_ ) );
NAND2_X1 _12518_ ( .A1(_02505_ ), .A2(fanout_net_37 ), .ZN(_04778_ ) );
OAI211_X1 _12519_ ( .A(_04778_ ), .B(_04056_ ), .C1(fanout_net_37 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04779_ ) );
NAND3_X1 _12520_ ( .A1(_04777_ ), .A2(_04779_ ), .A3(_04029_ ), .ZN(_04780_ ) );
MUX2_X1 _12521_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04781_ ) );
MUX2_X1 _12522_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04782_ ) );
MUX2_X1 _12523_ ( .A(_04781_ ), .B(_04782_ ), .S(_04021_ ), .Z(_04783_ ) );
OAI211_X1 _12524_ ( .A(_04018_ ), .B(_04780_ ), .C1(_04783_ ), .C2(_04030_ ), .ZN(_04784_ ) );
OR2_X1 _12525_ ( .A1(fanout_net_37 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04785_ ) );
OAI211_X1 _12526_ ( .A(_04785_ ), .B(_04056_ ), .C1(_04493_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04786_ ) );
NAND2_X1 _12527_ ( .A1(_02515_ ), .A2(fanout_net_37 ), .ZN(_04787_ ) );
OAI211_X1 _12528_ ( .A(_04787_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04788_ ) );
NAND3_X1 _12529_ ( .A1(_04786_ ), .A2(_04788_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04789_ ) );
MUX2_X1 _12530_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04790_ ) );
MUX2_X1 _12531_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04791_ ) );
MUX2_X1 _12532_ ( .A(_04790_ ), .B(_04791_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04792_ ) );
OAI211_X1 _12533_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04789_ ), .C1(_04792_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04793_ ) );
OAI211_X4 _12534_ ( .A(_04784_ ), .B(_04793_ ), .C1(_04047_ ), .C2(_02043_ ), .ZN(_04794_ ) );
NAND2_X2 _12535_ ( .A1(_04775_ ), .A2(_04794_ ), .ZN(_04795_ ) );
XNOR2_X1 _12536_ ( .A(_04795_ ), .B(_02525_ ), .ZN(_04796_ ) );
OR3_X1 _12537_ ( .A1(_04014_ ), .A2(\EX_LS_result_reg [4] ), .A3(_02327_ ), .ZN(_04797_ ) );
OR2_X1 _12538_ ( .A1(_04060_ ), .A2(\myreg.Reg[5][4] ), .ZN(_04798_ ) );
OAI211_X1 _12539_ ( .A(_04798_ ), .B(_04146_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[4][4] ), .ZN(_04799_ ) );
OR2_X1 _12540_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[6][4] ), .ZN(_04800_ ) );
OAI211_X1 _12541_ ( .A(_04800_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04025_ ), .C2(\myreg.Reg[7][4] ), .ZN(_04801_ ) );
NAND3_X1 _12542_ ( .A1(_04799_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04801_ ), .ZN(_04802_ ) );
MUX2_X1 _12543_ ( .A(\myreg.Reg[2][4] ), .B(\myreg.Reg[3][4] ), .S(fanout_net_37 ), .Z(_04803_ ) );
MUX2_X1 _12544_ ( .A(\myreg.Reg[0][4] ), .B(\myreg.Reg[1][4] ), .S(fanout_net_37 ), .Z(_04804_ ) );
MUX2_X1 _12545_ ( .A(_04803_ ), .B(_04804_ ), .S(_04022_ ), .Z(_04805_ ) );
OAI211_X1 _12546_ ( .A(_04018_ ), .B(_04802_ ), .C1(_04805_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04806_ ) );
NOR2_X1 _12547_ ( .A1(_04493_ ), .A2(\myreg.Reg[11][4] ), .ZN(_04807_ ) );
OAI21_X1 _12548_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_37 ), .B2(\myreg.Reg[10][4] ), .ZN(_04808_ ) );
NOR2_X1 _12549_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][4] ), .ZN(_04809_ ) );
OAI21_X1 _12550_ ( .A(_04022_ ), .B1(_04025_ ), .B2(\myreg.Reg[9][4] ), .ZN(_04810_ ) );
OAI221_X1 _12551_ ( .A(_04030_ ), .B1(_04807_ ), .B2(_04808_ ), .C1(_04809_ ), .C2(_04810_ ), .ZN(_04811_ ) );
MUX2_X1 _12552_ ( .A(\myreg.Reg[12][4] ), .B(\myreg.Reg[13][4] ), .S(fanout_net_37 ), .Z(_04812_ ) );
MUX2_X1 _12553_ ( .A(\myreg.Reg[14][4] ), .B(\myreg.Reg[15][4] ), .S(fanout_net_37 ), .Z(_04813_ ) );
MUX2_X1 _12554_ ( .A(_04812_ ), .B(_04813_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04814_ ) );
OAI211_X1 _12555_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04811_ ), .C1(_04814_ ), .C2(_04066_ ), .ZN(_04815_ ) );
OAI211_X4 _12556_ ( .A(_04806_ ), .B(_04815_ ), .C1(_04048_ ), .C2(_02093_ ), .ZN(_04816_ ) );
NAND2_X1 _12557_ ( .A1(_04797_ ), .A2(_04816_ ), .ZN(_04817_ ) );
XNOR2_X1 _12558_ ( .A(_04817_ ), .B(_02533_ ), .ZN(_04818_ ) );
AND2_X1 _12559_ ( .A1(_04796_ ), .A2(_04818_ ), .ZN(_04819_ ) );
AND4_X1 _12560_ ( .A1(_04631_ ), .A2(_04725_ ), .A3(_04774_ ), .A4(_04819_ ), .ZN(_04820_ ) );
NAND3_X1 _12561_ ( .A1(_04437_ ), .A2(_04535_ ), .A3(_04820_ ), .ZN(_04821_ ) );
NOR2_X1 _12562_ ( .A1(_03779_ ), .A2(\ID_EX_typ [1] ), .ZN(_04822_ ) );
AND2_X2 _12563_ ( .A1(_04822_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04823_ ) );
INV_X1 _12564_ ( .A(\ID_EX_typ [1] ), .ZN(_04824_ ) );
NOR2_X1 _12565_ ( .A1(_04824_ ), .A2(fanout_net_5 ), .ZN(_04825_ ) );
INV_X1 _12566_ ( .A(fanout_net_6 ), .ZN(_04826_ ) );
AND2_X2 _12567_ ( .A1(_04825_ ), .A2(_04826_ ), .ZN(_04827_ ) );
INV_X1 _12568_ ( .A(_04827_ ), .ZN(_04828_ ) );
AND2_X1 _12569_ ( .A1(_04001_ ), .A2(fanout_net_6 ), .ZN(_04829_ ) );
INV_X1 _12570_ ( .A(_04829_ ), .ZN(_04830_ ) );
OR2_X1 _12571_ ( .A1(_04316_ ), .A2(fanout_net_7 ), .ZN(_04831_ ) );
INV_X1 _12572_ ( .A(fanout_net_7 ), .ZN(_04832_ ) );
BUF_X4 _12573_ ( .A(_04832_ ), .Z(_04833_ ) );
BUF_X4 _12574_ ( .A(_04833_ ), .Z(_04834_ ) );
BUF_X2 _12575_ ( .A(_04834_ ), .Z(_04835_ ) );
OR2_X1 _12576_ ( .A1(_04835_ ), .A2(\ID_EX_imm [31] ), .ZN(_04836_ ) );
NAND2_X1 _12577_ ( .A1(_04831_ ), .A2(_04836_ ), .ZN(_04837_ ) );
INV_X1 _12578_ ( .A(_02928_ ), .ZN(_04838_ ) );
NAND2_X1 _12579_ ( .A1(_04837_ ), .A2(_04838_ ), .ZN(_04839_ ) );
NAND3_X1 _12580_ ( .A1(_04831_ ), .A2(_02928_ ), .A3(_04836_ ), .ZN(_04840_ ) );
NAND2_X1 _12581_ ( .A1(_04839_ ), .A2(_04840_ ), .ZN(_04841_ ) );
OR2_X1 _12582_ ( .A1(_04339_ ), .A2(fanout_net_7 ), .ZN(_04842_ ) );
NAND2_X1 _12583_ ( .A1(fanout_net_7 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04843_ ) );
AND3_X1 _12584_ ( .A1(_04842_ ), .A2(_04340_ ), .A3(_04843_ ), .ZN(_04844_ ) );
AOI21_X1 _12585_ ( .A(_04340_ ), .B1(_04842_ ), .B2(_04843_ ), .ZN(_04845_ ) );
OAI21_X1 _12586_ ( .A(_04841_ ), .B1(_04844_ ), .B2(_04845_ ), .ZN(_04846_ ) );
NAND3_X1 _12587_ ( .A1(_04270_ ), .A2(_04835_ ), .A3(_04289_ ), .ZN(_04847_ ) );
NAND2_X1 _12588_ ( .A1(fanout_net_7 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04848_ ) );
AND2_X1 _12589_ ( .A1(_04847_ ), .A2(_04848_ ), .ZN(_04849_ ) );
XNOR2_X1 _12590_ ( .A(_04849_ ), .B(_02900_ ), .ZN(_04850_ ) );
NAND3_X1 _12591_ ( .A1(_04245_ ), .A2(_04835_ ), .A3(_04267_ ), .ZN(_04851_ ) );
NAND2_X1 _12592_ ( .A1(fanout_net_7 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04852_ ) );
AND2_X2 _12593_ ( .A1(_04851_ ), .A2(_04852_ ), .ZN(_04853_ ) );
INV_X1 _12594_ ( .A(_02125_ ), .ZN(_04854_ ) );
XNOR2_X1 _12595_ ( .A(_04853_ ), .B(_04854_ ), .ZN(_04855_ ) );
NOR3_X1 _12596_ ( .A1(_04846_ ), .A2(_04850_ ), .A3(_04855_ ), .ZN(_04856_ ) );
OR2_X4 _12597_ ( .A1(_04050_ ), .A2(fanout_net_7 ), .ZN(_04857_ ) );
NAND2_X1 _12598_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [23] ), .ZN(_04858_ ) );
AND2_X4 _12599_ ( .A1(_04857_ ), .A2(_04858_ ), .ZN(_04859_ ) );
XNOR2_X2 _12600_ ( .A(_04859_ ), .B(_02179_ ), .ZN(_04860_ ) );
NAND3_X2 _12601_ ( .A1(_04091_ ), .A2(_04834_ ), .A3(_04111_ ), .ZN(_04861_ ) );
NAND2_X1 _12602_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [21] ), .ZN(_04862_ ) );
AND2_X4 _12603_ ( .A1(_04861_ ), .A2(_04862_ ), .ZN(_04863_ ) );
XNOR2_X2 _12604_ ( .A(_04863_ ), .B(_04113_ ), .ZN(_04864_ ) );
NAND3_X1 _12605_ ( .A1(_04054_ ), .A2(_04086_ ), .A3(_04834_ ), .ZN(_04865_ ) );
NAND2_X1 _12606_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [22] ), .ZN(_04866_ ) );
AND2_X4 _12607_ ( .A1(_04865_ ), .A2(_04866_ ), .ZN(_04867_ ) );
XNOR2_X2 _12608_ ( .A(_04867_ ), .B(_02155_ ), .ZN(_04868_ ) );
NOR3_X2 _12609_ ( .A1(_04860_ ), .A2(_04864_ ), .A3(_04868_ ), .ZN(_04869_ ) );
NAND3_X1 _12610_ ( .A1(_04116_ ), .A2(_04138_ ), .A3(_04834_ ), .ZN(_04870_ ) );
NAND2_X1 _12611_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [20] ), .ZN(_04871_ ) );
AND2_X4 _12612_ ( .A1(_04870_ ), .A2(_04871_ ), .ZN(_04872_ ) );
XNOR2_X1 _12613_ ( .A(_04872_ ), .B(_02202_ ), .ZN(_04873_ ) );
INV_X1 _12614_ ( .A(_04873_ ), .ZN(_04874_ ) );
NAND3_X1 _12615_ ( .A1(_04169_ ), .A2(_04188_ ), .A3(_04834_ ), .ZN(_04875_ ) );
NAND2_X1 _12616_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [18] ), .ZN(_04876_ ) );
AND2_X4 _12617_ ( .A1(_04875_ ), .A2(_04876_ ), .ZN(_04877_ ) );
XNOR2_X2 _12618_ ( .A(_04877_ ), .B(_02275_ ), .ZN(_04878_ ) );
NAND3_X2 _12619_ ( .A1(_04143_ ), .A2(_04834_ ), .A3(_04165_ ), .ZN(_04879_ ) );
NAND2_X1 _12620_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [19] ), .ZN(_04880_ ) );
AND2_X4 _12621_ ( .A1(_04879_ ), .A2(_04880_ ), .ZN(_04881_ ) );
XNOR2_X2 _12622_ ( .A(_04881_ ), .B(_02252_ ), .ZN(_04882_ ) );
NOR2_X1 _12623_ ( .A1(_04878_ ), .A2(_04882_ ), .ZN(_04883_ ) );
NAND3_X1 _12624_ ( .A1(_04869_ ), .A2(_04874_ ), .A3(_04883_ ), .ZN(_04884_ ) );
NAND3_X1 _12625_ ( .A1(_04220_ ), .A2(_04834_ ), .A3(_04239_ ), .ZN(_04885_ ) );
NAND2_X1 _12626_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [17] ), .ZN(_04886_ ) );
AND2_X4 _12627_ ( .A1(_04885_ ), .A2(_04886_ ), .ZN(_04887_ ) );
XNOR2_X2 _12628_ ( .A(_04887_ ), .B(_02299_ ), .ZN(_04888_ ) );
NAND3_X1 _12629_ ( .A1(_04193_ ), .A2(_04216_ ), .A3(_04835_ ), .ZN(_04889_ ) );
NAND2_X1 _12630_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [16] ), .ZN(_04890_ ) );
AND2_X4 _12631_ ( .A1(_04889_ ), .A2(_04890_ ), .ZN(_04891_ ) );
XNOR2_X1 _12632_ ( .A(_04891_ ), .B(_02322_ ), .ZN(_04892_ ) );
NOR3_X4 _12633_ ( .A1(_04884_ ), .A2(_04888_ ), .A3(_04892_ ), .ZN(_04893_ ) );
NAND2_X4 _12634_ ( .A1(_04628_ ), .A2(_04834_ ), .ZN(_04894_ ) );
NAND2_X1 _12635_ ( .A1(_02632_ ), .A2(fanout_net_7 ), .ZN(_04895_ ) );
NAND2_X4 _12636_ ( .A1(_04894_ ), .A2(_04895_ ), .ZN(_04896_ ) );
XNOR2_X2 _12637_ ( .A(_04896_ ), .B(_02631_ ), .ZN(_04897_ ) );
OR2_X4 _12638_ ( .A1(_04605_ ), .A2(fanout_net_7 ), .ZN(_04898_ ) );
NAND2_X1 _12639_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [15] ), .ZN(_04899_ ) );
AND2_X4 _12640_ ( .A1(_04898_ ), .A2(_04899_ ), .ZN(_04900_ ) );
NOR2_X4 _12641_ ( .A1(_04900_ ), .A2(_04606_ ), .ZN(_04901_ ) );
INV_X2 _12642_ ( .A(_04901_ ), .ZN(_04902_ ) );
NAND3_X1 _12643_ ( .A1(_04898_ ), .A2(_04606_ ), .A3(_04899_ ), .ZN(_04903_ ) );
AOI21_X4 _12644_ ( .A(_04897_ ), .B1(_04902_ ), .B2(_04903_ ), .ZN(_04904_ ) );
NAND3_X1 _12645_ ( .A1(_04536_ ), .A2(_04555_ ), .A3(_04834_ ), .ZN(_04905_ ) );
NAND2_X1 _12646_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [12] ), .ZN(_04906_ ) );
AND2_X4 _12647_ ( .A1(_04905_ ), .A2(_04906_ ), .ZN(_04907_ ) );
XNOR2_X2 _12648_ ( .A(_04907_ ), .B(_02560_ ), .ZN(_04908_ ) );
INV_X1 _12649_ ( .A(_04908_ ), .ZN(_04909_ ) );
NAND2_X4 _12650_ ( .A1(_04904_ ), .A2(_04909_ ), .ZN(_04910_ ) );
AOI21_X2 _12651_ ( .A(fanout_net_7 ), .B1(_04558_ ), .B2(_04577_ ), .ZN(_04911_ ) );
NOR2_X1 _12652_ ( .A1(_04833_ ), .A2(\ID_EX_imm [13] ), .ZN(_04912_ ) );
NOR2_X4 _12653_ ( .A1(_04911_ ), .A2(_04912_ ), .ZN(_04913_ ) );
INV_X1 _12654_ ( .A(_04579_ ), .ZN(_04914_ ) );
XNOR2_X2 _12655_ ( .A(_04913_ ), .B(_04914_ ), .ZN(_04915_ ) );
NOR2_X4 _12656_ ( .A1(_04910_ ), .A2(_04915_ ), .ZN(_04916_ ) );
NAND3_X1 _12657_ ( .A1(_04655_ ), .A2(_04674_ ), .A3(_04833_ ), .ZN(_04917_ ) );
NAND2_X1 _12658_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [10] ), .ZN(_04918_ ) );
AND2_X2 _12659_ ( .A1(_04917_ ), .A2(_04918_ ), .ZN(_04919_ ) );
XNOR2_X2 _12660_ ( .A(_04919_ ), .B(_02724_ ), .ZN(_04920_ ) );
NAND3_X1 _12661_ ( .A1(_04632_ ), .A2(_04833_ ), .A3(_04651_ ), .ZN(_04921_ ) );
NAND2_X1 _12662_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [11] ), .ZN(_04922_ ) );
AND2_X4 _12663_ ( .A1(_04921_ ), .A2(_04922_ ), .ZN(_04923_ ) );
XNOR2_X2 _12664_ ( .A(_04923_ ), .B(_02702_ ), .ZN(_04924_ ) );
NOR2_X4 _12665_ ( .A1(_04920_ ), .A2(_04924_ ), .ZN(_04925_ ) );
NAND3_X1 _12666_ ( .A1(_04702_ ), .A2(_04833_ ), .A3(_04721_ ), .ZN(_04926_ ) );
NAND2_X1 _12667_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [9] ), .ZN(_04927_ ) );
AND2_X4 _12668_ ( .A1(_04926_ ), .A2(_04927_ ), .ZN(_04928_ ) );
XNOR2_X2 _12669_ ( .A(_04928_ ), .B(_02678_ ), .ZN(_04929_ ) );
INV_X2 _12670_ ( .A(_04929_ ), .ZN(_04930_ ) );
NAND3_X1 _12671_ ( .A1(_04679_ ), .A2(_04834_ ), .A3(_04698_ ), .ZN(_04931_ ) );
NAND2_X1 _12672_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [8] ), .ZN(_04932_ ) );
AND2_X4 _12673_ ( .A1(_04931_ ), .A2(_04932_ ), .ZN(_04933_ ) );
XNOR2_X1 _12674_ ( .A(_04933_ ), .B(_02655_ ), .ZN(_04934_ ) );
INV_X1 _12675_ ( .A(_04934_ ), .ZN(_04935_ ) );
NAND4_X4 _12676_ ( .A1(_04916_ ), .A2(_04925_ ), .A3(_04930_ ), .A4(_04935_ ), .ZN(_04936_ ) );
OAI21_X2 _12677_ ( .A(_04833_ ), .B1(_04531_ ), .B2(_04532_ ), .ZN(_04937_ ) );
NAND2_X1 _12678_ ( .A1(fanout_net_7 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_04938_ ) );
AND2_X4 _12679_ ( .A1(_04937_ ), .A2(_04938_ ), .ZN(_04939_ ) );
INV_X1 _12680_ ( .A(_02352_ ), .ZN(_04940_ ) );
XNOR2_X2 _12681_ ( .A(_04939_ ), .B(_04940_ ), .ZN(_04941_ ) );
INV_X1 _12682_ ( .A(_04941_ ), .ZN(_04942_ ) );
NAND2_X4 _12683_ ( .A1(_04458_ ), .A2(_04832_ ), .ZN(_04943_ ) );
NAND2_X1 _12684_ ( .A1(_02400_ ), .A2(fanout_net_7 ), .ZN(_04944_ ) );
NAND2_X1 _12685_ ( .A1(_04943_ ), .A2(_04944_ ), .ZN(_04945_ ) );
NAND2_X1 _12686_ ( .A1(_04945_ ), .A2(_02399_ ), .ZN(_04946_ ) );
AND3_X4 _12687_ ( .A1(_04943_ ), .A2(_02399_ ), .A3(_04944_ ), .ZN(_04947_ ) );
AOI21_X4 _12688_ ( .A(_02399_ ), .B1(_04943_ ), .B2(_04944_ ), .ZN(_04948_ ) );
NOR2_X2 _12689_ ( .A1(_04947_ ), .A2(_04948_ ), .ZN(_04949_ ) );
INV_X1 _12690_ ( .A(_04486_ ), .ZN(_04950_ ) );
NAND3_X4 _12691_ ( .A1(_04464_ ), .A2(_04832_ ), .A3(_04484_ ), .ZN(_04951_ ) );
OR2_X1 _12692_ ( .A1(_04832_ ), .A2(\ID_EX_imm [0] ), .ZN(_04952_ ) );
AND3_X1 _12693_ ( .A1(_04950_ ), .A2(_04951_ ), .A3(_04952_ ), .ZN(_04953_ ) );
OAI21_X1 _12694_ ( .A(_04946_ ), .B1(_04949_ ), .B2(_04953_ ), .ZN(_04954_ ) );
NAND3_X1 _12695_ ( .A1(_04489_ ), .A2(_04833_ ), .A3(_04509_ ), .ZN(_04955_ ) );
NAND2_X1 _12696_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [2] ), .ZN(_04956_ ) );
AND2_X4 _12697_ ( .A1(_04955_ ), .A2(_04956_ ), .ZN(_04957_ ) );
XNOR2_X1 _12698_ ( .A(_04957_ ), .B(_02376_ ), .ZN(_04958_ ) );
INV_X2 _12699_ ( .A(_04958_ ), .ZN(_04959_ ) );
AND3_X2 _12700_ ( .A1(_04942_ ), .A2(_04954_ ), .A3(_04959_ ), .ZN(_04960_ ) );
INV_X1 _12701_ ( .A(_04957_ ), .ZN(_04961_ ) );
NOR3_X1 _12702_ ( .A1(_04941_ ), .A2(_04511_ ), .A3(_04961_ ), .ZN(_04962_ ) );
AOI21_X1 _12703_ ( .A(_04940_ ), .B1(_04937_ ), .B2(_04938_ ), .ZN(_04963_ ) );
OR3_X4 _12704_ ( .A1(_04960_ ), .A2(_04962_ ), .A3(_04963_ ), .ZN(_04964_ ) );
NAND3_X1 _12705_ ( .A1(_04752_ ), .A2(_04771_ ), .A3(_04833_ ), .ZN(_04965_ ) );
NAND2_X1 _12706_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [6] ), .ZN(_04966_ ) );
AND2_X4 _12707_ ( .A1(_04965_ ), .A2(_04966_ ), .ZN(_04967_ ) );
XNOR2_X2 _12708_ ( .A(_04967_ ), .B(_02530_ ), .ZN(_04968_ ) );
OR2_X4 _12709_ ( .A1(_04748_ ), .A2(fanout_net_7 ), .ZN(_04969_ ) );
NAND2_X1 _12710_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [7] ), .ZN(_04970_ ) );
AND2_X1 _12711_ ( .A1(_04969_ ), .A2(_04970_ ), .ZN(_04971_ ) );
OR2_X2 _12712_ ( .A1(_04971_ ), .A2(_04749_ ), .ZN(_04972_ ) );
NAND3_X1 _12713_ ( .A1(_04969_ ), .A2(_04749_ ), .A3(_04970_ ), .ZN(_04973_ ) );
AOI21_X1 _12714_ ( .A(_04968_ ), .B1(_04972_ ), .B2(_04973_ ), .ZN(_04974_ ) );
NAND2_X2 _12715_ ( .A1(_04795_ ), .A2(_04833_ ), .ZN(_04975_ ) );
NAND2_X1 _12716_ ( .A1(_02535_ ), .A2(\ID_EX_typ [4] ), .ZN(_04976_ ) );
NAND2_X4 _12717_ ( .A1(_04975_ ), .A2(_04976_ ), .ZN(_04977_ ) );
INV_X1 _12718_ ( .A(_02525_ ), .ZN(_04978_ ) );
XNOR2_X2 _12719_ ( .A(_04977_ ), .B(_04978_ ), .ZN(_04979_ ) );
INV_X2 _12720_ ( .A(_04979_ ), .ZN(_04980_ ) );
NAND3_X1 _12721_ ( .A1(_04797_ ), .A2(_04816_ ), .A3(_04833_ ), .ZN(_04981_ ) );
NAND2_X1 _12722_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [4] ), .ZN(_04982_ ) );
AND2_X2 _12723_ ( .A1(_04981_ ), .A2(_04982_ ), .ZN(_04983_ ) );
BUF_X8 _12724_ ( .A(_04983_ ), .Z(_04984_ ) );
XNOR2_X1 _12725_ ( .A(_04984_ ), .B(_02452_ ), .ZN(_04985_ ) );
INV_X1 _12726_ ( .A(_04985_ ), .ZN(_04986_ ) );
NAND4_X1 _12727_ ( .A1(_04964_ ), .A2(_04974_ ), .A3(_04980_ ), .A4(_04986_ ), .ZN(_04987_ ) );
INV_X1 _12728_ ( .A(_02530_ ), .ZN(_04988_ ) );
INV_X1 _12729_ ( .A(_04967_ ), .ZN(_04989_ ) );
AOI211_X1 _12730_ ( .A(_04988_ ), .B(_04989_ ), .C1(_04972_ ), .C2(_04973_ ), .ZN(_04990_ ) );
NAND3_X1 _12731_ ( .A1(_04980_ ), .A2(_02452_ ), .A3(_04984_ ), .ZN(_04991_ ) );
OAI21_X1 _12732_ ( .A(_04991_ ), .B1(_04978_ ), .B2(_04977_ ), .ZN(_04992_ ) );
AOI221_X1 _12733_ ( .A(_04990_ ), .B1(_02477_ ), .B2(_04971_ ), .C1(_04974_ ), .C2(_04992_ ), .ZN(_04993_ ) );
AOI21_X2 _12734_ ( .A(_04936_ ), .B1(_04987_ ), .B2(_04993_ ), .ZN(_04994_ ) );
INV_X1 _12735_ ( .A(_04925_ ), .ZN(_04995_ ) );
NAND3_X1 _12736_ ( .A1(_04926_ ), .A2(_02678_ ), .A3(_04927_ ), .ZN(_04996_ ) );
NAND3_X1 _12737_ ( .A1(_04930_ ), .A2(_02655_ ), .A3(_04933_ ), .ZN(_04997_ ) );
AOI21_X1 _12738_ ( .A(_04995_ ), .B1(_04996_ ), .B2(_04997_ ), .ZN(_04998_ ) );
AND3_X1 _12739_ ( .A1(_04921_ ), .A2(_02702_ ), .A3(_04922_ ), .ZN(_04999_ ) );
OR2_X2 _12740_ ( .A1(_04998_ ), .A2(_04999_ ), .ZN(_05000_ ) );
INV_X1 _12741_ ( .A(_04919_ ), .ZN(_05001_ ) );
NOR3_X1 _12742_ ( .A1(_04924_ ), .A2(_04676_ ), .A3(_05001_ ), .ZN(_05002_ ) );
OAI21_X1 _12743_ ( .A(_04916_ ), .B1(_05000_ ), .B2(_05002_ ), .ZN(_05003_ ) );
NOR2_X1 _12744_ ( .A1(_04913_ ), .A2(_04914_ ), .ZN(_05004_ ) );
INV_X1 _12745_ ( .A(_02561_ ), .ZN(_05005_ ) );
INV_X1 _12746_ ( .A(_04907_ ), .ZN(_05006_ ) );
NOR3_X1 _12747_ ( .A1(_04915_ ), .A2(_05005_ ), .A3(_05006_ ), .ZN(_05007_ ) );
OAI21_X1 _12748_ ( .A(_04904_ ), .B1(_05004_ ), .B2(_05007_ ), .ZN(_05008_ ) );
XNOR2_X1 _12749_ ( .A(_04900_ ), .B(_02609_ ), .ZN(_05009_ ) );
NAND2_X1 _12750_ ( .A1(_04896_ ), .A2(_02631_ ), .ZN(_05010_ ) );
OR2_X1 _12751_ ( .A1(_05009_ ), .A2(_05010_ ), .ZN(_05011_ ) );
NAND3_X1 _12752_ ( .A1(_04898_ ), .A2(_02609_ ), .A3(_04899_ ), .ZN(_05012_ ) );
NAND4_X1 _12753_ ( .A1(_05003_ ), .A2(_05008_ ), .A3(_05011_ ), .A4(_05012_ ), .ZN(_05013_ ) );
OAI21_X1 _12754_ ( .A(_04893_ ), .B1(_04994_ ), .B2(_05013_ ), .ZN(_05014_ ) );
INV_X1 _12755_ ( .A(_04860_ ), .ZN(_05015_ ) );
NAND3_X1 _12756_ ( .A1(_05015_ ), .A2(_02155_ ), .A3(_04867_ ), .ZN(_05016_ ) );
INV_X1 _12757_ ( .A(_04888_ ), .ZN(_05017_ ) );
AND3_X2 _12758_ ( .A1(_05017_ ), .A2(_02322_ ), .A3(_04891_ ), .ZN(_05018_ ) );
AND3_X1 _12759_ ( .A1(_04885_ ), .A2(_02299_ ), .A3(_04886_ ), .ZN(_05019_ ) );
OAI21_X1 _12760_ ( .A(_04883_ ), .B1(_05018_ ), .B2(_05019_ ), .ZN(_05020_ ) );
INV_X1 _12761_ ( .A(_04882_ ), .ZN(_05021_ ) );
NAND3_X1 _12762_ ( .A1(_05021_ ), .A2(_02275_ ), .A3(_04877_ ), .ZN(_05022_ ) );
NAND3_X1 _12763_ ( .A1(_04879_ ), .A2(_02252_ ), .A3(_04880_ ), .ZN(_05023_ ) );
NAND3_X1 _12764_ ( .A1(_05020_ ), .A2(_05022_ ), .A3(_05023_ ), .ZN(_05024_ ) );
NAND3_X1 _12765_ ( .A1(_05024_ ), .A2(_04874_ ), .A3(_04869_ ), .ZN(_05025_ ) );
AND2_X1 _12766_ ( .A1(_04863_ ), .A2(_04114_ ), .ZN(_05026_ ) );
NOR2_X1 _12767_ ( .A1(_04863_ ), .A2(_04114_ ), .ZN(_05027_ ) );
OAI211_X1 _12768_ ( .A(_02202_ ), .B(_04872_ ), .C1(_05026_ ), .C2(_05027_ ), .ZN(_05028_ ) );
NAND3_X1 _12769_ ( .A1(_04861_ ), .A2(_04113_ ), .A3(_04862_ ), .ZN(_05029_ ) );
AND2_X1 _12770_ ( .A1(_05028_ ), .A2(_05029_ ), .ZN(_05030_ ) );
NOR3_X1 _12771_ ( .A1(_05030_ ), .A2(_04860_ ), .A3(_04868_ ), .ZN(_05031_ ) );
AOI21_X1 _12772_ ( .A(_05031_ ), .B1(_02179_ ), .B2(_04859_ ), .ZN(_05032_ ) );
NAND4_X1 _12773_ ( .A1(_05014_ ), .A2(_05016_ ), .A3(_05025_ ), .A4(_05032_ ), .ZN(_05033_ ) );
NAND3_X1 _12774_ ( .A1(_04360_ ), .A2(_04362_ ), .A3(_04835_ ), .ZN(_05034_ ) );
NAND2_X1 _12775_ ( .A1(_02819_ ), .A2(\ID_EX_typ [4] ), .ZN(_05035_ ) );
NAND2_X1 _12776_ ( .A1(_05034_ ), .A2(_05035_ ), .ZN(_05036_ ) );
INV_X1 _12777_ ( .A(_04364_ ), .ZN(_05037_ ) );
NOR2_X1 _12778_ ( .A1(_05036_ ), .A2(_05037_ ), .ZN(_05038_ ) );
AOI21_X1 _12779_ ( .A(_04364_ ), .B1(_05034_ ), .B2(_05035_ ), .ZN(_05039_ ) );
NOR2_X1 _12780_ ( .A1(_05038_ ), .A2(_05039_ ), .ZN(_05040_ ) );
NAND3_X1 _12781_ ( .A1(_04366_ ), .A2(_04835_ ), .A3(_04385_ ), .ZN(_05041_ ) );
NAND2_X1 _12782_ ( .A1(_02865_ ), .A2(\ID_EX_typ [4] ), .ZN(_05042_ ) );
NAND2_X1 _12783_ ( .A1(_05041_ ), .A2(_05042_ ), .ZN(_05043_ ) );
INV_X1 _12784_ ( .A(_02864_ ), .ZN(_05044_ ) );
NOR2_X1 _12785_ ( .A1(_05043_ ), .A2(_05044_ ), .ZN(_05045_ ) );
AOI21_X1 _12786_ ( .A(_02864_ ), .B1(_05041_ ), .B2(_05042_ ), .ZN(_05046_ ) );
NOR2_X1 _12787_ ( .A1(_05045_ ), .A2(_05046_ ), .ZN(_05047_ ) );
NOR2_X1 _12788_ ( .A1(_05040_ ), .A2(_05047_ ), .ZN(_05048_ ) );
NAND3_X1 _12789_ ( .A1(_04389_ ), .A2(_04835_ ), .A3(_04408_ ), .ZN(_05049_ ) );
NAND2_X1 _12790_ ( .A1(_02788_ ), .A2(\ID_EX_typ [4] ), .ZN(_05050_ ) );
NAND2_X1 _12791_ ( .A1(_05049_ ), .A2(_05050_ ), .ZN(_05051_ ) );
INV_X1 _12792_ ( .A(_02787_ ), .ZN(_05052_ ) );
NOR2_X1 _12793_ ( .A1(_05051_ ), .A2(_05052_ ), .ZN(_05053_ ) );
AOI21_X1 _12794_ ( .A(_02787_ ), .B1(_05049_ ), .B2(_05050_ ), .ZN(_05054_ ) );
NOR2_X1 _12795_ ( .A1(_05053_ ), .A2(_05054_ ), .ZN(_05055_ ) );
INV_X1 _12796_ ( .A(_05055_ ), .ZN(_05056_ ) );
NAND3_X1 _12797_ ( .A1(_04412_ ), .A2(_04835_ ), .A3(_04431_ ), .ZN(_05057_ ) );
NAND2_X1 _12798_ ( .A1(_02867_ ), .A2(\ID_EX_typ [4] ), .ZN(_05058_ ) );
NAND2_X1 _12799_ ( .A1(_05057_ ), .A2(_05058_ ), .ZN(_05059_ ) );
XNOR2_X1 _12800_ ( .A(_05059_ ), .B(_02814_ ), .ZN(_05060_ ) );
INV_X1 _12801_ ( .A(_05060_ ), .ZN(_05061_ ) );
AND4_X2 _12802_ ( .A1(_05033_ ), .A2(_05048_ ), .A3(_05056_ ), .A4(_05061_ ), .ZN(_05062_ ) );
INV_X1 _12803_ ( .A(_05051_ ), .ZN(_05063_ ) );
NOR3_X1 _12804_ ( .A1(_05060_ ), .A2(_05052_ ), .A3(_05063_ ), .ZN(_05064_ ) );
AOI22_X1 _12805_ ( .A1(_05057_ ), .A2(_05058_ ), .B1(_02793_ ), .B2(_02813_ ), .ZN(_05065_ ) );
OAI21_X1 _12806_ ( .A(_05048_ ), .B1(_05064_ ), .B2(_05065_ ), .ZN(_05066_ ) );
INV_X1 _12807_ ( .A(_05040_ ), .ZN(_05067_ ) );
NAND3_X1 _12808_ ( .A1(_05067_ ), .A2(_02864_ ), .A3(_05043_ ), .ZN(_05068_ ) );
NAND2_X1 _12809_ ( .A1(_05036_ ), .A2(_04364_ ), .ZN(_05069_ ) );
NAND3_X1 _12810_ ( .A1(_05066_ ), .A2(_05068_ ), .A3(_05069_ ), .ZN(_05070_ ) );
OAI21_X2 _12811_ ( .A(_04856_ ), .B1(_05062_ ), .B2(_05070_ ), .ZN(_05071_ ) );
AND3_X1 _12812_ ( .A1(_04831_ ), .A2(_04838_ ), .A3(_04836_ ), .ZN(_05072_ ) );
AOI21_X1 _12813_ ( .A(_02090_ ), .B1(_04842_ ), .B2(_04843_ ), .ZN(_05073_ ) );
AND2_X1 _12814_ ( .A1(_04841_ ), .A2(_05073_ ), .ZN(_05074_ ) );
AOI21_X1 _12815_ ( .A(_04854_ ), .B1(_04851_ ), .B2(_04852_ ), .ZN(_05075_ ) );
AND2_X1 _12816_ ( .A1(_04849_ ), .A2(_02894_ ), .ZN(_05076_ ) );
AOI21_X1 _12817_ ( .A(_02894_ ), .B1(_04847_ ), .B2(_04848_ ), .ZN(_05077_ ) );
OAI21_X1 _12818_ ( .A(_05075_ ), .B1(_05076_ ), .B2(_05077_ ), .ZN(_05078_ ) );
OAI21_X1 _12819_ ( .A(_05078_ ), .B1(_02900_ ), .B2(_04849_ ), .ZN(_05079_ ) );
NOR2_X1 _12820_ ( .A1(_04844_ ), .A2(_04845_ ), .ZN(_05080_ ) );
AOI21_X1 _12821_ ( .A(_04838_ ), .B1(_04831_ ), .B2(_04836_ ), .ZN(_05081_ ) );
NOR3_X1 _12822_ ( .A1(_05080_ ), .A2(_05072_ ), .A3(_05081_ ), .ZN(_05082_ ) );
AOI211_X1 _12823_ ( .A(_05072_ ), .B(_05074_ ), .C1(_05079_ ), .C2(_05082_ ), .ZN(_05083_ ) );
AND2_X2 _12824_ ( .A1(_05071_ ), .A2(_05083_ ), .ZN(_05084_ ) );
MUX2_X1 _12825_ ( .A(_04828_ ), .B(_04830_ ), .S(_05084_ ), .Z(_05085_ ) );
AND3_X1 _12826_ ( .A1(_04607_ ), .A2(_02631_ ), .A3(_04628_ ), .ZN(_05086_ ) );
AND2_X1 _12827_ ( .A1(_04722_ ), .A2(_02678_ ), .ZN(_05087_ ) );
AND3_X2 _12828_ ( .A1(_04724_ ), .A2(_02655_ ), .A3(_04699_ ), .ZN(_05088_ ) );
OAI21_X1 _12829_ ( .A(_04678_ ), .B1(_05087_ ), .B2(_05088_ ), .ZN(_05089_ ) );
AND2_X1 _12830_ ( .A1(_04675_ ), .A2(_02724_ ), .ZN(_05090_ ) );
AND2_X2 _12831_ ( .A1(_04654_ ), .A2(_05090_ ), .ZN(_05091_ ) );
AOI21_X1 _12832_ ( .A(_05091_ ), .B1(_02702_ ), .B2(_04652_ ), .ZN(_05092_ ) );
AND2_X2 _12833_ ( .A1(_05089_ ), .A2(_05092_ ), .ZN(_05093_ ) );
INV_X1 _12834_ ( .A(_05093_ ), .ZN(_05094_ ) );
AND2_X2 _12835_ ( .A1(_05094_ ), .A2(_04631_ ), .ZN(_05095_ ) );
NAND2_X1 _12836_ ( .A1(_04556_ ), .A2(_02561_ ), .ZN(_05096_ ) );
NOR3_X1 _12837_ ( .A1(_04580_ ), .A2(_04581_ ), .A3(_05096_ ), .ZN(_05097_ ) );
OR2_X1 _12838_ ( .A1(_05097_ ), .A2(_04580_ ), .ZN(_05098_ ) );
AND3_X1 _12839_ ( .A1(_05098_ ), .A2(_04607_ ), .A3(_04630_ ), .ZN(_05099_ ) );
OR2_X4 _12840_ ( .A1(_05095_ ), .A2(_05099_ ), .ZN(_05100_ ) );
AOI211_X1 _12841_ ( .A(_05086_ ), .B(_05100_ ), .C1(_02609_ ), .C2(_04605_ ), .ZN(_05101_ ) );
AOI21_X1 _12842_ ( .A(_04486_ ), .B1(_04484_ ), .B2(_04464_ ), .ZN(_05102_ ) );
OAI21_X1 _12843_ ( .A(_04459_ ), .B1(_04462_ ), .B2(_05102_ ), .ZN(_05103_ ) );
NAND2_X1 _12844_ ( .A1(_05103_ ), .A2(_04512_ ), .ZN(_05104_ ) );
AOI21_X1 _12845_ ( .A(_04511_ ), .B1(_04489_ ), .B2(_04509_ ), .ZN(_05105_ ) );
INV_X1 _12846_ ( .A(_05105_ ), .ZN(_05106_ ) );
OAI211_X1 _12847_ ( .A(_05104_ ), .B(_05106_ ), .C1(_04940_ ), .C2(_04533_ ), .ZN(_05107_ ) );
NAND2_X1 _12848_ ( .A1(_04940_ ), .A2(_04533_ ), .ZN(_05108_ ) );
AND2_X1 _12849_ ( .A1(_04774_ ), .A2(_04819_ ), .ZN(_05109_ ) );
NAND3_X1 _12850_ ( .A1(_05107_ ), .A2(_05108_ ), .A3(_05109_ ), .ZN(_05110_ ) );
AND3_X1 _12851_ ( .A1(_04750_ ), .A2(_02530_ ), .A3(_04772_ ), .ZN(_05111_ ) );
NAND3_X1 _12852_ ( .A1(_04796_ ), .A2(_02452_ ), .A3(_04817_ ), .ZN(_05112_ ) );
OAI21_X1 _12853_ ( .A(_05112_ ), .B1(_04978_ ), .B2(_04795_ ), .ZN(_05113_ ) );
AOI221_X4 _12854_ ( .A(_05111_ ), .B1(_02477_ ), .B2(_04748_ ), .C1(_05113_ ), .C2(_04774_ ), .ZN(_05114_ ) );
AND2_X1 _12855_ ( .A1(_05110_ ), .A2(_05114_ ), .ZN(_05115_ ) );
INV_X1 _12856_ ( .A(_05115_ ), .ZN(_05116_ ) );
NAND3_X1 _12857_ ( .A1(_05116_ ), .A2(_04631_ ), .A3(_04725_ ), .ZN(_05117_ ) );
AND2_X1 _12858_ ( .A1(_05101_ ), .A2(_05117_ ), .ZN(_05118_ ) );
INV_X1 _12859_ ( .A(_04437_ ), .ZN(_05119_ ) );
OR2_X2 _12860_ ( .A1(_05118_ ), .A2(_05119_ ), .ZN(_05120_ ) );
NOR2_X1 _12861_ ( .A1(_04112_ ), .A2(_04113_ ), .ZN(_05121_ ) );
AND2_X1 _12862_ ( .A1(_04112_ ), .A2(_04113_ ), .ZN(_05122_ ) );
INV_X1 _12863_ ( .A(_05122_ ), .ZN(_05123_ ) );
NAND2_X1 _12864_ ( .A1(_04139_ ), .A2(_02202_ ), .ZN(_05124_ ) );
AOI21_X1 _12865_ ( .A(_05121_ ), .B1(_05123_ ), .B2(_05124_ ), .ZN(_05125_ ) );
NAND3_X1 _12866_ ( .A1(_05125_ ), .A2(_04052_ ), .A3(_04089_ ), .ZN(_05126_ ) );
NOR2_X1 _12867_ ( .A1(_04240_ ), .A2(_02299_ ), .ZN(_05127_ ) );
AND2_X1 _12868_ ( .A1(_04240_ ), .A2(_02299_ ), .ZN(_05128_ ) );
INV_X1 _12869_ ( .A(_05128_ ), .ZN(_05129_ ) );
NAND2_X1 _12870_ ( .A1(_04217_ ), .A2(_02322_ ), .ZN(_05130_ ) );
AOI21_X1 _12871_ ( .A(_05127_ ), .B1(_05129_ ), .B2(_05130_ ), .ZN(_05131_ ) );
AND3_X1 _12872_ ( .A1(_05131_ ), .A2(_04168_ ), .A3(_04191_ ), .ZN(_05132_ ) );
AOI21_X1 _12873_ ( .A(_04167_ ), .B1(_04143_ ), .B2(_04165_ ), .ZN(_05133_ ) );
AND3_X1 _12874_ ( .A1(_04168_ ), .A2(_02275_ ), .A3(_04189_ ), .ZN(_05134_ ) );
NOR3_X4 _12875_ ( .A1(_05132_ ), .A2(_05133_ ), .A3(_05134_ ), .ZN(_05135_ ) );
INV_X1 _12876_ ( .A(_04142_ ), .ZN(_05136_ ) );
OAI21_X1 _12877_ ( .A(_05126_ ), .B1(_05135_ ), .B2(_05136_ ), .ZN(_05137_ ) );
AND3_X1 _12878_ ( .A1(_02179_ ), .A2(_04049_ ), .A3(_04016_ ), .ZN(_05138_ ) );
AND3_X1 _12879_ ( .A1(_04052_ ), .A2(_02155_ ), .A3(_04087_ ), .ZN(_05139_ ) );
NOR3_X2 _12880_ ( .A1(_05137_ ), .A2(_05138_ ), .A3(_05139_ ), .ZN(_05140_ ) );
INV_X1 _12881_ ( .A(_04436_ ), .ZN(_05141_ ) );
NOR2_X1 _12882_ ( .A1(_05140_ ), .A2(_05141_ ), .ZN(_05142_ ) );
NOR2_X1 _12883_ ( .A1(_04386_ ), .A2(_05044_ ), .ZN(_05143_ ) );
NAND2_X1 _12884_ ( .A1(_04365_ ), .A2(_05143_ ), .ZN(_05144_ ) );
OAI21_X1 _12885_ ( .A(_05144_ ), .B1(_05037_ ), .B2(_04363_ ), .ZN(_05145_ ) );
AND3_X1 _12886_ ( .A1(_02815_ ), .A2(_04412_ ), .A3(_04431_ ), .ZN(_05146_ ) );
NOR2_X1 _12887_ ( .A1(_04409_ ), .A2(_05052_ ), .ZN(_05147_ ) );
AOI21_X1 _12888_ ( .A(_05146_ ), .B1(_04433_ ), .B2(_05147_ ), .ZN(_05148_ ) );
INV_X1 _12889_ ( .A(_05148_ ), .ZN(_05149_ ) );
AOI21_X1 _12890_ ( .A(_05145_ ), .B1(_04388_ ), .B2(_05149_ ), .ZN(_05150_ ) );
INV_X1 _12891_ ( .A(_04342_ ), .ZN(_05151_ ) );
NOR2_X1 _12892_ ( .A1(_05150_ ), .A2(_05151_ ), .ZN(_05152_ ) );
NOR2_X1 _12893_ ( .A1(_04268_ ), .A2(_04854_ ), .ZN(_05153_ ) );
NAND2_X1 _12894_ ( .A1(_04291_ ), .A2(_05153_ ), .ZN(_05154_ ) );
NOR2_X1 _12895_ ( .A1(_04290_ ), .A2(_02900_ ), .ZN(_05155_ ) );
INV_X1 _12896_ ( .A(_05155_ ), .ZN(_05156_ ) );
NAND2_X1 _12897_ ( .A1(_05154_ ), .A2(_05156_ ), .ZN(_05157_ ) );
AND3_X1 _12898_ ( .A1(_05157_ ), .A2(_04317_ ), .A3(_04341_ ), .ZN(_05158_ ) );
NOR2_X1 _12899_ ( .A1(_04339_ ), .A2(_02090_ ), .ZN(_05159_ ) );
NAND2_X1 _12900_ ( .A1(_04317_ ), .A2(_05159_ ), .ZN(_05160_ ) );
OAI21_X1 _12901_ ( .A(_05160_ ), .B1(_04838_ ), .B2(_04316_ ), .ZN(_05161_ ) );
NOR4_X4 _12902_ ( .A1(_05142_ ), .A2(_05152_ ), .A3(_05158_ ), .A4(_05161_ ), .ZN(_05162_ ) );
AND2_X2 _12903_ ( .A1(_04822_ ), .A2(fanout_net_6 ), .ZN(_05163_ ) );
AND3_X1 _12904_ ( .A1(_05120_ ), .A2(_05162_ ), .A3(_05163_ ), .ZN(_05164_ ) );
AND2_X1 _12905_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_5 ), .ZN(_05165_ ) );
AND2_X2 _12906_ ( .A1(_05165_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05166_ ) );
INV_X1 _12907_ ( .A(_05166_ ), .ZN(_05167_ ) );
AOI21_X1 _12908_ ( .A(_05167_ ), .B1(_05120_ ), .B2(_05162_ ), .ZN(_05168_ ) );
NOR3_X2 _12909_ ( .A1(_05164_ ), .A2(_05168_ ), .A3(_04823_ ), .ZN(_05169_ ) );
AOI221_X2 _12910_ ( .A(_04002_ ), .B1(_04821_ ), .B2(_04823_ ), .C1(_05085_ ), .C2(_05169_ ), .ZN(_05170_ ) );
INV_X1 _12911_ ( .A(_04002_ ), .ZN(_05171_ ) );
AND4_X1 _12912_ ( .A1(_04631_ ), .A2(_05109_ ), .A3(_04725_ ), .A4(_04535_ ), .ZN(_05172_ ) );
AOI21_X1 _12913_ ( .A(_05171_ ), .B1(_04437_ ), .B2(_05172_ ), .ZN(_05173_ ) );
NOR2_X4 _12914_ ( .A1(_05170_ ), .A2(_05173_ ), .ZN(_05174_ ) );
BUF_X8 _12915_ ( .A(_05174_ ), .Z(_05175_ ) );
MUX2_X1 _12916_ ( .A(_03891_ ), .B(_04000_ ), .S(_05175_ ), .Z(_05176_ ) );
INV_X1 _12917_ ( .A(\ID_EX_typ [3] ), .ZN(_05177_ ) );
BUF_X4 _12918_ ( .A(_05177_ ), .Z(_05178_ ) );
MUX2_X2 _12919_ ( .A(_03872_ ), .B(_05176_ ), .S(_05178_ ), .Z(_05179_ ) );
INV_X2 _12920_ ( .A(_03777_ ), .ZN(_05180_ ) );
BUF_X4 _12921_ ( .A(_05180_ ), .Z(_05181_ ) );
BUF_X4 _12922_ ( .A(_05181_ ), .Z(_05182_ ) );
NAND2_X1 _12923_ ( .A1(_05179_ ), .A2(_05182_ ), .ZN(_05183_ ) );
BUF_X2 _12924_ ( .A(_03778_ ), .Z(_05184_ ) );
OAI21_X1 _12925_ ( .A(_05184_ ), .B1(_04000_ ), .B2(fanout_net_5 ), .ZN(_05185_ ) );
BUF_X4 _12926_ ( .A(_03779_ ), .Z(_05186_ ) );
AOI21_X1 _12927_ ( .A(_05186_ ), .B1(_02933_ ), .B2(_02902_ ), .ZN(_05187_ ) );
OR2_X1 _12928_ ( .A1(_05185_ ), .A2(_05187_ ), .ZN(_05188_ ) );
AOI21_X1 _12929_ ( .A(_03801_ ), .B1(_05183_ ), .B2(_05188_ ), .ZN(_00122_ ) );
BUF_X4 _12930_ ( .A(_05177_ ), .Z(_05189_ ) );
AND4_X1 _12931_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_05190_ ) );
AND4_X1 _12932_ ( .A1(\ID_EX_pc [13] ), .A2(_05190_ ), .A3(\ID_EX_pc [12] ), .A4(_03880_ ), .ZN(_05191_ ) );
AND2_X2 _12933_ ( .A1(_03879_ ), .A2(_05191_ ), .ZN(_05192_ ) );
AND4_X1 _12934_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_05193_ ) );
AND2_X1 _12935_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_05194_ ) );
AND4_X1 _12936_ ( .A1(\ID_EX_pc [21] ), .A2(_05193_ ), .A3(\ID_EX_pc [20] ), .A4(_05194_ ), .ZN(_05195_ ) );
AND2_X1 _12937_ ( .A1(_05192_ ), .A2(_05195_ ), .ZN(_05196_ ) );
AND3_X1 _12938_ ( .A1(_05196_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_05197_ ) );
NAND2_X1 _12939_ ( .A1(_05197_ ), .A2(\ID_EX_pc [28] ), .ZN(_05198_ ) );
XNOR2_X1 _12940_ ( .A(_05198_ ), .B(\ID_EX_pc [29] ), .ZN(_05199_ ) );
OAI21_X1 _12941_ ( .A(_05199_ ), .B1(_05170_ ), .B2(_05173_ ), .ZN(_05200_ ) );
INV_X4 _12942_ ( .A(_05174_ ), .ZN(_05201_ ) );
BUF_X2 _12943_ ( .A(_05201_ ), .Z(_05202_ ) );
NAND2_X1 _12944_ ( .A1(_03994_ ), .A2(_03995_ ), .ZN(_05203_ ) );
NOR2_X1 _12945_ ( .A1(_03997_ ), .A2(_03892_ ), .ZN(_05204_ ) );
XNOR2_X1 _12946_ ( .A(_05203_ ), .B(_05204_ ), .ZN(_05205_ ) );
OAI211_X1 _12947_ ( .A(_05189_ ), .B(_05200_ ), .C1(_05202_ ), .C2(_05205_ ), .ZN(_05206_ ) );
BUF_X4 _12948_ ( .A(_05181_ ), .Z(_05207_ ) );
BUF_X4 _12949_ ( .A(_05178_ ), .Z(_05208_ ) );
XNOR2_X1 _12950_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_05209_ ) );
XNOR2_X1 _12951_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_05210_ ) );
XNOR2_X1 _12952_ ( .A(fanout_net_4 ), .B(\ID_EX_csr [1] ), .ZN(_05211_ ) );
XNOR2_X1 _12953_ ( .A(fanout_net_3 ), .B(\ID_EX_csr [0] ), .ZN(_05212_ ) );
AND4_X1 _12954_ ( .A1(_05209_ ), .A2(_05210_ ), .A3(_05211_ ), .A4(_05212_ ), .ZN(_05213_ ) );
XNOR2_X1 _12955_ ( .A(\EX_LS_dest_csreg_mem [9] ), .B(\ID_EX_csr [9] ), .ZN(_05214_ ) );
INV_X1 _12956_ ( .A(_01943_ ), .ZN(_05215_ ) );
NOR3_X1 _12957_ ( .A1(_03809_ ), .A2(_01924_ ), .A3(_05215_ ), .ZN(_05216_ ) );
AND4_X1 _12958_ ( .A1(_03820_ ), .A2(_05213_ ), .A3(_05214_ ), .A4(_05216_ ), .ZN(_05217_ ) );
XNOR2_X1 _12959_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_05218_ ) );
AND3_X1 _12960_ ( .A1(_03810_ ), .A2(_03804_ ), .A3(_05218_ ), .ZN(_05219_ ) );
AND4_X1 _12961_ ( .A1(_03822_ ), .A2(_05219_ ), .A3(_03826_ ), .A4(_03811_ ), .ZN(_05220_ ) );
AND2_X1 _12962_ ( .A1(_05217_ ), .A2(_05220_ ), .ZN(_05221_ ) );
INV_X1 _12963_ ( .A(_05221_ ), .ZN(_05222_ ) );
CLKBUF_X3 _12964_ ( .A(_03866_ ), .Z(_05223_ ) );
BUF_X2 _12965_ ( .A(_05223_ ), .Z(_05224_ ) );
NAND3_X1 _12966_ ( .A1(_03838_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_05224_ ), .ZN(_05225_ ) );
BUF_X2 _12967_ ( .A(_03848_ ), .Z(_05226_ ) );
BUF_X2 _12968_ ( .A(_03851_ ), .Z(_05227_ ) );
NAND3_X1 _12969_ ( .A1(_05226_ ), .A2(\mepc [29] ), .A3(_05227_ ), .ZN(_05228_ ) );
BUF_X2 _12970_ ( .A(_03855_ ), .Z(_05229_ ) );
AND3_X1 _12971_ ( .A1(_03848_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_05229_ ), .ZN(_05230_ ) );
AND3_X1 _12972_ ( .A1(_03860_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_05231_ ) );
AND3_X1 _12973_ ( .A1(_03832_ ), .A2(_03816_ ), .A3(\ID_EX_csr [4] ), .ZN(_05232_ ) );
AND2_X1 _12974_ ( .A1(_05231_ ), .A2(_05232_ ), .ZN(_05233_ ) );
AND2_X1 _12975_ ( .A1(_05233_ ), .A2(_03850_ ), .ZN(_05234_ ) );
AND3_X1 _12976_ ( .A1(_03837_ ), .A2(\mtvec [29] ), .A3(_03841_ ), .ZN(_05235_ ) );
NOR3_X1 _12977_ ( .A1(_05230_ ), .A2(_05234_ ), .A3(_05235_ ), .ZN(_05236_ ) );
NAND4_X1 _12978_ ( .A1(_05222_ ), .A2(_05225_ ), .A3(_05228_ ), .A4(_05236_ ), .ZN(_05237_ ) );
BUF_X4 _12979_ ( .A(_05217_ ), .Z(_05238_ ) );
INV_X1 _12980_ ( .A(\EX_LS_result_csreg_mem [29] ), .ZN(_05239_ ) );
BUF_X4 _12981_ ( .A(_05220_ ), .Z(_05240_ ) );
NAND3_X1 _12982_ ( .A1(_05238_ ), .A2(_05239_ ), .A3(_05240_ ), .ZN(_05241_ ) );
AND2_X1 _12983_ ( .A1(_05237_ ), .A2(_05241_ ), .ZN(_05242_ ) );
OAI211_X1 _12984_ ( .A(_05206_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05242_ ), .ZN(_05243_ ) );
MUX2_X1 _12985_ ( .A(_05205_ ), .B(_02970_ ), .S(fanout_net_5 ), .Z(_05244_ ) );
BUF_X2 _12986_ ( .A(_05180_ ), .Z(_05245_ ) );
OR2_X1 _12987_ ( .A1(_05244_ ), .A2(_05245_ ), .ZN(_05246_ ) );
AOI21_X1 _12988_ ( .A(_03801_ ), .B1(_05243_ ), .B2(_05246_ ), .ZN(_00123_ ) );
BUF_X4 _12989_ ( .A(_05181_ ), .Z(_05247_ ) );
BUF_X4 _12990_ ( .A(_05178_ ), .Z(_05248_ ) );
INV_X1 _12991_ ( .A(_03871_ ), .ZN(_05249_ ) );
AND2_X1 _12992_ ( .A1(_03861_ ), .A2(_05229_ ), .ZN(_05250_ ) );
INV_X1 _12993_ ( .A(_05250_ ), .ZN(_05251_ ) );
BUF_X2 _12994_ ( .A(_03847_ ), .Z(_05252_ ) );
NAND3_X1 _12995_ ( .A1(_05252_ ), .A2(\mepc [20] ), .A3(_03851_ ), .ZN(_05253_ ) );
NAND3_X1 _12996_ ( .A1(_05252_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_05229_ ), .ZN(_05254_ ) );
BUF_X2 _12997_ ( .A(_03836_ ), .Z(_05255_ ) );
NAND3_X1 _12998_ ( .A1(_05255_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_03866_ ), .ZN(_05256_ ) );
NAND3_X1 _12999_ ( .A1(_05255_ ), .A2(\mtvec [20] ), .A3(_03841_ ), .ZN(_05257_ ) );
AND4_X1 _13000_ ( .A1(_05253_ ), .A2(_05254_ ), .A3(_05256_ ), .A4(_05257_ ), .ZN(_05258_ ) );
NAND4_X1 _13001_ ( .A1(_05249_ ), .A2(_03863_ ), .A3(_05251_ ), .A4(_05258_ ), .ZN(_05259_ ) );
INV_X1 _13002_ ( .A(\EX_LS_result_csreg_mem [20] ), .ZN(_05260_ ) );
NAND3_X1 _13003_ ( .A1(_03814_ ), .A2(_03829_ ), .A3(_05260_ ), .ZN(_05261_ ) );
AND2_X1 _13004_ ( .A1(_05259_ ), .A2(_05261_ ), .ZN(_05262_ ) );
BUF_X2 _13005_ ( .A(_05175_ ), .Z(_05263_ ) );
XOR2_X1 _13006_ ( .A(_03967_ ), .B(_03972_ ), .Z(_05264_ ) );
AND2_X1 _13007_ ( .A1(_05263_ ), .A2(_05264_ ), .ZN(_05265_ ) );
BUF_X4 _13008_ ( .A(_05175_ ), .Z(_05266_ ) );
NAND3_X1 _13009_ ( .A1(_03879_ ), .A2(_05191_ ), .A3(_05194_ ), .ZN(_05267_ ) );
INV_X1 _13010_ ( .A(\ID_EX_pc [20] ), .ZN(_05268_ ) );
XNOR2_X1 _13011_ ( .A(_05267_ ), .B(_05268_ ), .ZN(_05269_ ) );
OAI21_X1 _13012_ ( .A(_05189_ ), .B1(_05266_ ), .B2(_05269_ ), .ZN(_05270_ ) );
OAI221_X1 _13013_ ( .A(_05247_ ), .B1(_05248_ ), .B2(_05262_ ), .C1(_05265_ ), .C2(_05270_ ), .ZN(_05271_ ) );
AND2_X2 _13014_ ( .A1(_03778_ ), .A2(fanout_net_5 ), .ZN(_05272_ ) );
AND3_X1 _13015_ ( .A1(_02941_ ), .A2(_02938_ ), .A3(_05272_ ), .ZN(_05273_ ) );
BUF_X4 _13016_ ( .A(_03780_ ), .Z(_05274_ ) );
AOI21_X1 _13017_ ( .A(_05273_ ), .B1(_05274_ ), .B2(_05264_ ), .ZN(_05275_ ) );
AOI21_X1 _13018_ ( .A(_03801_ ), .B1(_05271_ ), .B2(_05275_ ), .ZN(_00124_ ) );
NAND3_X1 _13019_ ( .A1(_03955_ ), .A2(_03956_ ), .A3(_03957_ ), .ZN(_05276_ ) );
NAND2_X1 _13020_ ( .A1(_05276_ ), .A2(_03964_ ), .ZN(_05277_ ) );
AND2_X1 _13021_ ( .A1(_05277_ ), .A2(_03896_ ), .ZN(_05278_ ) );
NOR2_X1 _13022_ ( .A1(_05278_ ), .A2(_03959_ ), .ZN(_05279_ ) );
XNOR2_X1 _13023_ ( .A(_05279_ ), .B(_03895_ ), .ZN(_05280_ ) );
AOI21_X1 _13024_ ( .A(\ID_EX_typ [3] ), .B1(_05263_ ), .B2(_05280_ ), .ZN(_05281_ ) );
NAND3_X1 _13025_ ( .A1(_03879_ ), .A2(\ID_EX_pc [18] ), .A3(_05191_ ), .ZN(_05282_ ) );
INV_X1 _13026_ ( .A(\ID_EX_pc [19] ), .ZN(_05283_ ) );
XNOR2_X1 _13027_ ( .A(_05282_ ), .B(_05283_ ), .ZN(_05284_ ) );
OAI21_X1 _13028_ ( .A(_05281_ ), .B1(_05266_ ), .B2(_05284_ ), .ZN(_05285_ ) );
AND2_X1 _13029_ ( .A1(_03837_ ), .A2(_03841_ ), .ZN(_05286_ ) );
BUF_X2 _13030_ ( .A(_05229_ ), .Z(_05287_ ) );
AOI22_X1 _13031_ ( .A1(_05286_ ), .A2(\mtvec [19] ), .B1(_03861_ ), .B2(_05287_ ), .ZN(_05288_ ) );
BUF_X2 _13032_ ( .A(_05252_ ), .Z(_05289_ ) );
NAND3_X1 _13033_ ( .A1(_05289_ ), .A2(\mepc [19] ), .A3(_05227_ ), .ZN(_05290_ ) );
BUF_X2 _13034_ ( .A(_03856_ ), .Z(_05291_ ) );
NAND3_X1 _13035_ ( .A1(_05289_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_05291_ ), .ZN(_05292_ ) );
NAND3_X1 _13036_ ( .A1(_03864_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_03867_ ), .ZN(_05293_ ) );
NAND4_X1 _13037_ ( .A1(_05288_ ), .A2(_05290_ ), .A3(_05292_ ), .A4(_05293_ ), .ZN(_05294_ ) );
NAND2_X1 _13038_ ( .A1(_05249_ ), .A2(_05294_ ), .ZN(_05295_ ) );
NAND3_X1 _13039_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(\EX_LS_result_csreg_mem [19] ), .ZN(_05296_ ) );
AND2_X1 _13040_ ( .A1(_05295_ ), .A2(_05296_ ), .ZN(_05297_ ) );
INV_X1 _13041_ ( .A(_05297_ ), .ZN(_05298_ ) );
OAI211_X1 _13042_ ( .A(_05285_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05298_ ), .ZN(_05299_ ) );
BUF_X4 _13043_ ( .A(_03779_ ), .Z(_05300_ ) );
NOR3_X1 _13044_ ( .A1(_02949_ ), .A2(_05300_ ), .A3(_05181_ ), .ZN(_05301_ ) );
AOI21_X1 _13045_ ( .A(_05301_ ), .B1(_05274_ ), .B2(_05280_ ), .ZN(_05302_ ) );
AOI21_X1 _13046_ ( .A(_03801_ ), .B1(_05299_ ), .B2(_05302_ ), .ZN(_00125_ ) );
INV_X1 _13047_ ( .A(\ID_EX_pc [18] ), .ZN(_05303_ ) );
XNOR2_X1 _13048_ ( .A(_05192_ ), .B(_05303_ ), .ZN(_05304_ ) );
XOR2_X1 _13049_ ( .A(_05277_ ), .B(_03896_ ), .Z(_05305_ ) );
MUX2_X1 _13050_ ( .A(_05304_ ), .B(_05305_ ), .S(_05175_ ), .Z(_05306_ ) );
OR2_X2 _13051_ ( .A1(_05306_ ), .A2(\ID_EX_typ [3] ), .ZN(_05307_ ) );
BUF_X2 _13052_ ( .A(_03814_ ), .Z(_05308_ ) );
BUF_X2 _13053_ ( .A(_03829_ ), .Z(_05309_ ) );
NAND3_X1 _13054_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [18] ), .ZN(_05310_ ) );
BUF_X2 _13055_ ( .A(_05252_ ), .Z(_05311_ ) );
BUF_X2 _13056_ ( .A(_05311_ ), .Z(_05312_ ) );
BUF_X2 _13057_ ( .A(_03851_ ), .Z(_05313_ ) );
BUF_X2 _13058_ ( .A(_05313_ ), .Z(_05314_ ) );
NAND3_X1 _13059_ ( .A1(_05312_ ), .A2(\mepc [18] ), .A3(_05314_ ), .ZN(_05315_ ) );
BUF_X2 _13060_ ( .A(_05255_ ), .Z(_05316_ ) );
BUF_X2 _13061_ ( .A(_05316_ ), .Z(_05317_ ) );
NAND3_X1 _13062_ ( .A1(_05317_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_05224_ ), .ZN(_05318_ ) );
NAND3_X1 _13063_ ( .A1(_03838_ ), .A2(\mtvec [18] ), .A3(_03842_ ), .ZN(_05319_ ) );
NAND3_X1 _13064_ ( .A1(_05315_ ), .A2(_05318_ ), .A3(_05319_ ), .ZN(_05320_ ) );
AND3_X1 _13065_ ( .A1(_05226_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_05291_ ), .ZN(_05321_ ) );
NOR3_X1 _13066_ ( .A1(_05320_ ), .A2(_05250_ ), .A3(_05321_ ), .ZN(_05322_ ) );
OAI21_X1 _13067_ ( .A(_05310_ ), .B1(_05322_ ), .B2(_03871_ ), .ZN(_05323_ ) );
OAI211_X1 _13068_ ( .A(_05307_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05323_ ), .ZN(_05324_ ) );
BUF_X4 _13069_ ( .A(_05272_ ), .Z(_05325_ ) );
BUF_X4 _13070_ ( .A(_03780_ ), .Z(_05326_ ) );
AOI22_X1 _13071_ ( .A1(_02950_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05305_ ), .ZN(_05327_ ) );
AOI21_X1 _13072_ ( .A(_03801_ ), .B1(_05324_ ), .B2(_05327_ ), .ZN(_00126_ ) );
AND2_X1 _13073_ ( .A1(_03955_ ), .A2(_03956_ ), .ZN(_05328_ ) );
NOR2_X1 _13074_ ( .A1(_05328_ ), .A2(_03963_ ), .ZN(_05329_ ) );
XNOR2_X1 _13075_ ( .A(_05329_ ), .B(_03957_ ), .ZN(_05330_ ) );
AOI21_X1 _13076_ ( .A(\ID_EX_typ [3] ), .B1(_05263_ ), .B2(_05330_ ), .ZN(_05331_ ) );
AND3_X1 _13077_ ( .A1(_03880_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_05332_ ) );
AND2_X1 _13078_ ( .A1(_03879_ ), .A2(_05332_ ), .ZN(_05333_ ) );
NAND3_X1 _13079_ ( .A1(_05333_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05334_ ) );
INV_X1 _13080_ ( .A(\ID_EX_pc [16] ), .ZN(_05335_ ) );
NOR2_X1 _13081_ ( .A1(_05334_ ), .A2(_05335_ ), .ZN(_05336_ ) );
XNOR2_X1 _13082_ ( .A(_05336_ ), .B(\ID_EX_pc [17] ), .ZN(_05337_ ) );
OAI21_X1 _13083_ ( .A(_05331_ ), .B1(_05266_ ), .B2(_05337_ ), .ZN(_05338_ ) );
AND3_X1 _13084_ ( .A1(_03837_ ), .A2(\mtvec [17] ), .A3(_03841_ ), .ZN(_05339_ ) );
AOI21_X1 _13085_ ( .A(_05339_ ), .B1(_05238_ ), .B2(_05240_ ), .ZN(_05340_ ) );
AND3_X1 _13086_ ( .A1(_05252_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_05229_ ), .ZN(_05341_ ) );
BUF_X4 _13087_ ( .A(_05234_ ), .Z(_05342_ ) );
AND2_X2 _13088_ ( .A1(_05233_ ), .A2(_05229_ ), .ZN(_05343_ ) );
NOR3_X1 _13089_ ( .A1(_05341_ ), .A2(_05342_ ), .A3(_05343_ ), .ZN(_05344_ ) );
NAND3_X1 _13090_ ( .A1(_05311_ ), .A2(\mepc [17] ), .A3(_05313_ ), .ZN(_05345_ ) );
CLKBUF_X2 _13091_ ( .A(_05255_ ), .Z(_05346_ ) );
NAND3_X1 _13092_ ( .A1(_05346_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_05223_ ), .ZN(_05347_ ) );
AND2_X1 _13093_ ( .A1(_05345_ ), .A2(_05347_ ), .ZN(_05348_ ) );
NAND3_X1 _13094_ ( .A1(_05340_ ), .A2(_05344_ ), .A3(_05348_ ), .ZN(_05349_ ) );
INV_X1 _13095_ ( .A(\EX_LS_result_csreg_mem [17] ), .ZN(_05350_ ) );
NAND3_X1 _13096_ ( .A1(_05238_ ), .A2(_05350_ ), .A3(_05240_ ), .ZN(_05351_ ) );
AND2_X1 _13097_ ( .A1(_05349_ ), .A2(_05351_ ), .ZN(_05352_ ) );
OAI211_X1 _13098_ ( .A(_05338_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05352_ ), .ZN(_05353_ ) );
NOR3_X1 _13099_ ( .A1(_02952_ ), .A2(_05300_ ), .A3(_05181_ ), .ZN(_05354_ ) );
AOI21_X1 _13100_ ( .A(_05354_ ), .B1(_05274_ ), .B2(_05330_ ), .ZN(_05355_ ) );
AOI21_X1 _13101_ ( .A(_03801_ ), .B1(_05353_ ), .B2(_05355_ ), .ZN(_00127_ ) );
NOR2_X1 _13102_ ( .A1(_03870_ ), .A2(_03862_ ), .ZN(_05356_ ) );
AND3_X1 _13103_ ( .A1(_05252_ ), .A2(\mepc [16] ), .A3(_03851_ ), .ZN(_05357_ ) );
AND3_X1 _13104_ ( .A1(_05255_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_03866_ ), .ZN(_05358_ ) );
NOR2_X1 _13105_ ( .A1(_05357_ ), .A2(_05358_ ), .ZN(_05359_ ) );
NAND3_X1 _13106_ ( .A1(_05252_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_05229_ ), .ZN(_05360_ ) );
NAND3_X1 _13107_ ( .A1(_03837_ ), .A2(\mtvec [16] ), .A3(_03841_ ), .ZN(_05361_ ) );
AND2_X1 _13108_ ( .A1(_05360_ ), .A2(_05361_ ), .ZN(_05362_ ) );
NAND4_X1 _13109_ ( .A1(_05356_ ), .A2(_05251_ ), .A3(_05359_ ), .A4(_05362_ ), .ZN(_05363_ ) );
INV_X1 _13110_ ( .A(\EX_LS_result_csreg_mem [16] ), .ZN(_05364_ ) );
NAND3_X1 _13111_ ( .A1(_03814_ ), .A2(_03829_ ), .A3(_05364_ ), .ZN(_05365_ ) );
AND2_X1 _13112_ ( .A1(_05363_ ), .A2(_05365_ ), .ZN(_05366_ ) );
XNOR2_X1 _13113_ ( .A(_05334_ ), .B(\ID_EX_pc [16] ), .ZN(_05367_ ) );
XOR2_X1 _13114_ ( .A(_03955_ ), .B(_03956_ ), .Z(_05368_ ) );
MUX2_X1 _13115_ ( .A(_05367_ ), .B(_05368_ ), .S(_05174_ ), .Z(_05369_ ) );
MUX2_X1 _13116_ ( .A(_05366_ ), .B(_05369_ ), .S(_05178_ ), .Z(_05370_ ) );
NAND2_X1 _13117_ ( .A1(_05370_ ), .A2(_05182_ ), .ZN(_05371_ ) );
NOR4_X1 _13118_ ( .A1(_02953_ ), .A2(_02943_ ), .A3(_05186_ ), .A4(_05180_ ), .ZN(_05372_ ) );
AOI21_X1 _13119_ ( .A(_05372_ ), .B1(_05274_ ), .B2(_05368_ ), .ZN(_05373_ ) );
AOI21_X1 _13120_ ( .A(_03801_ ), .B1(_05371_ ), .B2(_05373_ ), .ZN(_00128_ ) );
AND3_X1 _13121_ ( .A1(_05311_ ), .A2(\mepc [15] ), .A3(_05313_ ), .ZN(_05374_ ) );
AND3_X1 _13122_ ( .A1(_03848_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_03856_ ), .ZN(_05375_ ) );
AND3_X1 _13123_ ( .A1(_05346_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_05223_ ), .ZN(_05376_ ) );
NOR3_X1 _13124_ ( .A1(_05374_ ), .A2(_05375_ ), .A3(_05376_ ), .ZN(_05377_ ) );
AOI22_X1 _13125_ ( .A1(_05286_ ), .A2(\mtvec [15] ), .B1(_03861_ ), .B2(_05291_ ), .ZN(_05378_ ) );
AOI22_X1 _13126_ ( .A1(_05377_ ), .A2(_05378_ ), .B1(_03830_ ), .B2(_03815_ ), .ZN(_05379_ ) );
AND3_X1 _13127_ ( .A1(_03814_ ), .A2(_03829_ ), .A3(\EX_LS_result_csreg_mem [15] ), .ZN(_05380_ ) );
NOR2_X1 _13128_ ( .A1(_05379_ ), .A2(_05380_ ), .ZN(_05381_ ) );
INV_X1 _13129_ ( .A(_05381_ ), .ZN(_05382_ ) );
NAND3_X1 _13130_ ( .A1(_03879_ ), .A2(\ID_EX_pc [14] ), .A3(_05332_ ), .ZN(_05383_ ) );
XNOR2_X1 _13131_ ( .A(_05383_ ), .B(\ID_EX_pc [15] ), .ZN(_05384_ ) );
INV_X1 _13132_ ( .A(_03941_ ), .ZN(_05385_ ) );
OAI21_X1 _13133_ ( .A(_03944_ ), .B1(_03930_ ), .B2(_03938_ ), .ZN(_05386_ ) );
AOI21_X1 _13134_ ( .A(_05385_ ), .B1(_05386_ ), .B2(_03948_ ), .ZN(_05387_ ) );
NOR2_X1 _13135_ ( .A1(_05387_ ), .A2(_03952_ ), .ZN(_05388_ ) );
XNOR2_X1 _13136_ ( .A(_05388_ ), .B(_03940_ ), .ZN(_05389_ ) );
MUX2_X1 _13137_ ( .A(_05384_ ), .B(_05389_ ), .S(_05174_ ), .Z(_05390_ ) );
MUX2_X1 _13138_ ( .A(_05382_ ), .B(_05390_ ), .S(_05178_ ), .Z(_05391_ ) );
NAND2_X1 _13139_ ( .A1(_05391_ ), .A2(_05182_ ), .ZN(_05392_ ) );
NOR3_X1 _13140_ ( .A1(_02963_ ), .A2(_05300_ ), .A3(_05180_ ), .ZN(_05393_ ) );
AOI21_X1 _13141_ ( .A(_05393_ ), .B1(_05274_ ), .B2(_05389_ ), .ZN(_05394_ ) );
AOI21_X1 _13142_ ( .A(_03801_ ), .B1(_05392_ ), .B2(_05394_ ), .ZN(_00129_ ) );
BUF_X4 _13143_ ( .A(_03800_ ), .Z(_05395_ ) );
AND2_X1 _13144_ ( .A1(_05356_ ), .A2(_05251_ ), .ZN(_05396_ ) );
AND3_X1 _13145_ ( .A1(_05311_ ), .A2(\mepc [14] ), .A3(_05313_ ), .ZN(_05397_ ) );
AND3_X1 _13146_ ( .A1(_05346_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_05223_ ), .ZN(_05398_ ) );
NOR2_X1 _13147_ ( .A1(_05397_ ), .A2(_05398_ ), .ZN(_05399_ ) );
NAND3_X1 _13148_ ( .A1(_03838_ ), .A2(\mtvec [14] ), .A3(_03842_ ), .ZN(_05400_ ) );
AND3_X1 _13149_ ( .A1(_05311_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_03856_ ), .ZN(_05401_ ) );
INV_X1 _13150_ ( .A(_05401_ ), .ZN(_05402_ ) );
NAND4_X1 _13151_ ( .A1(_05396_ ), .A2(_05399_ ), .A3(_05400_ ), .A4(_05402_ ), .ZN(_05403_ ) );
INV_X1 _13152_ ( .A(\EX_LS_result_csreg_mem [14] ), .ZN(_05404_ ) );
NAND3_X1 _13153_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(_05404_ ), .ZN(_05405_ ) );
AND2_X1 _13154_ ( .A1(_05403_ ), .A2(_05405_ ), .ZN(_05406_ ) );
INV_X1 _13155_ ( .A(\ID_EX_pc [14] ), .ZN(_05407_ ) );
XNOR2_X1 _13156_ ( .A(_05333_ ), .B(_05407_ ), .ZN(_05408_ ) );
AND3_X1 _13157_ ( .A1(_05386_ ), .A2(_05385_ ), .A3(_03948_ ), .ZN(_05409_ ) );
NOR2_X1 _13158_ ( .A1(_05409_ ), .A2(_05387_ ), .ZN(_05410_ ) );
MUX2_X1 _13159_ ( .A(_05408_ ), .B(_05410_ ), .S(_05174_ ), .Z(_05411_ ) );
MUX2_X1 _13160_ ( .A(_05406_ ), .B(_05411_ ), .S(_05178_ ), .Z(_05412_ ) );
NAND2_X1 _13161_ ( .A1(_05412_ ), .A2(_05182_ ), .ZN(_05413_ ) );
AOI22_X1 _13162_ ( .A1(_02964_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05410_ ), .ZN(_05414_ ) );
AOI21_X1 _13163_ ( .A(_05395_ ), .B1(_05413_ ), .B2(_05414_ ), .ZN(_00130_ ) );
AND2_X1 _13164_ ( .A1(_03939_ ), .A2(_03942_ ), .ZN(_05415_ ) );
NOR2_X1 _13165_ ( .A1(_05415_ ), .A2(_03946_ ), .ZN(_05416_ ) );
XNOR2_X1 _13166_ ( .A(_05416_ ), .B(_03943_ ), .ZN(_05417_ ) );
AOI21_X1 _13167_ ( .A(\ID_EX_typ [3] ), .B1(_05263_ ), .B2(_05417_ ), .ZN(_05418_ ) );
AND2_X1 _13168_ ( .A1(_03881_ ), .A2(\ID_EX_pc [12] ), .ZN(_05419_ ) );
XNOR2_X1 _13169_ ( .A(_05419_ ), .B(\ID_EX_pc [13] ), .ZN(_05420_ ) );
OAI21_X1 _13170_ ( .A(_05418_ ), .B1(_05266_ ), .B2(_05420_ ), .ZN(_05421_ ) );
NAND3_X1 _13171_ ( .A1(_05255_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_03866_ ), .ZN(_05422_ ) );
NAND3_X1 _13172_ ( .A1(_03847_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_03855_ ), .ZN(_05423_ ) );
NAND3_X1 _13173_ ( .A1(_03847_ ), .A2(\mepc [13] ), .A3(_03851_ ), .ZN(_05424_ ) );
NAND3_X1 _13174_ ( .A1(_05255_ ), .A2(\mtvec [13] ), .A3(_03840_ ), .ZN(_05425_ ) );
AND4_X1 _13175_ ( .A1(_05422_ ), .A2(_05423_ ), .A3(_05424_ ), .A4(_05425_ ), .ZN(_05426_ ) );
NAND3_X1 _13176_ ( .A1(_05249_ ), .A2(_03863_ ), .A3(_05426_ ), .ZN(_05427_ ) );
INV_X1 _13177_ ( .A(\EX_LS_result_csreg_mem [13] ), .ZN(_05428_ ) );
NAND3_X1 _13178_ ( .A1(_03814_ ), .A2(_03829_ ), .A3(_05428_ ), .ZN(_05429_ ) );
AND2_X1 _13179_ ( .A1(_05427_ ), .A2(_05429_ ), .ZN(_05430_ ) );
OAI211_X1 _13180_ ( .A(_05421_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05430_ ), .ZN(_05431_ ) );
NOR3_X1 _13181_ ( .A1(_02967_ ), .A2(_05300_ ), .A3(_05180_ ), .ZN(_05432_ ) );
AOI21_X1 _13182_ ( .A(_05432_ ), .B1(_05274_ ), .B2(_05417_ ), .ZN(_05433_ ) );
AOI21_X1 _13183_ ( .A(_05395_ ), .B1(_05431_ ), .B2(_05433_ ), .ZN(_00131_ ) );
INV_X1 _13184_ ( .A(\EX_LS_result_csreg_mem [12] ), .ZN(_05434_ ) );
AND3_X1 _13185_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(_05434_ ), .ZN(_05435_ ) );
AND3_X1 _13186_ ( .A1(_05289_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_05287_ ), .ZN(_05436_ ) );
BUF_X2 _13187_ ( .A(_05252_ ), .Z(_05437_ ) );
AND3_X1 _13188_ ( .A1(_05437_ ), .A2(\mepc [12] ), .A3(_05227_ ), .ZN(_05438_ ) );
CLKBUF_X2 _13189_ ( .A(_03840_ ), .Z(_05439_ ) );
AND3_X1 _13190_ ( .A1(_05316_ ), .A2(\mtvec [12] ), .A3(_05439_ ), .ZN(_05440_ ) );
AND3_X1 _13191_ ( .A1(_03864_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_03867_ ), .ZN(_05441_ ) );
NOR4_X1 _13192_ ( .A1(_05436_ ), .A2(_05438_ ), .A3(_05440_ ), .A4(_05441_ ), .ZN(_05442_ ) );
AOI21_X1 _13193_ ( .A(_05435_ ), .B1(_05396_ ), .B2(_05442_ ), .ZN(_05443_ ) );
INV_X1 _13194_ ( .A(\ID_EX_pc [12] ), .ZN(_05444_ ) );
XNOR2_X1 _13195_ ( .A(_03881_ ), .B(_05444_ ), .ZN(_05445_ ) );
XOR2_X1 _13196_ ( .A(_03939_ ), .B(_03942_ ), .Z(_05446_ ) );
MUX2_X1 _13197_ ( .A(_05445_ ), .B(_05446_ ), .S(_05174_ ), .Z(_05447_ ) );
MUX2_X1 _13198_ ( .A(_05443_ ), .B(_05447_ ), .S(_05177_ ), .Z(_05448_ ) );
NAND2_X1 _13199_ ( .A1(_05448_ ), .A2(_05182_ ), .ZN(_05449_ ) );
AND3_X1 _13200_ ( .A1(_02968_ ), .A2(_02965_ ), .A3(_05272_ ), .ZN(_05450_ ) );
AOI21_X1 _13201_ ( .A(_05450_ ), .B1(_05274_ ), .B2(_05446_ ), .ZN(_05451_ ) );
AOI21_X1 _13202_ ( .A(_05395_ ), .B1(_05449_ ), .B2(_05451_ ), .ZN(_00132_ ) );
INV_X1 _13203_ ( .A(_03925_ ), .ZN(_05452_ ) );
NAND2_X1 _13204_ ( .A1(_03923_ ), .A2(_03929_ ), .ZN(_05453_ ) );
AOI21_X1 _13205_ ( .A(_05452_ ), .B1(_05453_ ), .B2(_03936_ ), .ZN(_05454_ ) );
NOR2_X1 _13206_ ( .A1(_05454_ ), .A2(_03931_ ), .ZN(_05455_ ) );
XNOR2_X1 _13207_ ( .A(_05455_ ), .B(_03924_ ), .ZN(_05456_ ) );
AOI21_X1 _13208_ ( .A(\ID_EX_typ [3] ), .B1(_05263_ ), .B2(_05456_ ), .ZN(_05457_ ) );
AND2_X1 _13209_ ( .A1(_03879_ ), .A2(\ID_EX_pc [10] ), .ZN(_05458_ ) );
XNOR2_X1 _13210_ ( .A(_05458_ ), .B(\ID_EX_pc [11] ), .ZN(_05459_ ) );
OAI21_X1 _13211_ ( .A(_05457_ ), .B1(_05266_ ), .B2(_05459_ ), .ZN(_05460_ ) );
NAND3_X1 _13212_ ( .A1(_05317_ ), .A2(\mtvec [11] ), .A3(_03842_ ), .ZN(_05461_ ) );
AND3_X1 _13213_ ( .A1(_05437_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_05287_ ), .ZN(_05462_ ) );
NOR3_X1 _13214_ ( .A1(_05462_ ), .A2(_05342_ ), .A3(_05343_ ), .ZN(_05463_ ) );
NAND3_X1 _13215_ ( .A1(_05226_ ), .A2(\mepc [11] ), .A3(_05227_ ), .ZN(_05464_ ) );
NAND3_X1 _13216_ ( .A1(_03838_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_05224_ ), .ZN(_05465_ ) );
AND2_X1 _13217_ ( .A1(_05464_ ), .A2(_05465_ ), .ZN(_05466_ ) );
NAND4_X1 _13218_ ( .A1(_05222_ ), .A2(_05461_ ), .A3(_05463_ ), .A4(_05466_ ), .ZN(_05467_ ) );
BUF_X2 _13219_ ( .A(_05238_ ), .Z(_05468_ ) );
INV_X1 _13220_ ( .A(\EX_LS_result_csreg_mem [11] ), .ZN(_05469_ ) );
BUF_X2 _13221_ ( .A(_05240_ ), .Z(_05470_ ) );
NAND3_X1 _13222_ ( .A1(_05468_ ), .A2(_05469_ ), .A3(_05470_ ), .ZN(_05471_ ) );
AND2_X1 _13223_ ( .A1(_05467_ ), .A2(_05471_ ), .ZN(_05472_ ) );
OAI211_X1 _13224_ ( .A(_05460_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05472_ ), .ZN(_05473_ ) );
AOI21_X1 _13225_ ( .A(_02732_ ), .B1(_02539_ ), .B2(_02682_ ), .ZN(_05474_ ) );
AND3_X1 _13226_ ( .A1(_02722_ ), .A2(_02723_ ), .A3(_02725_ ), .ZN(_05475_ ) );
NOR3_X1 _13227_ ( .A1(_05474_ ), .A2(_02735_ ), .A3(_05475_ ), .ZN(_05476_ ) );
NOR2_X1 _13228_ ( .A1(_05476_ ), .A2(_02735_ ), .ZN(_05477_ ) );
XNOR2_X1 _13229_ ( .A(_05477_ ), .B(_02704_ ), .ZN(_05478_ ) );
AOI22_X1 _13230_ ( .A1(_05478_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05456_ ), .ZN(_05479_ ) );
AOI21_X1 _13231_ ( .A(_05395_ ), .B1(_05473_ ), .B2(_05479_ ), .ZN(_00133_ ) );
NAND3_X1 _13232_ ( .A1(_05196_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_05480_ ) );
XNOR2_X1 _13233_ ( .A(_05480_ ), .B(\ID_EX_pc [28] ), .ZN(_05481_ ) );
OAI21_X1 _13234_ ( .A(_05481_ ), .B1(_05170_ ), .B2(_05173_ ), .ZN(_05482_ ) );
XNOR2_X1 _13235_ ( .A(_03992_ ), .B(_03993_ ), .ZN(_05483_ ) );
OAI211_X1 _13236_ ( .A(_05189_ ), .B(_05482_ ), .C1(_05202_ ), .C2(_05483_ ), .ZN(_05484_ ) );
NOR2_X1 _13237_ ( .A1(_05222_ ), .A2(\EX_LS_result_csreg_mem [28] ), .ZN(_05485_ ) );
AND3_X1 _13238_ ( .A1(_05289_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_05287_ ), .ZN(_05486_ ) );
AND3_X1 _13239_ ( .A1(_03864_ ), .A2(\mtvec [28] ), .A3(_05439_ ), .ZN(_05487_ ) );
NOR3_X1 _13240_ ( .A1(_05486_ ), .A2(_05342_ ), .A3(_05487_ ), .ZN(_05488_ ) );
NAND3_X1 _13241_ ( .A1(_05289_ ), .A2(\mepc [28] ), .A3(_05227_ ), .ZN(_05489_ ) );
NAND3_X1 _13242_ ( .A1(_03864_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_03867_ ), .ZN(_05490_ ) );
NAND2_X1 _13243_ ( .A1(_05489_ ), .A2(_05490_ ), .ZN(_05491_ ) );
BUF_X2 _13244_ ( .A(_05217_ ), .Z(_05492_ ) );
BUF_X2 _13245_ ( .A(_05220_ ), .Z(_05493_ ) );
AOI21_X1 _13246_ ( .A(_05491_ ), .B1(_05492_ ), .B2(_05493_ ), .ZN(_05494_ ) );
AOI21_X1 _13247_ ( .A(_05485_ ), .B1(_05488_ ), .B2(_05494_ ), .ZN(_05495_ ) );
OAI211_X1 _13248_ ( .A(_05484_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05495_ ), .ZN(_05496_ ) );
OAI21_X1 _13249_ ( .A(fanout_net_5 ), .B1(_02971_ ), .B2(_02873_ ), .ZN(_05497_ ) );
BUF_X4 _13250_ ( .A(_05180_ ), .Z(_05498_ ) );
BUF_X4 _13251_ ( .A(_05186_ ), .Z(_05499_ ) );
AOI21_X1 _13252_ ( .A(_05498_ ), .B1(_05483_ ), .B2(_05499_ ), .ZN(_05500_ ) );
NAND2_X1 _13253_ ( .A1(_05497_ ), .A2(_05500_ ), .ZN(_05501_ ) );
AOI21_X1 _13254_ ( .A(_05395_ ), .B1(_05496_ ), .B2(_05501_ ), .ZN(_00134_ ) );
INV_X1 _13255_ ( .A(\ID_EX_pc [10] ), .ZN(_05502_ ) );
XNOR2_X1 _13256_ ( .A(_03879_ ), .B(_05502_ ), .ZN(_05503_ ) );
AND3_X1 _13257_ ( .A1(_05453_ ), .A2(_05452_ ), .A3(_03936_ ), .ZN(_05504_ ) );
NOR2_X1 _13258_ ( .A1(_05504_ ), .A2(_05454_ ), .ZN(_05505_ ) );
MUX2_X1 _13259_ ( .A(_05503_ ), .B(_05505_ ), .S(_05175_ ), .Z(_05506_ ) );
OR2_X2 _13260_ ( .A1(_05506_ ), .A2(\ID_EX_typ [3] ), .ZN(_05507_ ) );
AOI22_X1 _13261_ ( .A1(_05286_ ), .A2(\mtvec [10] ), .B1(_03861_ ), .B2(_05287_ ), .ZN(_05508_ ) );
NAND3_X1 _13262_ ( .A1(_05289_ ), .A2(\mepc [10] ), .A3(_05227_ ), .ZN(_05509_ ) );
NAND3_X1 _13263_ ( .A1(_05289_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_05287_ ), .ZN(_05510_ ) );
NAND3_X1 _13264_ ( .A1(_03864_ ), .A2(\mycsreg.CSReg[0][10] ), .A3(_03867_ ), .ZN(_05511_ ) );
NAND4_X1 _13265_ ( .A1(_05508_ ), .A2(_05509_ ), .A3(_05510_ ), .A4(_05511_ ), .ZN(_05512_ ) );
NAND2_X1 _13266_ ( .A1(_05249_ ), .A2(_05512_ ), .ZN(_05513_ ) );
NAND3_X1 _13267_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(\EX_LS_result_csreg_mem [10] ), .ZN(_05514_ ) );
AND2_X1 _13268_ ( .A1(_05513_ ), .A2(_05514_ ), .ZN(_05515_ ) );
INV_X1 _13269_ ( .A(_05515_ ), .ZN(_05516_ ) );
OAI211_X1 _13270_ ( .A(_05507_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05516_ ), .ZN(_05517_ ) );
XNOR2_X1 _13271_ ( .A(_05474_ ), .B(_02726_ ), .ZN(_05518_ ) );
AOI22_X1 _13272_ ( .A1(_05518_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05505_ ), .ZN(_05519_ ) );
AOI21_X1 _13273_ ( .A(_05395_ ), .B1(_05517_ ), .B2(_05519_ ), .ZN(_00135_ ) );
AND3_X1 _13274_ ( .A1(_05311_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_03856_ ), .ZN(_05520_ ) );
INV_X1 _13275_ ( .A(_05520_ ), .ZN(_05521_ ) );
AOI22_X1 _13276_ ( .A1(_05286_ ), .A2(\mtvec [9] ), .B1(_03861_ ), .B2(_05287_ ), .ZN(_05522_ ) );
NAND3_X1 _13277_ ( .A1(_05226_ ), .A2(\mepc [9] ), .A3(_05227_ ), .ZN(_05523_ ) );
AND3_X1 _13278_ ( .A1(_05346_ ), .A2(\mycsreg.CSReg[0][9] ), .A3(_05223_ ), .ZN(_05524_ ) );
INV_X1 _13279_ ( .A(_05524_ ), .ZN(_05525_ ) );
NAND4_X1 _13280_ ( .A1(_05521_ ), .A2(_05522_ ), .A3(_05523_ ), .A4(_05525_ ), .ZN(_05526_ ) );
NAND2_X1 _13281_ ( .A1(_05526_ ), .A2(_05249_ ), .ZN(_05527_ ) );
NAND3_X1 _13282_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(\EX_LS_result_csreg_mem [9] ), .ZN(_05528_ ) );
AND2_X1 _13283_ ( .A1(_05527_ ), .A2(_05528_ ), .ZN(_05529_ ) );
INV_X1 _13284_ ( .A(_05529_ ), .ZN(_05530_ ) );
AND2_X1 _13285_ ( .A1(_03923_ ), .A2(_03927_ ), .ZN(_05531_ ) );
NOR2_X1 _13286_ ( .A1(_05531_ ), .A2(_03934_ ), .ZN(_05532_ ) );
XNOR2_X1 _13287_ ( .A(_05532_ ), .B(_03928_ ), .ZN(_05533_ ) );
AND2_X1 _13288_ ( .A1(_05263_ ), .A2(_05533_ ), .ZN(_05534_ ) );
XNOR2_X1 _13289_ ( .A(_03878_ ), .B(\ID_EX_pc [9] ), .ZN(_05535_ ) );
OAI21_X1 _13290_ ( .A(_05189_ ), .B1(_05266_ ), .B2(_05535_ ), .ZN(_05536_ ) );
OAI221_X1 _13291_ ( .A(_05247_ ), .B1(_05248_ ), .B2(_05530_ ), .C1(_05534_ ), .C2(_05536_ ), .ZN(_05537_ ) );
NAND2_X1 _13292_ ( .A1(_02539_ ), .A2(_02656_ ), .ZN(_05538_ ) );
AND2_X1 _13293_ ( .A1(_05538_ ), .A2(_02731_ ), .ZN(_05539_ ) );
XNOR2_X1 _13294_ ( .A(_05539_ ), .B(_02730_ ), .ZN(_05540_ ) );
NOR3_X1 _13295_ ( .A1(_05540_ ), .A2(_05300_ ), .A3(_05180_ ), .ZN(_05541_ ) );
AOI21_X1 _13296_ ( .A(_05541_ ), .B1(_05274_ ), .B2(_05533_ ), .ZN(_05542_ ) );
AOI21_X1 _13297_ ( .A(_05395_ ), .B1(_05537_ ), .B2(_05542_ ), .ZN(_00136_ ) );
BUF_X4 _13298_ ( .A(_05181_ ), .Z(_05543_ ) );
INV_X1 _13299_ ( .A(\EX_LS_result_csreg_mem [8] ), .ZN(_05544_ ) );
AND3_X1 _13300_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(_05544_ ), .ZN(_05545_ ) );
AND3_X1 _13301_ ( .A1(_03864_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_03867_ ), .ZN(_05546_ ) );
INV_X1 _13302_ ( .A(_05546_ ), .ZN(_05547_ ) );
NAND3_X1 _13303_ ( .A1(_05312_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_05291_ ), .ZN(_05548_ ) );
NAND2_X1 _13304_ ( .A1(_05547_ ), .A2(_05548_ ), .ZN(_05549_ ) );
AND3_X1 _13305_ ( .A1(_05226_ ), .A2(\mepc [8] ), .A3(_05314_ ), .ZN(_05550_ ) );
AND3_X1 _13306_ ( .A1(_03838_ ), .A2(\mtvec [8] ), .A3(_03842_ ), .ZN(_05551_ ) );
NOR3_X1 _13307_ ( .A1(_05549_ ), .A2(_05550_ ), .A3(_05551_ ), .ZN(_05552_ ) );
AOI21_X1 _13308_ ( .A(_05545_ ), .B1(_05396_ ), .B2(_05552_ ), .ZN(_05553_ ) );
XOR2_X1 _13309_ ( .A(_03923_ ), .B(_03927_ ), .Z(_05554_ ) );
AND2_X1 _13310_ ( .A1(_05263_ ), .A2(_05554_ ), .ZN(_05555_ ) );
XNOR2_X1 _13311_ ( .A(_03877_ ), .B(\ID_EX_pc [8] ), .ZN(_05556_ ) );
OAI21_X1 _13312_ ( .A(_05189_ ), .B1(_05266_ ), .B2(_05556_ ), .ZN(_05557_ ) );
OAI221_X1 _13313_ ( .A(_05543_ ), .B1(_05189_ ), .B2(_05553_ ), .C1(_05555_ ), .C2(_05557_ ), .ZN(_05558_ ) );
XOR2_X1 _13314_ ( .A(_02539_ ), .B(_02656_ ), .Z(_05559_ ) );
AOI22_X1 _13315_ ( .A1(_05559_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05554_ ), .ZN(_05560_ ) );
AOI21_X1 _13316_ ( .A(_05395_ ), .B1(_05558_ ), .B2(_05560_ ), .ZN(_00137_ ) );
NAND3_X1 _13317_ ( .A1(_05311_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_03856_ ), .ZN(_05561_ ) );
NAND3_X1 _13318_ ( .A1(_05311_ ), .A2(\mepc [7] ), .A3(_05313_ ), .ZN(_05562_ ) );
NAND3_X1 _13319_ ( .A1(_05316_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_05223_ ), .ZN(_05563_ ) );
NAND3_X1 _13320_ ( .A1(_05346_ ), .A2(\mtvec [7] ), .A3(_05439_ ), .ZN(_05564_ ) );
NAND4_X1 _13321_ ( .A1(_05561_ ), .A2(_05562_ ), .A3(_05563_ ), .A4(_05564_ ), .ZN(_05565_ ) );
AOI21_X1 _13322_ ( .A(_05565_ ), .B1(_05468_ ), .B2(_05470_ ), .ZN(_05566_ ) );
INV_X1 _13323_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_05567_ ) );
AND3_X1 _13324_ ( .A1(_05468_ ), .A2(_05567_ ), .A3(_05470_ ), .ZN(_05568_ ) );
NOR2_X1 _13325_ ( .A1(_05566_ ), .A2(_05568_ ), .ZN(_05569_ ) );
XNOR2_X1 _13326_ ( .A(\ID_EX_pc [7] ), .B(\ID_EX_imm [7] ), .ZN(_05570_ ) );
XNOR2_X1 _13327_ ( .A(_03919_ ), .B(_05570_ ), .ZN(_05571_ ) );
AND2_X1 _13328_ ( .A1(_05263_ ), .A2(_05571_ ), .ZN(_05572_ ) );
XNOR2_X1 _13329_ ( .A(_03876_ ), .B(\ID_EX_pc [7] ), .ZN(_05573_ ) );
OAI21_X1 _13330_ ( .A(_05189_ ), .B1(_05266_ ), .B2(_05573_ ), .ZN(_05574_ ) );
OAI221_X1 _13331_ ( .A(_05543_ ), .B1(_05189_ ), .B2(_05569_ ), .C1(_05572_ ), .C2(_05574_ ), .ZN(_05575_ ) );
NOR3_X1 _13332_ ( .A1(_02431_ ), .A2(_02526_ ), .A3(_02455_ ), .ZN(_05576_ ) );
OAI21_X1 _13333_ ( .A(_02500_ ), .B1(_05576_ ), .B2(_02537_ ), .ZN(_05577_ ) );
NAND2_X1 _13334_ ( .A1(_05577_ ), .A2(_02531_ ), .ZN(_05578_ ) );
XNOR2_X1 _13335_ ( .A(_05578_ ), .B(_02529_ ), .ZN(_05579_ ) );
AOI22_X1 _13336_ ( .A1(_05579_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05571_ ), .ZN(_05580_ ) );
AOI21_X1 _13337_ ( .A(_05395_ ), .B1(_05575_ ), .B2(_05580_ ), .ZN(_00138_ ) );
INV_X1 _13338_ ( .A(\ID_EX_pc [6] ), .ZN(_05581_ ) );
XNOR2_X1 _13339_ ( .A(_03875_ ), .B(_05581_ ), .ZN(_05582_ ) );
XOR2_X1 _13340_ ( .A(_03915_ ), .B(_03916_ ), .Z(_05583_ ) );
MUX2_X1 _13341_ ( .A(_05582_ ), .B(_05583_ ), .S(_05175_ ), .Z(_05584_ ) );
AND2_X2 _13342_ ( .A1(_05584_ ), .A2(_05178_ ), .ZN(_05585_ ) );
NAND3_X1 _13343_ ( .A1(_05226_ ), .A2(\mepc [6] ), .A3(_05314_ ), .ZN(_05586_ ) );
NAND3_X1 _13344_ ( .A1(_03838_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_05224_ ), .ZN(_05587_ ) );
NAND2_X1 _13345_ ( .A1(_05586_ ), .A2(_05587_ ), .ZN(_05588_ ) );
AOI21_X1 _13346_ ( .A(_05588_ ), .B1(_05492_ ), .B2(_05493_ ), .ZN(_05589_ ) );
AND3_X1 _13347_ ( .A1(_05226_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_05291_ ), .ZN(_05590_ ) );
AND3_X1 _13348_ ( .A1(_03864_ ), .A2(\mtvec [6] ), .A3(_05439_ ), .ZN(_05591_ ) );
NOR3_X1 _13349_ ( .A1(_05590_ ), .A2(_05342_ ), .A3(_05591_ ), .ZN(_05592_ ) );
NAND2_X1 _13350_ ( .A1(_05589_ ), .A2(_05592_ ), .ZN(_05593_ ) );
INV_X1 _13351_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_05594_ ) );
NAND3_X1 _13352_ ( .A1(_05468_ ), .A2(_05594_ ), .A3(_05470_ ), .ZN(_05595_ ) );
AND3_X1 _13353_ ( .A1(_05593_ ), .A2(\ID_EX_typ [3] ), .A3(_05595_ ), .ZN(_05596_ ) );
OAI21_X1 _13354_ ( .A(_05182_ ), .B1(_05585_ ), .B2(_05596_ ), .ZN(_05597_ ) );
OR3_X1 _13355_ ( .A1(_05576_ ), .A2(_02500_ ), .A3(_02537_ ), .ZN(_05598_ ) );
AND2_X1 _13356_ ( .A1(_05598_ ), .A2(_05577_ ), .ZN(_05599_ ) );
AOI22_X1 _13357_ ( .A1(_05599_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05583_ ), .ZN(_05600_ ) );
AOI21_X1 _13358_ ( .A(_05395_ ), .B1(_05597_ ), .B2(_05600_ ), .ZN(_00139_ ) );
BUF_X4 _13359_ ( .A(_03800_ ), .Z(_05601_ ) );
INV_X1 _13360_ ( .A(\ID_EX_pc [5] ), .ZN(_05602_ ) );
XNOR2_X1 _13361_ ( .A(_03874_ ), .B(_05602_ ), .ZN(_05603_ ) );
AOI21_X1 _13362_ ( .A(\ID_EX_typ [3] ), .B1(_05201_ ), .B2(_05603_ ), .ZN(_05604_ ) );
XOR2_X1 _13363_ ( .A(\ID_EX_pc [5] ), .B(\ID_EX_imm [5] ), .Z(_05605_ ) );
XNOR2_X1 _13364_ ( .A(_03911_ ), .B(_05605_ ), .ZN(_05606_ ) );
OAI21_X1 _13365_ ( .A(_05604_ ), .B1(_05202_ ), .B2(_05606_ ), .ZN(_05607_ ) );
AND3_X1 _13366_ ( .A1(_03848_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_03856_ ), .ZN(_05608_ ) );
AND3_X1 _13367_ ( .A1(_05346_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_05223_ ), .ZN(_05609_ ) );
NOR2_X1 _13368_ ( .A1(_05608_ ), .A2(_05609_ ), .ZN(_05610_ ) );
AND3_X1 _13369_ ( .A1(_05226_ ), .A2(\mepc [5] ), .A3(_05314_ ), .ZN(_05611_ ) );
AND3_X1 _13370_ ( .A1(_03837_ ), .A2(\mtvec [5] ), .A3(_03841_ ), .ZN(_05612_ ) );
NOR2_X1 _13371_ ( .A1(_05611_ ), .A2(_05612_ ), .ZN(_05613_ ) );
NAND4_X1 _13372_ ( .A1(_05249_ ), .A2(_03863_ ), .A3(_05610_ ), .A4(_05613_ ), .ZN(_05614_ ) );
INV_X1 _13373_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_05615_ ) );
NAND3_X1 _13374_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(_05615_ ), .ZN(_05616_ ) );
AND2_X1 _13375_ ( .A1(_05614_ ), .A2(_05616_ ), .ZN(_05617_ ) );
OAI211_X1 _13376_ ( .A(_05607_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05617_ ), .ZN(_05618_ ) );
NOR2_X1 _13377_ ( .A1(_05606_ ), .A2(_03781_ ), .ZN(_05619_ ) );
AOI21_X1 _13378_ ( .A(_02453_ ), .B1(_02432_ ), .B2(_02451_ ), .ZN(_05620_ ) );
NOR2_X1 _13379_ ( .A1(_02456_ ), .A2(_05620_ ), .ZN(_05621_ ) );
XNOR2_X1 _13380_ ( .A(_05621_ ), .B(_02527_ ), .ZN(_05622_ ) );
AOI21_X1 _13381_ ( .A(_05619_ ), .B1(_05622_ ), .B2(_05325_ ), .ZN(_05623_ ) );
AOI21_X1 _13382_ ( .A(_05601_ ), .B1(_05618_ ), .B2(_05623_ ), .ZN(_00140_ ) );
INV_X1 _13383_ ( .A(\ID_EX_pc [4] ), .ZN(_05624_ ) );
XNOR2_X1 _13384_ ( .A(_03873_ ), .B(_05624_ ), .ZN(_05625_ ) );
AOI21_X1 _13385_ ( .A(\ID_EX_typ [3] ), .B1(_05201_ ), .B2(_05625_ ), .ZN(_05626_ ) );
OR2_X1 _13386_ ( .A1(_03907_ ), .A2(_03908_ ), .ZN(_05627_ ) );
XOR2_X1 _13387_ ( .A(_05627_ ), .B(_03898_ ), .Z(_05628_ ) );
INV_X1 _13388_ ( .A(_05628_ ), .ZN(_05629_ ) );
OAI21_X1 _13389_ ( .A(_05626_ ), .B1(_05202_ ), .B2(_05629_ ), .ZN(_05630_ ) );
NAND3_X1 _13390_ ( .A1(_03847_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_05229_ ), .ZN(_05631_ ) );
NAND3_X1 _13391_ ( .A1(_03847_ ), .A2(\mepc [4] ), .A3(_03851_ ), .ZN(_05632_ ) );
NAND3_X1 _13392_ ( .A1(_05255_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_03866_ ), .ZN(_05633_ ) );
NAND3_X1 _13393_ ( .A1(_05255_ ), .A2(\mtvec [4] ), .A3(_03841_ ), .ZN(_05634_ ) );
AND4_X1 _13394_ ( .A1(_05631_ ), .A2(_05632_ ), .A3(_05633_ ), .A4(_05634_ ), .ZN(_05635_ ) );
NAND3_X1 _13395_ ( .A1(_05249_ ), .A2(_03863_ ), .A3(_05635_ ), .ZN(_05636_ ) );
INV_X1 _13396_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_05637_ ) );
NAND3_X1 _13397_ ( .A1(_03814_ ), .A2(_03829_ ), .A3(_05637_ ), .ZN(_05638_ ) );
AND2_X1 _13398_ ( .A1(_05636_ ), .A2(_05638_ ), .ZN(_05639_ ) );
OAI211_X1 _13399_ ( .A(_05630_ ), .B(_05207_ ), .C1(_05208_ ), .C2(_05639_ ), .ZN(_05640_ ) );
XNOR2_X1 _13400_ ( .A(_02431_ ), .B(_02454_ ), .ZN(_05641_ ) );
AOI22_X1 _13401_ ( .A1(_05641_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05628_ ), .ZN(_05642_ ) );
AOI21_X1 _13402_ ( .A(_05601_ ), .B1(_05640_ ), .B2(_05642_ ), .ZN(_00141_ ) );
XOR2_X1 _13403_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .Z(_05643_ ) );
NAND2_X1 _13404_ ( .A1(_03905_ ), .A2(_03906_ ), .ZN(_05644_ ) );
XNOR2_X1 _13405_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_imm [3] ), .ZN(_05645_ ) );
XNOR2_X1 _13406_ ( .A(_05644_ ), .B(_05645_ ), .ZN(_05646_ ) );
MUX2_X1 _13407_ ( .A(_05643_ ), .B(_05646_ ), .S(_05175_ ), .Z(_05647_ ) );
OR2_X2 _13408_ ( .A1(_05647_ ), .A2(\ID_EX_typ [3] ), .ZN(_05648_ ) );
INV_X1 _13409_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_05649_ ) );
AND3_X1 _13410_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(_05649_ ), .ZN(_05650_ ) );
NAND3_X1 _13411_ ( .A1(_05316_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_03867_ ), .ZN(_05651_ ) );
NAND3_X1 _13412_ ( .A1(_05437_ ), .A2(\mepc [3] ), .A3(_05313_ ), .ZN(_05652_ ) );
NAND3_X1 _13413_ ( .A1(_05312_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_05291_ ), .ZN(_05653_ ) );
NAND3_X1 _13414_ ( .A1(_05317_ ), .A2(\mtvec [3] ), .A3(_03842_ ), .ZN(_05654_ ) );
AND4_X1 _13415_ ( .A1(_05651_ ), .A2(_05652_ ), .A3(_05653_ ), .A4(_05654_ ), .ZN(_05655_ ) );
AOI21_X1 _13416_ ( .A(_05650_ ), .B1(_05356_ ), .B2(_05655_ ), .ZN(_05656_ ) );
OAI211_X1 _13417_ ( .A(_05648_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05656_ ), .ZN(_05657_ ) );
OAI21_X1 _13418_ ( .A(_02427_ ), .B1(_02377_ ), .B2(_04511_ ), .ZN(_05658_ ) );
XNOR2_X1 _13419_ ( .A(_05658_ ), .B(_02353_ ), .ZN(_05659_ ) );
AOI22_X1 _13420_ ( .A1(_05659_ ), .A2(_05325_ ), .B1(_05326_ ), .B2(_05646_ ), .ZN(_05660_ ) );
AOI21_X1 _13421_ ( .A(_05601_ ), .B1(_05657_ ), .B2(_05660_ ), .ZN(_00142_ ) );
OR3_X1 _13422_ ( .A1(_03903_ ), .A2(_03904_ ), .A3(_03900_ ), .ZN(_05661_ ) );
AND2_X1 _13423_ ( .A1(_05661_ ), .A2(_03905_ ), .ZN(_05662_ ) );
AOI21_X1 _13424_ ( .A(\ID_EX_typ [3] ), .B1(_05263_ ), .B2(_05662_ ), .ZN(_05663_ ) );
INV_X1 _13425_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05664_ ) );
OAI21_X1 _13426_ ( .A(_05663_ ), .B1(_05664_ ), .B2(_05266_ ), .ZN(_05665_ ) );
NAND3_X1 _13427_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [2] ), .ZN(_05666_ ) );
NAND3_X1 _13428_ ( .A1(_05289_ ), .A2(\mepc [2] ), .A3(_05227_ ), .ZN(_05667_ ) );
NAND2_X1 _13429_ ( .A1(_05251_ ), .A2(_05667_ ), .ZN(_05668_ ) );
AND3_X1 _13430_ ( .A1(_05437_ ), .A2(\mycsreg.CSReg[3][2] ), .A3(_05287_ ), .ZN(_05669_ ) );
AND3_X1 _13431_ ( .A1(_05317_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_05224_ ), .ZN(_05670_ ) );
AND3_X1 _13432_ ( .A1(_03864_ ), .A2(\mtvec [2] ), .A3(_05439_ ), .ZN(_05671_ ) );
NOR4_X1 _13433_ ( .A1(_05668_ ), .A2(_05669_ ), .A3(_05670_ ), .A4(_05671_ ), .ZN(_05672_ ) );
OAI21_X1 _13434_ ( .A(_05666_ ), .B1(_05672_ ), .B2(_03871_ ), .ZN(_05673_ ) );
OAI211_X1 _13435_ ( .A(_05665_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05673_ ), .ZN(_05674_ ) );
OR3_X1 _13436_ ( .A1(_02425_ ), .A2(_02426_ ), .A3(_02378_ ), .ZN(_05675_ ) );
AND2_X1 _13437_ ( .A1(_05675_ ), .A2(_02427_ ), .ZN(_05676_ ) );
AOI22_X1 _13438_ ( .A1(_05676_ ), .A2(_05272_ ), .B1(_03780_ ), .B2(_05662_ ), .ZN(_05677_ ) );
AOI21_X1 _13439_ ( .A(_05601_ ), .B1(_05674_ ), .B2(_05677_ ), .ZN(_00143_ ) );
XOR2_X1 _13440_ ( .A(_03901_ ), .B(_03902_ ), .Z(_05678_ ) );
AOI21_X1 _13441_ ( .A(\ID_EX_typ [3] ), .B1(_05175_ ), .B2(_05678_ ), .ZN(_05679_ ) );
INV_X1 _13442_ ( .A(\ID_EX_pc [1] ), .ZN(_05680_ ) );
OAI21_X1 _13443_ ( .A(_05679_ ), .B1(_05680_ ), .B2(_05266_ ), .ZN(_05681_ ) );
NAND3_X1 _13444_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [1] ), .ZN(_05682_ ) );
NAND3_X1 _13445_ ( .A1(_05312_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_05291_ ), .ZN(_05683_ ) );
NAND3_X1 _13446_ ( .A1(_05312_ ), .A2(\mepc [1] ), .A3(_05314_ ), .ZN(_05684_ ) );
NAND3_X1 _13447_ ( .A1(_05317_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_05224_ ), .ZN(_05685_ ) );
NAND3_X1 _13448_ ( .A1(_05317_ ), .A2(\mtvec [1] ), .A3(_03842_ ), .ZN(_05686_ ) );
AND4_X1 _13449_ ( .A1(_05683_ ), .A2(_05684_ ), .A3(_05685_ ), .A4(_05686_ ), .ZN(_05687_ ) );
OAI21_X1 _13450_ ( .A(_05682_ ), .B1(_05687_ ), .B2(_03871_ ), .ZN(_05688_ ) );
OAI211_X1 _13451_ ( .A(_05681_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05688_ ), .ZN(_05689_ ) );
XOR2_X1 _13452_ ( .A(_02401_ ), .B(_02424_ ), .Z(_05690_ ) );
AOI22_X1 _13453_ ( .A1(_05690_ ), .A2(_05272_ ), .B1(_03780_ ), .B2(_05678_ ), .ZN(_05691_ ) );
AOI21_X1 _13454_ ( .A(_05601_ ), .B1(_05689_ ), .B2(_05691_ ), .ZN(_00144_ ) );
NAND3_X1 _13455_ ( .A1(_05192_ ), .A2(\ID_EX_pc [26] ), .A3(_05195_ ), .ZN(_05692_ ) );
XNOR2_X1 _13456_ ( .A(_05692_ ), .B(\ID_EX_pc [27] ), .ZN(_05693_ ) );
AOI21_X1 _13457_ ( .A(\ID_EX_typ [3] ), .B1(_05201_ ), .B2(_05693_ ), .ZN(_05694_ ) );
NOR2_X1 _13458_ ( .A1(_05222_ ), .A2(\EX_LS_result_csreg_mem [27] ), .ZN(_05695_ ) );
AND3_X1 _13459_ ( .A1(_05437_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_05287_ ), .ZN(_05696_ ) );
AND3_X1 _13460_ ( .A1(_05316_ ), .A2(\mtvec [27] ), .A3(_05439_ ), .ZN(_05697_ ) );
NOR3_X1 _13461_ ( .A1(_05696_ ), .A2(_05342_ ), .A3(_05697_ ), .ZN(_05698_ ) );
NAND3_X1 _13462_ ( .A1(_05437_ ), .A2(\mepc [27] ), .A3(_05313_ ), .ZN(_05699_ ) );
NAND3_X1 _13463_ ( .A1(_03864_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_03867_ ), .ZN(_05700_ ) );
NAND2_X1 _13464_ ( .A1(_05699_ ), .A2(_05700_ ), .ZN(_05701_ ) );
AOI21_X1 _13465_ ( .A(_05701_ ), .B1(_05238_ ), .B2(_05240_ ), .ZN(_05702_ ) );
AOI21_X1 _13466_ ( .A(_05695_ ), .B1(_05698_ ), .B2(_05702_ ), .ZN(_05703_ ) );
INV_X1 _13467_ ( .A(_05703_ ), .ZN(_05704_ ) );
AOI211_X1 _13468_ ( .A(_05184_ ), .B(_05694_ ), .C1(\ID_EX_typ [3] ), .C2(_05704_ ), .ZN(_05705_ ) );
NAND2_X1 _13469_ ( .A1(_03986_ ), .A2(_03988_ ), .ZN(_05706_ ) );
NAND2_X1 _13470_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_05707_ ) );
NAND2_X1 _13471_ ( .A1(_05706_ ), .A2(_05707_ ), .ZN(_05708_ ) );
XNOR2_X1 _13472_ ( .A(_05708_ ), .B(_03987_ ), .ZN(_05709_ ) );
OAI211_X1 _13473_ ( .A(_05263_ ), .B(_05180_ ), .C1(_05178_ ), .C2(_05703_ ), .ZN(_05710_ ) );
AOI21_X1 _13474_ ( .A(_05709_ ), .B1(_05710_ ), .B2(_03781_ ), .ZN(_05711_ ) );
NOR2_X1 _13475_ ( .A1(_05705_ ), .A2(_05711_ ), .ZN(_05712_ ) );
BUF_X2 _13476_ ( .A(_03779_ ), .Z(_05713_ ) );
OR3_X1 _13477_ ( .A1(_02974_ ), .A2(_05713_ ), .A3(_05181_ ), .ZN(_05714_ ) );
AOI21_X1 _13478_ ( .A(_05601_ ), .B1(_05712_ ), .B2(_05714_ ), .ZN(_00145_ ) );
AND3_X1 _13479_ ( .A1(_05346_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_05223_ ), .ZN(_05715_ ) );
AOI21_X1 _13480_ ( .A(_05715_ ), .B1(_05238_ ), .B2(_05240_ ), .ZN(_05716_ ) );
NAND3_X1 _13481_ ( .A1(_05312_ ), .A2(\mepc [0] ), .A3(_05314_ ), .ZN(_05717_ ) );
AND3_X1 _13482_ ( .A1(_05311_ ), .A2(\mycsreg.CSReg[3][0] ), .A3(_03856_ ), .ZN(_05718_ ) );
AND3_X1 _13483_ ( .A1(_05346_ ), .A2(\mtvec [0] ), .A3(_05439_ ), .ZN(_05719_ ) );
NOR3_X1 _13484_ ( .A1(_05718_ ), .A2(_05343_ ), .A3(_05719_ ), .ZN(_05720_ ) );
NAND3_X1 _13485_ ( .A1(_05716_ ), .A2(_05717_ ), .A3(_05720_ ), .ZN(_05721_ ) );
INV_X1 _13486_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_05722_ ) );
NAND3_X1 _13487_ ( .A1(_05492_ ), .A2(_05722_ ), .A3(_05493_ ), .ZN(_05723_ ) );
AND2_X1 _13488_ ( .A1(_05721_ ), .A2(_05723_ ), .ZN(_05724_ ) );
XOR2_X1 _13489_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05725_ ) );
MUX2_X1 _13490_ ( .A(\ID_EX_pc [0] ), .B(_05725_ ), .S(_05174_ ), .Z(_05726_ ) );
MUX2_X2 _13491_ ( .A(_05724_ ), .B(_05726_ ), .S(_05177_ ), .Z(_05727_ ) );
AOI22_X1 _13492_ ( .A1(_05727_ ), .A2(_05182_ ), .B1(_05274_ ), .B2(_05725_ ), .ZN(_05728_ ) );
NOR2_X1 _13493_ ( .A1(_05728_ ), .A2(_03801_ ), .ZN(_00146_ ) );
NAND2_X1 _13494_ ( .A1(_05192_ ), .A2(_05195_ ), .ZN(_05729_ ) );
XNOR2_X1 _13495_ ( .A(_05729_ ), .B(\ID_EX_pc [26] ), .ZN(_05730_ ) );
AOI21_X1 _13496_ ( .A(\ID_EX_typ [3] ), .B1(_05201_ ), .B2(_05730_ ), .ZN(_05731_ ) );
XOR2_X1 _13497_ ( .A(_03986_ ), .B(_03988_ ), .Z(_05732_ ) );
INV_X1 _13498_ ( .A(_05732_ ), .ZN(_05733_ ) );
OAI21_X1 _13499_ ( .A(_05731_ ), .B1(_05202_ ), .B2(_05733_ ), .ZN(_05734_ ) );
NAND3_X1 _13500_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [26] ), .ZN(_05735_ ) );
NAND3_X1 _13501_ ( .A1(_05437_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_05287_ ), .ZN(_05736_ ) );
NAND3_X1 _13502_ ( .A1(_05437_ ), .A2(\mepc [26] ), .A3(_05313_ ), .ZN(_05737_ ) );
NAND3_X1 _13503_ ( .A1(_05316_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_03867_ ), .ZN(_05738_ ) );
NAND3_X1 _13504_ ( .A1(_05316_ ), .A2(\mtvec [26] ), .A3(_05439_ ), .ZN(_05739_ ) );
AND4_X1 _13505_ ( .A1(_05736_ ), .A2(_05737_ ), .A3(_05738_ ), .A4(_05739_ ), .ZN(_05740_ ) );
OAI21_X1 _13506_ ( .A(_05735_ ), .B1(_05740_ ), .B2(_03871_ ), .ZN(_05741_ ) );
OAI211_X1 _13507_ ( .A(_05734_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05741_ ), .ZN(_05742_ ) );
AOI22_X1 _13508_ ( .A1(_02976_ ), .A2(_05272_ ), .B1(_03780_ ), .B2(_05732_ ), .ZN(_05743_ ) );
AOI21_X1 _13509_ ( .A(_05601_ ), .B1(_05742_ ), .B2(_05743_ ), .ZN(_00147_ ) );
NAND3_X1 _13510_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [25] ), .ZN(_05744_ ) );
NAND3_X1 _13511_ ( .A1(_05289_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_05291_ ), .ZN(_05745_ ) );
NAND3_X1 _13512_ ( .A1(_05289_ ), .A2(\mepc [25] ), .A3(_05227_ ), .ZN(_05746_ ) );
NAND3_X1 _13513_ ( .A1(_05317_ ), .A2(\mtvec [25] ), .A3(_03842_ ), .ZN(_05747_ ) );
NAND3_X1 _13514_ ( .A1(_05317_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_05224_ ), .ZN(_05748_ ) );
AND4_X1 _13515_ ( .A1(_05745_ ), .A2(_05746_ ), .A3(_05747_ ), .A4(_05748_ ), .ZN(_05749_ ) );
OAI21_X1 _13516_ ( .A(_05744_ ), .B1(_05749_ ), .B2(_03871_ ), .ZN(_05750_ ) );
AND3_X1 _13517_ ( .A1(_05194_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05751_ ) );
AND2_X1 _13518_ ( .A1(_05192_ ), .A2(_05751_ ), .ZN(_05752_ ) );
AND3_X1 _13519_ ( .A1(_05752_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05753_ ) );
NAND2_X1 _13520_ ( .A1(_05753_ ), .A2(\ID_EX_pc [24] ), .ZN(_05754_ ) );
XNOR2_X1 _13521_ ( .A(_05754_ ), .B(\ID_EX_pc [25] ), .ZN(_05755_ ) );
AND2_X1 _13522_ ( .A1(_05202_ ), .A2(_05755_ ), .ZN(_05756_ ) );
OR2_X1 _13523_ ( .A1(_03974_ ), .A2(_03981_ ), .ZN(_05757_ ) );
AND2_X1 _13524_ ( .A1(_05757_ ), .A2(_03894_ ), .ZN(_05758_ ) );
OR2_X1 _13525_ ( .A1(_05758_ ), .A2(_03983_ ), .ZN(_05759_ ) );
XNOR2_X1 _13526_ ( .A(_05759_ ), .B(_03893_ ), .ZN(_05760_ ) );
OAI21_X1 _13527_ ( .A(_05178_ ), .B1(_05202_ ), .B2(_05760_ ), .ZN(_05761_ ) );
OAI221_X1 _13528_ ( .A(_05543_ ), .B1(_05189_ ), .B2(_05750_ ), .C1(_05756_ ), .C2(_05761_ ), .ZN(_05762_ ) );
NOR2_X1 _13529_ ( .A1(_05760_ ), .A2(_03781_ ), .ZN(_05763_ ) );
NOR3_X1 _13530_ ( .A1(_02978_ ), .A2(_05713_ ), .A3(_05181_ ), .ZN(_05764_ ) );
NOR2_X1 _13531_ ( .A1(_05763_ ), .A2(_05764_ ), .ZN(_05765_ ) );
AOI21_X1 _13532_ ( .A(_05601_ ), .B1(_05762_ ), .B2(_05765_ ), .ZN(_00148_ ) );
NAND3_X1 _13533_ ( .A1(_05752_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05766_ ) );
XNOR2_X1 _13534_ ( .A(_05766_ ), .B(\ID_EX_pc [24] ), .ZN(_05767_ ) );
AOI21_X1 _13535_ ( .A(\ID_EX_typ [3] ), .B1(_05201_ ), .B2(_05767_ ), .ZN(_05768_ ) );
XOR2_X1 _13536_ ( .A(_05757_ ), .B(_03894_ ), .Z(_05769_ ) );
INV_X1 _13537_ ( .A(_05769_ ), .ZN(_05770_ ) );
OAI21_X1 _13538_ ( .A(_05768_ ), .B1(_05202_ ), .B2(_05770_ ), .ZN(_05771_ ) );
OR2_X1 _13539_ ( .A1(_05222_ ), .A2(\EX_LS_result_csreg_mem [24] ), .ZN(_05772_ ) );
AND3_X1 _13540_ ( .A1(_05346_ ), .A2(\mtvec [24] ), .A3(_03841_ ), .ZN(_05773_ ) );
AOI21_X1 _13541_ ( .A(_05773_ ), .B1(_05238_ ), .B2(_05240_ ), .ZN(_05774_ ) );
AND3_X1 _13542_ ( .A1(_03848_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_03856_ ), .ZN(_05775_ ) );
NOR3_X1 _13543_ ( .A1(_05775_ ), .A2(_05342_ ), .A3(_05343_ ), .ZN(_05776_ ) );
NAND3_X1 _13544_ ( .A1(_05311_ ), .A2(\mepc [24] ), .A3(_05313_ ), .ZN(_05777_ ) );
NAND3_X1 _13545_ ( .A1(_05316_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_05223_ ), .ZN(_05778_ ) );
AND2_X1 _13546_ ( .A1(_05777_ ), .A2(_05778_ ), .ZN(_05779_ ) );
NAND3_X1 _13547_ ( .A1(_05774_ ), .A2(_05776_ ), .A3(_05779_ ), .ZN(_05780_ ) );
AND2_X1 _13548_ ( .A1(_05772_ ), .A2(_05780_ ), .ZN(_05781_ ) );
OAI211_X1 _13549_ ( .A(_05771_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05781_ ), .ZN(_05782_ ) );
AOI22_X1 _13550_ ( .A1(_05769_ ), .A2(_05326_ ), .B1(_02979_ ), .B2(_05272_ ), .ZN(_05783_ ) );
AOI21_X1 _13551_ ( .A(_05601_ ), .B1(_05782_ ), .B2(_05783_ ), .ZN(_00149_ ) );
NAND3_X1 _13552_ ( .A1(_05192_ ), .A2(\ID_EX_pc [22] ), .A3(_05751_ ), .ZN(_05784_ ) );
XNOR2_X1 _13553_ ( .A(_05784_ ), .B(\ID_EX_pc [23] ), .ZN(_05785_ ) );
OAI21_X1 _13554_ ( .A(_05785_ ), .B1(_05170_ ), .B2(_05173_ ), .ZN(_05786_ ) );
INV_X1 _13555_ ( .A(_03969_ ), .ZN(_05787_ ) );
OAI21_X1 _13556_ ( .A(_03973_ ), .B1(_03958_ ), .B2(_03966_ ), .ZN(_05788_ ) );
AOI21_X1 _13557_ ( .A(_05787_ ), .B1(_05788_ ), .B2(_03979_ ), .ZN(_05789_ ) );
OR2_X1 _13558_ ( .A1(_05789_ ), .A2(_03975_ ), .ZN(_05790_ ) );
XNOR2_X1 _13559_ ( .A(_05790_ ), .B(_03968_ ), .ZN(_05791_ ) );
OAI211_X1 _13560_ ( .A(_05189_ ), .B(_05786_ ), .C1(_05202_ ), .C2(_05791_ ), .ZN(_05792_ ) );
NAND3_X1 _13561_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [23] ), .ZN(_05793_ ) );
NAND3_X1 _13562_ ( .A1(_05312_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_05291_ ), .ZN(_05794_ ) );
NAND3_X1 _13563_ ( .A1(_05312_ ), .A2(\mepc [23] ), .A3(_05314_ ), .ZN(_05795_ ) );
NAND3_X1 _13564_ ( .A1(_05317_ ), .A2(\mtvec [23] ), .A3(_03842_ ), .ZN(_05796_ ) );
NAND3_X1 _13565_ ( .A1(_05317_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_05224_ ), .ZN(_05797_ ) );
AND4_X1 _13566_ ( .A1(_05794_ ), .A2(_05795_ ), .A3(_05796_ ), .A4(_05797_ ), .ZN(_05798_ ) );
OAI21_X1 _13567_ ( .A(_05793_ ), .B1(_05798_ ), .B2(_03871_ ), .ZN(_05799_ ) );
OAI211_X1 _13568_ ( .A(_05792_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05799_ ), .ZN(_05800_ ) );
MUX2_X1 _13569_ ( .A(_05791_ ), .B(_02986_ ), .S(fanout_net_5 ), .Z(_05801_ ) );
OR2_X1 _13570_ ( .A1(_05801_ ), .A2(_05245_ ), .ZN(_05802_ ) );
AOI21_X1 _13571_ ( .A(_05601_ ), .B1(_05800_ ), .B2(_05802_ ), .ZN(_00150_ ) );
INV_X1 _13572_ ( .A(\ID_EX_pc [22] ), .ZN(_05803_ ) );
XNOR2_X1 _13573_ ( .A(_05752_ ), .B(_05803_ ), .ZN(_05804_ ) );
AND3_X1 _13574_ ( .A1(_05788_ ), .A2(_05787_ ), .A3(_03979_ ), .ZN(_05805_ ) );
NOR2_X1 _13575_ ( .A1(_05805_ ), .A2(_05789_ ), .ZN(_05806_ ) );
MUX2_X1 _13576_ ( .A(_05804_ ), .B(_05806_ ), .S(_05175_ ), .Z(_05807_ ) );
OR2_X2 _13577_ ( .A1(_05807_ ), .A2(\ID_EX_typ [3] ), .ZN(_05808_ ) );
NAND3_X1 _13578_ ( .A1(_03848_ ), .A2(\mepc [22] ), .A3(_03851_ ), .ZN(_05809_ ) );
NAND3_X1 _13579_ ( .A1(_05346_ ), .A2(\mtvec [22] ), .A3(_05439_ ), .ZN(_05810_ ) );
NAND2_X1 _13580_ ( .A1(_05809_ ), .A2(_05810_ ), .ZN(_05811_ ) );
AND3_X1 _13581_ ( .A1(_03848_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_05229_ ), .ZN(_05812_ ) );
AND3_X1 _13582_ ( .A1(_03837_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_05223_ ), .ZN(_05813_ ) );
NOR3_X1 _13583_ ( .A1(_05811_ ), .A2(_05812_ ), .A3(_05813_ ), .ZN(_05814_ ) );
NAND4_X1 _13584_ ( .A1(_05249_ ), .A2(_05814_ ), .A3(_03863_ ), .A4(_05251_ ), .ZN(_05815_ ) );
INV_X1 _13585_ ( .A(\EX_LS_result_csreg_mem [22] ), .ZN(_05816_ ) );
NAND3_X1 _13586_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(_05816_ ), .ZN(_05817_ ) );
AND2_X1 _13587_ ( .A1(_05815_ ), .A2(_05817_ ), .ZN(_05818_ ) );
OAI211_X1 _13588_ ( .A(_05808_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05818_ ), .ZN(_05819_ ) );
AND3_X1 _13589_ ( .A1(_02987_ ), .A2(_02982_ ), .A3(_05272_ ), .ZN(_05820_ ) );
AOI21_X1 _13590_ ( .A(_05820_ ), .B1(_05274_ ), .B2(_05806_ ), .ZN(_05821_ ) );
AOI21_X1 _13591_ ( .A(_03800_ ), .B1(_05819_ ), .B2(_05821_ ), .ZN(_00151_ ) );
NOR2_X1 _13592_ ( .A1(_05267_ ), .A2(_05268_ ), .ZN(_05822_ ) );
INV_X1 _13593_ ( .A(\ID_EX_pc [21] ), .ZN(_05823_ ) );
XNOR2_X1 _13594_ ( .A(_05822_ ), .B(_05823_ ), .ZN(_05824_ ) );
AOI21_X1 _13595_ ( .A(\ID_EX_typ [3] ), .B1(_05201_ ), .B2(_05824_ ), .ZN(_05825_ ) );
OAI21_X1 _13596_ ( .A(_03972_ ), .B1(_03958_ ), .B2(_03966_ ), .ZN(_05826_ ) );
NAND2_X1 _13597_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_05827_ ) );
NAND2_X1 _13598_ ( .A1(_05826_ ), .A2(_05827_ ), .ZN(_05828_ ) );
XNOR2_X1 _13599_ ( .A(_05828_ ), .B(_03971_ ), .ZN(_05829_ ) );
OAI21_X1 _13600_ ( .A(_05825_ ), .B1(_05202_ ), .B2(_05829_ ), .ZN(_05830_ ) );
NAND3_X1 _13601_ ( .A1(_03837_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_03866_ ), .ZN(_05831_ ) );
NAND3_X1 _13602_ ( .A1(_05252_ ), .A2(\mepc [21] ), .A3(_03851_ ), .ZN(_05832_ ) );
NAND3_X1 _13603_ ( .A1(_05252_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_05229_ ), .ZN(_05833_ ) );
NAND3_X1 _13604_ ( .A1(_05255_ ), .A2(\mtvec [21] ), .A3(_03841_ ), .ZN(_05834_ ) );
AND4_X1 _13605_ ( .A1(_05831_ ), .A2(_05832_ ), .A3(_05833_ ), .A4(_05834_ ), .ZN(_05835_ ) );
NAND3_X1 _13606_ ( .A1(_05249_ ), .A2(_03863_ ), .A3(_05835_ ), .ZN(_05836_ ) );
INV_X1 _13607_ ( .A(\EX_LS_result_csreg_mem [21] ), .ZN(_05837_ ) );
AND3_X1 _13608_ ( .A1(_03814_ ), .A2(_03829_ ), .A3(_05837_ ), .ZN(_05838_ ) );
INV_X1 _13609_ ( .A(_05838_ ), .ZN(_05839_ ) );
AND2_X1 _13610_ ( .A1(_05836_ ), .A2(_05839_ ), .ZN(_05840_ ) );
OAI211_X1 _13611_ ( .A(_05830_ ), .B(_05247_ ), .C1(_05248_ ), .C2(_05840_ ), .ZN(_05841_ ) );
NOR3_X1 _13612_ ( .A1(_02940_ ), .A2(_05499_ ), .A3(_05181_ ), .ZN(_05842_ ) );
NOR2_X1 _13613_ ( .A1(_05829_ ), .A2(_03781_ ), .ZN(_05843_ ) );
NOR2_X1 _13614_ ( .A1(_05842_ ), .A2(_05843_ ), .ZN(_05844_ ) );
AOI21_X1 _13615_ ( .A(_03800_ ), .B1(_05841_ ), .B2(_05844_ ), .ZN(_00152_ ) );
OAI21_X1 _13616_ ( .A(_03999_ ), .B1(_03996_ ), .B2(_03997_ ), .ZN(_05845_ ) );
NAND2_X1 _13617_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_05846_ ) );
AND2_X1 _13618_ ( .A1(_05845_ ), .A2(_05846_ ), .ZN(_05847_ ) );
XNOR2_X1 _13619_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_05848_ ) );
XNOR2_X1 _13620_ ( .A(_05847_ ), .B(_05848_ ), .ZN(_05849_ ) );
MUX2_X1 _13621_ ( .A(_05849_ ), .B(_02930_ ), .S(fanout_net_5 ), .Z(_05850_ ) );
OR2_X1 _13622_ ( .A1(_05850_ ), .A2(_05245_ ), .ZN(_05851_ ) );
BUF_X4 _13623_ ( .A(_03778_ ), .Z(_05852_ ) );
NAND3_X1 _13624_ ( .A1(_05437_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_03856_ ), .ZN(_05853_ ) );
NAND3_X1 _13625_ ( .A1(_05437_ ), .A2(\mepc [31] ), .A3(_05313_ ), .ZN(_05854_ ) );
NAND3_X1 _13626_ ( .A1(_05316_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_03867_ ), .ZN(_05855_ ) );
NAND3_X1 _13627_ ( .A1(_05316_ ), .A2(\mtvec [31] ), .A3(_05439_ ), .ZN(_05856_ ) );
NAND4_X1 _13628_ ( .A1(_05853_ ), .A2(_05854_ ), .A3(_05855_ ), .A4(_05856_ ), .ZN(_05857_ ) );
OR2_X1 _13629_ ( .A1(_05221_ ), .A2(_05857_ ), .ZN(_05858_ ) );
OAI21_X1 _13630_ ( .A(_05858_ ), .B1(\EX_LS_result_csreg_mem [31] ), .B2(_05222_ ), .ZN(_05859_ ) );
INV_X1 _13631_ ( .A(\ID_EX_pc [30] ), .ZN(_05860_ ) );
NOR2_X1 _13632_ ( .A1(_03890_ ), .A2(_05860_ ), .ZN(_05861_ ) );
XNOR2_X1 _13633_ ( .A(_05861_ ), .B(\ID_EX_pc [31] ), .ZN(_05862_ ) );
MUX2_X1 _13634_ ( .A(_05862_ ), .B(_05849_ ), .S(_05175_ ), .Z(_05863_ ) );
MUX2_X2 _13635_ ( .A(_05859_ ), .B(_05863_ ), .S(_05178_ ), .Z(_05864_ ) );
OAI211_X1 _13636_ ( .A(_05851_ ), .B(_03790_ ), .C1(_05852_ ), .C2(_05864_ ), .ZN(_00153_ ) );
AND3_X1 _13637_ ( .A1(_03797_ ), .A2(\ID_EX_pc [31] ), .A3(_03799_ ), .ZN(_00154_ ) );
AND3_X1 _13638_ ( .A1(_03797_ ), .A2(\ID_EX_pc [30] ), .A3(_03799_ ), .ZN(_00155_ ) );
AND3_X1 _13639_ ( .A1(_03797_ ), .A2(\ID_EX_pc [21] ), .A3(_03799_ ), .ZN(_00156_ ) );
AND3_X1 _13640_ ( .A1(_03797_ ), .A2(\ID_EX_pc [20] ), .A3(_03799_ ), .ZN(_00157_ ) );
AND3_X1 _13641_ ( .A1(_03797_ ), .A2(\ID_EX_pc [19] ), .A3(_03799_ ), .ZN(_00158_ ) );
CLKBUF_X2 _13642_ ( .A(_03787_ ), .Z(_05865_ ) );
CLKBUF_X2 _13643_ ( .A(_03788_ ), .Z(_05866_ ) );
AND3_X1 _13644_ ( .A1(_05865_ ), .A2(\ID_EX_pc [18] ), .A3(_05866_ ), .ZN(_00159_ ) );
AND3_X1 _13645_ ( .A1(_05865_ ), .A2(\ID_EX_pc [17] ), .A3(_05866_ ), .ZN(_00160_ ) );
AND3_X1 _13646_ ( .A1(_05865_ ), .A2(\ID_EX_pc [16] ), .A3(_05866_ ), .ZN(_00161_ ) );
AND3_X1 _13647_ ( .A1(_05865_ ), .A2(\ID_EX_pc [15] ), .A3(_05866_ ), .ZN(_00162_ ) );
AND3_X1 _13648_ ( .A1(_05865_ ), .A2(\ID_EX_pc [14] ), .A3(_05866_ ), .ZN(_00163_ ) );
AND3_X1 _13649_ ( .A1(_05865_ ), .A2(\ID_EX_pc [13] ), .A3(_05866_ ), .ZN(_00164_ ) );
AND3_X1 _13650_ ( .A1(_05865_ ), .A2(\ID_EX_pc [12] ), .A3(_05866_ ), .ZN(_00165_ ) );
AND3_X1 _13651_ ( .A1(_05865_ ), .A2(\ID_EX_pc [29] ), .A3(_05866_ ), .ZN(_00166_ ) );
AND3_X1 _13652_ ( .A1(_05865_ ), .A2(\ID_EX_pc [11] ), .A3(_05866_ ), .ZN(_00167_ ) );
AND3_X1 _13653_ ( .A1(_05865_ ), .A2(\ID_EX_pc [10] ), .A3(_05866_ ), .ZN(_00168_ ) );
CLKBUF_X2 _13654_ ( .A(_03787_ ), .Z(_05867_ ) );
CLKBUF_X2 _13655_ ( .A(_03788_ ), .Z(_05868_ ) );
AND3_X1 _13656_ ( .A1(_05867_ ), .A2(\ID_EX_pc [9] ), .A3(_05868_ ), .ZN(_00169_ ) );
AND3_X1 _13657_ ( .A1(_05867_ ), .A2(\ID_EX_pc [8] ), .A3(_05868_ ), .ZN(_00170_ ) );
AND3_X1 _13658_ ( .A1(_05867_ ), .A2(\ID_EX_pc [7] ), .A3(_05868_ ), .ZN(_00171_ ) );
AND3_X1 _13659_ ( .A1(_05867_ ), .A2(\ID_EX_pc [6] ), .A3(_05868_ ), .ZN(_00172_ ) );
AND3_X1 _13660_ ( .A1(_05867_ ), .A2(\ID_EX_pc [5] ), .A3(_05868_ ), .ZN(_00173_ ) );
AND3_X1 _13661_ ( .A1(_05867_ ), .A2(\ID_EX_pc [4] ), .A3(_05868_ ), .ZN(_00174_ ) );
AND3_X1 _13662_ ( .A1(_05867_ ), .A2(\ID_EX_pc [3] ), .A3(_05868_ ), .ZN(_00175_ ) );
AND3_X1 _13663_ ( .A1(_05867_ ), .A2(\ID_EX_pc [2] ), .A3(_05868_ ), .ZN(_00176_ ) );
AND3_X1 _13664_ ( .A1(_05867_ ), .A2(\ID_EX_pc [28] ), .A3(_05868_ ), .ZN(_00177_ ) );
AND3_X1 _13665_ ( .A1(_05867_ ), .A2(\ID_EX_pc [1] ), .A3(_05868_ ), .ZN(_00178_ ) );
CLKBUF_X2 _13666_ ( .A(_03787_ ), .Z(_05869_ ) );
CLKBUF_X2 _13667_ ( .A(_03788_ ), .Z(_05870_ ) );
AND3_X1 _13668_ ( .A1(_05869_ ), .A2(\ID_EX_pc [0] ), .A3(_05870_ ), .ZN(_00179_ ) );
AND3_X1 _13669_ ( .A1(_05869_ ), .A2(\ID_EX_pc [27] ), .A3(_05870_ ), .ZN(_00180_ ) );
AND3_X1 _13670_ ( .A1(_05869_ ), .A2(\ID_EX_pc [26] ), .A3(_05870_ ), .ZN(_00181_ ) );
AND3_X1 _13671_ ( .A1(_05869_ ), .A2(\ID_EX_pc [25] ), .A3(_05870_ ), .ZN(_00182_ ) );
AND3_X1 _13672_ ( .A1(_05869_ ), .A2(\ID_EX_pc [24] ), .A3(_05870_ ), .ZN(_00183_ ) );
AND3_X1 _13673_ ( .A1(_05869_ ), .A2(\ID_EX_pc [23] ), .A3(_05870_ ), .ZN(_00184_ ) );
AND3_X1 _13674_ ( .A1(_05869_ ), .A2(\ID_EX_pc [22] ), .A3(_05870_ ), .ZN(_00185_ ) );
AND3_X1 _13675_ ( .A1(_05869_ ), .A2(\ID_EX_typ [7] ), .A3(_05870_ ), .ZN(_00186_ ) );
AND3_X1 _13676_ ( .A1(_01923_ ), .A2(_03748_ ), .A3(EXU_valid_LSU ), .ZN(_05871_ ) );
NAND3_X1 _13677_ ( .A1(_01998_ ), .A2(\myclint.rvalid ), .A3(_02001_ ), .ZN(_05872_ ) );
OAI21_X1 _13678_ ( .A(_05872_ ), .B1(_03714_ ), .B2(io_master_arready ), .ZN(_05873_ ) );
INV_X1 _13679_ ( .A(_01884_ ), .ZN(_05874_ ) );
BUF_X2 _13680_ ( .A(_05874_ ), .Z(_05875_ ) );
BUF_X2 _13681_ ( .A(_05875_ ), .Z(_05876_ ) );
BUF_X2 _13682_ ( .A(_05876_ ), .Z(_05877_ ) );
BUF_X4 _13683_ ( .A(_05877_ ), .Z(_05878_ ) );
BUF_X4 _13684_ ( .A(_05878_ ), .Z(_05879_ ) );
OAI211_X1 _13685_ ( .A(_05871_ ), .B(_03790_ ), .C1(_05873_ ), .C2(_05879_ ), .ZN(_05880_ ) );
INV_X1 _13686_ ( .A(io_master_awready ), .ZN(_05881_ ) );
AND4_X1 _13687_ ( .A1(\EX_LS_flag [1] ), .A2(_01871_ ), .A3(_05881_ ), .A4(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_05882_ ) );
INV_X1 _13688_ ( .A(\mylsu.state [4] ), .ZN(_05883_ ) );
INV_X1 _13689_ ( .A(\mylsu.state [0] ), .ZN(_05884_ ) );
AOI21_X1 _13690_ ( .A(_05882_ ), .B1(_05883_ ), .B2(_05884_ ), .ZN(_05885_ ) );
AND2_X1 _13691_ ( .A1(_03790_ ), .A2(EXU_valid_LSU ), .ZN(_05886_ ) );
INV_X1 _13692_ ( .A(_05886_ ), .ZN(_05887_ ) );
OAI221_X1 _13693_ ( .A(_05880_ ), .B1(_03775_ ), .B2(_03800_ ), .C1(_05885_ ), .C2(_05887_ ), .ZN(_00187_ ) );
AND3_X1 _13694_ ( .A1(_05869_ ), .A2(\ID_EX_typ [6] ), .A3(_05870_ ), .ZN(_00188_ ) );
AND3_X1 _13695_ ( .A1(_05869_ ), .A2(\ID_EX_typ [5] ), .A3(_05870_ ), .ZN(_00189_ ) );
AND3_X1 _13696_ ( .A1(_03796_ ), .A2(\ID_EX_typ [4] ), .A3(_03798_ ), .ZN(_00190_ ) );
AND3_X1 _13697_ ( .A1(_03796_ ), .A2(\ID_EX_typ [3] ), .A3(_03798_ ), .ZN(_00191_ ) );
AND3_X1 _13698_ ( .A1(_03796_ ), .A2(fanout_net_6 ), .A3(_03798_ ), .ZN(_00192_ ) );
AND3_X1 _13699_ ( .A1(_03796_ ), .A2(\ID_EX_typ [1] ), .A3(_03798_ ), .ZN(_00193_ ) );
AND3_X1 _13700_ ( .A1(_03796_ ), .A2(fanout_net_5 ), .A3(_03798_ ), .ZN(_00194_ ) );
AND2_X1 _13701_ ( .A1(_01989_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_05888_ ) );
CLKBUF_X2 _13702_ ( .A(_05888_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _13703_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .ZN(_05889_ ) );
BUF_X2 _13704_ ( .A(_05889_ ), .Z(_05890_ ) );
AND3_X1 _13705_ ( .A1(_01989_ ), .A2(_05890_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00242_ ) );
CLKBUF_X2 _13706_ ( .A(_03636_ ), .Z(_05891_ ) );
BUF_X2 _13707_ ( .A(_05891_ ), .Z(_05892_ ) );
AND3_X1 _13708_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05892_ ), .A3(fanout_net_8 ), .ZN(_00243_ ) );
AND3_X1 _13709_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_12 ), .A3(_03655_ ), .ZN(_00244_ ) );
AND3_X1 _13710_ ( .A1(_03796_ ), .A2(\EX_LS_pc [2] ), .A3(_03798_ ), .ZN(_00282_ ) );
AND2_X1 _13711_ ( .A1(_03790_ ), .A2(fanout_net_44 ), .ZN(_00283_ ) );
INV_X1 _13712_ ( .A(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_05893_ ) );
AND3_X1 _13713_ ( .A1(_03787_ ), .A2(_05893_ ), .A3(_03788_ ), .ZN(_05894_ ) );
NOR2_X1 _13714_ ( .A1(fanout_net_44 ), .A2(\mylsu.state [1] ), .ZN(_05895_ ) );
NAND2_X1 _13715_ ( .A1(_05894_ ), .A2(_05895_ ), .ZN(_05896_ ) );
NOR2_X1 _13716_ ( .A1(_02013_ ), .A2(_02015_ ), .ZN(_05897_ ) );
AOI21_X1 _13717_ ( .A(_03748_ ), .B1(_05897_ ), .B2(_01870_ ), .ZN(_05898_ ) );
NOR3_X1 _13718_ ( .A1(_03732_ ), .A2(_05898_ ), .A3(_03740_ ), .ZN(_05899_ ) );
AOI21_X1 _13719_ ( .A(_05896_ ), .B1(_05899_ ), .B2(_01941_ ), .ZN(_00296_ ) );
INV_X1 _13720_ ( .A(_01941_ ), .ZN(_05900_ ) );
AOI21_X1 _13721_ ( .A(_05900_ ), .B1(_05215_ ), .B2(_05898_ ), .ZN(_05901_ ) );
AOI21_X1 _13722_ ( .A(_05896_ ), .B1(_05901_ ), .B2(_03745_ ), .ZN(_00297_ ) );
NAND3_X1 _13723_ ( .A1(_05897_ ), .A2(\EX_LS_flag [2] ), .A3(_01923_ ), .ZN(_05902_ ) );
NOR2_X1 _13724_ ( .A1(_05902_ ), .A2(_05896_ ), .ZN(_00298_ ) );
AOI21_X1 _13725_ ( .A(_05896_ ), .B1(_03734_ ), .B2(_01941_ ), .ZN(_00299_ ) );
AOI21_X1 _13726_ ( .A(_05896_ ), .B1(_03745_ ), .B2(_05902_ ), .ZN(_00300_ ) );
NAND2_X1 _13727_ ( .A1(_01926_ ), .A2(_01940_ ), .ZN(_05903_ ) );
INV_X1 _13728_ ( .A(_01945_ ), .ZN(_05904_ ) );
NOR3_X1 _13729_ ( .A1(_02015_ ), .A2(_01943_ ), .A3(_03748_ ), .ZN(_05905_ ) );
OAI21_X1 _13730_ ( .A(_05905_ ), .B1(_02013_ ), .B2(\EX_LS_flag [1] ), .ZN(_05906_ ) );
AND3_X1 _13731_ ( .A1(_05903_ ), .A2(_05904_ ), .A3(_05906_ ), .ZN(_05907_ ) );
NOR4_X1 _13732_ ( .A1(_05907_ ), .A2(_03793_ ), .A3(_01950_ ), .A4(_03740_ ), .ZN(_05908_ ) );
AND3_X1 _13733_ ( .A1(_05908_ ), .A2(_03790_ ), .A3(_05895_ ), .ZN(_00301_ ) );
INV_X1 _13734_ ( .A(_00283_ ), .ZN(_05909_ ) );
AND4_X1 _13735_ ( .A1(EXU_valid_LSU ), .A2(_03787_ ), .A3(_03788_ ), .A4(_05895_ ), .ZN(_05910_ ) );
NOR2_X1 _13736_ ( .A1(_01871_ ), .A2(\EX_LS_flag [1] ), .ZN(_05911_ ) );
OAI21_X1 _13737_ ( .A(_05910_ ), .B1(_05911_ ), .B2(_03735_ ), .ZN(_05912_ ) );
OAI21_X1 _13738_ ( .A(_05909_ ), .B1(_01945_ ), .B2(_05912_ ), .ZN(_00302_ ) );
CLKBUF_X2 _13739_ ( .A(_01918_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _13740_ ( .A(_01885_ ), .Z(_05913_ ) );
NOR3_X1 _13741_ ( .A1(_05913_ ), .A2(fanout_net_4 ), .A3(_03793_ ), .ZN(_05914_ ) );
INV_X1 _13742_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_05915_ ) );
INV_X1 _13743_ ( .A(_01888_ ), .ZN(_05916_ ) );
AOI211_X1 _13744_ ( .A(_05914_ ), .B(_05879_ ), .C1(_05915_ ), .C2(_05916_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _13745_ ( .A1(_05913_ ), .A2(fanout_net_3 ), .A3(_03793_ ), .ZN(_05917_ ) );
INV_X1 _13746_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_05918_ ) );
AOI211_X1 _13747_ ( .A(_05917_ ), .B(_05879_ ), .C1(_05918_ ), .C2(_05916_ ), .ZN(\io_master_araddr [0] ) );
BUF_X4 _13748_ ( .A(_05879_ ), .Z(_05919_ ) );
OR3_X1 _13749_ ( .A1(_05913_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(_03793_ ), .ZN(_05920_ ) );
BUF_X4 _13750_ ( .A(_01888_ ), .Z(_05921_ ) );
OAI21_X1 _13751_ ( .A(_05920_ ), .B1(\mylsu.araddr_tmp [15] ), .B2(_05921_ ), .ZN(_05922_ ) );
BUF_X4 _13752_ ( .A(_01883_ ), .Z(_05923_ ) );
BUF_X4 _13753_ ( .A(_05923_ ), .Z(_05924_ ) );
BUF_X4 _13754_ ( .A(_05924_ ), .Z(_05925_ ) );
OAI22_X1 _13755_ ( .A1(_05919_ ), .A2(_05922_ ), .B1(_03459_ ), .B2(_05925_ ), .ZN(\io_master_araddr [15] ) );
AND2_X1 _13756_ ( .A1(_01888_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .ZN(_05926_ ) );
AOI21_X1 _13757_ ( .A(_05926_ ), .B1(\mylsu.araddr_tmp [14] ), .B2(_05916_ ), .ZN(_05927_ ) );
OAI22_X1 _13758_ ( .A1(_05919_ ), .A2(_05927_ ), .B1(_01830_ ), .B2(_05925_ ), .ZN(\io_master_araddr [14] ) );
OR3_X1 _13759_ ( .A1(_05913_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(_03793_ ), .ZN(_05928_ ) );
OAI21_X1 _13760_ ( .A(_05928_ ), .B1(\mylsu.araddr_tmp [5] ), .B2(_05921_ ), .ZN(_05929_ ) );
OAI22_X1 _13761_ ( .A1(_05919_ ), .A2(_05929_ ), .B1(_03389_ ), .B2(_05925_ ), .ZN(\io_master_araddr [5] ) );
OR3_X1 _13762_ ( .A1(_05913_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(_03793_ ), .ZN(_05930_ ) );
OAI21_X1 _13763_ ( .A(_05930_ ), .B1(\mylsu.araddr_tmp [4] ), .B2(_05921_ ), .ZN(_05931_ ) );
BUF_X4 _13764_ ( .A(_01993_ ), .Z(_05932_ ) );
OAI22_X1 _13765_ ( .A1(_05919_ ), .A2(_05931_ ), .B1(_05892_ ), .B2(_05932_ ), .ZN(\io_master_araddr [4] ) );
OR3_X1 _13766_ ( .A1(_05913_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(_03793_ ), .ZN(_05933_ ) );
OAI21_X1 _13767_ ( .A(_05933_ ), .B1(\mylsu.araddr_tmp [3] ), .B2(_05921_ ), .ZN(_05934_ ) );
OAI22_X1 _13768_ ( .A1(_05919_ ), .A2(_05934_ ), .B1(_03655_ ), .B2(_05932_ ), .ZN(\io_master_araddr [3] ) );
INV_X1 _13769_ ( .A(_01897_ ), .ZN(\io_master_araddr [31] ) );
INV_X1 _13770_ ( .A(_01893_ ), .ZN(\io_master_araddr [30] ) );
INV_X1 _13771_ ( .A(_01974_ ), .ZN(\io_master_araddr [29] ) );
INV_X1 _13772_ ( .A(_01957_ ), .ZN(\io_master_araddr [28] ) );
INV_X1 _13773_ ( .A(_01978_ ), .ZN(\io_master_araddr [27] ) );
INV_X1 _13774_ ( .A(_01961_ ), .ZN(\io_master_araddr [26] ) );
INV_X1 _13775_ ( .A(_01901_ ), .ZN(\io_master_araddr [24] ) );
OR3_X1 _13776_ ( .A1(_05913_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(_03792_ ), .ZN(_05935_ ) );
OAI21_X1 _13777_ ( .A(_05935_ ), .B1(\mylsu.araddr_tmp [13] ), .B2(_05921_ ), .ZN(_05936_ ) );
OAI22_X1 _13778_ ( .A1(_05919_ ), .A2(_05936_ ), .B1(_01838_ ), .B2(_05932_ ), .ZN(\io_master_araddr [13] ) );
OAI221_X1 _13779_ ( .A(\IF_ID_pc [12] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01890_ ), .C2(_01891_ ), .ZN(_05937_ ) );
INV_X1 _13780_ ( .A(_01876_ ), .ZN(_05938_ ) );
OR3_X1 _13781_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(_03792_ ), .ZN(_05939_ ) );
OAI211_X1 _13782_ ( .A(_05938_ ), .B(_05939_ ), .C1(\mylsu.araddr_tmp [12] ), .C2(_01888_ ), .ZN(_05940_ ) );
OAI21_X1 _13783_ ( .A(_05937_ ), .B1(\io_master_arburst [0] ), .B2(_05940_ ), .ZN(\io_master_araddr [12] ) );
OR3_X1 _13784_ ( .A1(_05913_ ), .A2(\EX_LS_dest_csreg_mem [11] ), .A3(_03792_ ), .ZN(_05941_ ) );
OAI21_X1 _13785_ ( .A(_05941_ ), .B1(\mylsu.araddr_tmp [11] ), .B2(_05921_ ), .ZN(_05942_ ) );
OAI22_X1 _13786_ ( .A1(_05919_ ), .A2(_05942_ ), .B1(_01741_ ), .B2(_05932_ ), .ZN(\io_master_araddr [11] ) );
OR3_X1 _13787_ ( .A1(_05913_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(_03792_ ), .ZN(_05943_ ) );
OAI21_X1 _13788_ ( .A(_05943_ ), .B1(\mylsu.araddr_tmp [10] ), .B2(_05921_ ), .ZN(_05944_ ) );
OAI22_X1 _13789_ ( .A1(_05919_ ), .A2(_05944_ ), .B1(_03446_ ), .B2(_05932_ ), .ZN(\io_master_araddr [10] ) );
OR3_X1 _13790_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [9] ), .A3(_03792_ ), .ZN(_05945_ ) );
OAI21_X1 _13791_ ( .A(_05945_ ), .B1(\mylsu.araddr_tmp [9] ), .B2(_05921_ ), .ZN(_05946_ ) );
OAI22_X1 _13792_ ( .A1(_05919_ ), .A2(_05946_ ), .B1(_01686_ ), .B2(_05932_ ), .ZN(\io_master_araddr [9] ) );
OR3_X1 _13793_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [8] ), .A3(_03792_ ), .ZN(_05947_ ) );
OAI21_X1 _13794_ ( .A(_05947_ ), .B1(\mylsu.araddr_tmp [8] ), .B2(_05921_ ), .ZN(_05948_ ) );
OAI22_X1 _13795_ ( .A1(_05919_ ), .A2(_05948_ ), .B1(_03407_ ), .B2(_05932_ ), .ZN(\io_master_araddr [8] ) );
NOR3_X1 _13796_ ( .A1(_05913_ ), .A2(_03802_ ), .A3(_03793_ ), .ZN(_05949_ ) );
AOI21_X1 _13797_ ( .A(_05949_ ), .B1(_05916_ ), .B2(\mylsu.araddr_tmp [7] ), .ZN(_05950_ ) );
OAI22_X1 _13798_ ( .A1(_05879_ ), .A2(_05950_ ), .B1(_03404_ ), .B2(_05932_ ), .ZN(\io_master_araddr [7] ) );
OR3_X1 _13799_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [6] ), .A3(_03792_ ), .ZN(_05951_ ) );
OAI21_X1 _13800_ ( .A(_05951_ ), .B1(\mylsu.araddr_tmp [6] ), .B2(_05921_ ), .ZN(_05952_ ) );
OAI22_X1 _13801_ ( .A1(_05879_ ), .A2(_05952_ ), .B1(_01808_ ), .B2(_05932_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _13802_ ( .A1(_01885_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(_03792_ ), .ZN(_05953_ ) );
OAI211_X1 _13803_ ( .A(_05938_ ), .B(_05953_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01888_ ), .ZN(_05954_ ) );
NOR2_X1 _13804_ ( .A1(_01869_ ), .A2(_05954_ ), .ZN(_05955_ ) );
BUF_X4 _13805_ ( .A(_05955_ ), .Z(_05956_ ) );
BUF_X4 _13806_ ( .A(_05956_ ), .Z(_05957_ ) );
BUF_X2 _13807_ ( .A(_05957_ ), .Z(\io_master_araddr [2] ) );
CLKBUF_X2 _13808_ ( .A(_01884_ ), .Z(\io_master_arid [1] ) );
NOR3_X1 _13809_ ( .A1(\io_master_arburst [0] ), .A2(_01933_ ), .A3(_01876_ ), .ZN(\io_master_arsize [2] ) );
NOR3_X1 _13810_ ( .A1(\io_master_arburst [0] ), .A2(_01932_ ), .A3(_01876_ ), .ZN(\io_master_arsize [0] ) );
INV_X1 _13811_ ( .A(\EX_LS_typ [2] ), .ZN(_05958_ ) );
OAI22_X1 _13812_ ( .A1(_01867_ ), .A2(_01868_ ), .B1(_05958_ ), .B2(_01876_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _13813_ ( .A(_01953_ ), .B(_01990_ ), .C1(_01998_ ), .C2(_02001_ ), .ZN(io_master_arvalid ) );
AND2_X1 _13814_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ) );
AND2_X1 _13815_ ( .A1(_01944_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_05959_ ) );
BUF_X4 _13816_ ( .A(_05959_ ), .Z(_05960_ ) );
BUF_X4 _13817_ ( .A(_05960_ ), .Z(_05961_ ) );
MUX2_X1 _13818_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_05961_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _13819_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_05961_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _13820_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_05961_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _13821_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_05961_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _13822_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_05961_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _13823_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_05961_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _13824_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_05961_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _13825_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_05961_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _13826_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_05961_ ), .Z(\io_master_awaddr [15] ) );
BUF_X4 _13827_ ( .A(_05960_ ), .Z(_05962_ ) );
MUX2_X1 _13828_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_05962_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _13829_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_05962_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _13830_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_05962_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _13831_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_05962_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _13832_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_05962_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _13833_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_05962_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _13834_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_05962_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _13835_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_05962_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _13836_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_05962_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _13837_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_05962_ ), .Z(\io_master_awaddr [6] ) );
BUF_X4 _13838_ ( .A(_05960_ ), .Z(_05963_ ) );
MUX2_X1 _13839_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_05963_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _13840_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_05963_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _13841_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_05963_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _13842_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_05963_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _13843_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_05963_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _13844_ ( .A(\mylsu.awaddr_tmp [1] ), .B(fanout_net_4 ), .S(_05963_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _13845_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_3 ), .S(_05963_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _13846_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_05963_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _13847_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_05963_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _13848_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_05963_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _13849_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_05960_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _13850_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_05960_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _13851_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_05960_ ), .Z(\io_master_awaddr [22] ) );
AND3_X1 _13852_ ( .A1(_01949_ ), .A2(\EX_LS_typ [1] ), .A3(_01936_ ), .ZN(\io_master_awsize [0] ) );
NAND2_X1 _13853_ ( .A1(_01949_ ), .A2(_01936_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _13854_ ( .A1(_01941_ ), .A2(_01951_ ), .A3(_05961_ ), .ZN(_05964_ ) );
NAND2_X1 _13855_ ( .A1(_05964_ ), .A2(_05883_ ), .ZN(io_master_awvalid ) );
INV_X1 _13856_ ( .A(\mylsu.state [2] ), .ZN(_05965_ ) );
INV_X1 _13857_ ( .A(\mylsu.state [1] ), .ZN(_05966_ ) );
NAND4_X1 _13858_ ( .A1(_05964_ ), .A2(_05965_ ), .A3(_05883_ ), .A4(_05966_ ), .ZN(io_master_bready ) );
NOR3_X1 _13859_ ( .A1(_01875_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_05967_ ) );
INV_X1 _13860_ ( .A(fanout_net_44 ), .ZN(_05968_ ) );
BUF_X2 _13861_ ( .A(_05968_ ), .Z(_05969_ ) );
NOR2_X1 _13862_ ( .A1(_03711_ ), .A2(\io_master_rid [0] ), .ZN(_05970_ ) );
NAND4_X1 _13863_ ( .A1(_05970_ ), .A2(io_master_rlast ), .A3(_03709_ ), .A4(_03710_ ), .ZN(_05971_ ) );
AOI21_X1 _13864_ ( .A(_05878_ ), .B1(_03708_ ), .B2(_05971_ ), .ZN(_05972_ ) );
AOI21_X1 _13865_ ( .A(_05969_ ), .B1(_05972_ ), .B2(_03725_ ), .ZN(_05973_ ) );
NAND2_X1 _13866_ ( .A1(\io_master_bid [1] ), .A2(\io_master_bid [0] ), .ZN(_05974_ ) );
OR3_X1 _13867_ ( .A1(_05974_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bid [2] ), .ZN(_05975_ ) );
NOR2_X1 _13868_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_05976_ ) );
NAND2_X1 _13869_ ( .A1(_05976_ ), .A2(io_master_bvalid ), .ZN(_05977_ ) );
NOR2_X1 _13870_ ( .A1(_05975_ ), .A2(_05977_ ), .ZN(_05978_ ) );
INV_X1 _13871_ ( .A(_05978_ ), .ZN(_05979_ ) );
AOI211_X1 _13872_ ( .A(_05967_ ), .B(_05973_ ), .C1(\mylsu.state [1] ), .C2(_05979_ ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _13873_ ( .A(_01995_ ), .B(_01994_ ), .C1(_01998_ ), .C2(_02001_ ), .ZN(io_master_rready ) );
MUX2_X1 _13874_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_3 ), .Z(_05980_ ) );
CLKBUF_X2 _13875_ ( .A(_03818_ ), .Z(_05981_ ) );
AND2_X1 _13876_ ( .A1(_05980_ ), .A2(_05981_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _13877_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_3 ), .Z(_05982_ ) );
AND2_X1 _13878_ ( .A1(_05982_ ), .A2(_05981_ ), .ZN(\io_master_wdata [14] ) );
NOR3_X1 _13879_ ( .A1(_05615_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _13880_ ( .A1(_05637_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [4] ) );
NOR3_X1 _13881_ ( .A1(_05649_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [3] ) );
INV_X1 _13882_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_05983_ ) );
NOR3_X1 _13883_ ( .A1(_05983_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [2] ) );
INV_X1 _13884_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_05984_ ) );
NOR3_X1 _13885_ ( .A1(_05984_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [1] ) );
NOR3_X1 _13886_ ( .A1(_05722_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _13887_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_3 ), .Z(_05985_ ) );
AND2_X1 _13888_ ( .A1(_05985_ ), .A2(_05981_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _13889_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_3 ), .Z(_05986_ ) );
AND2_X1 _13890_ ( .A1(_05986_ ), .A2(_05981_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _13891_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_3 ), .Z(_05987_ ) );
AND2_X1 _13892_ ( .A1(_05987_ ), .A2(_05981_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _13893_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_3 ), .Z(_05988_ ) );
AND2_X1 _13894_ ( .A1(_05988_ ), .A2(_05981_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _13895_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_3 ), .Z(_05989_ ) );
AND2_X1 _13896_ ( .A1(_05989_ ), .A2(_05981_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _13897_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_3 ), .Z(_05990_ ) );
AND2_X1 _13898_ ( .A1(_05990_ ), .A2(_05981_ ), .ZN(\io_master_wdata [8] ) );
NOR3_X1 _13899_ ( .A1(_05567_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [7] ) );
NOR3_X1 _13900_ ( .A1(_05594_ ), .A2(fanout_net_3 ), .A3(fanout_net_4 ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _13901_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_3 ), .Z(_05991_ ) );
MUX2_X1 _13902_ ( .A(_05991_ ), .B(_05980_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _13903_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_3 ), .Z(_05992_ ) );
MUX2_X1 _13904_ ( .A(_05992_ ), .B(_05982_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [30] ) );
MUX2_X1 _13905_ ( .A(_05837_ ), .B(_05428_ ), .S(fanout_net_3 ), .Z(_05993_ ) );
NOR2_X1 _13906_ ( .A1(_03818_ ), .A2(fanout_net_3 ), .ZN(_05994_ ) );
INV_X1 _13907_ ( .A(_05994_ ), .ZN(_05995_ ) );
OAI22_X1 _13908_ ( .A1(_05993_ ), .A2(fanout_net_4 ), .B1(_05995_ ), .B2(_05615_ ), .ZN(\io_master_wdata [21] ) );
MUX2_X1 _13909_ ( .A(_05260_ ), .B(_05434_ ), .S(fanout_net_3 ), .Z(_05996_ ) );
OAI22_X1 _13910_ ( .A1(_05996_ ), .A2(fanout_net_4 ), .B1(_05995_ ), .B2(_05637_ ), .ZN(\io_master_wdata [20] ) );
INV_X1 _13911_ ( .A(\EX_LS_result_csreg_mem [19] ), .ZN(_05997_ ) );
MUX2_X1 _13912_ ( .A(_05997_ ), .B(_05469_ ), .S(fanout_net_3 ), .Z(_05998_ ) );
OAI22_X1 _13913_ ( .A1(_05998_ ), .A2(fanout_net_4 ), .B1(_05995_ ), .B2(_05649_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _13914_ ( .A(_03818_ ), .B1(_03771_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_05999_ ) );
NOR2_X1 _13915_ ( .A1(fanout_net_3 ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_06000_ ) );
OAI22_X1 _13916_ ( .A1(_05995_ ), .A2(_05983_ ), .B1(_05999_ ), .B2(_06000_ ), .ZN(\io_master_wdata [18] ) );
INV_X1 _13917_ ( .A(\EX_LS_result_csreg_mem [9] ), .ZN(_06001_ ) );
MUX2_X1 _13918_ ( .A(_05350_ ), .B(_06001_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06002_ ) );
OAI22_X1 _13919_ ( .A1(_06002_ ), .A2(fanout_net_4 ), .B1(_05995_ ), .B2(_05984_ ), .ZN(\io_master_wdata [17] ) );
MUX2_X1 _13920_ ( .A(_05364_ ), .B(_05544_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06003_ ) );
OAI22_X1 _13921_ ( .A1(_06003_ ), .A2(fanout_net_4 ), .B1(_05995_ ), .B2(_05722_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _13922_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06004_ ) );
MUX2_X1 _13923_ ( .A(_06004_ ), .B(_05985_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _13924_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06005_ ) );
MUX2_X1 _13925_ ( .A(_06005_ ), .B(_05986_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _13926_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06006_ ) );
MUX2_X1 _13927_ ( .A(_06006_ ), .B(_05987_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _13928_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06007_ ) );
MUX2_X1 _13929_ ( .A(_06007_ ), .B(_05988_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _13930_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06008_ ) );
MUX2_X1 _13931_ ( .A(_06008_ ), .B(_05989_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _13932_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06009_ ) );
MUX2_X1 _13933_ ( .A(_06009_ ), .B(_05990_ ), .S(fanout_net_4 ), .Z(\io_master_wdata [24] ) );
INV_X1 _13934_ ( .A(\EX_LS_result_csreg_mem [23] ), .ZN(_06010_ ) );
INV_X1 _13935_ ( .A(\EX_LS_result_csreg_mem [15] ), .ZN(_06011_ ) );
MUX2_X1 _13936_ ( .A(_06010_ ), .B(_06011_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06012_ ) );
OAI22_X1 _13937_ ( .A1(_06012_ ), .A2(fanout_net_4 ), .B1(_05995_ ), .B2(_05567_ ), .ZN(\io_master_wdata [23] ) );
MUX2_X1 _13938_ ( .A(_05816_ ), .B(_05404_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06013_ ) );
OAI22_X1 _13939_ ( .A1(_06013_ ), .A2(fanout_net_4 ), .B1(_05995_ ), .B2(_05594_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _13940_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06014_ ) );
AND2_X1 _13941_ ( .A1(_06014_ ), .A2(_05981_ ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _13942_ ( .A1(_03771_ ), .A2(_05981_ ), .A3(\EX_LS_typ [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _13943_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06015_ ) );
MUX2_X1 _13944_ ( .A(_06015_ ), .B(_06014_ ), .S(fanout_net_4 ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _13945_ ( .A1(_03818_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_06016_ ) );
NAND3_X1 _13946_ ( .A1(_03771_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_typ [0] ), .ZN(_06017_ ) );
OAI211_X1 _13947_ ( .A(_06016_ ), .B(_06017_ ), .C1(_01931_ ), .C2(_05958_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _13948_ ( .A1(_05964_ ), .A2(_05965_ ), .ZN(io_master_wvalid ) );
MUX2_X1 _13949_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _13950_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _13951_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _13952_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
INV_X1 _13953_ ( .A(_01952_ ), .ZN(_06018_ ) );
NOR2_X1 _13954_ ( .A1(_05897_ ), .A2(exception_quest_IDU ), .ZN(_06019_ ) );
NOR2_X1 _13955_ ( .A1(_06018_ ), .A2(_06019_ ), .ZN(_06020_ ) );
BUF_X4 _13956_ ( .A(_06020_ ), .Z(_06021_ ) );
MUX2_X1 _13957_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _13958_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _13959_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _13960_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _13961_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _13962_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _13963_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _13964_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _13965_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _13966_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_06021_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _13967_ ( .A(_06020_ ), .Z(_06022_ ) );
MUX2_X1 _13968_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _13969_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _13970_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _13971_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _13972_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _13973_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _13974_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _13975_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _13976_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _13977_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_06022_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _13978_ ( .A(_06020_ ), .Z(_06023_ ) );
MUX2_X1 _13979_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _13980_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _13981_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _13982_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _13983_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _13984_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _13985_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _13986_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _13987_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _13988_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_06023_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _13989_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_06020_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _13990_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_06020_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
OAI21_X1 _13991_ ( .A(_02017_ ), .B1(_06018_ ), .B2(_02016_ ), .ZN(_06024_ ) );
XNOR2_X1 _13992_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06025_ ) );
XNOR2_X1 _13993_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06026_ ) );
XNOR2_X1 _13994_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06027_ ) );
XNOR2_X1 _13995_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06028_ ) );
NAND4_X1 _13996_ ( .A1(_06025_ ), .A2(_06026_ ), .A3(_06027_ ), .A4(_06028_ ), .ZN(_06029_ ) );
XNOR2_X1 _13997_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_06030_ ) );
XNOR2_X1 _13998_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_06031_ ) );
XNOR2_X1 _13999_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_06032_ ) );
XNOR2_X1 _14000_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_06033_ ) );
NAND4_X1 _14001_ ( .A1(_06030_ ), .A2(_06031_ ), .A3(_06032_ ), .A4(_06033_ ), .ZN(_06034_ ) );
XNOR2_X1 _14002_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06035_ ) );
XNOR2_X1 _14003_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06036_ ) );
XNOR2_X1 _14004_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06037_ ) );
XNOR2_X1 _14005_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06038_ ) );
NAND4_X1 _14006_ ( .A1(_06035_ ), .A2(_06036_ ), .A3(_06037_ ), .A4(_06038_ ), .ZN(_06039_ ) );
XNOR2_X1 _14007_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06040_ ) );
XNOR2_X1 _14008_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06041_ ) );
XNOR2_X1 _14009_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06042_ ) );
XNOR2_X1 _14010_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06043_ ) );
NAND4_X1 _14011_ ( .A1(_06040_ ), .A2(_06041_ ), .A3(_06042_ ), .A4(_06043_ ), .ZN(_06044_ ) );
NOR4_X1 _14012_ ( .A1(_06029_ ), .A2(_06034_ ), .A3(_06039_ ), .A4(_06044_ ), .ZN(_06045_ ) );
XNOR2_X1 _14013_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06046_ ) );
XNOR2_X1 _14014_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06047_ ) );
XNOR2_X1 _14015_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06048_ ) );
XNOR2_X1 _14016_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06049_ ) );
XNOR2_X1 _14017_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06050_ ) );
AND4_X1 _14018_ ( .A1(_06047_ ), .A2(_06048_ ), .A3(_06049_ ), .A4(_06050_ ), .ZN(_06051_ ) );
XNOR2_X1 _14019_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06052_ ) );
XNOR2_X1 _14020_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06053_ ) );
AND2_X1 _14021_ ( .A1(_06052_ ), .A2(_06053_ ), .ZN(_06054_ ) );
XNOR2_X1 _14022_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06055_ ) );
AND4_X1 _14023_ ( .A1(_06046_ ), .A2(_06051_ ), .A3(_06054_ ), .A4(_06055_ ), .ZN(_06056_ ) );
XNOR2_X1 _14024_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06057_ ) );
XNOR2_X1 _14025_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06058_ ) );
XNOR2_X1 _14026_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06059_ ) );
XNOR2_X1 _14027_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06060_ ) );
AND4_X1 _14028_ ( .A1(_06057_ ), .A2(_06058_ ), .A3(_06059_ ), .A4(_06060_ ), .ZN(_06061_ ) );
XNOR2_X1 _14029_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06062_ ) );
XNOR2_X1 _14030_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06063_ ) );
XNOR2_X1 _14031_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06064_ ) );
XNOR2_X1 _14032_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06065_ ) );
AND4_X1 _14033_ ( .A1(_06062_ ), .A2(_06063_ ), .A3(_06064_ ), .A4(_06065_ ), .ZN(_06066_ ) );
NAND4_X1 _14034_ ( .A1(_06045_ ), .A2(_06056_ ), .A3(_06061_ ), .A4(_06066_ ), .ZN(_06067_ ) );
OR3_X1 _14035_ ( .A1(_06067_ ), .A2(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(_02017_ ), .ZN(_06068_ ) );
NAND2_X1 _14036_ ( .A1(_06024_ ), .A2(_06068_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14037_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_06069_ ) );
NOR2_X1 _14038_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06070_ ) );
NAND2_X1 _14039_ ( .A1(_06070_ ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06071_ ) );
NOR2_X1 _14040_ ( .A1(_06071_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06072_ ) );
NAND2_X1 _14041_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06073_ ) );
NOR3_X1 _14042_ ( .A1(_06073_ ), .A2(\LS_WB_waddr_csreg [11] ), .A3(\LS_WB_waddr_csreg [10] ), .ZN(_06074_ ) );
NOR2_X1 _14043_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_06075_ ) );
AND3_X1 _14044_ ( .A1(_06072_ ), .A2(_06074_ ), .A3(_06075_ ), .ZN(_06076_ ) );
NOR3_X1 _14045_ ( .A1(reset ), .A2(excp_written ), .A3(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_B ), .ZN(_06077_ ) );
AND4_X1 _14046_ ( .A1(_06069_ ), .A2(_06076_ ), .A3(\LS_WB_waddr_csreg [0] ), .A4(_06077_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14047_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .A3(\LS_WB_waddr_csreg [5] ), .A4(\LS_WB_waddr_csreg [4] ), .ZN(_06078_ ) );
NOR4_X1 _14048_ ( .A1(\LS_WB_waddr_csreg [1] ), .A2(\LS_WB_waddr_csreg [0] ), .A3(\LS_WB_waddr_csreg [3] ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_06079_ ) );
AND4_X1 _14049_ ( .A1(_06077_ ), .A2(_06078_ ), .A3(_06079_ ), .A4(_06074_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _14050_ ( .A1(_06078_ ), .A2(_06074_ ), .ZN(_06080_ ) );
NAND3_X1 _14051_ ( .A1(_06077_ ), .A2(_06069_ ), .A3(\LS_WB_waddr_csreg [0] ), .ZN(_06081_ ) );
INV_X1 _14052_ ( .A(\LS_WB_waddr_csreg [2] ), .ZN(_06082_ ) );
NOR4_X1 _14053_ ( .A1(_06080_ ), .A2(_06081_ ), .A3(\LS_WB_waddr_csreg [3] ), .A4(_06082_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND3_X1 _14054_ ( .A1(_01459_ ), .A2(\LS_WB_wen_csreg [7] ), .A3(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06083_ ) );
NOR4_X1 _14055_ ( .A1(_06069_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(\LS_WB_waddr_csreg [3] ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_06084_ ) );
NAND3_X1 _14056_ ( .A1(_06072_ ), .A2(_06074_ ), .A3(_06084_ ), .ZN(_06085_ ) );
AOI21_X1 _14057_ ( .A(_06083_ ), .B1(_06085_ ), .B2(_02004_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NAND2_X1 _14058_ ( .A1(_05690_ ), .A2(_02934_ ), .ZN(_06086_ ) );
AND2_X1 _14059_ ( .A1(_02931_ ), .A2(_03782_ ), .ZN(_06087_ ) );
BUF_X4 _14060_ ( .A(_06087_ ), .Z(_06088_ ) );
INV_X1 _14061_ ( .A(_06088_ ), .ZN(_06089_ ) );
BUF_X4 _14062_ ( .A(_06089_ ), .Z(_06090_ ) );
BUF_X4 _14063_ ( .A(_06090_ ), .Z(_06091_ ) );
OAI21_X1 _14064_ ( .A(_06086_ ), .B1(_03865_ ), .B2(_06091_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _14065_ ( .A(_04486_ ), .B(\ID_EX_imm [0] ), .ZN(_06092_ ) );
BUF_X4 _14066_ ( .A(_06088_ ), .Z(_06093_ ) );
BUF_X4 _14067_ ( .A(_06093_ ), .Z(_06094_ ) );
AOI22_X1 _14068_ ( .A1(_06092_ ), .A2(_02935_ ), .B1(_03805_ ), .B2(_06094_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND2_X2 _14069_ ( .A1(_03258_ ), .A2(\ID_EX_typ [7] ), .ZN(_06095_ ) );
INV_X1 _14070_ ( .A(_06095_ ), .ZN(_06096_ ) );
BUF_X4 _14071_ ( .A(_06096_ ), .Z(_06097_ ) );
AND2_X1 _14072_ ( .A1(_05518_ ), .A2(_06097_ ), .ZN(_06098_ ) );
BUF_X4 _14073_ ( .A(_06089_ ), .Z(_06099_ ) );
MUX2_X1 _14074_ ( .A(\ID_EX_csr [10] ), .B(_06098_ ), .S(_06099_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
NOR4_X1 _14075_ ( .A1(_03259_ ), .A2(_03791_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [9] ), .ZN(_06100_ ) );
AOI21_X1 _14076_ ( .A(_06100_ ), .B1(_05540_ ), .B2(_02935_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR2_X1 _14077_ ( .A1(_05559_ ), .A2(_06095_ ), .ZN(_06101_ ) );
MUX2_X1 _14078_ ( .A(\ID_EX_csr [8] ), .B(_06101_ ), .S(_06099_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _14079_ ( .A1(_05579_ ), .A2(_02934_ ), .ZN(_06102_ ) );
OAI21_X1 _14080_ ( .A(_06102_ ), .B1(_03806_ ), .B2(_06091_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
AOI21_X1 _14081_ ( .A(_02931_ ), .B1(_05598_ ), .B2(_05577_ ), .ZN(_06103_ ) );
BUF_X4 _14082_ ( .A(_06088_ ), .Z(_06104_ ) );
BUF_X4 _14083_ ( .A(_06104_ ), .Z(_06105_ ) );
AOI21_X1 _14084_ ( .A(_06103_ ), .B1(_03844_ ), .B2(_06105_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14085_ ( .A1(_05622_ ), .A2(_02934_ ), .ZN(_06106_ ) );
OAI21_X1 _14086_ ( .A(_06106_ ), .B1(_03816_ ), .B2(_06091_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _14087_ ( .A1(_05641_ ), .A2(_02934_ ), .ZN(_06107_ ) );
OAI21_X1 _14088_ ( .A(_06107_ ), .B1(_03824_ ), .B2(_06091_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _14089_ ( .A1(_05659_ ), .A2(_02934_ ), .ZN(_06108_ ) );
OAI21_X1 _14090_ ( .A(_06108_ ), .B1(_03821_ ), .B2(_06091_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _14091_ ( .A1(_05675_ ), .A2(_02934_ ), .A3(_02427_ ), .ZN(_06109_ ) );
OAI21_X1 _14092_ ( .A(_06109_ ), .B1(_03853_ ), .B2(_06091_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
NAND2_X1 _14093_ ( .A1(_05478_ ), .A2(_02934_ ), .ZN(_06110_ ) );
OAI21_X1 _14094_ ( .A(_06110_ ), .B1(_03834_ ), .B2(_06091_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X4 _14095_ ( .A(_06093_ ), .Z(_06111_ ) );
INV_X1 _14096_ ( .A(_05840_ ), .ZN(_06112_ ) );
AOI22_X1 _14097_ ( .A1(_06112_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02206_ ), .ZN(_06113_ ) );
NAND3_X1 _14098_ ( .A1(_02205_ ), .A2(_02227_ ), .A3(_05186_ ), .ZN(_06114_ ) );
AND2_X1 _14099_ ( .A1(_06113_ ), .A2(_06114_ ), .ZN(_06115_ ) );
NOR2_X1 _14100_ ( .A1(_04824_ ), .A2(fanout_net_6 ), .ZN(_06116_ ) );
INV_X1 _14101_ ( .A(_06116_ ), .ZN(_06117_ ) );
AOI211_X1 _14102_ ( .A(_06117_ ), .B(_05838_ ), .C1(_05356_ ), .C2(_05835_ ), .ZN(_06118_ ) );
OAI21_X1 _14103_ ( .A(_06111_ ), .B1(_06115_ ), .B2(_06118_ ), .ZN(_06119_ ) );
MUX2_X1 _14104_ ( .A(_05823_ ), .B(_04112_ ), .S(_06097_ ), .Z(_06120_ ) );
OAI21_X1 _14105_ ( .A(_06119_ ), .B1(_06105_ ), .B2(_06120_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
INV_X1 _14106_ ( .A(_05262_ ), .ZN(_06121_ ) );
AOI22_X1 _14107_ ( .A1(_06121_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02203_ ), .ZN(_06122_ ) );
NAND3_X1 _14108_ ( .A1(_02182_ ), .A2(_02201_ ), .A3(_05186_ ), .ZN(_06123_ ) );
AND2_X1 _14109_ ( .A1(_06122_ ), .A2(_06123_ ), .ZN(_06124_ ) );
BUF_X4 _14110_ ( .A(_06116_ ), .Z(_06125_ ) );
AND3_X1 _14111_ ( .A1(_05259_ ), .A2(_06125_ ), .A3(_05261_ ), .ZN(_06126_ ) );
OAI21_X1 _14112_ ( .A(_06111_ ), .B1(_06124_ ), .B2(_06126_ ), .ZN(_06127_ ) );
MUX2_X1 _14113_ ( .A(_05268_ ), .B(_04139_ ), .S(_06097_ ), .Z(_06128_ ) );
OAI21_X1 _14114_ ( .A(_06127_ ), .B1(_06105_ ), .B2(_06128_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
AOI21_X1 _14115_ ( .A(_06117_ ), .B1(_05295_ ), .B2(_05296_ ), .ZN(_06129_ ) );
AOI22_X1 _14116_ ( .A1(_05297_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02253_ ), .ZN(_06130_ ) );
NAND3_X1 _14117_ ( .A1(_02250_ ), .A2(_02251_ ), .A3(_05300_ ), .ZN(_06131_ ) );
AOI211_X1 _14118_ ( .A(_06090_ ), .B(_06129_ ), .C1(_06130_ ), .C2(_06131_ ), .ZN(_06132_ ) );
BUF_X4 _14119_ ( .A(_06096_ ), .Z(_06133_ ) );
MUX2_X1 _14120_ ( .A(_05283_ ), .B(_04166_ ), .S(_06133_ ), .Z(_06134_ ) );
AOI21_X1 _14121_ ( .A(_06132_ ), .B1(_06134_ ), .B2(_06091_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
BUF_X4 _14122_ ( .A(_06125_ ), .Z(_06135_ ) );
BUF_X4 _14123_ ( .A(_06088_ ), .Z(_06136_ ) );
NAND3_X1 _14124_ ( .A1(_05323_ ), .A2(_06135_ ), .A3(_06136_ ), .ZN(_06137_ ) );
BUF_X4 _14125_ ( .A(_04826_ ), .Z(_06138_ ) );
OAI221_X1 _14126_ ( .A(_06093_ ), .B1(_05713_ ), .B2(\ID_EX_imm [18] ), .C1(_05323_ ), .C2(_06138_ ), .ZN(_06139_ ) );
AND3_X1 _14127_ ( .A1(_02255_ ), .A2(_05713_ ), .A3(_02274_ ), .ZN(_06140_ ) );
MUX2_X1 _14128_ ( .A(_05303_ ), .B(_04189_ ), .S(_06097_ ), .Z(_06141_ ) );
OAI221_X1 _14129_ ( .A(_06137_ ), .B1(_06139_ ), .B2(_06140_ ), .C1(_06141_ ), .C2(_06094_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
AND3_X1 _14130_ ( .A1(_03848_ ), .A2(\mepc [17] ), .A3(_03851_ ), .ZN(_06142_ ) );
AND3_X1 _14131_ ( .A1(_03837_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_03866_ ), .ZN(_06143_ ) );
NOR4_X1 _14132_ ( .A1(_05341_ ), .A2(_06142_ ), .A3(_06143_ ), .A4(_05339_ ), .ZN(_06144_ ) );
AND3_X1 _14133_ ( .A1(_05356_ ), .A2(_05251_ ), .A3(_06144_ ), .ZN(_06145_ ) );
AND3_X1 _14134_ ( .A1(_03815_ ), .A2(_03830_ ), .A3(_05350_ ), .ZN(_06146_ ) );
NOR3_X1 _14135_ ( .A1(_06145_ ), .A2(_06117_ ), .A3(_06146_ ), .ZN(_06147_ ) );
INV_X1 _14136_ ( .A(_05352_ ), .ZN(_06148_ ) );
AOI22_X1 _14137_ ( .A1(_06148_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02300_ ), .ZN(_06149_ ) );
NAND3_X1 _14138_ ( .A1(_02279_ ), .A2(_02298_ ), .A3(_05186_ ), .ZN(_06150_ ) );
AOI21_X1 _14139_ ( .A(_06147_ ), .B1(_06149_ ), .B2(_06150_ ), .ZN(_06151_ ) );
BUF_X4 _14140_ ( .A(_06088_ ), .Z(_06152_ ) );
NAND2_X1 _14141_ ( .A1(_06151_ ), .A2(_06152_ ), .ZN(_06153_ ) );
NAND4_X1 _14142_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06154_ ) );
OAI211_X1 _14143_ ( .A(_06099_ ), .B(_06154_ ), .C1(_04240_ ), .C2(_06095_ ), .ZN(_06155_ ) );
AND2_X1 _14144_ ( .A1(_06153_ ), .A2(_06155_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
BUF_X4 _14145_ ( .A(_06088_ ), .Z(_06156_ ) );
INV_X1 _14146_ ( .A(_05366_ ), .ZN(_06157_ ) );
AOI22_X1 _14147_ ( .A1(_06157_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02323_ ), .ZN(_06158_ ) );
NAND3_X1 _14148_ ( .A1(_02302_ ), .A2(_02321_ ), .A3(_05186_ ), .ZN(_06159_ ) );
AND2_X1 _14149_ ( .A1(_06158_ ), .A2(_06159_ ), .ZN(_06160_ ) );
AND3_X1 _14150_ ( .A1(_05363_ ), .A2(_06116_ ), .A3(_05365_ ), .ZN(_06161_ ) );
OAI21_X1 _14151_ ( .A(_06156_ ), .B1(_06160_ ), .B2(_06161_ ), .ZN(_06162_ ) );
MUX2_X1 _14152_ ( .A(_05335_ ), .B(_04217_ ), .S(_06097_ ), .Z(_06163_ ) );
OAI21_X1 _14153_ ( .A(_06162_ ), .B1(_06105_ ), .B2(_06163_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
BUF_X4 _14154_ ( .A(_06090_ ), .Z(_06164_ ) );
AOI21_X1 _14155_ ( .A(_06095_ ), .B1(_04584_ ), .B2(_04604_ ), .ZN(_06165_ ) );
CLKBUF_X2 _14156_ ( .A(_03258_ ), .Z(_06166_ ) );
AND3_X1 _14157_ ( .A1(_06166_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_typ [7] ), .ZN(_06167_ ) );
OAI21_X1 _14158_ ( .A(_06164_ ), .B1(_06165_ ), .B2(_06167_ ), .ZN(_06168_ ) );
AND3_X1 _14159_ ( .A1(_05492_ ), .A2(_06011_ ), .A3(_05493_ ), .ZN(_06169_ ) );
AND3_X1 _14160_ ( .A1(_03838_ ), .A2(\mtvec [15] ), .A3(_03842_ ), .ZN(_06170_ ) );
NOR4_X1 _14161_ ( .A1(_05374_ ), .A2(_05375_ ), .A3(_05343_ ), .A4(_06170_ ), .ZN(_06171_ ) );
AOI21_X1 _14162_ ( .A(_05376_ ), .B1(_05468_ ), .B2(_05470_ ), .ZN(_06172_ ) );
AOI21_X1 _14163_ ( .A(_06169_ ), .B1(_06171_ ), .B2(_06172_ ), .ZN(_06173_ ) );
AOI21_X1 _14164_ ( .A(fanout_net_5 ), .B1(_02589_ ), .B2(_02608_ ), .ZN(_06174_ ) );
AND2_X1 _14165_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [15] ), .ZN(_06175_ ) );
OAI221_X1 _14166_ ( .A(_06136_ ), .B1(_06138_ ), .B2(_06173_ ), .C1(_06174_ ), .C2(_06175_ ), .ZN(_06176_ ) );
NAND3_X1 _14167_ ( .A1(_05312_ ), .A2(\mepc [15] ), .A3(_05314_ ), .ZN(_06177_ ) );
NOR3_X1 _14168_ ( .A1(_05375_ ), .A2(_05343_ ), .A3(_06170_ ), .ZN(_06178_ ) );
NAND3_X1 _14169_ ( .A1(_06172_ ), .A2(_06177_ ), .A3(_06178_ ), .ZN(_06179_ ) );
NAND3_X1 _14170_ ( .A1(_05468_ ), .A2(_06011_ ), .A3(_05470_ ), .ZN(_06180_ ) );
NAND4_X1 _14171_ ( .A1(_06179_ ), .A2(_06135_ ), .A3(_06180_ ), .A4(_06136_ ), .ZN(_06181_ ) );
NAND3_X1 _14172_ ( .A1(_06168_ ), .A2(_06176_ ), .A3(_06181_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
NAND2_X1 _14173_ ( .A1(_05403_ ), .A2(_05405_ ), .ZN(_06182_ ) );
AOI22_X1 _14174_ ( .A1(_06182_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02632_ ), .ZN(_06183_ ) );
NAND3_X1 _14175_ ( .A1(_02611_ ), .A2(_02630_ ), .A3(_05186_ ), .ZN(_06184_ ) );
AND2_X1 _14176_ ( .A1(_06183_ ), .A2(_06184_ ), .ZN(_06185_ ) );
AND3_X1 _14177_ ( .A1(_05403_ ), .A2(_06116_ ), .A3(_05405_ ), .ZN(_06186_ ) );
OAI21_X1 _14178_ ( .A(_06156_ ), .B1(_06185_ ), .B2(_06186_ ), .ZN(_06187_ ) );
MUX2_X1 _14179_ ( .A(_05407_ ), .B(_04628_ ), .S(_06097_ ), .Z(_06188_ ) );
OAI21_X1 _14180_ ( .A(_06187_ ), .B1(_06105_ ), .B2(_06188_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OAI22_X1 _14181_ ( .A1(_05430_ ), .A2(_04826_ ), .B1(_03779_ ), .B2(\ID_EX_imm [13] ), .ZN(_06189_ ) );
AOI21_X1 _14182_ ( .A(_06189_ ), .B1(_05186_ ), .B2(_04914_ ), .ZN(_06190_ ) );
NAND3_X1 _14183_ ( .A1(_05427_ ), .A2(_06116_ ), .A3(_05429_ ), .ZN(_06191_ ) );
INV_X1 _14184_ ( .A(_06191_ ), .ZN(_06192_ ) );
OR3_X1 _14185_ ( .A1(_06190_ ), .A2(_06089_ ), .A3(_06192_ ), .ZN(_06193_ ) );
NAND4_X1 _14186_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06194_ ) );
OAI211_X1 _14187_ ( .A(_06099_ ), .B(_06194_ ), .C1(_04578_ ), .C2(_06095_ ), .ZN(_06195_ ) );
AND2_X1 _14188_ ( .A1(_06193_ ), .A2(_06195_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _14189_ ( .A1(_05226_ ), .A2(\mepc [12] ), .A3(_05227_ ), .ZN(_06196_ ) );
NAND3_X1 _14190_ ( .A1(_03838_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_05224_ ), .ZN(_06197_ ) );
NAND2_X1 _14191_ ( .A1(_06196_ ), .A2(_06197_ ), .ZN(_06198_ ) );
AOI21_X1 _14192_ ( .A(_06198_ ), .B1(_05492_ ), .B2(_05493_ ), .ZN(_06199_ ) );
INV_X1 _14193_ ( .A(_05440_ ), .ZN(_06200_ ) );
NOR3_X1 _14194_ ( .A1(_05436_ ), .A2(_05342_ ), .A3(_05343_ ), .ZN(_06201_ ) );
NAND3_X1 _14195_ ( .A1(_06199_ ), .A2(_06200_ ), .A3(_06201_ ), .ZN(_06202_ ) );
AND3_X1 _14196_ ( .A1(_05492_ ), .A2(_05434_ ), .A3(_05493_ ), .ZN(_06203_ ) );
INV_X1 _14197_ ( .A(_06203_ ), .ZN(_06204_ ) );
NAND2_X1 _14198_ ( .A1(_06202_ ), .A2(_06204_ ), .ZN(_06205_ ) );
AOI22_X1 _14199_ ( .A1(_06205_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02562_ ), .ZN(_06206_ ) );
BUF_X4 _14200_ ( .A(_06088_ ), .Z(_06207_ ) );
OAI211_X1 _14201_ ( .A(_06206_ ), .B(_06207_ ), .C1(fanout_net_5 ), .C2(_02561_ ), .ZN(_06208_ ) );
NAND4_X1 _14202_ ( .A1(_06202_ ), .A2(_06135_ ), .A3(_06204_ ), .A4(_06104_ ), .ZN(_06209_ ) );
MUX2_X1 _14203_ ( .A(_05444_ ), .B(_04556_ ), .S(_06133_ ), .Z(_06210_ ) );
BUF_X4 _14204_ ( .A(_06093_ ), .Z(_06211_ ) );
OAI211_X1 _14205_ ( .A(_06208_ ), .B(_06209_ ), .C1(_06210_ ), .C2(_06211_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
NAND3_X1 _14206_ ( .A1(_03872_ ), .A2(_06135_ ), .A3(_06136_ ), .ZN(_06212_ ) );
AND3_X1 _14207_ ( .A1(_02046_ ), .A2(_05713_ ), .A3(_02089_ ), .ZN(_06213_ ) );
OAI221_X1 _14208_ ( .A(_06093_ ), .B1(_05713_ ), .B2(\ID_EX_imm [30] ), .C1(_03872_ ), .C2(_06138_ ), .ZN(_06214_ ) );
AND4_X1 _14209_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06215_ ) );
BUF_X4 _14210_ ( .A(_06097_ ), .Z(_06216_ ) );
AOI21_X1 _14211_ ( .A(_06215_ ), .B1(_04339_ ), .B2(_06216_ ), .ZN(_06217_ ) );
OAI221_X1 _14212_ ( .A(_06212_ ), .B1(_06213_ ), .B2(_06214_ ), .C1(_06217_ ), .C2(_06094_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
AND3_X1 _14213_ ( .A1(_04632_ ), .A2(_04651_ ), .A3(_06097_ ), .ZN(_06218_ ) );
AND3_X1 _14214_ ( .A1(_06166_ ), .A2(\ID_EX_pc [11] ), .A3(\ID_EX_typ [7] ), .ZN(_06219_ ) );
OAI21_X1 _14215_ ( .A(_06164_ ), .B1(_06218_ ), .B2(_06219_ ), .ZN(_06220_ ) );
NAND2_X1 _14216_ ( .A1(_05467_ ), .A2(_05471_ ), .ZN(_06221_ ) );
AOI22_X1 _14217_ ( .A1(_06221_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02703_ ), .ZN(_06222_ ) );
OAI211_X1 _14218_ ( .A(_06222_ ), .B(_06136_ ), .C1(fanout_net_5 ), .C2(_02702_ ), .ZN(_06223_ ) );
NAND4_X1 _14219_ ( .A1(_05467_ ), .A2(_06135_ ), .A3(_05471_ ), .A4(_06136_ ), .ZN(_06224_ ) );
NAND3_X1 _14220_ ( .A1(_06220_ ), .A2(_06223_ ), .A3(_06224_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _14221_ ( .A(_06117_ ), .B1(_05513_ ), .B2(_05514_ ), .ZN(_06225_ ) );
AOI22_X1 _14222_ ( .A1(_05515_ ), .A2(fanout_net_6 ), .B1(fanout_net_5 ), .B2(_02725_ ), .ZN(_06226_ ) );
NAND3_X1 _14223_ ( .A1(_02722_ ), .A2(_02723_ ), .A3(_05300_ ), .ZN(_06227_ ) );
AOI211_X1 _14224_ ( .A(_06090_ ), .B(_06225_ ), .C1(_06226_ ), .C2(_06227_ ), .ZN(_06228_ ) );
MUX2_X1 _14225_ ( .A(_05502_ ), .B(_04675_ ), .S(_06133_ ), .Z(_06229_ ) );
AOI21_X1 _14226_ ( .A(_06228_ ), .B1(_06229_ ), .B2(_06091_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
AOI21_X1 _14227_ ( .A(_06117_ ), .B1(_05527_ ), .B2(_05528_ ), .ZN(_06230_ ) );
AOI21_X1 _14228_ ( .A(_06230_ ), .B1(fanout_net_5 ), .B2(\ID_EX_imm [9] ), .ZN(_06231_ ) );
OAI21_X1 _14229_ ( .A(_06231_ ), .B1(fanout_net_5 ), .B2(_04723_ ), .ZN(_06232_ ) );
OAI211_X1 _14230_ ( .A(_06232_ ), .B(_06111_ ), .C1(_06138_ ), .C2(_05530_ ), .ZN(_06233_ ) );
BUF_X4 _14231_ ( .A(_06090_ ), .Z(_06234_ ) );
OR4_X1 _14232_ ( .A1(\ID_EX_pc [9] ), .A2(_03259_ ), .A3(_03791_ ), .A4(_03782_ ), .ZN(_06235_ ) );
INV_X1 _14233_ ( .A(_04722_ ), .ZN(_06236_ ) );
OAI211_X1 _14234_ ( .A(_06234_ ), .B(_06235_ ), .C1(_06236_ ), .C2(_06095_ ), .ZN(_06237_ ) );
NAND2_X1 _14235_ ( .A1(_06233_ ), .A2(_06237_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _14236_ ( .A(fanout_net_5 ), .B1(_02635_ ), .B2(_02654_ ), .ZN(_06238_ ) );
AND2_X1 _14237_ ( .A1(fanout_net_5 ), .A2(\ID_EX_imm [8] ), .ZN(_06239_ ) );
OAI221_X1 _14238_ ( .A(_06104_ ), .B1(_06238_ ), .B2(_06239_ ), .C1(_05553_ ), .C2(_06138_ ), .ZN(_06240_ ) );
AND3_X1 _14239_ ( .A1(_05468_ ), .A2(_05544_ ), .A3(_05470_ ), .ZN(_06241_ ) );
NOR2_X1 _14240_ ( .A1(_05342_ ), .A2(_05343_ ), .ZN(_06242_ ) );
INV_X1 _14241_ ( .A(_05550_ ), .ZN(_06243_ ) );
INV_X1 _14242_ ( .A(_05551_ ), .ZN(_06244_ ) );
AND4_X1 _14243_ ( .A1(_06242_ ), .A2(_05548_ ), .A3(_06243_ ), .A4(_06244_ ), .ZN(_06245_ ) );
AOI21_X1 _14244_ ( .A(_05546_ ), .B1(_05468_ ), .B2(_05470_ ), .ZN(_06246_ ) );
AOI21_X1 _14245_ ( .A(_06241_ ), .B1(_06245_ ), .B2(_06246_ ), .ZN(_06247_ ) );
NAND3_X1 _14246_ ( .A1(_06247_ ), .A2(_06135_ ), .A3(_06136_ ), .ZN(_06248_ ) );
AND3_X1 _14247_ ( .A1(_06166_ ), .A2(\ID_EX_pc [8] ), .A3(\ID_EX_typ [7] ), .ZN(_06249_ ) );
INV_X1 _14248_ ( .A(_04699_ ), .ZN(_06250_ ) );
AOI21_X1 _14249_ ( .A(_06249_ ), .B1(_06250_ ), .B2(_06216_ ), .ZN(_06251_ ) );
OAI211_X1 _14250_ ( .A(_06240_ ), .B(_06248_ ), .C1(_06251_ ), .C2(_06211_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
AND2_X1 _14251_ ( .A1(_05561_ ), .A2(_05563_ ), .ZN(_06252_ ) );
AND2_X1 _14252_ ( .A1(_05562_ ), .A2(_05564_ ), .ZN(_06253_ ) );
AOI22_X1 _14253_ ( .A1(_06252_ ), .A2(_06253_ ), .B1(_03829_ ), .B2(_03814_ ), .ZN(_06254_ ) );
AND3_X1 _14254_ ( .A1(_03814_ ), .A2(_03829_ ), .A3(\EX_LS_result_csreg_mem [7] ), .ZN(_06255_ ) );
OR2_X1 _14255_ ( .A1(_06254_ ), .A2(_06255_ ), .ZN(_06256_ ) );
AOI22_X1 _14256_ ( .A1(_06256_ ), .A2(_06116_ ), .B1(fanout_net_5 ), .B2(\ID_EX_imm [7] ), .ZN(_06257_ ) );
OAI21_X1 _14257_ ( .A(_06257_ ), .B1(fanout_net_5 ), .B2(_04749_ ), .ZN(_06258_ ) );
OAI211_X1 _14258_ ( .A(_06258_ ), .B(_06111_ ), .C1(_06138_ ), .C2(_05569_ ), .ZN(_06259_ ) );
NAND3_X1 _14259_ ( .A1(_04727_ ), .A2(_04747_ ), .A3(_06133_ ), .ZN(_06260_ ) );
OAI211_X1 _14260_ ( .A(_06260_ ), .B(_06234_ ), .C1(\ID_EX_pc [7] ), .C2(_06216_ ), .ZN(_06261_ ) );
NAND2_X1 _14261_ ( .A1(_06259_ ), .A2(_06261_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
AND3_X1 _14262_ ( .A1(_05492_ ), .A2(_05594_ ), .A3(_05493_ ), .ZN(_06262_ ) );
AOI21_X1 _14263_ ( .A(_06262_ ), .B1(_05592_ ), .B2(_05589_ ), .ZN(_06263_ ) );
AOI21_X1 _14264_ ( .A(\ID_EX_typ [0] ), .B1(_02479_ ), .B2(_02498_ ), .ZN(_06264_ ) );
AND2_X1 _14265_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [6] ), .ZN(_06265_ ) );
OAI221_X1 _14266_ ( .A(_06104_ ), .B1(_06138_ ), .B2(_06263_ ), .C1(_06264_ ), .C2(_06265_ ), .ZN(_06266_ ) );
NAND4_X1 _14267_ ( .A1(_05593_ ), .A2(_06135_ ), .A3(_05595_ ), .A4(_06104_ ), .ZN(_06267_ ) );
MUX2_X1 _14268_ ( .A(_05581_ ), .B(_04772_ ), .S(_06133_ ), .Z(_06268_ ) );
OAI211_X1 _14269_ ( .A(_06266_ ), .B(_06267_ ), .C1(_06268_ ), .C2(_06211_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
AOI21_X1 _14270_ ( .A(_05609_ ), .B1(_05238_ ), .B2(_05240_ ), .ZN(_06269_ ) );
NAND3_X1 _14271_ ( .A1(_05226_ ), .A2(\mepc [5] ), .A3(_05314_ ), .ZN(_06270_ ) );
NOR3_X1 _14272_ ( .A1(_05608_ ), .A2(_05342_ ), .A3(_05612_ ), .ZN(_06271_ ) );
NAND3_X1 _14273_ ( .A1(_06269_ ), .A2(_06270_ ), .A3(_06271_ ), .ZN(_06272_ ) );
NAND3_X1 _14274_ ( .A1(_05238_ ), .A2(_05615_ ), .A3(_05240_ ), .ZN(_06273_ ) );
AND2_X1 _14275_ ( .A1(_06272_ ), .A2(_06273_ ), .ZN(_06274_ ) );
OAI22_X1 _14276_ ( .A1(_06274_ ), .A2(_06138_ ), .B1(_03779_ ), .B2(\ID_EX_imm [5] ), .ZN(_06275_ ) );
AOI21_X1 _14277_ ( .A(_06275_ ), .B1(_05499_ ), .B2(_04978_ ), .ZN(_06276_ ) );
NAND3_X1 _14278_ ( .A1(_06272_ ), .A2(_06125_ ), .A3(_06273_ ), .ZN(_06277_ ) );
INV_X1 _14279_ ( .A(_06277_ ), .ZN(_06278_ ) );
OAI21_X1 _14280_ ( .A(_06156_ ), .B1(_06276_ ), .B2(_06278_ ), .ZN(_06279_ ) );
AND4_X1 _14281_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06280_ ) );
AOI21_X1 _14282_ ( .A(_06280_ ), .B1(_04795_ ), .B2(_06216_ ), .ZN(_06281_ ) );
OAI21_X1 _14283_ ( .A(_06279_ ), .B1(_06105_ ), .B2(_06281_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
AND4_X1 _14284_ ( .A1(_05624_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06282_ ) );
AOI211_X1 _14285_ ( .A(_06093_ ), .B(_06282_ ), .C1(_04817_ ), .C2(_06133_ ), .ZN(_06283_ ) );
NAND2_X1 _14286_ ( .A1(_05636_ ), .A2(_05638_ ), .ZN(_06284_ ) );
NAND3_X1 _14287_ ( .A1(_05636_ ), .A2(_06116_ ), .A3(_05638_ ), .ZN(_06285_ ) );
NAND2_X1 _14288_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [4] ), .ZN(_06286_ ) );
AND2_X1 _14289_ ( .A1(_06285_ ), .A2(_06286_ ), .ZN(_06287_ ) );
NAND2_X1 _14290_ ( .A1(_02452_ ), .A2(_03779_ ), .ZN(_06288_ ) );
AOI221_X4 _14291_ ( .A(_06089_ ), .B1(fanout_net_6 ), .B2(_06284_ ), .C1(_06287_ ), .C2(_06288_ ), .ZN(_06289_ ) );
OR2_X1 _14292_ ( .A1(_06283_ ), .A2(_06289_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _14293_ ( .A1(_05652_ ), .A2(_05651_ ), .ZN(_06290_ ) );
AOI21_X1 _14294_ ( .A(_06290_ ), .B1(_05238_ ), .B2(_05240_ ), .ZN(_06291_ ) );
INV_X1 _14295_ ( .A(_05342_ ), .ZN(_06292_ ) );
NAND4_X1 _14296_ ( .A1(_06291_ ), .A2(_06292_ ), .A3(_05654_ ), .A4(_05653_ ), .ZN(_06293_ ) );
NAND3_X1 _14297_ ( .A1(_05492_ ), .A2(_05649_ ), .A3(_05493_ ), .ZN(_06294_ ) );
NAND2_X1 _14298_ ( .A1(_06293_ ), .A2(_06294_ ), .ZN(_06295_ ) );
AOI22_X1 _14299_ ( .A1(_04940_ ), .A2(_05713_ ), .B1(fanout_net_6 ), .B2(_06295_ ), .ZN(_06296_ ) );
OAI211_X1 _14300_ ( .A(_06296_ ), .B(_06207_ ), .C1(_05499_ ), .C2(\ID_EX_imm [3] ), .ZN(_06297_ ) );
NAND4_X1 _14301_ ( .A1(_06293_ ), .A2(_06135_ ), .A3(_06294_ ), .A4(_06104_ ), .ZN(_06298_ ) );
AND3_X1 _14302_ ( .A1(_06166_ ), .A2(\ID_EX_pc [3] ), .A3(\ID_EX_typ [7] ), .ZN(_06299_ ) );
AOI21_X1 _14303_ ( .A(_06299_ ), .B1(_04533_ ), .B2(_06216_ ), .ZN(_06300_ ) );
OAI211_X1 _14304_ ( .A(_06297_ ), .B(_06298_ ), .C1(_06300_ ), .C2(_06211_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
NAND3_X1 _14305_ ( .A1(_03838_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_05224_ ), .ZN(_06301_ ) );
NAND2_X1 _14306_ ( .A1(_05667_ ), .A2(_06301_ ), .ZN(_06302_ ) );
NOR3_X1 _14307_ ( .A1(_06302_ ), .A2(_05669_ ), .A3(_05343_ ), .ZN(_06303_ ) );
AOI21_X1 _14308_ ( .A(_05671_ ), .B1(_05492_ ), .B2(_05493_ ), .ZN(_06304_ ) );
NAND2_X1 _14309_ ( .A1(_06303_ ), .A2(_06304_ ), .ZN(_06305_ ) );
NAND3_X1 _14310_ ( .A1(_05492_ ), .A2(_05983_ ), .A3(_05493_ ), .ZN(_06306_ ) );
NAND2_X1 _14311_ ( .A1(_06305_ ), .A2(_06306_ ), .ZN(_06307_ ) );
AOI22_X1 _14312_ ( .A1(_04511_ ), .A2(_05713_ ), .B1(fanout_net_6 ), .B2(_06307_ ), .ZN(_06308_ ) );
OAI211_X1 _14313_ ( .A(_06308_ ), .B(_06207_ ), .C1(_05499_ ), .C2(\ID_EX_imm [2] ), .ZN(_06309_ ) );
NAND4_X1 _14314_ ( .A1(_06305_ ), .A2(_06135_ ), .A3(_06306_ ), .A4(_06104_ ), .ZN(_06310_ ) );
INV_X1 _14315_ ( .A(\ID_EX_pc [2] ), .ZN(_06311_ ) );
MUX2_X1 _14316_ ( .A(_06311_ ), .B(_04510_ ), .S(_06097_ ), .Z(_06312_ ) );
OAI211_X1 _14317_ ( .A(_06309_ ), .B(_06310_ ), .C1(_06312_ ), .C2(_06211_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
INV_X1 _14318_ ( .A(_05242_ ), .ZN(_06313_ ) );
AOI22_X1 _14319_ ( .A1(_06313_ ), .A2(fanout_net_6 ), .B1(\ID_EX_typ [0] ), .B2(_02895_ ), .ZN(_06314_ ) );
OAI211_X1 _14320_ ( .A(_06314_ ), .B(_06207_ ), .C1(\ID_EX_typ [0] ), .C2(_02894_ ), .ZN(_06315_ ) );
NAND4_X1 _14321_ ( .A1(_05237_ ), .A2(_06125_ ), .A3(_05241_ ), .A4(_06104_ ), .ZN(_06316_ ) );
AND3_X1 _14322_ ( .A1(_06166_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_typ [7] ), .ZN(_06317_ ) );
AOI21_X1 _14323_ ( .A(_06317_ ), .B1(_04290_ ), .B2(_06216_ ), .ZN(_06318_ ) );
OAI211_X1 _14324_ ( .A(_06315_ ), .B(_06316_ ), .C1(_06105_ ), .C2(_06318_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
AND3_X1 _14325_ ( .A1(_04438_ ), .A2(_04457_ ), .A3(_06097_ ), .ZN(_06319_ ) );
AND3_X1 _14326_ ( .A1(_06166_ ), .A2(\ID_EX_pc [1] ), .A3(\ID_EX_typ [7] ), .ZN(_06320_ ) );
OAI21_X1 _14327_ ( .A(_06164_ ), .B1(_06319_ ), .B2(_06320_ ), .ZN(_06321_ ) );
NAND3_X1 _14328_ ( .A1(_05468_ ), .A2(_05984_ ), .A3(_05470_ ), .ZN(_06322_ ) );
NAND4_X1 _14329_ ( .A1(_05683_ ), .A2(_05684_ ), .A3(_05685_ ), .A4(_05686_ ), .ZN(_06323_ ) );
OAI21_X1 _14330_ ( .A(_06322_ ), .B1(_05221_ ), .B2(_06323_ ), .ZN(_06324_ ) );
AOI22_X1 _14331_ ( .A1(_06324_ ), .A2(fanout_net_6 ), .B1(\ID_EX_typ [0] ), .B2(_02400_ ), .ZN(_06325_ ) );
OAI211_X1 _14332_ ( .A(_06325_ ), .B(_06136_ ), .C1(_02399_ ), .C2(\ID_EX_typ [0] ), .ZN(_06326_ ) );
OR2_X1 _14333_ ( .A1(_05221_ ), .A2(_06323_ ), .ZN(_06327_ ) );
NAND4_X1 _14334_ ( .A1(_06327_ ), .A2(_06135_ ), .A3(_06322_ ), .A4(_06207_ ), .ZN(_06328_ ) );
NAND3_X1 _14335_ ( .A1(_06321_ ), .A2(_06326_ ), .A3(_06328_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
NAND3_X1 _14336_ ( .A1(_04464_ ), .A2(_04484_ ), .A3(_06133_ ), .ZN(_06329_ ) );
OAI211_X1 _14337_ ( .A(_06329_ ), .B(_06234_ ), .C1(\ID_EX_pc [0] ), .C2(_06216_ ), .ZN(_06330_ ) );
AND3_X1 _14338_ ( .A1(_05312_ ), .A2(\mepc [0] ), .A3(_05314_ ), .ZN(_06331_ ) );
NOR3_X1 _14339_ ( .A1(_06331_ ), .A2(_05718_ ), .A3(_05715_ ), .ZN(_06332_ ) );
AOI22_X1 _14340_ ( .A1(_05286_ ), .A2(\mtvec [0] ), .B1(_03861_ ), .B2(_05291_ ), .ZN(_06333_ ) );
AOI21_X1 _14341_ ( .A(_03871_ ), .B1(_06332_ ), .B2(_06333_ ), .ZN(_06334_ ) );
AND3_X1 _14342_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [0] ), .ZN(_06335_ ) );
OAI21_X1 _14343_ ( .A(_06125_ ), .B1(_06334_ ), .B2(_06335_ ), .ZN(_06336_ ) );
NAND2_X1 _14344_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [0] ), .ZN(_06337_ ) );
NAND2_X1 _14345_ ( .A1(_06336_ ), .A2(_06337_ ), .ZN(_06338_ ) );
AND3_X1 _14346_ ( .A1(_02403_ ), .A2(_05186_ ), .A3(_02423_ ), .ZN(_06339_ ) );
OAI221_X1 _14347_ ( .A(_06152_ ), .B1(_06138_ ), .B2(_05724_ ), .C1(_06338_ ), .C2(_06339_ ), .ZN(_06340_ ) );
NAND2_X1 _14348_ ( .A1(_06330_ ), .A2(_06340_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
INV_X1 _14349_ ( .A(_05495_ ), .ZN(_06341_ ) );
AOI22_X1 _14350_ ( .A1(_06341_ ), .A2(fanout_net_6 ), .B1(_05300_ ), .B2(_04854_ ), .ZN(_06342_ ) );
OAI211_X1 _14351_ ( .A(_06342_ ), .B(_06207_ ), .C1(_05499_ ), .C2(\ID_EX_imm [28] ), .ZN(_06343_ ) );
INV_X1 _14352_ ( .A(_05485_ ), .ZN(_06344_ ) );
NAND2_X1 _14353_ ( .A1(_05494_ ), .A2(_05488_ ), .ZN(_06345_ ) );
NAND4_X1 _14354_ ( .A1(_06344_ ), .A2(_06125_ ), .A3(_06345_ ), .A4(_06104_ ), .ZN(_06346_ ) );
AND3_X1 _14355_ ( .A1(_06166_ ), .A2(\ID_EX_pc [28] ), .A3(\ID_EX_typ [7] ), .ZN(_06347_ ) );
AOI21_X1 _14356_ ( .A(_06347_ ), .B1(_04268_ ), .B2(_06216_ ), .ZN(_06348_ ) );
OAI211_X1 _14357_ ( .A(_06343_ ), .B(_06346_ ), .C1(_06105_ ), .C2(_06348_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
AOI22_X1 _14358_ ( .A1(_05704_ ), .A2(fanout_net_6 ), .B1(_05300_ ), .B2(_05037_ ), .ZN(_06349_ ) );
OAI211_X1 _14359_ ( .A(_06349_ ), .B(_06207_ ), .C1(_05499_ ), .C2(\ID_EX_imm [27] ), .ZN(_06350_ ) );
INV_X1 _14360_ ( .A(_05695_ ), .ZN(_06351_ ) );
NAND2_X1 _14361_ ( .A1(_05702_ ), .A2(_05698_ ), .ZN(_06352_ ) );
NAND4_X1 _14362_ ( .A1(_06351_ ), .A2(_06125_ ), .A3(_06352_ ), .A4(_06093_ ), .ZN(_06353_ ) );
AND3_X1 _14363_ ( .A1(_06166_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_06354_ ) );
AOI21_X1 _14364_ ( .A(_06354_ ), .B1(_04363_ ), .B2(_06216_ ), .ZN(_06355_ ) );
OAI211_X1 _14365_ ( .A(_06350_ ), .B(_06353_ ), .C1(_06105_ ), .C2(_06355_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
NAND4_X1 _14366_ ( .A1(_05736_ ), .A2(_05737_ ), .A3(_05738_ ), .A4(_05739_ ), .ZN(_06356_ ) );
OR2_X1 _14367_ ( .A1(_05221_ ), .A2(_06356_ ), .ZN(_06357_ ) );
OAI21_X1 _14368_ ( .A(_06357_ ), .B1(\EX_LS_result_csreg_mem [26] ), .B2(_05222_ ), .ZN(_06358_ ) );
AOI22_X1 _14369_ ( .A1(_05044_ ), .A2(_05713_ ), .B1(fanout_net_6 ), .B2(_06358_ ), .ZN(_06359_ ) );
OAI211_X1 _14370_ ( .A(_06359_ ), .B(_06207_ ), .C1(_05499_ ), .C2(\ID_EX_imm [26] ), .ZN(_06360_ ) );
OR3_X1 _14371_ ( .A1(_06358_ ), .A2(_06117_ ), .A3(_06089_ ), .ZN(_06361_ ) );
AND3_X1 _14372_ ( .A1(_03258_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_06362_ ) );
AOI21_X1 _14373_ ( .A(_06362_ ), .B1(_04386_ ), .B2(_06133_ ), .ZN(_06363_ ) );
OAI211_X1 _14374_ ( .A(_06360_ ), .B(_06361_ ), .C1(_06105_ ), .C2(_06363_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
OR2_X1 _14375_ ( .A1(_05222_ ), .A2(\EX_LS_result_csreg_mem [25] ), .ZN(_06364_ ) );
AND2_X1 _14376_ ( .A1(_05745_ ), .A2(_05746_ ), .ZN(_06365_ ) );
NAND4_X1 _14377_ ( .A1(_05222_ ), .A2(_05747_ ), .A3(_05748_ ), .A4(_06365_ ), .ZN(_06366_ ) );
NAND2_X1 _14378_ ( .A1(_06364_ ), .A2(_06366_ ), .ZN(_06367_ ) );
AOI22_X1 _14379_ ( .A1(_06367_ ), .A2(fanout_net_6 ), .B1(\ID_EX_typ [0] ), .B2(_02867_ ), .ZN(_06368_ ) );
OAI211_X1 _14380_ ( .A(_06368_ ), .B(_06207_ ), .C1(\ID_EX_typ [0] ), .C2(_02815_ ), .ZN(_06369_ ) );
NAND4_X1 _14381_ ( .A1(_06364_ ), .A2(_06366_ ), .A3(_06125_ ), .A4(_06093_ ), .ZN(_06370_ ) );
AND3_X1 _14382_ ( .A1(_06166_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06371_ ) );
AOI21_X1 _14383_ ( .A(_06371_ ), .B1(_04432_ ), .B2(_06216_ ), .ZN(_06372_ ) );
OAI211_X1 _14384_ ( .A(_06369_ ), .B(_06370_ ), .C1(_06372_ ), .C2(_06094_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
INV_X1 _14385_ ( .A(_05781_ ), .ZN(_06373_ ) );
AOI22_X1 _14386_ ( .A1(_06373_ ), .A2(fanout_net_6 ), .B1(_05300_ ), .B2(_05052_ ), .ZN(_06374_ ) );
OAI211_X1 _14387_ ( .A(_06374_ ), .B(_06207_ ), .C1(_05499_ ), .C2(\ID_EX_imm [24] ), .ZN(_06375_ ) );
NAND4_X1 _14388_ ( .A1(_05772_ ), .A2(_06125_ ), .A3(_05780_ ), .A4(_06093_ ), .ZN(_06376_ ) );
AND3_X1 _14389_ ( .A1(_03258_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_typ [7] ), .ZN(_06377_ ) );
AOI21_X1 _14390_ ( .A(_06377_ ), .B1(_04409_ ), .B2(_06133_ ), .ZN(_06378_ ) );
OAI211_X1 _14391_ ( .A(_06375_ ), .B(_06376_ ), .C1(_06211_ ), .C2(_06378_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _14392_ ( .A(_06095_ ), .B1(_04016_ ), .B2(_04049_ ), .ZN(_06379_ ) );
AND3_X1 _14393_ ( .A1(_06166_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_typ [7] ), .ZN(_06380_ ) );
OAI21_X1 _14394_ ( .A(_06164_ ), .B1(_06379_ ), .B2(_06380_ ), .ZN(_06381_ ) );
NAND3_X1 _14395_ ( .A1(_05468_ ), .A2(_06010_ ), .A3(_05470_ ), .ZN(_06382_ ) );
NAND4_X1 _14396_ ( .A1(_05794_ ), .A2(_05795_ ), .A3(_05796_ ), .A4(_05797_ ), .ZN(_06383_ ) );
OAI21_X1 _14397_ ( .A(_06382_ ), .B1(_05221_ ), .B2(_06383_ ), .ZN(_06384_ ) );
AOI22_X1 _14398_ ( .A1(_06384_ ), .A2(fanout_net_6 ), .B1(\ID_EX_typ [0] ), .B2(_02177_ ), .ZN(_06385_ ) );
OAI211_X1 _14399_ ( .A(_06385_ ), .B(_06136_ ), .C1(_02179_ ), .C2(\ID_EX_typ [0] ), .ZN(_06386_ ) );
OR3_X1 _14400_ ( .A1(_06384_ ), .A2(_06117_ ), .A3(_06090_ ), .ZN(_06387_ ) );
NAND3_X1 _14401_ ( .A1(_06381_ ), .A2(_06386_ ), .A3(_06387_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
AOI22_X1 _14402_ ( .A1(_05818_ ), .A2(_06116_ ), .B1(\ID_EX_typ [0] ), .B2(\ID_EX_imm [22] ), .ZN(_06388_ ) );
OAI21_X1 _14403_ ( .A(_06388_ ), .B1(\ID_EX_typ [0] ), .B2(_04088_ ), .ZN(_06389_ ) );
OAI211_X1 _14404_ ( .A(_06389_ ), .B(_06111_ ), .C1(_06138_ ), .C2(_05818_ ), .ZN(_06390_ ) );
NAND4_X1 _14405_ ( .A1(_05803_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06391_ ) );
INV_X1 _14406_ ( .A(_04087_ ), .ZN(_06392_ ) );
OAI211_X1 _14407_ ( .A(_06234_ ), .B(_06391_ ), .C1(_06392_ ), .C2(_06095_ ), .ZN(_06393_ ) );
NAND2_X1 _14408_ ( .A1(_06390_ ), .A2(_06393_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
AOI22_X1 _14409_ ( .A1(_04838_ ), .A2(_05713_ ), .B1(fanout_net_6 ), .B2(_05859_ ), .ZN(_06394_ ) );
OAI211_X1 _14410_ ( .A(_06394_ ), .B(_06104_ ), .C1(_05499_ ), .C2(\ID_EX_imm [31] ), .ZN(_06395_ ) );
OR2_X1 _14411_ ( .A1(_05222_ ), .A2(\EX_LS_result_csreg_mem [31] ), .ZN(_06396_ ) );
NAND4_X1 _14412_ ( .A1(_06396_ ), .A2(_06125_ ), .A3(_05858_ ), .A4(_06093_ ), .ZN(_06397_ ) );
AND3_X1 _14413_ ( .A1(_03258_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06398_ ) );
AOI21_X1 _14414_ ( .A(_06398_ ), .B1(_04316_ ), .B2(_06133_ ), .ZN(_06399_ ) );
OAI211_X1 _14415_ ( .A(_06395_ ), .B(_06397_ ), .C1(_06211_ ), .C2(_06399_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
NAND3_X1 _14416_ ( .A1(_05836_ ), .A2(_05839_ ), .A3(_06156_ ), .ZN(_06400_ ) );
NOR3_X1 _14417_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06401_ ) );
AND2_X1 _14418_ ( .A1(\ID_EX_typ [3] ), .A2(fanout_net_6 ), .ZN(_06402_ ) );
AND2_X1 _14419_ ( .A1(_06401_ ), .A2(_06402_ ), .ZN(_06403_ ) );
BUF_X4 _14420_ ( .A(_06403_ ), .Z(_06404_ ) );
INV_X1 _14421_ ( .A(_06404_ ), .ZN(_06405_ ) );
BUF_X2 _14422_ ( .A(_06405_ ), .Z(_06406_ ) );
NOR3_X1 _14423_ ( .A1(_04824_ ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06407_ ) );
AND2_X2 _14424_ ( .A1(_06407_ ), .A2(_06402_ ), .ZN(_06408_ ) );
INV_X1 _14425_ ( .A(_06408_ ), .ZN(_06409_ ) );
BUF_X4 _14426_ ( .A(_06409_ ), .Z(_06410_ ) );
OAI22_X1 _14427_ ( .A1(_05829_ ), .A2(_06406_ ), .B1(_02206_ ), .B2(_06410_ ), .ZN(_06411_ ) );
INV_X1 _14428_ ( .A(_05118_ ), .ZN(_06412_ ) );
NAND2_X1 _14429_ ( .A1(_06412_ ), .A2(_04243_ ), .ZN(_06413_ ) );
AND2_X1 _14430_ ( .A1(_06413_ ), .A2(_05135_ ), .ZN(_06414_ ) );
INV_X1 _14431_ ( .A(_04141_ ), .ZN(_06415_ ) );
OR2_X1 _14432_ ( .A1(_06414_ ), .A2(_06415_ ), .ZN(_06416_ ) );
AND2_X1 _14433_ ( .A1(_06416_ ), .A2(_05124_ ), .ZN(_06417_ ) );
XNOR2_X1 _14434_ ( .A(_06417_ ), .B(_04115_ ), .ZN(_06418_ ) );
AND3_X1 _14435_ ( .A1(_04001_ ), .A2(\ID_EX_typ [3] ), .A3(_04826_ ), .ZN(_06419_ ) );
AND2_X1 _14436_ ( .A1(_06419_ ), .A2(_04835_ ), .ZN(_06420_ ) );
BUF_X2 _14437_ ( .A(_06420_ ), .Z(_06421_ ) );
BUF_X4 _14438_ ( .A(_06421_ ), .Z(_06422_ ) );
AOI21_X1 _14439_ ( .A(_06411_ ), .B1(_06418_ ), .B2(_06422_ ), .ZN(_06423_ ) );
NOR2_X1 _14440_ ( .A1(_03782_ ), .A2(\ID_EX_typ [6] ), .ZN(_06424_ ) );
AND2_X2 _14441_ ( .A1(_06424_ ), .A2(_03259_ ), .ZN(_06425_ ) );
INV_X1 _14442_ ( .A(_06425_ ), .ZN(_06426_ ) );
BUF_X4 _14443_ ( .A(_06426_ ), .Z(_06427_ ) );
BUF_X4 _14444_ ( .A(_06427_ ), .Z(_06428_ ) );
OAI21_X1 _14445_ ( .A(_05498_ ), .B1(_06423_ ), .B2(_06428_ ), .ZN(_06429_ ) );
AND2_X1 _14446_ ( .A1(_05165_ ), .A2(fanout_net_6 ), .ZN(_06430_ ) );
BUF_X4 _14447_ ( .A(_06430_ ), .Z(_06431_ ) );
BUF_X4 _14448_ ( .A(_06431_ ), .Z(_06432_ ) );
NAND2_X4 _14449_ ( .A1(_04951_ ), .A2(_04952_ ), .ZN(_06433_ ) );
AND2_X2 _14450_ ( .A1(_04945_ ), .A2(_06433_ ), .ZN(_06434_ ) );
BUF_X4 _14451_ ( .A(_04957_ ), .Z(_06435_ ) );
AND2_X4 _14452_ ( .A1(_06434_ ), .A2(_06435_ ), .ZN(_06436_ ) );
INV_X1 _14453_ ( .A(_04939_ ), .ZN(_06437_ ) );
AND2_X4 _14454_ ( .A1(_06436_ ), .A2(_06437_ ), .ZN(_06438_ ) );
AND2_X4 _14455_ ( .A1(_06438_ ), .A2(_04984_ ), .ZN(_06439_ ) );
INV_X1 _14456_ ( .A(_04977_ ), .ZN(_06440_ ) );
OAI21_X4 _14457_ ( .A(_04967_ ), .B1(_06439_ ), .B2(_06440_ ), .ZN(_06441_ ) );
INV_X1 _14458_ ( .A(_04971_ ), .ZN(_06442_ ) );
NOR2_X1 _14459_ ( .A1(_06441_ ), .A2(_06442_ ), .ZN(_06443_ ) );
NOR4_X1 _14460_ ( .A1(_06439_ ), .A2(_04971_ ), .A3(_04967_ ), .A4(_06440_ ), .ZN(_06444_ ) );
NOR2_X1 _14461_ ( .A1(_06443_ ), .A2(_06444_ ), .ZN(_06445_ ) );
NOR2_X1 _14462_ ( .A1(_06445_ ), .A2(_04838_ ), .ZN(_06446_ ) );
INV_X1 _14463_ ( .A(_04933_ ), .ZN(_06447_ ) );
OR3_X4 _14464_ ( .A1(_06441_ ), .A2(_06442_ ), .A3(_06447_ ), .ZN(_06448_ ) );
INV_X1 _14465_ ( .A(_04928_ ), .ZN(_06449_ ) );
NOR2_X1 _14466_ ( .A1(_06448_ ), .A2(_06449_ ), .ZN(_06450_ ) );
NOR3_X1 _14467_ ( .A1(_06443_ ), .A2(_04928_ ), .A3(_04933_ ), .ZN(_06451_ ) );
NOR3_X2 _14468_ ( .A1(_06448_ ), .A2(_06449_ ), .A3(_05001_ ), .ZN(_06452_ ) );
AND2_X2 _14469_ ( .A1(_06452_ ), .A2(_04923_ ), .ZN(_06453_ ) );
NOR3_X1 _14470_ ( .A1(_06450_ ), .A2(_04923_ ), .A3(_04919_ ), .ZN(_06454_ ) );
OAI221_X1 _14471_ ( .A(_06446_ ), .B1(_06450_ ), .B2(_06451_ ), .C1(_06453_ ), .C2(_06454_ ), .ZN(_06455_ ) );
NAND3_X1 _14472_ ( .A1(_04898_ ), .A2(_04899_ ), .A3(_04896_ ), .ZN(_06456_ ) );
NOR3_X1 _14473_ ( .A1(_06456_ ), .A2(_04913_ ), .A3(_05006_ ), .ZN(_06457_ ) );
AND4_X1 _14474_ ( .A1(_04863_ ), .A2(_04859_ ), .A3(_04872_ ), .A4(_04867_ ), .ZN(_06458_ ) );
AND4_X1 _14475_ ( .A1(_04880_ ), .A2(_04879_ ), .A3(_04875_ ), .A4(_04876_ ), .ZN(_06459_ ) );
AND3_X1 _14476_ ( .A1(_06459_ ), .A2(_04887_ ), .A3(_04891_ ), .ZN(_06460_ ) );
AOI22_X1 _14477_ ( .A1(_04842_ ), .A2(_04843_ ), .B1(_05041_ ), .B2(_05042_ ), .ZN(_06461_ ) );
AND3_X1 _14478_ ( .A1(_06461_ ), .A2(_05036_ ), .A3(_04837_ ), .ZN(_06462_ ) );
INV_X1 _14479_ ( .A(_05059_ ), .ZN(_06463_ ) );
NOR4_X1 _14480_ ( .A1(_05063_ ), .A2(_06463_ ), .A3(_04849_ ), .A4(_04853_ ), .ZN(_06464_ ) );
NAND4_X1 _14481_ ( .A1(_06458_ ), .A2(_06460_ ), .A3(_06462_ ), .A4(_06464_ ), .ZN(_06465_ ) );
AND4_X1 _14482_ ( .A1(_04923_ ), .A2(_06452_ ), .A3(_06457_ ), .A4(_06465_ ), .ZN(_06466_ ) );
NOR2_X2 _14483_ ( .A1(_06455_ ), .A2(_06466_ ), .ZN(_06467_ ) );
OR4_X1 _14484_ ( .A1(_04863_ ), .A2(_04859_ ), .A3(_04872_ ), .A4(_04867_ ), .ZN(_06468_ ) );
OR2_X1 _14485_ ( .A1(_04887_ ), .A2(_04891_ ), .ZN(_06469_ ) );
OR3_X1 _14486_ ( .A1(_06469_ ), .A2(_04881_ ), .A3(_04877_ ), .ZN(_06470_ ) );
OR2_X2 _14487_ ( .A1(_06468_ ), .A2(_06470_ ), .ZN(_06471_ ) );
NAND2_X1 _14488_ ( .A1(_05006_ ), .A2(_04913_ ), .ZN(_06472_ ) );
NOR4_X1 _14489_ ( .A1(_06471_ ), .A2(_04900_ ), .A3(_04896_ ), .A4(_06472_ ), .ZN(_06473_ ) );
AND2_X1 _14490_ ( .A1(_04842_ ), .A2(_04843_ ), .ZN(_06474_ ) );
NAND4_X1 _14491_ ( .A1(_05063_ ), .A2(_06463_ ), .A3(_04849_ ), .A4(_04853_ ), .ZN(_06475_ ) );
NOR4_X1 _14492_ ( .A1(_06475_ ), .A2(_04837_ ), .A3(_05036_ ), .A4(_05043_ ), .ZN(_06476_ ) );
AND3_X1 _14493_ ( .A1(_06473_ ), .A2(_06474_ ), .A3(_06476_ ), .ZN(_06477_ ) );
MUX2_X2 _14494_ ( .A(_06477_ ), .B(_06457_ ), .S(_06453_ ), .Z(_06478_ ) );
AND2_X4 _14495_ ( .A1(_06467_ ), .A2(_06478_ ), .ZN(_06479_ ) );
XNOR2_X1 _14496_ ( .A(_06439_ ), .B(_04977_ ), .ZN(_06480_ ) );
AND2_X2 _14497_ ( .A1(_06479_ ), .A2(_06480_ ), .ZN(_06481_ ) );
INV_X1 _14498_ ( .A(_06481_ ), .ZN(_06482_ ) );
XNOR2_X1 _14499_ ( .A(_06438_ ), .B(_04984_ ), .ZN(_06483_ ) );
NOR2_X1 _14500_ ( .A1(_06483_ ), .A2(_04977_ ), .ZN(_06484_ ) );
INV_X1 _14501_ ( .A(_06484_ ), .ZN(_06485_ ) );
INV_X1 _14502_ ( .A(_06483_ ), .ZN(_06486_ ) );
BUF_X4 _14503_ ( .A(_04945_ ), .Z(_06487_ ) );
BUF_X4 _14504_ ( .A(_06487_ ), .Z(_06488_ ) );
BUF_X4 _14505_ ( .A(_06488_ ), .Z(_06489_ ) );
BUF_X4 _14506_ ( .A(_06433_ ), .Z(_06490_ ) );
XNOR2_X1 _14507_ ( .A(_06489_ ), .B(_06490_ ), .ZN(_06491_ ) );
BUF_X4 _14508_ ( .A(_04961_ ), .Z(_06492_ ) );
BUF_X4 _14509_ ( .A(_06492_ ), .Z(_06493_ ) );
BUF_X4 _14510_ ( .A(_06493_ ), .Z(_06494_ ) );
NOR2_X1 _14511_ ( .A1(_06491_ ), .A2(_06494_ ), .ZN(_06495_ ) );
INV_X1 _14512_ ( .A(_06495_ ), .ZN(_06496_ ) );
XNOR2_X1 _14513_ ( .A(_06436_ ), .B(_04939_ ), .ZN(_06497_ ) );
INV_X1 _14514_ ( .A(_06497_ ), .ZN(_06498_ ) );
BUF_X2 _14515_ ( .A(_06498_ ), .Z(_06499_ ) );
NAND4_X1 _14516_ ( .A1(_06467_ ), .A2(_06478_ ), .A3(_06496_ ), .A4(_06499_ ), .ZN(_06500_ ) );
AOI22_X1 _14517_ ( .A1(_06482_ ), .A2(_06485_ ), .B1(_06486_ ), .B2(_06500_ ), .ZN(_06501_ ) );
BUF_X4 _14518_ ( .A(_06492_ ), .Z(_06502_ ) );
BUF_X4 _14519_ ( .A(_04943_ ), .Z(_06503_ ) );
BUF_X4 _14520_ ( .A(_04944_ ), .Z(_06504_ ) );
BUF_X2 _14521_ ( .A(_04951_ ), .Z(_06505_ ) );
BUF_X2 _14522_ ( .A(_06505_ ), .Z(_06506_ ) );
BUF_X2 _14523_ ( .A(_04952_ ), .Z(_06507_ ) );
BUF_X2 _14524_ ( .A(_06507_ ), .Z(_06508_ ) );
AND3_X1 _14525_ ( .A1(_05052_ ), .A2(_06506_ ), .A3(_06508_ ), .ZN(_06509_ ) );
AOI21_X1 _14526_ ( .A(_02179_ ), .B1(_06506_ ), .B2(_06508_ ), .ZN(_06510_ ) );
OAI211_X1 _14527_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06509_ ), .C2(_06510_ ), .ZN(_06511_ ) );
BUF_X4 _14528_ ( .A(_06487_ ), .Z(_06512_ ) );
BUF_X4 _14529_ ( .A(_06512_ ), .Z(_06513_ ) );
AND3_X1 _14530_ ( .A1(_04088_ ), .A2(_06506_ ), .A3(_06508_ ), .ZN(_06514_ ) );
AOI21_X1 _14531_ ( .A(_04113_ ), .B1(_06506_ ), .B2(_06508_ ), .ZN(_06515_ ) );
OAI21_X1 _14532_ ( .A(_06513_ ), .B1(_06514_ ), .B2(_06515_ ), .ZN(_06516_ ) );
AOI21_X1 _14533_ ( .A(_06502_ ), .B1(_06511_ ), .B2(_06516_ ), .ZN(_06517_ ) );
BUF_X4 _14534_ ( .A(_06435_ ), .Z(_06518_ ) );
BUF_X4 _14535_ ( .A(_06518_ ), .Z(_06519_ ) );
CLKBUF_X2 _14536_ ( .A(_04952_ ), .Z(_06520_ ) );
BUF_X2 _14537_ ( .A(_06520_ ), .Z(_06521_ ) );
CLKBUF_X2 _14538_ ( .A(_06521_ ), .Z(_06522_ ) );
AND3_X1 _14539_ ( .A1(_04854_ ), .A2(_06506_ ), .A3(_06522_ ), .ZN(_06523_ ) );
CLKBUF_X2 _14540_ ( .A(_04951_ ), .Z(_06524_ ) );
BUF_X2 _14541_ ( .A(_06524_ ), .Z(_06525_ ) );
CLKBUF_X2 _14542_ ( .A(_06525_ ), .Z(_06526_ ) );
AOI21_X1 _14543_ ( .A(_04364_ ), .B1(_06526_ ), .B2(_06522_ ), .ZN(_06527_ ) );
OAI211_X1 _14544_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06523_ ), .C2(_06527_ ), .ZN(_06528_ ) );
AND3_X1 _14545_ ( .A1(_05044_ ), .A2(_06525_ ), .A3(_06521_ ), .ZN(_06529_ ) );
AOI21_X1 _14546_ ( .A(_02815_ ), .B1(_06506_ ), .B2(_06508_ ), .ZN(_06530_ ) );
OAI21_X1 _14547_ ( .A(_06513_ ), .B1(_06529_ ), .B2(_06530_ ), .ZN(_06531_ ) );
AOI21_X1 _14548_ ( .A(_06519_ ), .B1(_06528_ ), .B2(_06531_ ), .ZN(_06532_ ) );
NOR2_X1 _14549_ ( .A1(_06517_ ), .A2(_06532_ ), .ZN(_06533_ ) );
AND2_X1 _14550_ ( .A1(_06490_ ), .A2(_02928_ ), .ZN(_06534_ ) );
INV_X1 _14551_ ( .A(_06534_ ), .ZN(_06535_ ) );
AND3_X1 _14552_ ( .A1(_06525_ ), .A2(_02090_ ), .A3(_06521_ ), .ZN(_06536_ ) );
AOI21_X1 _14553_ ( .A(_02894_ ), .B1(_06506_ ), .B2(_06508_ ), .ZN(_06537_ ) );
OR2_X1 _14554_ ( .A1(_06536_ ), .A2(_06537_ ), .ZN(_06538_ ) );
MUX2_X1 _14555_ ( .A(_06535_ ), .B(_06538_ ), .S(_06488_ ), .Z(_06539_ ) );
NOR2_X1 _14556_ ( .A1(_06539_ ), .A2(_06493_ ), .ZN(_06540_ ) );
BUF_X4 _14557_ ( .A(_04939_ ), .Z(_06541_ ) );
BUF_X4 _14558_ ( .A(_06541_ ), .Z(_06542_ ) );
MUX2_X1 _14559_ ( .A(_06533_ ), .B(_06540_ ), .S(_06542_ ), .Z(_06543_ ) );
BUF_X2 _14560_ ( .A(_04984_ ), .Z(_06544_ ) );
BUF_X2 _14561_ ( .A(_06544_ ), .Z(_06545_ ) );
BUF_X2 _14562_ ( .A(_06545_ ), .Z(_06546_ ) );
BUF_X2 _14563_ ( .A(_06546_ ), .Z(_06547_ ) );
AND2_X1 _14564_ ( .A1(_06543_ ), .A2(_06547_ ), .ZN(_06548_ ) );
OAI21_X1 _14565_ ( .A(_06432_ ), .B1(_06501_ ), .B2(_06548_ ), .ZN(_06549_ ) );
NOR2_X1 _14566_ ( .A1(fanout_net_6 ), .A2(\ID_EX_typ [1] ), .ZN(_06550_ ) );
INV_X1 _14567_ ( .A(_06550_ ), .ZN(_06551_ ) );
NOR2_X1 _14568_ ( .A1(_04823_ ), .A2(_06551_ ), .ZN(_06552_ ) );
INV_X1 _14569_ ( .A(_06552_ ), .ZN(_06553_ ) );
BUF_X2 _14570_ ( .A(_06553_ ), .Z(_06554_ ) );
AND2_X1 _14571_ ( .A1(_04929_ ), .A2(_04934_ ), .ZN(_06555_ ) );
INV_X1 _14572_ ( .A(_06555_ ), .ZN(_06556_ ) );
AND4_X1 _14573_ ( .A1(_02530_ ), .A2(_04972_ ), .A3(_04973_ ), .A4(_04989_ ), .ZN(_06557_ ) );
AND3_X2 _14574_ ( .A1(_04972_ ), .A2(_04973_ ), .A3(_04968_ ), .ZN(_06558_ ) );
AND2_X1 _14575_ ( .A1(_04977_ ), .A2(_02525_ ), .ZN(_06559_ ) );
NOR2_X1 _14576_ ( .A1(_04984_ ), .A2(_02533_ ), .ZN(_06560_ ) );
AOI21_X1 _14577_ ( .A(_06559_ ), .B1(_04979_ ), .B2(_06560_ ), .ZN(_06561_ ) );
INV_X1 _14578_ ( .A(_06561_ ), .ZN(_06562_ ) );
AOI221_X2 _14579_ ( .A(_06557_ ), .B1(_02477_ ), .B2(_06442_ ), .C1(_06558_ ), .C2(_06562_ ), .ZN(_06563_ ) );
NOR2_X4 _14580_ ( .A1(_06433_ ), .A2(_04950_ ), .ZN(_06564_ ) );
INV_X2 _14581_ ( .A(_06564_ ), .ZN(_06565_ ) );
NOR3_X4 _14582_ ( .A1(_06565_ ), .A2(_04947_ ), .A3(_04948_ ), .ZN(_06566_ ) );
INV_X2 _14583_ ( .A(_06566_ ), .ZN(_06567_ ) );
INV_X1 _14584_ ( .A(_04947_ ), .ZN(_06568_ ) );
AOI21_X4 _14585_ ( .A(_04959_ ), .B1(_06567_ ), .B2(_06568_ ), .ZN(_06569_ ) );
AND2_X1 _14586_ ( .A1(_04939_ ), .A2(_02352_ ), .ZN(_06570_ ) );
NOR2_X1 _14587_ ( .A1(_04957_ ), .A2(_04511_ ), .ZN(_06571_ ) );
OR3_X4 _14588_ ( .A1(_06569_ ), .A2(_06570_ ), .A3(_06571_ ), .ZN(_06572_ ) );
NOR2_X1 _14589_ ( .A1(_04939_ ), .A2(_02352_ ), .ZN(_06573_ ) );
INV_X1 _14590_ ( .A(_06573_ ), .ZN(_06574_ ) );
AND2_X2 _14591_ ( .A1(_04979_ ), .A2(_04985_ ), .ZN(_06575_ ) );
NAND4_X4 _14592_ ( .A1(_06572_ ), .A2(_06574_ ), .A3(_06558_ ), .A4(_06575_ ), .ZN(_06576_ ) );
AOI21_X2 _14593_ ( .A(_06556_ ), .B1(_06563_ ), .B2(_06576_ ), .ZN(_06577_ ) );
AND2_X2 _14594_ ( .A1(_04908_ ), .A2(_04915_ ), .ZN(_06578_ ) );
AND3_X2 _14595_ ( .A1(_05009_ ), .A2(_04897_ ), .A3(_06578_ ), .ZN(_06579_ ) );
AND2_X1 _14596_ ( .A1(_04924_ ), .A2(_04920_ ), .ZN(_06580_ ) );
NAND3_X2 _14597_ ( .A1(_06577_ ), .A2(_06579_ ), .A3(_06580_ ), .ZN(_06581_ ) );
NOR2_X1 _14598_ ( .A1(_04933_ ), .A2(_04700_ ), .ZN(_06582_ ) );
AND2_X1 _14599_ ( .A1(_04929_ ), .A2(_06582_ ), .ZN(_06583_ ) );
AOI21_X2 _14600_ ( .A(_06583_ ), .B1(_02678_ ), .B2(_06449_ ), .ZN(_06584_ ) );
INV_X1 _14601_ ( .A(_04924_ ), .ZN(_06585_ ) );
INV_X1 _14602_ ( .A(_04920_ ), .ZN(_06586_ ) );
NOR3_X1 _14603_ ( .A1(_06584_ ), .A2(_06585_ ), .A3(_06586_ ), .ZN(_06587_ ) );
NOR2_X1 _14604_ ( .A1(_04919_ ), .A2(_04676_ ), .ZN(_06588_ ) );
NAND2_X1 _14605_ ( .A1(_04924_ ), .A2(_06588_ ), .ZN(_06589_ ) );
OAI21_X1 _14606_ ( .A(_06589_ ), .B1(_04653_ ), .B2(_04923_ ), .ZN(_06590_ ) );
OAI21_X1 _14607_ ( .A(_06579_ ), .B1(_06587_ ), .B2(_06590_ ), .ZN(_06591_ ) );
NOR2_X1 _14608_ ( .A1(_04896_ ), .A2(_04629_ ), .ZN(_06592_ ) );
NAND3_X1 _14609_ ( .A1(_04902_ ), .A2(_04903_ ), .A3(_06592_ ), .ZN(_06593_ ) );
NOR2_X1 _14610_ ( .A1(_04913_ ), .A2(_04579_ ), .ZN(_06594_ ) );
NOR3_X1 _14611_ ( .A1(_06594_ ), .A2(_05005_ ), .A3(_04907_ ), .ZN(_06595_ ) );
AOI21_X1 _14612_ ( .A(_06595_ ), .B1(_04579_ ), .B2(_04913_ ), .ZN(_06596_ ) );
INV_X1 _14613_ ( .A(_06596_ ), .ZN(_06597_ ) );
NAND3_X1 _14614_ ( .A1(_06597_ ), .A2(_05009_ ), .A3(_04897_ ), .ZN(_06598_ ) );
AND4_X2 _14615_ ( .A1(_04902_ ), .A2(_06591_ ), .A3(_06593_ ), .A4(_06598_ ), .ZN(_06599_ ) );
AND2_X4 _14616_ ( .A1(_06581_ ), .A2(_06599_ ), .ZN(_06600_ ) );
INV_X4 _14617_ ( .A(_06600_ ), .ZN(_06601_ ) );
AND2_X1 _14618_ ( .A1(_04888_ ), .A2(_04892_ ), .ZN(_06602_ ) );
NAND4_X2 _14619_ ( .A1(_06601_ ), .A2(_04882_ ), .A3(_04878_ ), .A4(_06602_ ), .ZN(_06603_ ) );
NOR2_X1 _14620_ ( .A1(_04891_ ), .A2(_04218_ ), .ZN(_06604_ ) );
INV_X1 _14621_ ( .A(_06604_ ), .ZN(_06605_ ) );
AND2_X1 _14622_ ( .A1(_04887_ ), .A2(_04241_ ), .ZN(_06606_ ) );
NOR2_X1 _14623_ ( .A1(_04887_ ), .A2(_04241_ ), .ZN(_06607_ ) );
NOR3_X1 _14624_ ( .A1(_06605_ ), .A2(_06606_ ), .A3(_06607_ ), .ZN(_06608_ ) );
OAI211_X1 _14625_ ( .A(_04882_ ), .B(_04878_ ), .C1(_06608_ ), .C2(_06607_ ), .ZN(_06609_ ) );
OR2_X1 _14626_ ( .A1(_04881_ ), .A2(_04167_ ), .ZN(_06610_ ) );
INV_X1 _14627_ ( .A(_04877_ ), .ZN(_06611_ ) );
NAND3_X1 _14628_ ( .A1(_04882_ ), .A2(_02275_ ), .A3(_06611_ ), .ZN(_06612_ ) );
AND3_X1 _14629_ ( .A1(_06609_ ), .A2(_06610_ ), .A3(_06612_ ), .ZN(_06613_ ) );
AOI21_X1 _14630_ ( .A(_04874_ ), .B1(_06603_ ), .B2(_06613_ ), .ZN(_06614_ ) );
NOR2_X1 _14631_ ( .A1(_04872_ ), .A2(_04140_ ), .ZN(_06615_ ) );
OR2_X1 _14632_ ( .A1(_06614_ ), .A2(_06615_ ), .ZN(_06616_ ) );
AOI21_X1 _14633_ ( .A(_06554_ ), .B1(_06616_ ), .B2(_04864_ ), .ZN(_06617_ ) );
OAI21_X1 _14634_ ( .A(_06617_ ), .B1(_04864_ ), .B2(_06616_ ), .ZN(_06618_ ) );
BUF_X4 _14635_ ( .A(_06544_ ), .Z(_06619_ ) );
AND2_X1 _14636_ ( .A1(_04825_ ), .A2(fanout_net_6 ), .ZN(_06620_ ) );
NAND3_X1 _14637_ ( .A1(_06543_ ), .A2(_06619_ ), .A3(_06620_ ), .ZN(_06621_ ) );
INV_X1 _14638_ ( .A(_05163_ ), .ZN(_06622_ ) );
BUF_X2 _14639_ ( .A(_06518_ ), .Z(_06623_ ) );
INV_X1 _14640_ ( .A(_04945_ ), .ZN(_06624_ ) );
BUF_X2 _14641_ ( .A(_06624_ ), .Z(_06625_ ) );
BUF_X2 _14642_ ( .A(_06625_ ), .Z(_06626_ ) );
BUF_X2 _14643_ ( .A(_06626_ ), .Z(_06627_ ) );
BUF_X2 _14644_ ( .A(_06506_ ), .Z(_06628_ ) );
BUF_X2 _14645_ ( .A(_06508_ ), .Z(_06629_ ) );
AOI21_X1 _14646_ ( .A(_02525_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06630_ ) );
AND3_X1 _14647_ ( .A1(_02533_ ), .A2(_06628_ ), .A3(_06629_ ), .ZN(_06631_ ) );
NOR3_X1 _14648_ ( .A1(_06627_ ), .A2(_06630_ ), .A3(_06631_ ), .ZN(_06632_ ) );
AND3_X1 _14649_ ( .A1(_04511_ ), .A2(_06526_ ), .A3(_06522_ ), .ZN(_06633_ ) );
BUF_X2 _14650_ ( .A(_06488_ ), .Z(_06634_ ) );
AOI21_X1 _14651_ ( .A(_02352_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06635_ ) );
NOR3_X1 _14652_ ( .A1(_06633_ ), .A2(_06634_ ), .A3(_06635_ ), .ZN(_06636_ ) );
OAI21_X1 _14653_ ( .A(_06623_ ), .B1(_06632_ ), .B2(_06636_ ), .ZN(_06637_ ) );
AOI21_X1 _14654_ ( .A(_02399_ ), .B1(_06526_ ), .B2(_06522_ ), .ZN(_06638_ ) );
NOR2_X1 _14655_ ( .A1(_04953_ ), .A2(_06638_ ), .ZN(_06639_ ) );
BUF_X2 _14656_ ( .A(_06513_ ), .Z(_06640_ ) );
NAND3_X1 _14657_ ( .A1(_06639_ ), .A2(_06493_ ), .A3(_06640_ ), .ZN(_06641_ ) );
NAND2_X1 _14658_ ( .A1(_06637_ ), .A2(_06641_ ), .ZN(_06642_ ) );
BUF_X2 _14659_ ( .A(_06437_ ), .Z(_06643_ ) );
NAND2_X1 _14660_ ( .A1(_06642_ ), .A2(_06643_ ), .ZN(_06644_ ) );
INV_X1 _14661_ ( .A(_04984_ ), .ZN(_06645_ ) );
AOI21_X1 _14662_ ( .A(_06622_ ), .B1(_06644_ ), .B2(_06645_ ), .ZN(_06646_ ) );
BUF_X4 _14663_ ( .A(_06519_ ), .Z(_06647_ ) );
AND3_X1 _14664_ ( .A1(_04629_ ), .A2(_06526_ ), .A3(_06522_ ), .ZN(_06648_ ) );
INV_X1 _14665_ ( .A(_06648_ ), .ZN(_06649_ ) );
AOI21_X1 _14666_ ( .A(_02609_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06650_ ) );
INV_X1 _14667_ ( .A(_06650_ ), .ZN(_06651_ ) );
NAND3_X1 _14668_ ( .A1(_06649_ ), .A2(_06627_ ), .A3(_06651_ ), .ZN(_06652_ ) );
AOI21_X1 _14669_ ( .A(_02299_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06653_ ) );
INV_X1 _14670_ ( .A(_06653_ ), .ZN(_06654_ ) );
OAI211_X1 _14671_ ( .A(_06654_ ), .B(_06489_ ), .C1(_02322_ ), .C2(_06490_ ), .ZN(_06655_ ) );
AOI21_X1 _14672_ ( .A(_06647_ ), .B1(_06652_ ), .B2(_06655_ ), .ZN(_06656_ ) );
AND3_X1 _14673_ ( .A1(_04190_ ), .A2(_06526_ ), .A3(_06522_ ), .ZN(_06657_ ) );
AOI21_X1 _14674_ ( .A(_02252_ ), .B1(_06526_ ), .B2(_06508_ ), .ZN(_06658_ ) );
OAI211_X1 _14675_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06657_ ), .C2(_06658_ ), .ZN(_06659_ ) );
AND3_X1 _14676_ ( .A1(_04140_ ), .A2(_06506_ ), .A3(_06508_ ), .ZN(_06660_ ) );
OAI21_X1 _14677_ ( .A(_06634_ ), .B1(_06660_ ), .B2(_06515_ ), .ZN(_06661_ ) );
AND3_X1 _14678_ ( .A1(_06659_ ), .A2(_06623_ ), .A3(_06661_ ), .ZN(_06662_ ) );
OAI21_X1 _14679_ ( .A(_06643_ ), .B1(_06656_ ), .B2(_06662_ ), .ZN(_06663_ ) );
BUF_X4 _14680_ ( .A(_06503_ ), .Z(_06664_ ) );
BUF_X4 _14681_ ( .A(_06504_ ), .Z(_06665_ ) );
AND3_X1 _14682_ ( .A1(_04988_ ), .A2(_06526_ ), .A3(_06522_ ), .ZN(_06666_ ) );
AOI21_X1 _14683_ ( .A(_02477_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06667_ ) );
OAI211_X1 _14684_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06666_ ), .C2(_06667_ ), .ZN(_06668_ ) );
AND3_X1 _14685_ ( .A1(_04700_ ), .A2(_06526_ ), .A3(_06522_ ), .ZN(_06669_ ) );
AOI21_X1 _14686_ ( .A(_02678_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06670_ ) );
OAI21_X1 _14687_ ( .A(_06489_ ), .B1(_06669_ ), .B2(_06670_ ), .ZN(_06671_ ) );
NAND2_X1 _14688_ ( .A1(_06668_ ), .A2(_06671_ ), .ZN(_06672_ ) );
BUF_X4 _14689_ ( .A(_06502_ ), .Z(_06673_ ) );
NAND2_X1 _14690_ ( .A1(_06672_ ), .A2(_06673_ ), .ZN(_06674_ ) );
AND3_X1 _14691_ ( .A1(_04676_ ), .A2(_06526_ ), .A3(_06522_ ), .ZN(_06675_ ) );
AOI21_X1 _14692_ ( .A(_02702_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06676_ ) );
OR3_X1 _14693_ ( .A1(_06675_ ), .A2(_06676_ ), .A3(_06513_ ), .ZN(_06677_ ) );
AOI21_X1 _14694_ ( .A(_04579_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_06678_ ) );
INV_X1 _14695_ ( .A(_06678_ ), .ZN(_06679_ ) );
OAI211_X1 _14696_ ( .A(_06679_ ), .B(_06489_ ), .C1(_02561_ ), .C2(_06490_ ), .ZN(_06680_ ) );
NAND3_X1 _14697_ ( .A1(_06677_ ), .A2(_06647_ ), .A3(_06680_ ), .ZN(_06681_ ) );
NAND3_X1 _14698_ ( .A1(_06674_ ), .A2(_06681_ ), .A3(_06542_ ), .ZN(_06682_ ) );
NAND3_X1 _14699_ ( .A1(_06663_ ), .A2(_06682_ ), .A3(_06545_ ), .ZN(_06683_ ) );
NAND2_X1 _14700_ ( .A1(_06646_ ), .A2(_06683_ ), .ZN(_06684_ ) );
OAI211_X1 _14701_ ( .A(_06621_ ), .B(_06684_ ), .C1(_05026_ ), .C2(_04828_ ), .ZN(_06685_ ) );
BUF_X4 _14702_ ( .A(_04823_ ), .Z(_06686_ ) );
BUF_X4 _14703_ ( .A(_05166_ ), .Z(_06687_ ) );
AOI221_X4 _14704_ ( .A(_06685_ ), .B1(_05027_ ), .B2(_06686_ ), .C1(_04864_ ), .C2(_06687_ ), .ZN(_06688_ ) );
NAND3_X1 _14705_ ( .A1(_06549_ ), .A2(_06618_ ), .A3(_06688_ ), .ZN(_06689_ ) );
INV_X1 _14706_ ( .A(_06420_ ), .ZN(_06690_ ) );
NAND3_X1 _14707_ ( .A1(_06690_ ), .A2(_06405_ ), .A3(_06409_ ), .ZN(_06691_ ) );
AND4_X1 _14708_ ( .A1(\ID_EX_typ [3] ), .A2(_04826_ ), .A3(_04824_ ), .A4(\ID_EX_typ [0] ), .ZN(_06692_ ) );
MUX2_X1 _14709_ ( .A(_06692_ ), .B(_06419_ ), .S(\ID_EX_typ [4] ), .Z(_06693_ ) );
NOR2_X1 _14710_ ( .A1(_06691_ ), .A2(_06693_ ), .ZN(_06694_ ) );
NOR2_X1 _14711_ ( .A1(_06694_ ), .A2(_06426_ ), .ZN(_06695_ ) );
BUF_X4 _14712_ ( .A(_06695_ ), .Z(_06696_ ) );
INV_X1 _14713_ ( .A(_06696_ ), .ZN(_06697_ ) );
BUF_X4 _14714_ ( .A(_06697_ ), .Z(_06698_ ) );
AOI21_X1 _14715_ ( .A(_06429_ ), .B1(_06689_ ), .B2(_06698_ ), .ZN(_06699_ ) );
OAI21_X1 _14716_ ( .A(_06234_ ), .B1(_05824_ ), .B2(_05543_ ), .ZN(_06700_ ) );
OAI21_X1 _14717_ ( .A(_06400_ ), .B1(_06699_ ), .B2(_06700_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
NAND3_X1 _14718_ ( .A1(_05259_ ), .A2(_05261_ ), .A3(_06156_ ), .ZN(_06701_ ) );
NAND3_X1 _14719_ ( .A1(_06413_ ), .A2(_06415_ ), .A3(_05135_ ), .ZN(_06702_ ) );
NAND3_X1 _14720_ ( .A1(_06416_ ), .A2(_06422_ ), .A3(_06702_ ), .ZN(_06703_ ) );
BUF_X4 _14721_ ( .A(_06408_ ), .Z(_06704_ ) );
AOI22_X1 _14722_ ( .A1(_05264_ ), .A2(_06404_ ), .B1(\ID_EX_imm [20] ), .B2(_06704_ ), .ZN(_06705_ ) );
AOI21_X1 _14723_ ( .A(_06427_ ), .B1(_06703_ ), .B2(_06705_ ), .ZN(_06706_ ) );
OR2_X1 _14724_ ( .A1(_06706_ ), .A2(_05184_ ), .ZN(_06707_ ) );
BUF_X2 _14725_ ( .A(_06479_ ), .Z(_06708_ ) );
AND2_X1 _14726_ ( .A1(_06708_ ), .A2(_06498_ ), .ZN(_06709_ ) );
BUF_X4 _14727_ ( .A(_06673_ ), .Z(_06710_ ) );
OAI21_X1 _14728_ ( .A(_06709_ ), .B1(_06710_ ), .B2(_06434_ ), .ZN(_06711_ ) );
AOI22_X1 _14729_ ( .A1(_06711_ ), .A2(_06486_ ), .B1(_06485_ ), .B2(_06482_ ), .ZN(_06712_ ) );
NAND2_X1 _14730_ ( .A1(_06433_ ), .A2(_05044_ ), .ZN(_06713_ ) );
NAND3_X1 _14731_ ( .A1(_06525_ ), .A2(_05037_ ), .A3(_06521_ ), .ZN(_06714_ ) );
AND3_X1 _14732_ ( .A1(_06625_ ), .A2(_06713_ ), .A3(_06714_ ), .ZN(_06715_ ) );
NOR2_X1 _14733_ ( .A1(_06433_ ), .A2(_02815_ ), .ZN(_06716_ ) );
AOI21_X1 _14734_ ( .A(_02787_ ), .B1(_06525_ ), .B2(_06521_ ), .ZN(_06717_ ) );
NOR3_X1 _14735_ ( .A1(_06625_ ), .A2(_06716_ ), .A3(_06717_ ), .ZN(_06718_ ) );
NOR3_X1 _14736_ ( .A1(_06715_ ), .A2(_06718_ ), .A3(_06519_ ), .ZN(_06719_ ) );
AND3_X1 _14737_ ( .A1(_04051_ ), .A2(_06525_ ), .A3(_06521_ ), .ZN(_06720_ ) );
AOI21_X1 _14738_ ( .A(_02155_ ), .B1(_06525_ ), .B2(_06521_ ), .ZN(_06721_ ) );
OAI211_X1 _14739_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06720_ ), .C2(_06721_ ), .ZN(_06722_ ) );
AND3_X1 _14740_ ( .A1(_04114_ ), .A2(_06525_ ), .A3(_06521_ ), .ZN(_06723_ ) );
AOI21_X1 _14741_ ( .A(_02202_ ), .B1(_06525_ ), .B2(_06521_ ), .ZN(_06724_ ) );
OAI21_X1 _14742_ ( .A(_06512_ ), .B1(_06723_ ), .B2(_06724_ ), .ZN(_06725_ ) );
AOI21_X1 _14743_ ( .A(_06502_ ), .B1(_06722_ ), .B2(_06725_ ), .ZN(_06726_ ) );
NOR2_X1 _14744_ ( .A1(_06719_ ), .A2(_06726_ ), .ZN(_06727_ ) );
NAND2_X1 _14745_ ( .A1(_06433_ ), .A2(_04854_ ), .ZN(_06728_ ) );
NAND3_X1 _14746_ ( .A1(_06525_ ), .A2(_02900_ ), .A3(_06521_ ), .ZN(_06729_ ) );
AND2_X1 _14747_ ( .A1(_06728_ ), .A2(_06729_ ), .ZN(_06730_ ) );
MUX2_X1 _14748_ ( .A(_02928_ ), .B(_04340_ ), .S(_06433_ ), .Z(_06731_ ) );
MUX2_X1 _14749_ ( .A(_06730_ ), .B(_06731_ ), .S(_06625_ ), .Z(_06732_ ) );
AND2_X1 _14750_ ( .A1(_06732_ ), .A2(_06623_ ), .ZN(_06733_ ) );
MUX2_X1 _14751_ ( .A(_06727_ ), .B(_06733_ ), .S(_06542_ ), .Z(_06734_ ) );
AND2_X1 _14752_ ( .A1(_06734_ ), .A2(_06547_ ), .ZN(_06735_ ) );
OAI21_X1 _14753_ ( .A(_06432_ ), .B1(_06712_ ), .B2(_06735_ ), .ZN(_06736_ ) );
NOR2_X1 _14754_ ( .A1(_06614_ ), .A2(_06554_ ), .ZN(_06737_ ) );
AND2_X4 _14755_ ( .A1(_06603_ ), .A2(_06613_ ), .ZN(_06738_ ) );
INV_X4 _14756_ ( .A(_06738_ ), .ZN(_06739_ ) );
OAI21_X1 _14757_ ( .A(_06737_ ), .B1(_04873_ ), .B2(_06739_ ), .ZN(_06740_ ) );
BUF_X2 _14758_ ( .A(_06620_ ), .Z(_06741_ ) );
BUF_X2 _14759_ ( .A(_06741_ ), .Z(_06742_ ) );
NAND3_X1 _14760_ ( .A1(_06734_ ), .A2(_06547_ ), .A3(_06742_ ), .ZN(_06743_ ) );
NOR2_X1 _14761_ ( .A1(_06433_ ), .A2(_02399_ ), .ZN(_06744_ ) );
AOI21_X1 _14762_ ( .A(_02376_ ), .B1(_06524_ ), .B2(_06520_ ), .ZN(_06745_ ) );
OAI21_X1 _14763_ ( .A(_06626_ ), .B1(_06744_ ), .B2(_06745_ ), .ZN(_06746_ ) );
AND3_X1 _14764_ ( .A1(_04940_ ), .A2(_06524_ ), .A3(_06520_ ), .ZN(_06747_ ) );
AOI21_X1 _14765_ ( .A(_02452_ ), .B1(_06524_ ), .B2(_06520_ ), .ZN(_06748_ ) );
OAI21_X1 _14766_ ( .A(_06513_ ), .B1(_06747_ ), .B2(_06748_ ), .ZN(_06749_ ) );
NAND3_X1 _14767_ ( .A1(_06746_ ), .A2(_06623_ ), .A3(_06749_ ), .ZN(_06750_ ) );
AOI21_X1 _14768_ ( .A(_04950_ ), .B1(_06506_ ), .B2(_06508_ ), .ZN(_06751_ ) );
NAND3_X1 _14769_ ( .A1(_06751_ ), .A2(_06493_ ), .A3(_06640_ ), .ZN(_06752_ ) );
AOI21_X1 _14770_ ( .A(_06542_ ), .B1(_06750_ ), .B2(_06752_ ), .ZN(_06753_ ) );
INV_X1 _14771_ ( .A(_06753_ ), .ZN(_06754_ ) );
BUF_X4 _14772_ ( .A(_06645_ ), .Z(_06755_ ) );
AOI21_X1 _14773_ ( .A(_06622_ ), .B1(_06754_ ), .B2(_06755_ ), .ZN(_06756_ ) );
AND3_X1 _14774_ ( .A1(_04606_ ), .A2(_06505_ ), .A3(_06507_ ), .ZN(_06757_ ) );
AOI21_X1 _14775_ ( .A(_02322_ ), .B1(_06505_ ), .B2(_06507_ ), .ZN(_06758_ ) );
OR3_X1 _14776_ ( .A1(_06625_ ), .A2(_06757_ ), .A3(_06758_ ), .ZN(_06759_ ) );
AND3_X1 _14777_ ( .A1(_04914_ ), .A2(_06524_ ), .A3(_06520_ ), .ZN(_06760_ ) );
AOI21_X1 _14778_ ( .A(_02631_ ), .B1(_06505_ ), .B2(_06507_ ), .ZN(_06761_ ) );
OR3_X1 _14779_ ( .A1(_06760_ ), .A2(_06512_ ), .A3(_06761_ ), .ZN(_06762_ ) );
NAND3_X1 _14780_ ( .A1(_06759_ ), .A2(_06762_ ), .A3(_06494_ ), .ZN(_06763_ ) );
AND3_X1 _14781_ ( .A1(_04241_ ), .A2(_06524_ ), .A3(_06520_ ), .ZN(_06764_ ) );
AOI21_X1 _14782_ ( .A(_02275_ ), .B1(_06505_ ), .B2(_06507_ ), .ZN(_06765_ ) );
OAI211_X1 _14783_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06764_ ), .C2(_06765_ ), .ZN(_06766_ ) );
AND3_X1 _14784_ ( .A1(_04167_ ), .A2(_06505_ ), .A3(_06507_ ), .ZN(_06767_ ) );
OAI21_X1 _14785_ ( .A(_06640_ ), .B1(_06767_ ), .B2(_06724_ ), .ZN(_06768_ ) );
NAND2_X1 _14786_ ( .A1(_06766_ ), .A2(_06768_ ), .ZN(_06769_ ) );
BUF_X4 _14787_ ( .A(_06647_ ), .Z(_06770_ ) );
NAND2_X1 _14788_ ( .A1(_06769_ ), .A2(_06770_ ), .ZN(_06771_ ) );
AND2_X1 _14789_ ( .A1(_06763_ ), .A2(_06771_ ), .ZN(_06772_ ) );
AND3_X1 _14790_ ( .A1(_04653_ ), .A2(_06524_ ), .A3(_06520_ ), .ZN(_06773_ ) );
AOI21_X1 _14791_ ( .A(_02561_ ), .B1(_06505_ ), .B2(_06507_ ), .ZN(_06774_ ) );
OR3_X1 _14792_ ( .A1(_06625_ ), .A2(_06773_ ), .A3(_06774_ ), .ZN(_06775_ ) );
BUF_X2 _14793_ ( .A(_06519_ ), .Z(_06776_ ) );
AND3_X1 _14794_ ( .A1(_04723_ ), .A2(_06505_ ), .A3(_06507_ ), .ZN(_06777_ ) );
AOI21_X1 _14795_ ( .A(_02724_ ), .B1(_06505_ ), .B2(_06507_ ), .ZN(_06778_ ) );
OR3_X1 _14796_ ( .A1(_06777_ ), .A2(_06778_ ), .A3(_06512_ ), .ZN(_06779_ ) );
AND3_X1 _14797_ ( .A1(_06775_ ), .A2(_06776_ ), .A3(_06779_ ), .ZN(_06780_ ) );
AND3_X1 _14798_ ( .A1(_04749_ ), .A2(_06524_ ), .A3(_06520_ ), .ZN(_06781_ ) );
AOI21_X1 _14799_ ( .A(_02655_ ), .B1(_06505_ ), .B2(_06507_ ), .ZN(_06782_ ) );
NOR3_X1 _14800_ ( .A1(_06626_ ), .A2(_06781_ ), .A3(_06782_ ), .ZN(_06783_ ) );
AND3_X1 _14801_ ( .A1(_04978_ ), .A2(_06524_ ), .A3(_06520_ ), .ZN(_06784_ ) );
AOI21_X1 _14802_ ( .A(_02530_ ), .B1(_06524_ ), .B2(_06520_ ), .ZN(_06785_ ) );
NOR3_X1 _14803_ ( .A1(_06784_ ), .A2(_06488_ ), .A3(_06785_ ), .ZN(_06786_ ) );
NOR3_X1 _14804_ ( .A1(_06783_ ), .A2(_06786_ ), .A3(_06776_ ), .ZN(_06787_ ) );
NOR2_X1 _14805_ ( .A1(_06780_ ), .A2(_06787_ ), .ZN(_06788_ ) );
BUF_X4 _14806_ ( .A(_06542_ ), .Z(_06789_ ) );
BUF_X4 _14807_ ( .A(_06789_ ), .Z(_06790_ ) );
MUX2_X1 _14808_ ( .A(_06772_ ), .B(_06788_ ), .S(_06790_ ), .Z(_06791_ ) );
OAI21_X1 _14809_ ( .A(_06756_ ), .B1(_06791_ ), .B2(_06755_ ), .ZN(_06792_ ) );
AND2_X1 _14810_ ( .A1(_04873_ ), .A2(_06687_ ), .ZN(_06793_ ) );
INV_X1 _14811_ ( .A(_04823_ ), .ZN(_06794_ ) );
BUF_X2 _14812_ ( .A(_06794_ ), .Z(_06795_ ) );
NOR3_X1 _14813_ ( .A1(_04872_ ), .A2(_04140_ ), .A3(_06795_ ), .ZN(_06796_ ) );
BUF_X2 _14814_ ( .A(_04828_ ), .Z(_06797_ ) );
AOI21_X1 _14815_ ( .A(_06797_ ), .B1(_04872_ ), .B2(_04140_ ), .ZN(_06798_ ) );
NOR3_X1 _14816_ ( .A1(_06793_ ), .A2(_06796_ ), .A3(_06798_ ), .ZN(_06799_ ) );
AND3_X1 _14817_ ( .A1(_06743_ ), .A2(_06792_ ), .A3(_06799_ ), .ZN(_06800_ ) );
NAND3_X1 _14818_ ( .A1(_06736_ ), .A2(_06740_ ), .A3(_06800_ ), .ZN(_06801_ ) );
AOI21_X1 _14819_ ( .A(_06707_ ), .B1(_06801_ ), .B2(_06698_ ), .ZN(_06802_ ) );
NAND2_X1 _14820_ ( .A1(_05269_ ), .A2(_05852_ ), .ZN(_06803_ ) );
NAND2_X1 _14821_ ( .A1(_06803_ ), .A2(_06164_ ), .ZN(_06804_ ) );
OAI21_X1 _14822_ ( .A(_06701_ ), .B1(_06802_ ), .B2(_06804_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OR2_X1 _14823_ ( .A1(_05297_ ), .A2(_06090_ ), .ZN(_06805_ ) );
AND2_X1 _14824_ ( .A1(_04189_ ), .A2(_02275_ ), .ZN(_06806_ ) );
AND2_X1 _14825_ ( .A1(_04217_ ), .A2(_02322_ ), .ZN(_06807_ ) );
AOI21_X1 _14826_ ( .A(_06807_ ), .B1(_06412_ ), .B2(_04219_ ), .ZN(_06808_ ) );
OAI21_X1 _14827_ ( .A(_05129_ ), .B1(_06808_ ), .B2(_05127_ ), .ZN(_06809_ ) );
AOI21_X1 _14828_ ( .A(_06806_ ), .B1(_06809_ ), .B2(_04191_ ), .ZN(_06810_ ) );
XNOR2_X1 _14829_ ( .A(_06810_ ), .B(_04168_ ), .ZN(_06811_ ) );
NAND2_X1 _14830_ ( .A1(_06811_ ), .A2(_06422_ ), .ZN(_06812_ ) );
AOI22_X1 _14831_ ( .A1(_05280_ ), .A2(_06404_ ), .B1(\ID_EX_imm [19] ), .B2(_06704_ ), .ZN(_06813_ ) );
AOI21_X1 _14832_ ( .A(_06427_ ), .B1(_06812_ ), .B2(_06813_ ), .ZN(_06814_ ) );
OR2_X1 _14833_ ( .A1(_06814_ ), .A2(_03778_ ), .ZN(_06815_ ) );
OAI21_X1 _14834_ ( .A(_06513_ ), .B1(_06633_ ), .B2(_06635_ ), .ZN(_06816_ ) );
OAI21_X1 _14835_ ( .A(_06816_ ), .B1(_06639_ ), .B2(_06634_ ), .ZN(_06817_ ) );
NOR2_X1 _14836_ ( .A1(_06817_ ), .A2(_06673_ ), .ZN(_06818_ ) );
BUF_X4 _14837_ ( .A(_06437_ ), .Z(_06819_ ) );
BUF_X4 _14838_ ( .A(_06819_ ), .Z(_06820_ ) );
AND2_X1 _14839_ ( .A1(_06818_ ), .A2(_06820_ ), .ZN(_06821_ ) );
OAI21_X1 _14840_ ( .A(_05163_ ), .B1(_06821_ ), .B2(_06545_ ), .ZN(_06822_ ) );
NOR3_X1 _14841_ ( .A1(_06626_ ), .A2(_06666_ ), .A3(_06667_ ), .ZN(_06823_ ) );
NOR3_X1 _14842_ ( .A1(_06631_ ), .A2(_06513_ ), .A3(_06630_ ), .ZN(_06824_ ) );
NOR2_X1 _14843_ ( .A1(_06823_ ), .A2(_06824_ ), .ZN(_06825_ ) );
NAND2_X1 _14844_ ( .A1(_06825_ ), .A2(_06673_ ), .ZN(_06826_ ) );
OAI211_X1 _14845_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06669_ ), .C2(_06670_ ), .ZN(_06827_ ) );
OAI21_X1 _14846_ ( .A(_06634_ ), .B1(_06675_ ), .B2(_06676_ ), .ZN(_06828_ ) );
NAND2_X1 _14847_ ( .A1(_06827_ ), .A2(_06828_ ), .ZN(_06829_ ) );
NAND2_X1 _14848_ ( .A1(_06829_ ), .A2(_06647_ ), .ZN(_06830_ ) );
NAND3_X1 _14849_ ( .A1(_06826_ ), .A2(_06790_ ), .A3(_06830_ ), .ZN(_06831_ ) );
BUF_X2 _14850_ ( .A(_06645_ ), .Z(_06832_ ) );
OR3_X1 _14851_ ( .A1(_06627_ ), .A2(_06657_ ), .A3(_06658_ ), .ZN(_06833_ ) );
AND3_X1 _14852_ ( .A1(_04218_ ), .A2(_06526_ ), .A3(_06522_ ), .ZN(_06834_ ) );
INV_X1 _14853_ ( .A(_06834_ ), .ZN(_06835_ ) );
NAND3_X1 _14854_ ( .A1(_06835_ ), .A2(_06627_ ), .A3(_06654_ ), .ZN(_06836_ ) );
NAND2_X1 _14855_ ( .A1(_06833_ ), .A2(_06836_ ), .ZN(_06837_ ) );
NAND2_X1 _14856_ ( .A1(_06837_ ), .A2(_06770_ ), .ZN(_06838_ ) );
AND3_X1 _14857_ ( .A1(_05005_ ), .A2(_06628_ ), .A3(_06629_ ), .ZN(_06839_ ) );
OAI211_X1 _14858_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06839_ ), .C2(_06678_ ), .ZN(_06840_ ) );
OAI21_X1 _14859_ ( .A(_06640_ ), .B1(_06648_ ), .B2(_06650_ ), .ZN(_06841_ ) );
NAND3_X1 _14860_ ( .A1(_06840_ ), .A2(_06494_ ), .A3(_06841_ ), .ZN(_06842_ ) );
NAND2_X1 _14861_ ( .A1(_06838_ ), .A2(_06842_ ), .ZN(_06843_ ) );
BUF_X2 _14862_ ( .A(_06643_ ), .Z(_06844_ ) );
AOI21_X1 _14863_ ( .A(_06832_ ), .B1(_06843_ ), .B2(_06844_ ), .ZN(_06845_ ) );
AOI21_X1 _14864_ ( .A(_06822_ ), .B1(_06831_ ), .B2(_06845_ ), .ZN(_06846_ ) );
OAI211_X1 _14865_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06536_ ), .C2(_06537_ ), .ZN(_06847_ ) );
OAI21_X1 _14866_ ( .A(_06488_ ), .B1(_06523_ ), .B2(_06527_ ), .ZN(_06848_ ) );
NAND3_X1 _14867_ ( .A1(_06847_ ), .A2(_06848_ ), .A3(_06519_ ), .ZN(_06849_ ) );
NAND4_X1 _14868_ ( .A1(_06502_ ), .A2(_02928_ ), .A3(_06634_ ), .A4(_06490_ ), .ZN(_06850_ ) );
NAND2_X1 _14869_ ( .A1(_06849_ ), .A2(_06850_ ), .ZN(_06851_ ) );
NAND2_X1 _14870_ ( .A1(_06851_ ), .A2(_06541_ ), .ZN(_06852_ ) );
NOR3_X1 _14871_ ( .A1(_06626_ ), .A2(_06660_ ), .A3(_06658_ ), .ZN(_06853_ ) );
NOR3_X1 _14872_ ( .A1(_06514_ ), .A2(_06488_ ), .A3(_06515_ ), .ZN(_06854_ ) );
OR3_X1 _14873_ ( .A1(_06853_ ), .A2(_06854_ ), .A3(_06492_ ), .ZN(_06855_ ) );
NOR3_X1 _14874_ ( .A1(_06626_ ), .A2(_06509_ ), .A3(_06510_ ), .ZN(_06856_ ) );
NOR3_X1 _14875_ ( .A1(_06529_ ), .A2(_06512_ ), .A3(_06530_ ), .ZN(_06857_ ) );
OR3_X1 _14876_ ( .A1(_06856_ ), .A2(_06857_ ), .A3(_06518_ ), .ZN(_06858_ ) );
NAND2_X1 _14877_ ( .A1(_06855_ ), .A2(_06858_ ), .ZN(_06859_ ) );
OAI21_X1 _14878_ ( .A(_06852_ ), .B1(_06859_ ), .B2(_06542_ ), .ZN(_06860_ ) );
AND2_X1 _14879_ ( .A1(_06860_ ), .A2(_06544_ ), .ZN(_06861_ ) );
AND2_X4 _14880_ ( .A1(_06481_ ), .A2(_06483_ ), .ZN(_06862_ ) );
XNOR2_X1 _14881_ ( .A(_06434_ ), .B(_06518_ ), .ZN(_06863_ ) );
AND4_X1 _14882_ ( .A1(_06498_ ), .A2(_06479_ ), .A3(_06863_ ), .A4(_06480_ ), .ZN(_06864_ ) );
OR3_X1 _14883_ ( .A1(_06862_ ), .A2(_06861_ ), .A3(_06864_ ), .ZN(_06865_ ) );
AOI221_X4 _14884_ ( .A(_06846_ ), .B1(_06741_ ), .B2(_06861_ ), .C1(_06865_ ), .C2(_06431_ ), .ZN(_06866_ ) );
NAND2_X1 _14885_ ( .A1(_06601_ ), .A2(_06602_ ), .ZN(_06867_ ) );
AOI21_X1 _14886_ ( .A(_06607_ ), .B1(_04888_ ), .B2(_06604_ ), .ZN(_06868_ ) );
AND2_X1 _14887_ ( .A1(_06867_ ), .A2(_06868_ ), .ZN(_06869_ ) );
INV_X1 _14888_ ( .A(_04878_ ), .ZN(_06870_ ) );
OR2_X1 _14889_ ( .A1(_06869_ ), .A2(_06870_ ), .ZN(_06871_ ) );
OR2_X1 _14890_ ( .A1(_04877_ ), .A2(_04190_ ), .ZN(_06872_ ) );
NAND2_X1 _14891_ ( .A1(_06871_ ), .A2(_06872_ ), .ZN(_06873_ ) );
AOI21_X1 _14892_ ( .A(_06554_ ), .B1(_06873_ ), .B2(_04882_ ), .ZN(_06874_ ) );
OAI21_X1 _14893_ ( .A(_06874_ ), .B1(_04882_ ), .B2(_06873_ ), .ZN(_06875_ ) );
NOR3_X1 _14894_ ( .A1(_04881_ ), .A2(_04167_ ), .A3(_06795_ ), .ZN(_06876_ ) );
AOI21_X1 _14895_ ( .A(_06797_ ), .B1(_04881_ ), .B2(_04167_ ), .ZN(_06877_ ) );
OR2_X1 _14896_ ( .A1(_06876_ ), .A2(_06877_ ), .ZN(_06878_ ) );
BUF_X4 _14897_ ( .A(_06687_ ), .Z(_06879_ ) );
AOI21_X1 _14898_ ( .A(_06878_ ), .B1(_04882_ ), .B2(_06879_ ), .ZN(_06880_ ) );
NAND3_X1 _14899_ ( .A1(_06866_ ), .A2(_06875_ ), .A3(_06880_ ), .ZN(_06881_ ) );
AOI21_X1 _14900_ ( .A(_06815_ ), .B1(_06881_ ), .B2(_06698_ ), .ZN(_06882_ ) );
NAND2_X1 _14901_ ( .A1(_05284_ ), .A2(_05852_ ), .ZN(_06883_ ) );
NAND2_X1 _14902_ ( .A1(_06883_ ), .A2(_06164_ ), .ZN(_06884_ ) );
OAI21_X1 _14903_ ( .A(_06805_ ), .B1(_06882_ ), .B2(_06884_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
NAND2_X1 _14904_ ( .A1(_05323_ ), .A2(_06094_ ), .ZN(_06885_ ) );
BUF_X4 _14905_ ( .A(_06690_ ), .Z(_06886_ ) );
AOI21_X1 _14906_ ( .A(_06886_ ), .B1(_06809_ ), .B2(_04191_ ), .ZN(_06887_ ) );
OAI21_X1 _14907_ ( .A(_06887_ ), .B1(_04191_ ), .B2(_06809_ ), .ZN(_06888_ ) );
AOI22_X1 _14908_ ( .A1(_05305_ ), .A2(_06404_ ), .B1(\ID_EX_imm [18] ), .B2(_06704_ ), .ZN(_06889_ ) );
AOI21_X1 _14909_ ( .A(_06426_ ), .B1(_06888_ ), .B2(_06889_ ), .ZN(_06890_ ) );
OR2_X1 _14910_ ( .A1(_06890_ ), .A2(_03778_ ), .ZN(_06891_ ) );
INV_X1 _14911_ ( .A(_06490_ ), .ZN(_06892_ ) );
AND2_X1 _14912_ ( .A1(_06892_ ), .A2(_06488_ ), .ZN(_06893_ ) );
INV_X1 _14913_ ( .A(_06893_ ), .ZN(_06894_ ) );
NAND4_X1 _14914_ ( .A1(_06708_ ), .A2(_06894_ ), .A3(_06499_ ), .A4(_06863_ ), .ZN(_06895_ ) );
AOI22_X1 _14915_ ( .A1(_06482_ ), .A2(_06485_ ), .B1(_06486_ ), .B2(_06895_ ), .ZN(_06896_ ) );
AND3_X1 _14916_ ( .A1(_06731_ ), .A2(_06492_ ), .A3(_06634_ ), .ZN(_06897_ ) );
AOI22_X1 _14917_ ( .A1(_06713_ ), .A2(_06714_ ), .B1(_04943_ ), .B2(_04944_ ), .ZN(_06898_ ) );
AOI21_X1 _14918_ ( .A(_06487_ ), .B1(_06728_ ), .B2(_06729_ ), .ZN(_06899_ ) );
NOR3_X1 _14919_ ( .A1(_06898_ ), .A2(_06899_ ), .A3(_06492_ ), .ZN(_06900_ ) );
NOR2_X1 _14920_ ( .A1(_06897_ ), .A2(_06900_ ), .ZN(_06901_ ) );
NOR3_X1 _14921_ ( .A1(_06625_ ), .A2(_06720_ ), .A3(_06721_ ), .ZN(_06902_ ) );
NOR3_X1 _14922_ ( .A1(_06716_ ), .A2(_06512_ ), .A3(_06717_ ), .ZN(_06903_ ) );
OR3_X1 _14923_ ( .A1(_06902_ ), .A2(_06903_ ), .A3(_06518_ ), .ZN(_06904_ ) );
OAI211_X1 _14924_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06723_ ), .C2(_06724_ ), .ZN(_06905_ ) );
OAI21_X1 _14925_ ( .A(_06488_ ), .B1(_06767_ ), .B2(_06765_ ), .ZN(_06906_ ) );
NAND2_X1 _14926_ ( .A1(_06905_ ), .A2(_06906_ ), .ZN(_06907_ ) );
NAND2_X1 _14927_ ( .A1(_06907_ ), .A2(_06623_ ), .ZN(_06908_ ) );
NAND2_X1 _14928_ ( .A1(_06904_ ), .A2(_06908_ ), .ZN(_06909_ ) );
MUX2_X1 _14929_ ( .A(_06901_ ), .B(_06909_ ), .S(_06819_ ), .Z(_06910_ ) );
NOR2_X1 _14930_ ( .A1(_06910_ ), .A2(_06832_ ), .ZN(_06911_ ) );
OAI21_X1 _14931_ ( .A(_06432_ ), .B1(_06896_ ), .B2(_06911_ ), .ZN(_06912_ ) );
NOR3_X1 _14932_ ( .A1(_04877_ ), .A2(_04190_ ), .A3(_06795_ ), .ZN(_06913_ ) );
OAI21_X1 _14933_ ( .A(_06512_ ), .B1(_06744_ ), .B2(_06745_ ), .ZN(_06914_ ) );
OAI21_X1 _14934_ ( .A(_06914_ ), .B1(_06512_ ), .B2(_06751_ ), .ZN(_06915_ ) );
NOR2_X1 _14935_ ( .A1(_06915_ ), .A2(_06494_ ), .ZN(_06916_ ) );
AND2_X1 _14936_ ( .A1(_06916_ ), .A2(_06844_ ), .ZN(_06917_ ) );
OAI21_X1 _14937_ ( .A(_05163_ ), .B1(_06917_ ), .B2(_06546_ ), .ZN(_06918_ ) );
NOR3_X1 _14938_ ( .A1(_06625_ ), .A2(_06777_ ), .A3(_06778_ ), .ZN(_06919_ ) );
NOR3_X1 _14939_ ( .A1(_06781_ ), .A2(_06487_ ), .A3(_06782_ ), .ZN(_06920_ ) );
OAI21_X1 _14940_ ( .A(_06776_ ), .B1(_06919_ ), .B2(_06920_ ), .ZN(_06921_ ) );
NOR3_X1 _14941_ ( .A1(_06625_ ), .A2(_06784_ ), .A3(_06785_ ), .ZN(_06922_ ) );
NOR3_X1 _14942_ ( .A1(_06747_ ), .A2(_06512_ ), .A3(_06748_ ), .ZN(_06923_ ) );
OAI21_X1 _14943_ ( .A(_06494_ ), .B1(_06922_ ), .B2(_06923_ ), .ZN(_06924_ ) );
AND2_X1 _14944_ ( .A1(_06921_ ), .A2(_06924_ ), .ZN(_06925_ ) );
OR3_X1 _14945_ ( .A1(_06626_ ), .A2(_06764_ ), .A3(_06765_ ), .ZN(_06926_ ) );
OR3_X1 _14946_ ( .A1(_06757_ ), .A2(_06634_ ), .A3(_06758_ ), .ZN(_06927_ ) );
AND3_X1 _14947_ ( .A1(_06926_ ), .A2(_06647_ ), .A3(_06927_ ), .ZN(_06928_ ) );
OR3_X1 _14948_ ( .A1(_06624_ ), .A2(_06760_ ), .A3(_06761_ ), .ZN(_06929_ ) );
OR3_X1 _14949_ ( .A1(_06773_ ), .A2(_06487_ ), .A3(_06774_ ), .ZN(_06930_ ) );
AND3_X1 _14950_ ( .A1(_06929_ ), .A2(_06673_ ), .A3(_06930_ ), .ZN(_06931_ ) );
OR2_X1 _14951_ ( .A1(_06928_ ), .A2(_06931_ ), .ZN(_06932_ ) );
BUF_X4 _14952_ ( .A(_06820_ ), .Z(_06933_ ) );
MUX2_X1 _14953_ ( .A(_06925_ ), .B(_06932_ ), .S(_06933_ ), .Z(_06934_ ) );
AOI21_X1 _14954_ ( .A(_06918_ ), .B1(_06934_ ), .B2(_06547_ ), .ZN(_06935_ ) );
AOI211_X1 _14955_ ( .A(_06913_ ), .B(_06935_ ), .C1(_04878_ ), .C2(_06879_ ), .ZN(_06936_ ) );
AOI21_X1 _14956_ ( .A(_04828_ ), .B1(_04877_ ), .B2(_04190_ ), .ZN(_06937_ ) );
XNOR2_X1 _14957_ ( .A(_06869_ ), .B(_04878_ ), .ZN(_06938_ ) );
AOI221_X4 _14958_ ( .A(_06937_ ), .B1(_06741_ ), .B2(_06911_ ), .C1(_06938_ ), .C2(_06552_ ), .ZN(_06939_ ) );
NAND3_X1 _14959_ ( .A1(_06912_ ), .A2(_06936_ ), .A3(_06939_ ), .ZN(_06940_ ) );
AOI21_X1 _14960_ ( .A(_06891_ ), .B1(_06940_ ), .B2(_06698_ ), .ZN(_06941_ ) );
OAI21_X1 _14961_ ( .A(_06234_ ), .B1(_05304_ ), .B2(_05543_ ), .ZN(_06942_ ) );
OAI21_X1 _14962_ ( .A(_06885_ ), .B1(_06941_ ), .B2(_06942_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
INV_X1 _14963_ ( .A(_06146_ ), .ZN(_06943_ ) );
NAND2_X1 _14964_ ( .A1(_05356_ ), .A2(_05251_ ), .ZN(_06944_ ) );
INV_X1 _14965_ ( .A(_06144_ ), .ZN(_06945_ ) );
OAI211_X1 _14966_ ( .A(_06943_ ), .B(_06136_ ), .C1(_06944_ ), .C2(_06945_ ), .ZN(_06946_ ) );
XNOR2_X1 _14967_ ( .A(_06808_ ), .B(_04242_ ), .ZN(_06947_ ) );
NAND2_X1 _14968_ ( .A1(_06947_ ), .A2(_06422_ ), .ZN(_06948_ ) );
AOI22_X1 _14969_ ( .A1(_05330_ ), .A2(_06404_ ), .B1(\ID_EX_imm [17] ), .B2(_06704_ ), .ZN(_06949_ ) );
AOI21_X1 _14970_ ( .A(_06426_ ), .B1(_06948_ ), .B2(_06949_ ), .ZN(_06950_ ) );
OR2_X1 _14971_ ( .A1(_06950_ ), .A2(_03778_ ), .ZN(_06951_ ) );
AND3_X1 _14972_ ( .A1(_06708_ ), .A2(_06499_ ), .A3(_06863_ ), .ZN(_06952_ ) );
NAND2_X1 _14973_ ( .A1(_06952_ ), .A2(_06491_ ), .ZN(_06953_ ) );
AOI22_X1 _14974_ ( .A1(_06953_ ), .A2(_06486_ ), .B1(_06482_ ), .B2(_06485_ ), .ZN(_06954_ ) );
NOR3_X1 _14975_ ( .A1(_06626_ ), .A2(_06657_ ), .A3(_06653_ ), .ZN(_06955_ ) );
NOR3_X1 _14976_ ( .A1(_06660_ ), .A2(_06513_ ), .A3(_06658_ ), .ZN(_06956_ ) );
NOR3_X1 _14977_ ( .A1(_06955_ ), .A2(_06956_ ), .A3(_06493_ ), .ZN(_06957_ ) );
AOI21_X1 _14978_ ( .A(_06623_ ), .B1(_06511_ ), .B2(_06516_ ), .ZN(_06958_ ) );
OR2_X1 _14979_ ( .A1(_06957_ ), .A2(_06958_ ), .ZN(_06959_ ) );
NAND2_X1 _14980_ ( .A1(_06539_ ), .A2(_06673_ ), .ZN(_06960_ ) );
NAND2_X1 _14981_ ( .A1(_06528_ ), .A2(_06531_ ), .ZN(_06961_ ) );
NAND2_X1 _14982_ ( .A1(_06961_ ), .A2(_06647_ ), .ZN(_06962_ ) );
NAND2_X1 _14983_ ( .A1(_06960_ ), .A2(_06962_ ), .ZN(_06963_ ) );
MUX2_X1 _14984_ ( .A(_06959_ ), .B(_06963_ ), .S(_06789_ ), .Z(_06964_ ) );
NOR2_X1 _14985_ ( .A1(_06964_ ), .A2(_06755_ ), .ZN(_06965_ ) );
OAI21_X1 _14986_ ( .A(_06432_ ), .B1(_06954_ ), .B2(_06965_ ), .ZN(_06966_ ) );
AND3_X1 _14987_ ( .A1(_06639_ ), .A2(_06623_ ), .A3(_06640_ ), .ZN(_06967_ ) );
AND2_X1 _14988_ ( .A1(_06967_ ), .A2(_06643_ ), .ZN(_06968_ ) );
OAI21_X1 _14989_ ( .A(_05163_ ), .B1(_06968_ ), .B2(_06545_ ), .ZN(_06969_ ) );
AND3_X1 _14990_ ( .A1(_06677_ ), .A2(_06493_ ), .A3(_06680_ ), .ZN(_06970_ ) );
AND2_X1 _14991_ ( .A1(_06652_ ), .A2(_06655_ ), .ZN(_06971_ ) );
AOI21_X1 _14992_ ( .A(_06970_ ), .B1(_06770_ ), .B2(_06971_ ), .ZN(_06972_ ) );
AOI21_X1 _14993_ ( .A(_06832_ ), .B1(_06972_ ), .B2(_06933_ ), .ZN(_06973_ ) );
OR3_X1 _14994_ ( .A1(_06632_ ), .A2(_06636_ ), .A3(_06776_ ), .ZN(_06974_ ) );
BUF_X2 _14995_ ( .A(_06542_ ), .Z(_06975_ ) );
NAND2_X1 _14996_ ( .A1(_06672_ ), .A2(_06770_ ), .ZN(_06976_ ) );
NAND3_X1 _14997_ ( .A1(_06974_ ), .A2(_06975_ ), .A3(_06976_ ), .ZN(_06977_ ) );
AOI21_X1 _14998_ ( .A(_06969_ ), .B1(_06973_ ), .B2(_06977_ ), .ZN(_06978_ ) );
BUF_X4 _14999_ ( .A(_06686_ ), .Z(_06979_ ) );
AOI221_X4 _15000_ ( .A(_06978_ ), .B1(_06607_ ), .B2(_06979_ ), .C1(_04888_ ), .C2(_06879_ ), .ZN(_06980_ ) );
AOI21_X1 _15001_ ( .A(_06797_ ), .B1(_04887_ ), .B2(_04241_ ), .ZN(_06981_ ) );
INV_X1 _15002_ ( .A(_04892_ ), .ZN(_06982_ ) );
AOI21_X1 _15003_ ( .A(_06982_ ), .B1(_06581_ ), .B2(_06599_ ), .ZN(_06983_ ) );
OR3_X1 _15004_ ( .A1(_06983_ ), .A2(_04888_ ), .A3(_06604_ ), .ZN(_06984_ ) );
OAI21_X1 _15005_ ( .A(_04888_ ), .B1(_06983_ ), .B2(_06604_ ), .ZN(_06985_ ) );
AND3_X1 _15006_ ( .A1(_06984_ ), .A2(_06552_ ), .A3(_06985_ ), .ZN(_06986_ ) );
AOI211_X1 _15007_ ( .A(_06981_ ), .B(_06986_ ), .C1(_06742_ ), .C2(_06965_ ), .ZN(_06987_ ) );
NAND3_X1 _15008_ ( .A1(_06966_ ), .A2(_06980_ ), .A3(_06987_ ), .ZN(_06988_ ) );
AOI21_X1 _15009_ ( .A(_06951_ ), .B1(_06988_ ), .B2(_06698_ ), .ZN(_06989_ ) );
NAND2_X1 _15010_ ( .A1(_05337_ ), .A2(_05852_ ), .ZN(_06990_ ) );
NAND2_X1 _15011_ ( .A1(_06990_ ), .A2(_06164_ ), .ZN(_06991_ ) );
OAI21_X1 _15012_ ( .A(_06946_ ), .B1(_06989_ ), .B2(_06991_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _15013_ ( .A1(_05363_ ), .A2(_05365_ ), .A3(_06156_ ), .ZN(_06992_ ) );
AOI21_X1 _15014_ ( .A(_06690_ ), .B1(_06412_ ), .B2(_04219_ ), .ZN(_06993_ ) );
OAI21_X1 _15015_ ( .A(_06993_ ), .B1(_04219_ ), .B2(_06412_ ), .ZN(_06994_ ) );
BUF_X2 _15016_ ( .A(_06404_ ), .Z(_06995_ ) );
NAND2_X1 _15017_ ( .A1(_05368_ ), .A2(_06995_ ), .ZN(_06996_ ) );
CLKBUF_X2 _15018_ ( .A(_06402_ ), .Z(_06997_ ) );
NAND3_X1 _15019_ ( .A1(_06407_ ), .A2(\ID_EX_imm [16] ), .A3(_06997_ ), .ZN(_06998_ ) );
AND3_X1 _15020_ ( .A1(_06994_ ), .A2(_06996_ ), .A3(_06998_ ), .ZN(_06999_ ) );
OAI21_X1 _15021_ ( .A(_05498_ ), .B1(_06999_ ), .B2(_06428_ ), .ZN(_07000_ ) );
INV_X1 _15022_ ( .A(_06430_ ), .ZN(_07001_ ) );
BUF_X4 _15023_ ( .A(_07001_ ), .Z(_07002_ ) );
OAI211_X1 _15024_ ( .A(_06708_ ), .B(_06480_ ), .C1(_06755_ ), .C2(_06438_ ), .ZN(_07003_ ) );
OR3_X1 _15025_ ( .A1(_06624_ ), .A2(_06764_ ), .A3(_06758_ ), .ZN(_07004_ ) );
OR3_X1 _15026_ ( .A1(_06767_ ), .A2(_06487_ ), .A3(_06765_ ), .ZN(_07005_ ) );
AND3_X1 _15027_ ( .A1(_07004_ ), .A2(_07005_ ), .A3(_06435_ ), .ZN(_07006_ ) );
AOI21_X1 _15028_ ( .A(_06435_ ), .B1(_06722_ ), .B2(_06725_ ), .ZN(_07007_ ) );
NOR2_X1 _15029_ ( .A1(_07006_ ), .A2(_07007_ ), .ZN(_07008_ ) );
NOR2_X1 _15030_ ( .A1(_07008_ ), .A2(_06541_ ), .ZN(_07009_ ) );
OR3_X1 _15031_ ( .A1(_06715_ ), .A2(_06718_ ), .A3(_04961_ ), .ZN(_07010_ ) );
OAI21_X1 _15032_ ( .A(_07010_ ), .B1(_06732_ ), .B2(_06519_ ), .ZN(_07011_ ) );
AOI21_X1 _15033_ ( .A(_07009_ ), .B1(_06541_ ), .B2(_07011_ ), .ZN(_07012_ ) );
NAND2_X1 _15034_ ( .A1(_07012_ ), .A2(_06547_ ), .ZN(_07013_ ) );
AOI21_X1 _15035_ ( .A(_07002_ ), .B1(_07003_ ), .B2(_07013_ ), .ZN(_07014_ ) );
OAI21_X1 _15036_ ( .A(_06552_ ), .B1(_06600_ ), .B2(_06982_ ), .ZN(_07015_ ) );
AOI21_X1 _15037_ ( .A(_07015_ ), .B1(_06982_ ), .B2(_06600_ ), .ZN(_07016_ ) );
OAI21_X1 _15038_ ( .A(_06519_ ), .B1(_06783_ ), .B2(_06786_ ), .ZN(_07017_ ) );
NAND3_X1 _15039_ ( .A1(_06746_ ), .A2(_06502_ ), .A3(_06749_ ), .ZN(_07018_ ) );
AND3_X1 _15040_ ( .A1(_07017_ ), .A2(_06541_ ), .A3(_07018_ ), .ZN(_07019_ ) );
AND3_X1 _15041_ ( .A1(_06775_ ), .A2(_06492_ ), .A3(_06779_ ), .ZN(_07020_ ) );
AND2_X1 _15042_ ( .A1(_06759_ ), .A2(_06762_ ), .ZN(_07021_ ) );
AOI21_X1 _15043_ ( .A(_07020_ ), .B1(_06647_ ), .B2(_07021_ ), .ZN(_07022_ ) );
INV_X1 _15044_ ( .A(_07022_ ), .ZN(_07023_ ) );
AOI211_X1 _15045_ ( .A(_06645_ ), .B(_07019_ ), .C1(_07023_ ), .C2(_06820_ ), .ZN(_07024_ ) );
AND3_X1 _15046_ ( .A1(_06640_ ), .A2(_06623_ ), .A3(_06751_ ), .ZN(_07025_ ) );
AND3_X1 _15047_ ( .A1(_07025_ ), .A2(_06643_ ), .A3(_06645_ ), .ZN(_07026_ ) );
OAI21_X1 _15048_ ( .A(_05163_ ), .B1(_07024_ ), .B2(_07026_ ), .ZN(_07027_ ) );
OAI221_X1 _15049_ ( .A(_07027_ ), .B1(_06605_ ), .B2(_06795_ ), .C1(_06982_ ), .C2(_05167_ ), .ZN(_07028_ ) );
AND3_X1 _15050_ ( .A1(_07012_ ), .A2(_06619_ ), .A3(_06741_ ), .ZN(_07029_ ) );
AOI21_X1 _15051_ ( .A(_04828_ ), .B1(_04891_ ), .B2(_04218_ ), .ZN(_07030_ ) );
OR3_X1 _15052_ ( .A1(_07028_ ), .A2(_07029_ ), .A3(_07030_ ), .ZN(_07031_ ) );
OR3_X1 _15053_ ( .A1(_07014_ ), .A2(_07016_ ), .A3(_07031_ ), .ZN(_07032_ ) );
AOI21_X1 _15054_ ( .A(_07000_ ), .B1(_07032_ ), .B2(_06698_ ), .ZN(_07033_ ) );
OAI21_X1 _15055_ ( .A(_06234_ ), .B1(_05367_ ), .B2(_05543_ ), .ZN(_07034_ ) );
OAI21_X1 _15056_ ( .A(_06992_ ), .B1(_07033_ ), .B2(_07034_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OAI21_X1 _15057_ ( .A(_06156_ ), .B1(_05379_ ), .B2(_05380_ ), .ZN(_07035_ ) );
NAND4_X1 _15058_ ( .A1(_06708_ ), .A2(_06431_ ), .A3(_06483_ ), .A4(_06480_ ), .ZN(_07036_ ) );
AND2_X1 _15059_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_07037_ ) );
OR3_X1 _15060_ ( .A1(_06853_ ), .A2(_06854_ ), .A3(_06623_ ), .ZN(_07038_ ) );
NOR3_X1 _15061_ ( .A1(_06626_ ), .A2(_06834_ ), .A3(_06650_ ), .ZN(_07039_ ) );
NOR3_X1 _15062_ ( .A1(_06657_ ), .A2(_06513_ ), .A3(_06653_ ), .ZN(_07040_ ) );
OR3_X1 _15063_ ( .A1(_07039_ ), .A2(_07040_ ), .A3(_06502_ ), .ZN(_07041_ ) );
NAND3_X1 _15064_ ( .A1(_07038_ ), .A2(_07041_ ), .A3(_06933_ ), .ZN(_07042_ ) );
OAI21_X1 _15065_ ( .A(_06518_ ), .B1(_06856_ ), .B2(_06857_ ), .ZN(_07043_ ) );
NAND3_X1 _15066_ ( .A1(_06847_ ), .A2(_06848_ ), .A3(_06492_ ), .ZN(_07044_ ) );
NAND2_X1 _15067_ ( .A1(_07043_ ), .A2(_07044_ ), .ZN(_07045_ ) );
NAND2_X1 _15068_ ( .A1(_07045_ ), .A2(_06790_ ), .ZN(_07046_ ) );
AOI21_X1 _15069_ ( .A(_06755_ ), .B1(_07042_ ), .B2(_07046_ ), .ZN(_07047_ ) );
AND3_X1 _15070_ ( .A1(_06534_ ), .A2(_06518_ ), .A3(_06634_ ), .ZN(_07048_ ) );
AND3_X1 _15071_ ( .A1(_07048_ ), .A2(_06832_ ), .A3(_06933_ ), .ZN(_07049_ ) );
OAI21_X1 _15072_ ( .A(_07037_ ), .B1(_07047_ ), .B2(_07049_ ), .ZN(_07050_ ) );
MUX2_X1 _15073_ ( .A(_06817_ ), .B(_06825_ ), .S(_06623_ ), .Z(_07051_ ) );
BUF_X2 _15074_ ( .A(_06975_ ), .Z(_07052_ ) );
NAND2_X1 _15075_ ( .A1(_07051_ ), .A2(_07052_ ), .ZN(_07053_ ) );
BUF_X2 _15076_ ( .A(_06820_ ), .Z(_07054_ ) );
AOI21_X1 _15077_ ( .A(_06673_ ), .B1(_06840_ ), .B2(_06841_ ), .ZN(_07055_ ) );
AOI21_X1 _15078_ ( .A(_06647_ ), .B1(_06827_ ), .B2(_06828_ ), .ZN(_07056_ ) );
OAI21_X1 _15079_ ( .A(_07054_ ), .B1(_07055_ ), .B2(_07056_ ), .ZN(_07057_ ) );
AND2_X2 _15080_ ( .A1(_04984_ ), .A2(_05163_ ), .ZN(_07058_ ) );
BUF_X2 _15081_ ( .A(_07058_ ), .Z(_07059_ ) );
NAND3_X1 _15082_ ( .A1(_07053_ ), .A2(_07057_ ), .A3(_07059_ ), .ZN(_07060_ ) );
AOI22_X1 _15083_ ( .A1(_05009_ ), .A2(_05166_ ), .B1(_04903_ ), .B2(_04827_ ), .ZN(_07061_ ) );
OR3_X1 _15084_ ( .A1(_04900_ ), .A2(_04606_ ), .A3(_06794_ ), .ZN(_07062_ ) );
AND2_X1 _15085_ ( .A1(_07061_ ), .A2(_07062_ ), .ZN(_07063_ ) );
AND4_X1 _15086_ ( .A1(_07036_ ), .A2(_07050_ ), .A3(_07060_ ), .A4(_07063_ ), .ZN(_07064_ ) );
INV_X1 _15087_ ( .A(_06578_ ), .ZN(_07065_ ) );
AND2_X1 _15088_ ( .A1(_06577_ ), .A2(_06580_ ), .ZN(_07066_ ) );
INV_X1 _15089_ ( .A(_07066_ ), .ZN(_07067_ ) );
NOR2_X1 _15090_ ( .A1(_06587_ ), .A2(_06590_ ), .ZN(_07068_ ) );
AOI21_X1 _15091_ ( .A(_07065_ ), .B1(_07067_ ), .B2(_07068_ ), .ZN(_07069_ ) );
NOR2_X1 _15092_ ( .A1(_07069_ ), .A2(_06597_ ), .ZN(_07070_ ) );
INV_X1 _15093_ ( .A(_04897_ ), .ZN(_07071_ ) );
NOR2_X1 _15094_ ( .A1(_07070_ ), .A2(_07071_ ), .ZN(_07072_ ) );
OR3_X1 _15095_ ( .A1(_07072_ ), .A2(_05009_ ), .A3(_06592_ ), .ZN(_07073_ ) );
BUF_X2 _15096_ ( .A(_06552_ ), .Z(_07074_ ) );
OAI21_X1 _15097_ ( .A(_05009_ ), .B1(_07072_ ), .B2(_06592_ ), .ZN(_07075_ ) );
NAND3_X1 _15098_ ( .A1(_07073_ ), .A2(_07074_ ), .A3(_07075_ ), .ZN(_07076_ ) );
AOI21_X1 _15099_ ( .A(_06696_ ), .B1(_07064_ ), .B2(_07076_ ), .ZN(_07077_ ) );
AOI21_X1 _15100_ ( .A(_05094_ ), .B1(_05116_ ), .B2(_04725_ ), .ZN(_07078_ ) );
XNOR2_X1 _15101_ ( .A(_04578_ ), .B(_04914_ ), .ZN(_07079_ ) );
INV_X1 _15102_ ( .A(_07079_ ), .ZN(_07080_ ) );
NOR3_X1 _15103_ ( .A1(_07078_ ), .A2(_04557_ ), .A3(_07080_ ), .ZN(_07081_ ) );
OAI21_X1 _15104_ ( .A(_04630_ ), .B1(_07081_ ), .B2(_05098_ ), .ZN(_07082_ ) );
NAND2_X1 _15105_ ( .A1(_04628_ ), .A2(_02631_ ), .ZN(_07083_ ) );
NAND2_X1 _15106_ ( .A1(_07082_ ), .A2(_07083_ ), .ZN(_07084_ ) );
OAI21_X1 _15107_ ( .A(_06420_ ), .B1(_07084_ ), .B2(_04607_ ), .ZN(_07085_ ) );
AOI21_X1 _15108_ ( .A(_07085_ ), .B1(_04607_ ), .B2(_07084_ ), .ZN(_07086_ ) );
AOI21_X1 _15109_ ( .A(_07086_ ), .B1(\ID_EX_imm [15] ), .B2(_06704_ ), .ZN(_07087_ ) );
NAND2_X1 _15110_ ( .A1(_05389_ ), .A2(_06995_ ), .ZN(_07088_ ) );
AOI21_X1 _15111_ ( .A(_06427_ ), .B1(_07087_ ), .B2(_07088_ ), .ZN(_07089_ ) );
OR2_X1 _15112_ ( .A1(_07089_ ), .A2(_05184_ ), .ZN(_07090_ ) );
BUF_X4 _15113_ ( .A(_05181_ ), .Z(_07091_ ) );
OAI22_X1 _15114_ ( .A1(_07077_ ), .A2(_07090_ ), .B1(_07091_ ), .B2(_05384_ ), .ZN(_07092_ ) );
OAI21_X1 _15115_ ( .A(_07035_ ), .B1(_07092_ ), .B2(_06211_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
OR3_X1 _15116_ ( .A1(_07081_ ), .A2(_04630_ ), .A3(_05098_ ), .ZN(_07093_ ) );
AND3_X1 _15117_ ( .A1(_07093_ ), .A2(_06421_ ), .A3(_07082_ ), .ZN(_07094_ ) );
OR3_X1 _15118_ ( .A1(_05409_ ), .A2(_05387_ ), .A3(_06405_ ), .ZN(_07095_ ) );
OAI21_X1 _15119_ ( .A(_07095_ ), .B1(_02632_ ), .B2(_06410_ ), .ZN(_07096_ ) );
OAI21_X1 _15120_ ( .A(_06425_ ), .B1(_07094_ ), .B2(_07096_ ), .ZN(_07097_ ) );
INV_X4 _15121_ ( .A(_06479_ ), .ZN(_07098_ ) );
INV_X1 _15122_ ( .A(_06480_ ), .ZN(_07099_ ) );
AND2_X1 _15123_ ( .A1(_06893_ ), .A2(_06518_ ), .ZN(_07100_ ) );
AND2_X1 _15124_ ( .A1(_06497_ ), .A2(_07100_ ), .ZN(_07101_ ) );
OR4_X4 _15125_ ( .A1(_06486_ ), .A2(_07098_ ), .A3(_07099_ ), .A4(_07101_ ), .ZN(_07102_ ) );
AND3_X1 _15126_ ( .A1(_06731_ ), .A2(_06435_ ), .A3(_06488_ ), .ZN(_07103_ ) );
AND2_X1 _15127_ ( .A1(_07103_ ), .A2(_06437_ ), .ZN(_07104_ ) );
OR2_X1 _15128_ ( .A1(_07104_ ), .A2(_04984_ ), .ZN(_07105_ ) );
OR3_X1 _15129_ ( .A1(_06898_ ), .A2(_06899_ ), .A3(_06435_ ), .ZN(_07106_ ) );
OAI21_X1 _15130_ ( .A(_06518_ ), .B1(_06902_ ), .B2(_06903_ ), .ZN(_07107_ ) );
NAND2_X1 _15131_ ( .A1(_07106_ ), .A2(_07107_ ), .ZN(_07108_ ) );
NAND2_X1 _15132_ ( .A1(_07108_ ), .A2(_06541_ ), .ZN(_07109_ ) );
NOR3_X1 _15133_ ( .A1(_06625_ ), .A2(_06757_ ), .A3(_06761_ ), .ZN(_07110_ ) );
NOR3_X1 _15134_ ( .A1(_06764_ ), .A2(_06512_ ), .A3(_06758_ ), .ZN(_07111_ ) );
OR3_X1 _15135_ ( .A1(_07110_ ), .A2(_07111_ ), .A3(_06492_ ), .ZN(_07112_ ) );
NAND2_X1 _15136_ ( .A1(_06907_ ), .A2(_06492_ ), .ZN(_07113_ ) );
NAND3_X1 _15137_ ( .A1(_07112_ ), .A2(_06437_ ), .A3(_07113_ ), .ZN(_07114_ ) );
NAND3_X1 _15138_ ( .A1(_07109_ ), .A2(_04984_ ), .A3(_07114_ ), .ZN(_07115_ ) );
NAND2_X1 _15139_ ( .A1(_07105_ ), .A2(_07115_ ), .ZN(_07116_ ) );
AOI21_X1 _15140_ ( .A(_07001_ ), .B1(_07102_ ), .B2(_07116_ ), .ZN(_07117_ ) );
OAI21_X1 _15141_ ( .A(_06552_ ), .B1(_07070_ ), .B2(_07071_ ), .ZN(_07118_ ) );
AOI21_X1 _15142_ ( .A(_07118_ ), .B1(_07071_ ), .B2(_07070_ ), .ZN(_07119_ ) );
AND3_X1 _15143_ ( .A1(_06929_ ), .A2(_06435_ ), .A3(_06930_ ), .ZN(_07120_ ) );
NOR3_X1 _15144_ ( .A1(_06919_ ), .A2(_06920_ ), .A3(_06435_ ), .ZN(_07121_ ) );
OR3_X1 _15145_ ( .A1(_07120_ ), .A2(_06541_ ), .A3(_07121_ ), .ZN(_07122_ ) );
NOR2_X1 _15146_ ( .A1(_06922_ ), .A2(_06923_ ), .ZN(_07123_ ) );
MUX2_X1 _15147_ ( .A(_06915_ ), .B(_07123_ ), .S(_06518_ ), .Z(_07124_ ) );
OAI21_X1 _15148_ ( .A(_07122_ ), .B1(_06819_ ), .B2(_07124_ ), .ZN(_07125_ ) );
NAND2_X1 _15149_ ( .A1(_07125_ ), .A2(_07058_ ), .ZN(_07126_ ) );
OR3_X1 _15150_ ( .A1(_04896_ ), .A2(_04629_ ), .A3(_06794_ ), .ZN(_07127_ ) );
OAI211_X1 _15151_ ( .A(_07126_ ), .B(_07127_ ), .C1(_07071_ ), .C2(_05167_ ), .ZN(_07128_ ) );
AND3_X1 _15152_ ( .A1(_07105_ ), .A2(_07115_ ), .A3(_06620_ ), .ZN(_07129_ ) );
AOI21_X1 _15153_ ( .A(_04828_ ), .B1(_04896_ ), .B2(_04629_ ), .ZN(_07130_ ) );
OR3_X1 _15154_ ( .A1(_07128_ ), .A2(_07129_ ), .A3(_07130_ ), .ZN(_07131_ ) );
NOR3_X1 _15155_ ( .A1(_07117_ ), .A2(_07119_ ), .A3(_07131_ ), .ZN(_07132_ ) );
OAI21_X1 _15156_ ( .A(_07097_ ), .B1(_07132_ ), .B2(_06696_ ), .ZN(_07133_ ) );
MUX2_X2 _15157_ ( .A(_05408_ ), .B(_07133_ ), .S(_05180_ ), .Z(_07134_ ) );
MUX2_X1 _15158_ ( .A(_05406_ ), .B(_07134_ ), .S(_06099_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
NAND3_X1 _15159_ ( .A1(_05427_ ), .A2(_05429_ ), .A3(_06156_ ), .ZN(_07135_ ) );
OR2_X1 _15160_ ( .A1(_07078_ ), .A2(_04557_ ), .ZN(_07136_ ) );
AND2_X1 _15161_ ( .A1(_07136_ ), .A2(_05096_ ), .ZN(_07137_ ) );
OAI21_X1 _15162_ ( .A(_06421_ ), .B1(_07137_ ), .B2(_07080_ ), .ZN(_07138_ ) );
AOI21_X1 _15163_ ( .A(_07138_ ), .B1(_07080_ ), .B2(_07137_ ), .ZN(_07139_ ) );
AND2_X1 _15164_ ( .A1(_05417_ ), .A2(_06995_ ), .ZN(_07140_ ) );
AND3_X1 _15165_ ( .A1(_06407_ ), .A2(\ID_EX_imm [13] ), .A3(_06997_ ), .ZN(_07141_ ) );
NOR3_X1 _15166_ ( .A1(_07139_ ), .A2(_07140_ ), .A3(_07141_ ), .ZN(_07142_ ) );
OAI21_X1 _15167_ ( .A(_05498_ ), .B1(_07142_ ), .B2(_06428_ ), .ZN(_07143_ ) );
OAI211_X1 _15168_ ( .A(_06481_ ), .B(_06483_ ), .C1(_06496_ ), .C2(_06499_ ), .ZN(_07144_ ) );
OAI21_X1 _15169_ ( .A(_06789_ ), .B1(_06517_ ), .B2(_06532_ ), .ZN(_07145_ ) );
NAND3_X1 _15170_ ( .A1(_06835_ ), .A2(_06627_ ), .A3(_06651_ ), .ZN(_07146_ ) );
OAI211_X1 _15171_ ( .A(_06679_ ), .B(_06489_ ), .C1(_02631_ ), .C2(_06490_ ), .ZN(_07147_ ) );
AND3_X1 _15172_ ( .A1(_07146_ ), .A2(_07147_ ), .A3(_06647_ ), .ZN(_07148_ ) );
NOR3_X1 _15173_ ( .A1(_06955_ ), .A2(_06956_ ), .A3(_06776_ ), .ZN(_07149_ ) );
NOR2_X1 _15174_ ( .A1(_07148_ ), .A2(_07149_ ), .ZN(_07150_ ) );
OAI211_X1 _15175_ ( .A(_06619_ ), .B(_07145_ ), .C1(_07150_ ), .C2(_06975_ ), .ZN(_07151_ ) );
NAND3_X1 _15176_ ( .A1(_06540_ ), .A2(_06832_ ), .A3(_06933_ ), .ZN(_07152_ ) );
AND2_X1 _15177_ ( .A1(_07151_ ), .A2(_07152_ ), .ZN(_07153_ ) );
AOI21_X1 _15178_ ( .A(_07002_ ), .B1(_07144_ ), .B2(_07153_ ), .ZN(_07154_ ) );
AOI21_X1 _15179_ ( .A(_04909_ ), .B1(_07067_ ), .B2(_07068_ ), .ZN(_07155_ ) );
NOR2_X1 _15180_ ( .A1(_04907_ ), .A2(_05005_ ), .ZN(_07156_ ) );
OR3_X1 _15181_ ( .A1(_07155_ ), .A2(_04915_ ), .A3(_07156_ ), .ZN(_07157_ ) );
OAI21_X1 _15182_ ( .A(_04915_ ), .B1(_07155_ ), .B2(_07156_ ), .ZN(_07158_ ) );
AND3_X1 _15183_ ( .A1(_07157_ ), .A2(_07074_ ), .A3(_07158_ ), .ZN(_07159_ ) );
AND3_X1 _15184_ ( .A1(_04913_ ), .A2(_04579_ ), .A3(_06686_ ), .ZN(_07160_ ) );
INV_X1 _15185_ ( .A(_07058_ ), .ZN(_07161_ ) );
NAND2_X1 _15186_ ( .A1(_06642_ ), .A2(_06789_ ), .ZN(_07162_ ) );
NAND3_X1 _15187_ ( .A1(_06674_ ), .A2(_06681_ ), .A3(_06820_ ), .ZN(_07163_ ) );
AOI21_X1 _15188_ ( .A(_07161_ ), .B1(_07162_ ), .B2(_07163_ ), .ZN(_07164_ ) );
AOI211_X1 _15189_ ( .A(_07160_ ), .B(_07164_ ), .C1(_04915_ ), .C2(_06687_ ), .ZN(_07165_ ) );
INV_X1 _15190_ ( .A(_06620_ ), .ZN(_07166_ ) );
OAI221_X1 _15191_ ( .A(_07165_ ), .B1(_06594_ ), .B2(_06797_ ), .C1(_07166_ ), .C2(_07153_ ), .ZN(_07167_ ) );
OR3_X1 _15192_ ( .A1(_07154_ ), .A2(_07159_ ), .A3(_07167_ ), .ZN(_07168_ ) );
AOI21_X1 _15193_ ( .A(_07143_ ), .B1(_07168_ ), .B2(_06698_ ), .ZN(_07169_ ) );
NAND2_X1 _15194_ ( .A1(_05420_ ), .A2(_05852_ ), .ZN(_07170_ ) );
NAND2_X1 _15195_ ( .A1(_07170_ ), .A2(_06164_ ), .ZN(_07171_ ) );
OAI21_X1 _15196_ ( .A(_07135_ ), .B1(_07169_ ), .B2(_07171_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
AND3_X1 _15197_ ( .A1(_05356_ ), .A2(_05251_ ), .A3(_05442_ ), .ZN(_07172_ ) );
INV_X1 _15198_ ( .A(_07172_ ), .ZN(_07173_ ) );
INV_X1 _15199_ ( .A(_05435_ ), .ZN(_07174_ ) );
NAND3_X1 _15200_ ( .A1(_07173_ ), .A2(_07174_ ), .A3(_06156_ ), .ZN(_07175_ ) );
NOR3_X1 _15201_ ( .A1(_06719_ ), .A2(_06643_ ), .A3(_06726_ ), .ZN(_07176_ ) );
OR3_X1 _15202_ ( .A1(_06624_ ), .A2(_06760_ ), .A3(_06774_ ), .ZN(_07177_ ) );
OR3_X1 _15203_ ( .A1(_06757_ ), .A2(_06487_ ), .A3(_06761_ ), .ZN(_07178_ ) );
NAND3_X1 _15204_ ( .A1(_07177_ ), .A2(_07178_ ), .A3(_06519_ ), .ZN(_07179_ ) );
NAND3_X1 _15205_ ( .A1(_07004_ ), .A2(_07005_ ), .A3(_06502_ ), .ZN(_07180_ ) );
AND3_X1 _15206_ ( .A1(_07179_ ), .A2(_07180_ ), .A3(_06819_ ), .ZN(_07181_ ) );
OAI21_X1 _15207_ ( .A(_06544_ ), .B1(_07176_ ), .B2(_07181_ ), .ZN(_07182_ ) );
NAND4_X1 _15208_ ( .A1(_06732_ ), .A2(_06645_ ), .A3(_06643_ ), .A4(_06770_ ), .ZN(_07183_ ) );
AOI21_X1 _15209_ ( .A(_07166_ ), .B1(_07182_ ), .B2(_07183_ ), .ZN(_07184_ ) );
NOR3_X1 _15210_ ( .A1(_06434_ ), .A2(_06541_ ), .A3(_06493_ ), .ZN(_07185_ ) );
OR4_X1 _15211_ ( .A1(_06486_ ), .A2(_07098_ ), .A3(_07099_ ), .A4(_07185_ ), .ZN(_07186_ ) );
AND2_X1 _15212_ ( .A1(_07182_ ), .A2(_07183_ ), .ZN(_07187_ ) );
AOI21_X1 _15213_ ( .A(_07001_ ), .B1(_07186_ ), .B2(_07187_ ), .ZN(_07188_ ) );
NOR2_X1 _15214_ ( .A1(_06788_ ), .A2(_06790_ ), .ZN(_07189_ ) );
AND2_X1 _15215_ ( .A1(_06750_ ), .A2(_06752_ ), .ZN(_07190_ ) );
AOI21_X1 _15216_ ( .A(_07189_ ), .B1(_07052_ ), .B2(_07190_ ), .ZN(_07191_ ) );
AOI211_X1 _15217_ ( .A(_07184_ ), .B(_07188_ ), .C1(_07059_ ), .C2(_07191_ ), .ZN(_07192_ ) );
AND3_X1 _15218_ ( .A1(_07067_ ), .A2(_04909_ ), .A3(_07068_ ), .ZN(_07193_ ) );
OR3_X1 _15219_ ( .A1(_07193_ ), .A2(_07155_ ), .A3(_06553_ ), .ZN(_07194_ ) );
NAND2_X1 _15220_ ( .A1(_04908_ ), .A2(_06687_ ), .ZN(_07195_ ) );
NAND3_X1 _15221_ ( .A1(_05006_ ), .A2(_02561_ ), .A3(_06686_ ), .ZN(_07196_ ) );
BUF_X4 _15222_ ( .A(_04827_ ), .Z(_07197_ ) );
OAI21_X1 _15223_ ( .A(_07197_ ), .B1(_05006_ ), .B2(_02561_ ), .ZN(_07198_ ) );
AND3_X1 _15224_ ( .A1(_07195_ ), .A2(_07196_ ), .A3(_07198_ ), .ZN(_07199_ ) );
AND3_X1 _15225_ ( .A1(_07192_ ), .A2(_07194_ ), .A3(_07199_ ), .ZN(_07200_ ) );
NOR2_X1 _15226_ ( .A1(_07200_ ), .A2(_06696_ ), .ZN(_07201_ ) );
NAND2_X1 _15227_ ( .A1(_07078_ ), .A2(_04557_ ), .ZN(_07202_ ) );
NAND3_X1 _15228_ ( .A1(_07136_ ), .A2(_06422_ ), .A3(_07202_ ), .ZN(_07203_ ) );
AOI22_X1 _15229_ ( .A1(_05446_ ), .A2(_06995_ ), .B1(\ID_EX_imm [12] ), .B2(_06704_ ), .ZN(_07204_ ) );
AOI21_X1 _15230_ ( .A(_06427_ ), .B1(_07203_ ), .B2(_07204_ ), .ZN(_07205_ ) );
NOR3_X1 _15231_ ( .A1(_07201_ ), .A2(_05852_ ), .A3(_07205_ ), .ZN(_07206_ ) );
BUF_X4 _15232_ ( .A(_06090_ ), .Z(_07207_ ) );
OAI21_X1 _15233_ ( .A(_07207_ ), .B1(_05445_ ), .B2(_05543_ ), .ZN(_07208_ ) );
OAI21_X1 _15234_ ( .A(_07175_ ), .B1(_07206_ ), .B2(_07208_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
NAND2_X1 _15235_ ( .A1(_03872_ ), .A2(_06094_ ), .ZN(_07209_ ) );
INV_X1 _15236_ ( .A(_05047_ ), .ZN(_07210_ ) );
AND2_X1 _15237_ ( .A1(_04864_ ), .A2(_04873_ ), .ZN(_07211_ ) );
NAND4_X4 _15238_ ( .A1(_06739_ ), .A2(_04860_ ), .A3(_04868_ ), .A4(_07211_ ), .ZN(_07212_ ) );
INV_X1 _15239_ ( .A(_04868_ ), .ZN(_07213_ ) );
AOI21_X1 _15240_ ( .A(_05027_ ), .B1(_04864_ ), .B2(_06615_ ), .ZN(_07214_ ) );
NOR3_X1 _15241_ ( .A1(_05015_ ), .A2(_07213_ ), .A3(_07214_ ), .ZN(_07215_ ) );
NOR2_X1 _15242_ ( .A1(_04859_ ), .A2(_04051_ ), .ZN(_07216_ ) );
NOR2_X1 _15243_ ( .A1(_04867_ ), .A2(_04088_ ), .ZN(_07217_ ) );
AND2_X1 _15244_ ( .A1(_04860_ ), .A2(_07217_ ), .ZN(_07218_ ) );
NOR3_X1 _15245_ ( .A1(_07215_ ), .A2(_07216_ ), .A3(_07218_ ), .ZN(_07219_ ) );
AND2_X4 _15246_ ( .A1(_07212_ ), .A2(_07219_ ), .ZN(_07220_ ) );
INV_X2 _15247_ ( .A(_07220_ ), .ZN(_07221_ ) );
NAND3_X2 _15248_ ( .A1(_07221_ ), .A2(_05055_ ), .A3(_05060_ ), .ZN(_07222_ ) );
AND2_X1 _15249_ ( .A1(_05053_ ), .A2(_05060_ ), .ZN(_07223_ ) );
AOI21_X1 _15250_ ( .A(_07223_ ), .B1(_02815_ ), .B2(_06463_ ), .ZN(_07224_ ) );
AOI211_X2 _15251_ ( .A(_05067_ ), .B(_07210_ ), .C1(_07222_ ), .C2(_07224_ ), .ZN(_07225_ ) );
INV_X1 _15252_ ( .A(_05039_ ), .ZN(_07226_ ) );
AOI21_X1 _15253_ ( .A(_05038_ ), .B1(_05045_ ), .B2(_07226_ ), .ZN(_07227_ ) );
INV_X1 _15254_ ( .A(_07227_ ), .ZN(_07228_ ) );
OAI211_X2 _15255_ ( .A(_04850_ ), .B(_04855_ ), .C1(_07225_ ), .C2(_07228_ ), .ZN(_07229_ ) );
INV_X1 _15256_ ( .A(_05080_ ), .ZN(_07230_ ) );
AND2_X1 _15257_ ( .A1(_04853_ ), .A2(_02125_ ), .ZN(_07231_ ) );
AOI21_X1 _15258_ ( .A(_05076_ ), .B1(_04850_ ), .B2(_07231_ ), .ZN(_07232_ ) );
AND3_X1 _15259_ ( .A1(_07229_ ), .A2(_07230_ ), .A3(_07232_ ), .ZN(_07233_ ) );
AOI21_X1 _15260_ ( .A(_07230_ ), .B1(_07229_ ), .B2(_07232_ ), .ZN(_07234_ ) );
OR3_X2 _15261_ ( .A1(_07233_ ), .A2(_07234_ ), .A3(_06553_ ), .ZN(_07235_ ) );
AND2_X1 _15262_ ( .A1(_07104_ ), .A2(_06544_ ), .ZN(_07236_ ) );
NAND3_X1 _15263_ ( .A1(_06467_ ), .A2(_06478_ ), .A3(_06484_ ), .ZN(_07237_ ) );
NOR2_X1 _15264_ ( .A1(_07237_ ), .A2(_07101_ ), .ZN(_07238_ ) );
OR3_X1 _15265_ ( .A1(_06862_ ), .A2(_07236_ ), .A3(_07238_ ), .ZN(_07239_ ) );
NAND2_X1 _15266_ ( .A1(_07239_ ), .A2(_06431_ ), .ZN(_07240_ ) );
NAND3_X1 _15267_ ( .A1(_06926_ ), .A2(_06494_ ), .A3(_06927_ ), .ZN(_07241_ ) );
OAI211_X1 _15268_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06767_ ), .C2(_06724_ ), .ZN(_07242_ ) );
OAI21_X1 _15269_ ( .A(_06640_ ), .B1(_06723_ ), .B2(_06721_ ), .ZN(_07243_ ) );
NAND2_X1 _15270_ ( .A1(_07242_ ), .A2(_07243_ ), .ZN(_07244_ ) );
NAND2_X1 _15271_ ( .A1(_07244_ ), .A2(_06770_ ), .ZN(_07245_ ) );
NAND3_X1 _15272_ ( .A1(_07241_ ), .A2(_07245_ ), .A3(_06789_ ), .ZN(_07246_ ) );
OAI211_X1 _15273_ ( .A(_06640_ ), .B(_06729_ ), .C1(_06892_ ), .C2(_04340_ ), .ZN(_07247_ ) );
NAND2_X1 _15274_ ( .A1(_06728_ ), .A2(_06714_ ), .ZN(_07248_ ) );
BUF_X4 _15275_ ( .A(_06489_ ), .Z(_07249_ ) );
OAI211_X1 _15276_ ( .A(_07247_ ), .B(_06776_ ), .C1(_07248_ ), .C2(_07249_ ), .ZN(_07250_ ) );
NOR2_X1 _15277_ ( .A1(_06720_ ), .A2(_06717_ ), .ZN(_07251_ ) );
NAND2_X1 _15278_ ( .A1(_07251_ ), .A2(_06627_ ), .ZN(_07252_ ) );
OAI211_X1 _15279_ ( .A(_06713_ ), .B(_06489_ ), .C1(_02815_ ), .C2(_06490_ ), .ZN(_07253_ ) );
NAND2_X1 _15280_ ( .A1(_07252_ ), .A2(_07253_ ), .ZN(_07254_ ) );
OAI211_X1 _15281_ ( .A(_06820_ ), .B(_07250_ ), .C1(_07254_ ), .C2(_06770_ ), .ZN(_07255_ ) );
NAND3_X1 _15282_ ( .A1(_07246_ ), .A2(_06619_ ), .A3(_07255_ ), .ZN(_07256_ ) );
AND2_X1 _15283_ ( .A1(_07256_ ), .A2(_05163_ ), .ZN(_07257_ ) );
BUF_X2 _15284_ ( .A(_06619_ ), .Z(_07258_ ) );
OAI21_X1 _15285_ ( .A(_07257_ ), .B1(_07125_ ), .B2(_07258_ ), .ZN(_07259_ ) );
OAI21_X1 _15286_ ( .A(_07197_ ), .B1(_06474_ ), .B2(_04340_ ), .ZN(_07260_ ) );
AND3_X1 _15287_ ( .A1(_07104_ ), .A2(_06544_ ), .A3(_06620_ ), .ZN(_07261_ ) );
AOI221_X4 _15288_ ( .A(_07261_ ), .B1(_04844_ ), .B2(_06686_ ), .C1(_05080_ ), .C2(_05166_ ), .ZN(_07262_ ) );
AND4_X1 _15289_ ( .A1(_07240_ ), .A2(_07259_ ), .A3(_07260_ ), .A4(_07262_ ), .ZN(_07263_ ) );
AOI21_X1 _15290_ ( .A(_06696_ ), .B1(_07235_ ), .B2(_07263_ ), .ZN(_07264_ ) );
AOI22_X1 _15291_ ( .A1(_04000_ ), .A2(_06995_ ), .B1(\ID_EX_imm [30] ), .B2(_06704_ ), .ZN(_07265_ ) );
NAND2_X1 _15292_ ( .A1(_06412_ ), .A2(_04244_ ), .ZN(_07266_ ) );
NAND2_X1 _15293_ ( .A1(_07266_ ), .A2(_05140_ ), .ZN(_07267_ ) );
NAND2_X1 _15294_ ( .A1(_07267_ ), .A2(_04435_ ), .ZN(_07268_ ) );
NAND2_X1 _15295_ ( .A1(_07268_ ), .A2(_05150_ ), .ZN(_07269_ ) );
NAND2_X1 _15296_ ( .A1(_07269_ ), .A2(_04292_ ), .ZN(_07270_ ) );
NAND3_X1 _15297_ ( .A1(_07270_ ), .A2(_05156_ ), .A3(_05154_ ), .ZN(_07271_ ) );
AOI21_X1 _15298_ ( .A(_06886_ ), .B1(_07271_ ), .B2(_04341_ ), .ZN(_07272_ ) );
OAI21_X1 _15299_ ( .A(_07272_ ), .B1(_04341_ ), .B2(_07271_ ), .ZN(_07273_ ) );
AOI21_X1 _15300_ ( .A(_06427_ ), .B1(_07265_ ), .B2(_07273_ ), .ZN(_07274_ ) );
OR2_X1 _15301_ ( .A1(_07274_ ), .A2(_05184_ ), .ZN(_07275_ ) );
OAI22_X1 _15302_ ( .A1(_07264_ ), .A2(_07275_ ), .B1(_07091_ ), .B2(_03891_ ), .ZN(_07276_ ) );
OAI21_X1 _15303_ ( .A(_07209_ ), .B1(_07276_ ), .B2(_06211_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
AND2_X2 _15304_ ( .A1(_06480_ ), .A2(_06483_ ), .ZN(_07277_ ) );
OAI211_X1 _15305_ ( .A(_06708_ ), .B(_07277_ ), .C1(_06499_ ), .C2(_06863_ ), .ZN(_07278_ ) );
AOI21_X1 _15306_ ( .A(_06643_ ), .B1(_06855_ ), .B2(_06858_ ), .ZN(_07279_ ) );
OAI21_X1 _15307_ ( .A(_06502_ ), .B1(_07039_ ), .B2(_07040_ ), .ZN(_07280_ ) );
OAI211_X1 _15308_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06648_ ), .C2(_06678_ ), .ZN(_07281_ ) );
OAI21_X1 _15309_ ( .A(_06634_ ), .B1(_06839_ ), .B2(_06676_ ), .ZN(_07282_ ) );
NAND3_X1 _15310_ ( .A1(_07281_ ), .A2(_06519_ ), .A3(_07282_ ), .ZN(_07283_ ) );
AND3_X1 _15311_ ( .A1(_07280_ ), .A2(_06819_ ), .A3(_07283_ ), .ZN(_07284_ ) );
OAI21_X1 _15312_ ( .A(_06544_ ), .B1(_07279_ ), .B2(_07284_ ), .ZN(_07285_ ) );
AOI21_X1 _15313_ ( .A(_06541_ ), .B1(_06849_ ), .B2(_06850_ ), .ZN(_07286_ ) );
OR2_X1 _15314_ ( .A1(_07286_ ), .A2(_06544_ ), .ZN(_07287_ ) );
NAND2_X1 _15315_ ( .A1(_07285_ ), .A2(_07287_ ), .ZN(_07288_ ) );
AOI21_X1 _15316_ ( .A(_07002_ ), .B1(_07278_ ), .B2(_07288_ ), .ZN(_07289_ ) );
INV_X1 _15317_ ( .A(_06577_ ), .ZN(_07290_ ) );
AOI21_X1 _15318_ ( .A(_06586_ ), .B1(_07290_ ), .B2(_06584_ ), .ZN(_07291_ ) );
OR3_X1 _15319_ ( .A1(_07291_ ), .A2(_04924_ ), .A3(_06588_ ), .ZN(_07292_ ) );
OAI21_X1 _15320_ ( .A(_04924_ ), .B1(_07291_ ), .B2(_06588_ ), .ZN(_07293_ ) );
AND3_X1 _15321_ ( .A1(_07292_ ), .A2(_06552_ ), .A3(_07293_ ), .ZN(_07294_ ) );
AND3_X1 _15322_ ( .A1(_07285_ ), .A2(_06741_ ), .A3(_07287_ ), .ZN(_07295_ ) );
AOI21_X1 _15323_ ( .A(_04828_ ), .B1(_04923_ ), .B2(_04653_ ), .ZN(_07296_ ) );
NAND3_X1 _15324_ ( .A1(_06826_ ), .A2(_06643_ ), .A3(_06830_ ), .ZN(_07297_ ) );
OR3_X1 _15325_ ( .A1(_06817_ ), .A2(_06819_ ), .A3(_06493_ ), .ZN(_07298_ ) );
NAND2_X1 _15326_ ( .A1(_07297_ ), .A2(_07298_ ), .ZN(_07299_ ) );
NAND2_X1 _15327_ ( .A1(_07299_ ), .A2(_07058_ ), .ZN(_07300_ ) );
OR3_X1 _15328_ ( .A1(_04923_ ), .A2(_04653_ ), .A3(_06794_ ), .ZN(_07301_ ) );
OAI211_X1 _15329_ ( .A(_07300_ ), .B(_07301_ ), .C1(_06585_ ), .C2(_05167_ ), .ZN(_07302_ ) );
OR4_X1 _15330_ ( .A1(_07294_ ), .A2(_07295_ ), .A3(_07296_ ), .A4(_07302_ ), .ZN(_07303_ ) );
OAI21_X1 _15331_ ( .A(_06697_ ), .B1(_07289_ ), .B2(_07303_ ), .ZN(_07304_ ) );
INV_X1 _15332_ ( .A(_04701_ ), .ZN(_07305_ ) );
INV_X1 _15333_ ( .A(_04724_ ), .ZN(_07306_ ) );
AOI211_X1 _15334_ ( .A(_07305_ ), .B(_07306_ ), .C1(_05110_ ), .C2(_05114_ ), .ZN(_07307_ ) );
NOR3_X1 _15335_ ( .A1(_07307_ ), .A2(_05087_ ), .A3(_05088_ ), .ZN(_07308_ ) );
INV_X1 _15336_ ( .A(_04677_ ), .ZN(_07309_ ) );
NOR2_X1 _15337_ ( .A1(_07308_ ), .A2(_07309_ ), .ZN(_07310_ ) );
OR3_X1 _15338_ ( .A1(_07310_ ), .A2(_04654_ ), .A3(_05090_ ), .ZN(_07311_ ) );
OAI21_X1 _15339_ ( .A(_04654_ ), .B1(_07310_ ), .B2(_05090_ ), .ZN(_07312_ ) );
AND4_X1 _15340_ ( .A1(_04835_ ), .A2(_07311_ ), .A3(_06419_ ), .A4(_07312_ ), .ZN(_07313_ ) );
NAND2_X1 _15341_ ( .A1(_05456_ ), .A2(_06995_ ), .ZN(_07314_ ) );
OAI21_X1 _15342_ ( .A(_07314_ ), .B1(_02703_ ), .B2(_06410_ ), .ZN(_07315_ ) );
OAI21_X1 _15343_ ( .A(_06425_ ), .B1(_07313_ ), .B2(_07315_ ), .ZN(_07316_ ) );
AOI21_X1 _15344_ ( .A(_05184_ ), .B1(_07304_ ), .B2(_07316_ ), .ZN(_07317_ ) );
NOR2_X1 _15345_ ( .A1(_05459_ ), .A2(_05245_ ), .ZN(_07318_ ) );
OAI21_X1 _15346_ ( .A(_06164_ ), .B1(_07317_ ), .B2(_07318_ ), .ZN(_07319_ ) );
NAND3_X1 _15347_ ( .A1(_05467_ ), .A2(_05471_ ), .A3(_06111_ ), .ZN(_07320_ ) );
NAND2_X1 _15348_ ( .A1(_07319_ ), .A2(_07320_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OR2_X1 _15349_ ( .A1(_05515_ ), .A2(_06090_ ), .ZN(_07321_ ) );
AND4_X1 _15350_ ( .A1(_06894_ ), .A2(_06467_ ), .A3(_06478_ ), .A4(_06863_ ), .ZN(_07322_ ) );
OAI21_X1 _15351_ ( .A(_07277_ ), .B1(_06709_ ), .B2(_07322_ ), .ZN(_07323_ ) );
AND3_X1 _15352_ ( .A1(_06904_ ), .A2(_06975_ ), .A3(_06908_ ), .ZN(_07324_ ) );
NOR3_X1 _15353_ ( .A1(_07110_ ), .A2(_07111_ ), .A3(_06519_ ), .ZN(_07325_ ) );
OAI211_X1 _15354_ ( .A(_06503_ ), .B(_06504_ ), .C1(_06760_ ), .C2(_06774_ ), .ZN(_07326_ ) );
OAI21_X1 _15355_ ( .A(_06513_ ), .B1(_06773_ ), .B2(_06778_ ), .ZN(_07327_ ) );
AOI21_X1 _15356_ ( .A(_06502_ ), .B1(_07326_ ), .B2(_07327_ ), .ZN(_07328_ ) );
NOR3_X1 _15357_ ( .A1(_07325_ ), .A2(_06975_ ), .A3(_07328_ ), .ZN(_07329_ ) );
OAI21_X1 _15358_ ( .A(_07258_ ), .B1(_07324_ ), .B2(_07329_ ), .ZN(_07330_ ) );
OAI211_X1 _15359_ ( .A(_06832_ ), .B(_07054_ ), .C1(_06897_ ), .C2(_06900_ ), .ZN(_07331_ ) );
NAND3_X1 _15360_ ( .A1(_07323_ ), .A2(_07330_ ), .A3(_07331_ ), .ZN(_07332_ ) );
NAND2_X1 _15361_ ( .A1(_07332_ ), .A2(_06432_ ), .ZN(_07333_ ) );
AND3_X1 _15362_ ( .A1(_07290_ ), .A2(_06586_ ), .A3(_06584_ ), .ZN(_07334_ ) );
NOR3_X1 _15363_ ( .A1(_07334_ ), .A2(_07291_ ), .A3(_06553_ ), .ZN(_07335_ ) );
AOI21_X1 _15364_ ( .A(_07166_ ), .B1(_07330_ ), .B2(_07331_ ), .ZN(_07336_ ) );
AOI21_X1 _15365_ ( .A(_06797_ ), .B1(_04919_ ), .B2(_04676_ ), .ZN(_07337_ ) );
NAND3_X1 _15366_ ( .A1(_06924_ ), .A2(_06921_ ), .A3(_06844_ ), .ZN(_07338_ ) );
OAI21_X1 _15367_ ( .A(_06975_ ), .B1(_06915_ ), .B2(_06710_ ), .ZN(_07339_ ) );
NAND3_X1 _15368_ ( .A1(_07338_ ), .A2(_07059_ ), .A3(_07339_ ), .ZN(_07340_ ) );
NAND3_X1 _15369_ ( .A1(_05001_ ), .A2(_02724_ ), .A3(_06686_ ), .ZN(_07341_ ) );
OAI211_X1 _15370_ ( .A(_07340_ ), .B(_07341_ ), .C1(_06586_ ), .C2(_05167_ ), .ZN(_07342_ ) );
NOR4_X1 _15371_ ( .A1(_07335_ ), .A2(_07336_ ), .A3(_07337_ ), .A4(_07342_ ), .ZN(_07343_ ) );
AOI21_X1 _15372_ ( .A(_06696_ ), .B1(_07333_ ), .B2(_07343_ ), .ZN(_07344_ ) );
OAI21_X1 _15373_ ( .A(_06421_ ), .B1(_07308_ ), .B2(_07309_ ), .ZN(_07345_ ) );
AOI21_X1 _15374_ ( .A(_07345_ ), .B1(_07309_ ), .B2(_07308_ ), .ZN(_07346_ ) );
NOR3_X1 _15375_ ( .A1(_05504_ ), .A2(_05454_ ), .A3(_06405_ ), .ZN(_07347_ ) );
AND3_X1 _15376_ ( .A1(_06407_ ), .A2(\ID_EX_imm [10] ), .A3(_06997_ ), .ZN(_07348_ ) );
NOR3_X1 _15377_ ( .A1(_07346_ ), .A2(_07347_ ), .A3(_07348_ ), .ZN(_07349_ ) );
NOR2_X1 _15378_ ( .A1(_07349_ ), .A2(_06428_ ), .ZN(_07350_ ) );
NOR3_X1 _15379_ ( .A1(_07344_ ), .A2(_05852_ ), .A3(_07350_ ), .ZN(_07351_ ) );
OAI21_X1 _15380_ ( .A(_07207_ ), .B1(_05503_ ), .B2(_05543_ ), .ZN(_07352_ ) );
OAI21_X1 _15381_ ( .A(_07321_ ), .B1(_07351_ ), .B2(_07352_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
OR2_X1 _15382_ ( .A1(_05529_ ), .A2(_06090_ ), .ZN(_07353_ ) );
OR2_X1 _15383_ ( .A1(_05115_ ), .A2(_07305_ ), .ZN(_07354_ ) );
NAND2_X1 _15384_ ( .A1(_04699_ ), .A2(_02655_ ), .ZN(_07355_ ) );
AND3_X1 _15385_ ( .A1(_07354_ ), .A2(_07355_ ), .A3(_07306_ ), .ZN(_07356_ ) );
AOI21_X1 _15386_ ( .A(_07306_ ), .B1(_07354_ ), .B2(_07355_ ), .ZN(_07357_ ) );
NOR3_X1 _15387_ ( .A1(_07356_ ), .A2(_07357_ ), .A3(_06886_ ), .ZN(_07358_ ) );
AND2_X1 _15388_ ( .A1(_05533_ ), .A2(_06995_ ), .ZN(_07359_ ) );
AND3_X1 _15389_ ( .A1(_06407_ ), .A2(\ID_EX_imm [9] ), .A3(_06997_ ), .ZN(_07360_ ) );
NOR3_X1 _15390_ ( .A1(_07358_ ), .A2(_07359_ ), .A3(_07360_ ), .ZN(_07361_ ) );
OAI21_X1 _15391_ ( .A(_05498_ ), .B1(_07361_ ), .B2(_06428_ ), .ZN(_07362_ ) );
OAI21_X1 _15392_ ( .A(_06789_ ), .B1(_06957_ ), .B2(_06958_ ), .ZN(_07363_ ) );
AND3_X1 _15393_ ( .A1(_07146_ ), .A2(_07147_ ), .A3(_06673_ ), .ZN(_07364_ ) );
OAI211_X1 _15394_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06839_ ), .C2(_06676_ ), .ZN(_07365_ ) );
OAI21_X1 _15395_ ( .A(_07249_ ), .B1(_06675_ ), .B2(_06670_ ), .ZN(_07366_ ) );
AOI21_X1 _15396_ ( .A(_06673_ ), .B1(_07365_ ), .B2(_07366_ ), .ZN(_07367_ ) );
NOR2_X1 _15397_ ( .A1(_07364_ ), .A2(_07367_ ), .ZN(_07368_ ) );
OAI211_X1 _15398_ ( .A(_07363_ ), .B(_06619_ ), .C1(_07368_ ), .C2(_06975_ ), .ZN(_07369_ ) );
NAND4_X1 _15399_ ( .A1(_06960_ ), .A2(_06832_ ), .A3(_06844_ ), .A4(_06962_ ), .ZN(_07370_ ) );
AOI21_X1 _15400_ ( .A(_07166_ ), .B1(_07369_ ), .B2(_07370_ ), .ZN(_07371_ ) );
AND4_X1 _15401_ ( .A1(_06491_ ), .A2(_06467_ ), .A3(_06478_ ), .A4(_06863_ ), .ZN(_07372_ ) );
OAI21_X1 _15402_ ( .A(_07277_ ), .B1(_06709_ ), .B2(_07372_ ), .ZN(_07373_ ) );
AND2_X1 _15403_ ( .A1(_07369_ ), .A2(_07370_ ), .ZN(_07374_ ) );
AOI21_X1 _15404_ ( .A(_07002_ ), .B1(_07373_ ), .B2(_07374_ ), .ZN(_07375_ ) );
NAND3_X1 _15405_ ( .A1(_06974_ ), .A2(_07054_ ), .A3(_06976_ ), .ZN(_07376_ ) );
BUF_X4 _15406_ ( .A(_06776_ ), .Z(_07377_ ) );
NAND4_X1 _15407_ ( .A1(_06639_ ), .A2(_06790_ ), .A3(_07377_ ), .A4(_07249_ ), .ZN(_07378_ ) );
NAND2_X1 _15408_ ( .A1(_07376_ ), .A2(_07378_ ), .ZN(_07379_ ) );
AOI211_X1 _15409_ ( .A(_07371_ ), .B(_07375_ ), .C1(_07059_ ), .C2(_07379_ ), .ZN(_07380_ ) );
AOI21_X1 _15410_ ( .A(_04935_ ), .B1(_06563_ ), .B2(_06576_ ), .ZN(_07381_ ) );
INV_X1 _15411_ ( .A(_07381_ ), .ZN(_07382_ ) );
INV_X1 _15412_ ( .A(_06582_ ), .ZN(_07383_ ) );
NAND3_X1 _15413_ ( .A1(_07382_ ), .A2(_04930_ ), .A3(_07383_ ), .ZN(_07384_ ) );
OAI21_X1 _15414_ ( .A(_04929_ ), .B1(_07381_ ), .B2(_06582_ ), .ZN(_07385_ ) );
NAND3_X1 _15415_ ( .A1(_07384_ ), .A2(_07074_ ), .A3(_07385_ ), .ZN(_07386_ ) );
NAND2_X1 _15416_ ( .A1(_04929_ ), .A2(_06879_ ), .ZN(_07387_ ) );
NAND3_X1 _15417_ ( .A1(_06449_ ), .A2(_02678_ ), .A3(_06979_ ), .ZN(_07388_ ) );
OAI21_X1 _15418_ ( .A(_07197_ ), .B1(_06449_ ), .B2(_02678_ ), .ZN(_07389_ ) );
AND3_X1 _15419_ ( .A1(_07387_ ), .A2(_07388_ ), .A3(_07389_ ), .ZN(_07390_ ) );
NAND3_X1 _15420_ ( .A1(_07380_ ), .A2(_07386_ ), .A3(_07390_ ), .ZN(_07391_ ) );
AOI21_X1 _15421_ ( .A(_07362_ ), .B1(_07391_ ), .B2(_06698_ ), .ZN(_07392_ ) );
NAND2_X1 _15422_ ( .A1(_05535_ ), .A2(_05852_ ), .ZN(_07393_ ) );
NAND2_X1 _15423_ ( .A1(_07393_ ), .A2(_06234_ ), .ZN(_07394_ ) );
OAI21_X1 _15424_ ( .A(_07353_ ), .B1(_07392_ ), .B2(_07394_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _15425_ ( .A(_06886_ ), .B1(_05116_ ), .B2(_04701_ ), .ZN(_07395_ ) );
OAI21_X1 _15426_ ( .A(_07395_ ), .B1(_04701_ ), .B2(_05116_ ), .ZN(_07396_ ) );
AOI22_X1 _15427_ ( .A1(_05554_ ), .A2(_06995_ ), .B1(\ID_EX_imm [8] ), .B2(_06704_ ), .ZN(_07397_ ) );
AOI21_X1 _15428_ ( .A(_06427_ ), .B1(_07396_ ), .B2(_07397_ ), .ZN(_07398_ ) );
NOR2_X1 _15429_ ( .A1(_07398_ ), .A2(_05184_ ), .ZN(_07399_ ) );
OAI211_X1 _15430_ ( .A(_06481_ ), .B(_06483_ ), .C1(_07052_ ), .C2(_06436_ ), .ZN(_07400_ ) );
NOR2_X1 _15431_ ( .A1(_07008_ ), .A2(_06933_ ), .ZN(_07401_ ) );
NAND3_X1 _15432_ ( .A1(_07177_ ), .A2(_07178_ ), .A3(_06492_ ), .ZN(_07402_ ) );
OAI211_X1 _15433_ ( .A(_04943_ ), .B(_04944_ ), .C1(_06773_ ), .C2(_06778_ ), .ZN(_07403_ ) );
OAI21_X1 _15434_ ( .A(_06487_ ), .B1(_06777_ ), .B2(_06782_ ), .ZN(_07404_ ) );
NAND2_X1 _15435_ ( .A1(_07403_ ), .A2(_07404_ ), .ZN(_07405_ ) );
NAND2_X1 _15436_ ( .A1(_07405_ ), .A2(_06435_ ), .ZN(_07406_ ) );
AOI21_X1 _15437_ ( .A(_06975_ ), .B1(_07402_ ), .B2(_07406_ ), .ZN(_07407_ ) );
OAI21_X1 _15438_ ( .A(_06546_ ), .B1(_07401_ ), .B2(_07407_ ), .ZN(_07408_ ) );
OAI21_X1 _15439_ ( .A(_06755_ ), .B1(_07011_ ), .B2(_06790_ ), .ZN(_07409_ ) );
NAND2_X1 _15440_ ( .A1(_07408_ ), .A2(_07409_ ), .ZN(_07410_ ) );
AOI21_X1 _15441_ ( .A(_07002_ ), .B1(_07400_ ), .B2(_07410_ ), .ZN(_07411_ ) );
NAND3_X1 _15442_ ( .A1(_06563_ ), .A2(_06576_ ), .A3(_04935_ ), .ZN(_07412_ ) );
AND3_X1 _15443_ ( .A1(_07382_ ), .A2(_07074_ ), .A3(_07412_ ), .ZN(_07413_ ) );
NAND3_X1 _15444_ ( .A1(_06447_ ), .A2(_02655_ ), .A3(_06979_ ), .ZN(_07414_ ) );
AOI21_X1 _15445_ ( .A(_06789_ ), .B1(_07017_ ), .B2(_07018_ ), .ZN(_07415_ ) );
AND4_X1 _15446_ ( .A1(_06542_ ), .A2(_06776_ ), .A3(_07249_ ), .A4(_06751_ ), .ZN(_07416_ ) );
OAI21_X1 _15447_ ( .A(_07059_ ), .B1(_07415_ ), .B2(_07416_ ), .ZN(_07417_ ) );
NAND2_X1 _15448_ ( .A1(_04934_ ), .A2(_05166_ ), .ZN(_07418_ ) );
OAI21_X1 _15449_ ( .A(_04827_ ), .B1(_06447_ ), .B2(_02655_ ), .ZN(_07419_ ) );
AND3_X1 _15450_ ( .A1(_07417_ ), .A2(_07418_ ), .A3(_07419_ ), .ZN(_07420_ ) );
OAI211_X1 _15451_ ( .A(_07414_ ), .B(_07420_ ), .C1(_07410_ ), .C2(_07166_ ), .ZN(_07421_ ) );
NOR3_X1 _15452_ ( .A1(_07411_ ), .A2(_07413_ ), .A3(_07421_ ), .ZN(_07422_ ) );
OAI21_X1 _15453_ ( .A(_07399_ ), .B1(_07422_ ), .B2(_06696_ ), .ZN(_07423_ ) );
NAND2_X1 _15454_ ( .A1(_05556_ ), .A2(_05852_ ), .ZN(_07424_ ) );
NAND3_X1 _15455_ ( .A1(_07423_ ), .A2(_06091_ ), .A3(_07424_ ), .ZN(_07425_ ) );
NAND2_X1 _15456_ ( .A1(_05553_ ), .A2(_06094_ ), .ZN(_07426_ ) );
NAND2_X1 _15457_ ( .A1(_07425_ ), .A2(_07426_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
OAI21_X1 _15458_ ( .A(_06156_ ), .B1(_06254_ ), .B2(_06255_ ), .ZN(_07427_ ) );
AND3_X1 _15459_ ( .A1(_05107_ ), .A2(_05108_ ), .A3(_04819_ ), .ZN(_07428_ ) );
NOR2_X1 _15460_ ( .A1(_07428_ ), .A2(_05113_ ), .ZN(_07429_ ) );
OR2_X1 _15461_ ( .A1(_07429_ ), .A2(_04773_ ), .ZN(_07430_ ) );
NAND2_X1 _15462_ ( .A1(_04772_ ), .A2(_02530_ ), .ZN(_07431_ ) );
AND2_X1 _15463_ ( .A1(_07430_ ), .A2(_07431_ ), .ZN(_07432_ ) );
OAI21_X1 _15464_ ( .A(_06421_ ), .B1(_07432_ ), .B2(_04751_ ), .ZN(_07433_ ) );
AOI21_X1 _15465_ ( .A(_07433_ ), .B1(_04751_ ), .B2(_07432_ ), .ZN(_07434_ ) );
AND2_X1 _15466_ ( .A1(_05571_ ), .A2(_06995_ ), .ZN(_07435_ ) );
AND3_X1 _15467_ ( .A1(_06407_ ), .A2(\ID_EX_imm [7] ), .A3(_06997_ ), .ZN(_07436_ ) );
NOR3_X1 _15468_ ( .A1(_07434_ ), .A2(_07435_ ), .A3(_07436_ ), .ZN(_07437_ ) );
OAI21_X1 _15469_ ( .A(_05498_ ), .B1(_07437_ ), .B2(_06428_ ), .ZN(_07438_ ) );
AND3_X1 _15470_ ( .A1(_06481_ ), .A2(_06483_ ), .A3(_06499_ ), .ZN(_07439_ ) );
AND3_X1 _15471_ ( .A1(_07281_ ), .A2(_06493_ ), .A3(_07282_ ), .ZN(_07440_ ) );
OAI211_X1 _15472_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06675_ ), .C2(_06670_ ), .ZN(_07441_ ) );
OAI21_X1 _15473_ ( .A(_06640_ ), .B1(_06669_ ), .B2(_06667_ ), .ZN(_07442_ ) );
AND2_X1 _15474_ ( .A1(_07441_ ), .A2(_07442_ ), .ZN(_07443_ ) );
AOI211_X1 _15475_ ( .A(_06542_ ), .B(_07440_ ), .C1(_06770_ ), .C2(_07443_ ), .ZN(_07444_ ) );
AOI21_X1 _15476_ ( .A(_06820_ ), .B1(_07038_ ), .B2(_07041_ ), .ZN(_07445_ ) );
OR3_X1 _15477_ ( .A1(_07444_ ), .A2(_07445_ ), .A3(_06645_ ), .ZN(_07446_ ) );
MUX2_X1 _15478_ ( .A(_07048_ ), .B(_07045_ ), .S(_06819_ ), .Z(_07447_ ) );
NAND2_X1 _15479_ ( .A1(_07447_ ), .A2(_06755_ ), .ZN(_07448_ ) );
NAND2_X1 _15480_ ( .A1(_07446_ ), .A2(_07448_ ), .ZN(_07449_ ) );
OAI21_X1 _15481_ ( .A(_06432_ ), .B1(_07439_ ), .B2(_07449_ ), .ZN(_07450_ ) );
NAND2_X1 _15482_ ( .A1(_07449_ ), .A2(_06742_ ), .ZN(_07451_ ) );
OR3_X1 _15483_ ( .A1(_07051_ ), .A2(_07052_ ), .A3(_07161_ ), .ZN(_07452_ ) );
AND3_X1 _15484_ ( .A1(_07450_ ), .A2(_07451_ ), .A3(_07452_ ), .ZN(_07453_ ) );
NAND3_X1 _15485_ ( .A1(_06572_ ), .A2(_06574_ ), .A3(_06575_ ), .ZN(_07454_ ) );
NAND2_X1 _15486_ ( .A1(_07454_ ), .A2(_06561_ ), .ZN(_07455_ ) );
NAND2_X1 _15487_ ( .A1(_07455_ ), .A2(_04968_ ), .ZN(_07456_ ) );
XNOR2_X1 _15488_ ( .A(_04971_ ), .B(_02477_ ), .ZN(_07457_ ) );
OR2_X1 _15489_ ( .A1(_04967_ ), .A2(_04988_ ), .ZN(_07458_ ) );
AND3_X1 _15490_ ( .A1(_07456_ ), .A2(_07457_ ), .A3(_07458_ ), .ZN(_07459_ ) );
AOI21_X1 _15491_ ( .A(_07457_ ), .B1(_07456_ ), .B2(_07458_ ), .ZN(_07460_ ) );
OAI21_X1 _15492_ ( .A(_07074_ ), .B1(_07459_ ), .B2(_07460_ ), .ZN(_07461_ ) );
NAND3_X1 _15493_ ( .A1(_04972_ ), .A2(_04973_ ), .A3(_06879_ ), .ZN(_07462_ ) );
NAND3_X1 _15494_ ( .A1(_06442_ ), .A2(_02477_ ), .A3(_06979_ ), .ZN(_07463_ ) );
NAND2_X1 _15495_ ( .A1(_04973_ ), .A2(_07197_ ), .ZN(_07464_ ) );
AND3_X1 _15496_ ( .A1(_07462_ ), .A2(_07463_ ), .A3(_07464_ ), .ZN(_07465_ ) );
NAND3_X1 _15497_ ( .A1(_07453_ ), .A2(_07461_ ), .A3(_07465_ ), .ZN(_07466_ ) );
AOI21_X1 _15498_ ( .A(_07438_ ), .B1(_07466_ ), .B2(_06698_ ), .ZN(_07467_ ) );
NAND2_X1 _15499_ ( .A1(_05573_ ), .A2(_05184_ ), .ZN(_07468_ ) );
NAND2_X1 _15500_ ( .A1(_07468_ ), .A2(_06234_ ), .ZN(_07469_ ) );
OAI21_X1 _15501_ ( .A(_07427_ ), .B1(_07467_ ), .B2(_07469_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
NAND3_X1 _15502_ ( .A1(_05593_ ), .A2(_05595_ ), .A3(_06152_ ), .ZN(_07470_ ) );
NAND2_X1 _15503_ ( .A1(_07429_ ), .A2(_04773_ ), .ZN(_07471_ ) );
NAND3_X1 _15504_ ( .A1(_07430_ ), .A2(_06422_ ), .A3(_07471_ ), .ZN(_07472_ ) );
AOI22_X1 _15505_ ( .A1(_05583_ ), .A2(_06404_ ), .B1(\ID_EX_imm [6] ), .B2(_06408_ ), .ZN(_07473_ ) );
AOI21_X1 _15506_ ( .A(_06426_ ), .B1(_07472_ ), .B2(_07473_ ), .ZN(_07474_ ) );
OR2_X1 _15507_ ( .A1(_07474_ ), .A2(_03778_ ), .ZN(_07475_ ) );
OAI211_X1 _15508_ ( .A(_06709_ ), .B(_07277_ ), .C1(_06710_ ), .C2(_06894_ ), .ZN(_07476_ ) );
MUX2_X1 _15509_ ( .A(_07103_ ), .B(_07108_ ), .S(_06819_ ), .Z(_07477_ ) );
OR2_X1 _15510_ ( .A1(_07477_ ), .A2(_06546_ ), .ZN(_07478_ ) );
OR3_X1 _15511_ ( .A1(_06626_ ), .A2(_06781_ ), .A3(_06785_ ), .ZN(_07479_ ) );
OR3_X1 _15512_ ( .A1(_06777_ ), .A2(_06488_ ), .A3(_06782_ ), .ZN(_07480_ ) );
AOI21_X1 _15513_ ( .A(_06710_ ), .B1(_07479_ ), .B2(_07480_ ), .ZN(_07481_ ) );
AND3_X1 _15514_ ( .A1(_07326_ ), .A2(_06494_ ), .A3(_07327_ ), .ZN(_07482_ ) );
OAI21_X1 _15515_ ( .A(_07054_ ), .B1(_07481_ ), .B2(_07482_ ), .ZN(_07483_ ) );
NAND3_X1 _15516_ ( .A1(_07112_ ), .A2(_06790_ ), .A3(_07113_ ), .ZN(_07484_ ) );
NAND3_X1 _15517_ ( .A1(_07483_ ), .A2(_07484_ ), .A3(_06546_ ), .ZN(_07485_ ) );
NAND2_X1 _15518_ ( .A1(_07478_ ), .A2(_07485_ ), .ZN(_07486_ ) );
AOI21_X1 _15519_ ( .A(_07002_ ), .B1(_07476_ ), .B2(_07486_ ), .ZN(_07487_ ) );
AND3_X1 _15520_ ( .A1(_07478_ ), .A2(_06742_ ), .A3(_07485_ ), .ZN(_07488_ ) );
NOR3_X1 _15521_ ( .A1(_07124_ ), .A2(_07052_ ), .A3(_07161_ ), .ZN(_07489_ ) );
NOR3_X1 _15522_ ( .A1(_07487_ ), .A2(_07488_ ), .A3(_07489_ ), .ZN(_07490_ ) );
AOI21_X1 _15523_ ( .A(_06554_ ), .B1(_07455_ ), .B2(_04968_ ), .ZN(_07491_ ) );
OAI21_X1 _15524_ ( .A(_07491_ ), .B1(_04968_ ), .B2(_07455_ ), .ZN(_07492_ ) );
NAND2_X1 _15525_ ( .A1(_04968_ ), .A2(_06879_ ), .ZN(_07493_ ) );
NAND3_X1 _15526_ ( .A1(_04989_ ), .A2(_02530_ ), .A3(_06979_ ), .ZN(_07494_ ) );
OAI21_X1 _15527_ ( .A(_07197_ ), .B1(_04989_ ), .B2(_02530_ ), .ZN(_07495_ ) );
AND3_X1 _15528_ ( .A1(_07493_ ), .A2(_07494_ ), .A3(_07495_ ), .ZN(_07496_ ) );
NAND3_X1 _15529_ ( .A1(_07490_ ), .A2(_07492_ ), .A3(_07496_ ), .ZN(_07497_ ) );
BUF_X4 _15530_ ( .A(_06697_ ), .Z(_07498_ ) );
AOI21_X1 _15531_ ( .A(_07475_ ), .B1(_07497_ ), .B2(_07498_ ), .ZN(_07499_ ) );
OAI21_X1 _15532_ ( .A(_07207_ ), .B1(_05582_ ), .B2(_05543_ ), .ZN(_07500_ ) );
OAI21_X1 _15533_ ( .A(_07470_ ), .B1(_07499_ ), .B2(_07500_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
NAND3_X1 _15534_ ( .A1(_05614_ ), .A2(_05616_ ), .A3(_06152_ ), .ZN(_07501_ ) );
NAND3_X1 _15535_ ( .A1(_06407_ ), .A2(\ID_EX_imm [5] ), .A3(_06997_ ), .ZN(_07502_ ) );
OAI21_X1 _15536_ ( .A(_07502_ ), .B1(_05606_ ), .B2(_06406_ ), .ZN(_07503_ ) );
AND3_X1 _15537_ ( .A1(_05107_ ), .A2(_04818_ ), .A3(_05108_ ), .ZN(_07504_ ) );
AOI21_X1 _15538_ ( .A(_02533_ ), .B1(_04797_ ), .B2(_04816_ ), .ZN(_07505_ ) );
OAI21_X1 _15539_ ( .A(_04796_ ), .B1(_07504_ ), .B2(_07505_ ), .ZN(_07506_ ) );
AND2_X1 _15540_ ( .A1(_07506_ ), .A2(_06421_ ), .ZN(_07507_ ) );
OR3_X1 _15541_ ( .A1(_07504_ ), .A2(_07505_ ), .A3(_04796_ ), .ZN(_07508_ ) );
AOI21_X1 _15542_ ( .A(_07503_ ), .B1(_07507_ ), .B2(_07508_ ), .ZN(_07509_ ) );
OAI21_X1 _15543_ ( .A(_05498_ ), .B1(_07509_ ), .B2(_06428_ ), .ZN(_07510_ ) );
AND4_X1 _15544_ ( .A1(_06483_ ), .A2(_06481_ ), .A3(_06496_ ), .A4(_06498_ ), .ZN(_07511_ ) );
NAND2_X1 _15545_ ( .A1(_06543_ ), .A2(_06832_ ), .ZN(_07512_ ) );
NAND3_X1 _15546_ ( .A1(_07365_ ), .A2(_07366_ ), .A3(_06673_ ), .ZN(_07513_ ) );
OAI211_X1 _15547_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06669_ ), .C2(_06667_ ), .ZN(_07514_ ) );
OAI21_X1 _15548_ ( .A(_07249_ ), .B1(_06666_ ), .B2(_06630_ ), .ZN(_07515_ ) );
NAND2_X1 _15549_ ( .A1(_07514_ ), .A2(_07515_ ), .ZN(_07516_ ) );
OAI211_X1 _15550_ ( .A(_07513_ ), .B(_06820_ ), .C1(_07516_ ), .C2(_06494_ ), .ZN(_07517_ ) );
OAI211_X1 _15551_ ( .A(_06619_ ), .B(_07517_ ), .C1(_07150_ ), .C2(_06844_ ), .ZN(_07518_ ) );
NAND2_X1 _15552_ ( .A1(_07512_ ), .A2(_07518_ ), .ZN(_07519_ ) );
OAI21_X1 _15553_ ( .A(_06431_ ), .B1(_07511_ ), .B2(_07519_ ), .ZN(_07520_ ) );
NAND2_X1 _15554_ ( .A1(_07519_ ), .A2(_06742_ ), .ZN(_07521_ ) );
OAI211_X1 _15555_ ( .A(_07520_ ), .B(_07521_ ), .C1(_06644_ ), .C2(_07161_ ), .ZN(_07522_ ) );
NAND2_X1 _15556_ ( .A1(_06572_ ), .A2(_06574_ ), .ZN(_07523_ ) );
NOR2_X1 _15557_ ( .A1(_07523_ ), .A2(_04986_ ), .ZN(_07524_ ) );
INV_X1 _15558_ ( .A(_07524_ ), .ZN(_07525_ ) );
INV_X1 _15559_ ( .A(_06560_ ), .ZN(_07526_ ) );
NAND3_X1 _15560_ ( .A1(_07525_ ), .A2(_04980_ ), .A3(_07526_ ), .ZN(_07527_ ) );
OAI21_X1 _15561_ ( .A(_04979_ ), .B1(_07524_ ), .B2(_06560_ ), .ZN(_07528_ ) );
AND3_X1 _15562_ ( .A1(_07527_ ), .A2(_07074_ ), .A3(_07528_ ), .ZN(_07529_ ) );
NAND2_X1 _15563_ ( .A1(_04979_ ), .A2(_06879_ ), .ZN(_07530_ ) );
NAND3_X1 _15564_ ( .A1(_04977_ ), .A2(_02525_ ), .A3(_06979_ ), .ZN(_07531_ ) );
OAI21_X1 _15565_ ( .A(_07197_ ), .B1(_04977_ ), .B2(_02525_ ), .ZN(_07532_ ) );
NAND3_X1 _15566_ ( .A1(_07530_ ), .A2(_07531_ ), .A3(_07532_ ), .ZN(_07533_ ) );
OR3_X1 _15567_ ( .A1(_07522_ ), .A2(_07529_ ), .A3(_07533_ ), .ZN(_07534_ ) );
AOI21_X1 _15568_ ( .A(_07510_ ), .B1(_07534_ ), .B2(_07498_ ), .ZN(_07535_ ) );
OAI21_X1 _15569_ ( .A(_07207_ ), .B1(_05603_ ), .B2(_05543_ ), .ZN(_07536_ ) );
OAI21_X1 _15570_ ( .A(_07501_ ), .B1(_07535_ ), .B2(_07536_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
NAND3_X1 _15571_ ( .A1(_05636_ ), .A2(_05638_ ), .A3(_06152_ ), .ZN(_07537_ ) );
OAI211_X1 _15572_ ( .A(_06709_ ), .B(_07277_ ), .C1(_06710_ ), .C2(_06434_ ), .ZN(_07538_ ) );
NAND2_X1 _15573_ ( .A1(_06734_ ), .A2(_06832_ ), .ZN(_07539_ ) );
AND3_X1 _15574_ ( .A1(_07403_ ), .A2(_06502_ ), .A3(_07404_ ), .ZN(_07540_ ) );
NOR3_X1 _15575_ ( .A1(_06624_ ), .A2(_06784_ ), .A3(_06748_ ), .ZN(_07541_ ) );
NOR3_X1 _15576_ ( .A1(_06781_ ), .A2(_06487_ ), .A3(_06785_ ), .ZN(_07542_ ) );
NOR2_X1 _15577_ ( .A1(_07541_ ), .A2(_07542_ ), .ZN(_07543_ ) );
INV_X1 _15578_ ( .A(_07543_ ), .ZN(_07544_ ) );
AOI211_X1 _15579_ ( .A(_06541_ ), .B(_07540_ ), .C1(_07544_ ), .C2(_06647_ ), .ZN(_07545_ ) );
AOI21_X1 _15580_ ( .A(_06819_ ), .B1(_07179_ ), .B2(_07180_ ), .ZN(_07546_ ) );
OR3_X1 _15581_ ( .A1(_07545_ ), .A2(_06645_ ), .A3(_07546_ ), .ZN(_07547_ ) );
AND2_X1 _15582_ ( .A1(_07539_ ), .A2(_07547_ ), .ZN(_07548_ ) );
AOI21_X1 _15583_ ( .A(_07002_ ), .B1(_07538_ ), .B2(_07548_ ), .ZN(_07549_ ) );
OR2_X1 _15584_ ( .A1(_07548_ ), .A2(_07166_ ), .ZN(_07550_ ) );
AOI21_X1 _15585_ ( .A(_06553_ ), .B1(_07523_ ), .B2(_04986_ ), .ZN(_07551_ ) );
OAI21_X1 _15586_ ( .A(_07551_ ), .B1(_04986_ ), .B2(_07523_ ), .ZN(_07552_ ) );
OAI21_X1 _15587_ ( .A(_07197_ ), .B1(_06755_ ), .B2(_02452_ ), .ZN(_07553_ ) );
AND2_X1 _15588_ ( .A1(_06753_ ), .A2(_07058_ ), .ZN(_07554_ ) );
AOI221_X4 _15589_ ( .A(_07554_ ), .B1(_06560_ ), .B2(_06686_ ), .C1(_04985_ ), .C2(_05166_ ), .ZN(_07555_ ) );
NAND4_X1 _15590_ ( .A1(_07550_ ), .A2(_07552_ ), .A3(_07553_ ), .A4(_07555_ ), .ZN(_07556_ ) );
OAI21_X1 _15591_ ( .A(_06697_ ), .B1(_07549_ ), .B2(_07556_ ), .ZN(_07557_ ) );
AOI21_X1 _15592_ ( .A(_04818_ ), .B1(_05107_ ), .B2(_05108_ ), .ZN(_07558_ ) );
NOR3_X1 _15593_ ( .A1(_07504_ ), .A2(_07558_ ), .A3(_06886_ ), .ZN(_07559_ ) );
OAI22_X1 _15594_ ( .A1(_05629_ ), .A2(_06406_ ), .B1(_02453_ ), .B2(_06410_ ), .ZN(_07560_ ) );
OAI21_X1 _15595_ ( .A(_06425_ ), .B1(_07559_ ), .B2(_07560_ ), .ZN(_07561_ ) );
AND3_X1 _15596_ ( .A1(_07557_ ), .A2(_05245_ ), .A3(_07561_ ), .ZN(_07562_ ) );
OAI21_X1 _15597_ ( .A(_07207_ ), .B1(_05182_ ), .B2(_05625_ ), .ZN(_07563_ ) );
OAI21_X1 _15598_ ( .A(_07537_ ), .B1(_07562_ ), .B2(_07563_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _15599_ ( .A1(_05656_ ), .A2(_06094_ ), .ZN(_07564_ ) );
AND2_X1 _15600_ ( .A1(_05104_ ), .A2(_05106_ ), .ZN(_07565_ ) );
XNOR2_X1 _15601_ ( .A(_07565_ ), .B(_04534_ ), .ZN(_07566_ ) );
NAND2_X1 _15602_ ( .A1(_07566_ ), .A2(_06422_ ), .ZN(_07567_ ) );
AOI22_X1 _15603_ ( .A1(_05646_ ), .A2(_06404_ ), .B1(\ID_EX_imm [3] ), .B2(_06408_ ), .ZN(_07568_ ) );
AOI21_X1 _15604_ ( .A(_06426_ ), .B1(_07567_ ), .B2(_07568_ ), .ZN(_07569_ ) );
OR2_X1 _15605_ ( .A1(_07569_ ), .A2(_03778_ ), .ZN(_07570_ ) );
AND2_X1 _15606_ ( .A1(_07439_ ), .A2(_06863_ ), .ZN(_07571_ ) );
NAND2_X1 _15607_ ( .A1(_06860_ ), .A2(_06755_ ), .ZN(_07572_ ) );
NAND3_X1 _15608_ ( .A1(_07280_ ), .A2(_07052_ ), .A3(_07283_ ), .ZN(_07573_ ) );
NOR2_X1 _15609_ ( .A1(_06666_ ), .A2(_06630_ ), .ZN(_07574_ ) );
NOR2_X1 _15610_ ( .A1(_06631_ ), .A2(_06635_ ), .ZN(_07575_ ) );
MUX2_X1 _15611_ ( .A(_07574_ ), .B(_07575_ ), .S(_07249_ ), .Z(_07576_ ) );
MUX2_X1 _15612_ ( .A(_07443_ ), .B(_07576_ ), .S(_07377_ ), .Z(_07577_ ) );
OAI211_X1 _15613_ ( .A(_07258_ ), .B(_07573_ ), .C1(_07577_ ), .C2(_07052_ ), .ZN(_07578_ ) );
NAND2_X1 _15614_ ( .A1(_07572_ ), .A2(_07578_ ), .ZN(_07579_ ) );
OAI21_X1 _15615_ ( .A(_06432_ ), .B1(_07571_ ), .B2(_07579_ ), .ZN(_07580_ ) );
NAND2_X1 _15616_ ( .A1(_07579_ ), .A2(_06742_ ), .ZN(_07581_ ) );
AND3_X1 _15617_ ( .A1(_06818_ ), .A2(_06820_ ), .A3(_07058_ ), .ZN(_07582_ ) );
AOI221_X4 _15618_ ( .A(_07582_ ), .B1(_06570_ ), .B2(_06686_ ), .C1(_06574_ ), .C2(_04827_ ), .ZN(_07583_ ) );
NOR3_X1 _15619_ ( .A1(_06569_ ), .A2(_06571_ ), .A3(_06553_ ), .ZN(_07584_ ) );
OAI21_X1 _15620_ ( .A(_04941_ ), .B1(_07584_ ), .B2(_06879_ ), .ZN(_07585_ ) );
OAI211_X1 _15621_ ( .A(_04942_ ), .B(_07074_ ), .C1(_06569_ ), .C2(_06571_ ), .ZN(_07586_ ) );
AND3_X1 _15622_ ( .A1(_07583_ ), .A2(_07585_ ), .A3(_07586_ ), .ZN(_07587_ ) );
NAND3_X1 _15623_ ( .A1(_07580_ ), .A2(_07581_ ), .A3(_07587_ ), .ZN(_07588_ ) );
AOI21_X1 _15624_ ( .A(_07570_ ), .B1(_07588_ ), .B2(_07498_ ), .ZN(_07589_ ) );
OAI21_X1 _15625_ ( .A(_07207_ ), .B1(_05182_ ), .B2(_05643_ ), .ZN(_07590_ ) );
OAI21_X1 _15626_ ( .A(_07564_ ), .B1(_07589_ ), .B2(_07590_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
AOI21_X1 _15627_ ( .A(_06886_ ), .B1(_05103_ ), .B2(_04512_ ), .ZN(_07591_ ) );
OAI21_X1 _15628_ ( .A(_07591_ ), .B1(_04512_ ), .B2(_05103_ ), .ZN(_07592_ ) );
AOI22_X1 _15629_ ( .A1(_05662_ ), .A2(_06995_ ), .B1(\ID_EX_imm [2] ), .B2(_06704_ ), .ZN(_07593_ ) );
AOI21_X1 _15630_ ( .A(_06427_ ), .B1(_07592_ ), .B2(_07593_ ), .ZN(_07594_ ) );
NOR2_X1 _15631_ ( .A1(_07594_ ), .A2(_05184_ ), .ZN(_07595_ ) );
NAND2_X1 _15632_ ( .A1(_06910_ ), .A2(_06832_ ), .ZN(_07596_ ) );
OR3_X1 _15633_ ( .A1(_07325_ ), .A2(_06819_ ), .A3(_07328_ ), .ZN(_07597_ ) );
NOR3_X1 _15634_ ( .A1(_06784_ ), .A2(_06634_ ), .A3(_06748_ ), .ZN(_07598_ ) );
NOR2_X1 _15635_ ( .A1(_06747_ ), .A2(_06745_ ), .ZN(_07599_ ) );
AOI21_X1 _15636_ ( .A(_07598_ ), .B1(_06640_ ), .B2(_07599_ ), .ZN(_07600_ ) );
AND2_X1 _15637_ ( .A1(_07479_ ), .A2(_07480_ ), .ZN(_07601_ ) );
MUX2_X1 _15638_ ( .A(_07600_ ), .B(_07601_ ), .S(_06493_ ), .Z(_07602_ ) );
OAI211_X1 _15639_ ( .A(_06545_ ), .B(_07597_ ), .C1(_07602_ ), .C2(_06789_ ), .ZN(_07603_ ) );
AND3_X1 _15640_ ( .A1(_07596_ ), .A2(_06741_ ), .A3(_07603_ ), .ZN(_07604_ ) );
NAND4_X1 _15641_ ( .A1(_06862_ ), .A2(_06894_ ), .A3(_06499_ ), .A4(_06863_ ), .ZN(_07605_ ) );
NAND2_X1 _15642_ ( .A1(_07596_ ), .A2(_07603_ ), .ZN(_07606_ ) );
AOI21_X1 _15643_ ( .A(_07002_ ), .B1(_07605_ ), .B2(_07606_ ), .ZN(_07607_ ) );
AOI211_X1 _15644_ ( .A(_07604_ ), .B(_07607_ ), .C1(_06917_ ), .C2(_07059_ ), .ZN(_07608_ ) );
NAND3_X1 _15645_ ( .A1(_06567_ ), .A2(_06568_ ), .A3(_04959_ ), .ZN(_07609_ ) );
NAND2_X1 _15646_ ( .A1(_07609_ ), .A2(_06552_ ), .ZN(_07610_ ) );
OR2_X1 _15647_ ( .A1(_07610_ ), .A2(_06569_ ), .ZN(_07611_ ) );
AOI21_X1 _15648_ ( .A(_04828_ ), .B1(_07377_ ), .B2(_04511_ ), .ZN(_07612_ ) );
AOI221_X4 _15649_ ( .A(_07612_ ), .B1(_06571_ ), .B2(_06686_ ), .C1(_04958_ ), .C2(_06687_ ), .ZN(_07613_ ) );
AND3_X1 _15650_ ( .A1(_07608_ ), .A2(_07611_ ), .A3(_07613_ ), .ZN(_07614_ ) );
OAI21_X1 _15651_ ( .A(_07595_ ), .B1(_07614_ ), .B2(_06696_ ), .ZN(_07615_ ) );
NAND3_X1 _15652_ ( .A1(_06424_ ), .A2(\ID_EX_typ [7] ), .A3(_05664_ ), .ZN(_07616_ ) );
NAND3_X1 _15653_ ( .A1(_07615_ ), .A2(_06164_ ), .A3(_07616_ ), .ZN(_07617_ ) );
NAND2_X1 _15654_ ( .A1(_05673_ ), .A2(_06094_ ), .ZN(_07618_ ) );
NAND2_X1 _15655_ ( .A1(_07617_ ), .A2(_07618_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
NAND3_X1 _15656_ ( .A1(_05237_ ), .A2(_05241_ ), .A3(_06152_ ), .ZN(_07619_ ) );
OAI22_X1 _15657_ ( .A1(_05205_ ), .A2(_06405_ ), .B1(_02895_ ), .B2(_06410_ ), .ZN(_07620_ ) );
AOI21_X1 _15658_ ( .A(_05153_ ), .B1(_07269_ ), .B2(_04269_ ), .ZN(_07621_ ) );
XNOR2_X1 _15659_ ( .A(_07621_ ), .B(_04291_ ), .ZN(_07622_ ) );
AOI21_X1 _15660_ ( .A(_07620_ ), .B1(_06422_ ), .B2(_07622_ ), .ZN(_07623_ ) );
OAI21_X1 _15661_ ( .A(_05498_ ), .B1(_07623_ ), .B2(_06428_ ), .ZN(_07624_ ) );
INV_X1 _15662_ ( .A(_04855_ ), .ZN(_07625_ ) );
INV_X1 _15663_ ( .A(_07225_ ), .ZN(_07626_ ) );
AOI21_X1 _15664_ ( .A(_07625_ ), .B1(_07626_ ), .B2(_07227_ ), .ZN(_07627_ ) );
OR3_X1 _15665_ ( .A1(_07627_ ), .A2(_04850_ ), .A3(_07231_ ), .ZN(_07628_ ) );
OAI21_X1 _15666_ ( .A(_04850_ ), .B1(_07627_ ), .B2(_07231_ ), .ZN(_07629_ ) );
NAND3_X1 _15667_ ( .A1(_07628_ ), .A2(_07074_ ), .A3(_07629_ ), .ZN(_07630_ ) );
OAI211_X1 _15668_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06514_ ), .C2(_06510_ ), .ZN(_07631_ ) );
OAI21_X1 _15669_ ( .A(_07249_ ), .B1(_06509_ ), .B2(_06530_ ), .ZN(_07632_ ) );
NAND3_X1 _15670_ ( .A1(_07631_ ), .A2(_06710_ ), .A3(_07632_ ), .ZN(_07633_ ) );
OAI211_X1 _15671_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06529_ ), .C2(_06527_ ), .ZN(_07634_ ) );
NOR2_X1 _15672_ ( .A1(_06523_ ), .A2(_06537_ ), .ZN(_07635_ ) );
OAI21_X1 _15673_ ( .A(_07634_ ), .B1(_07635_ ), .B2(_06627_ ), .ZN(_07636_ ) );
OAI21_X1 _15674_ ( .A(_07633_ ), .B1(_07636_ ), .B2(_06710_ ), .ZN(_07637_ ) );
NAND2_X1 _15675_ ( .A1(_07637_ ), .A2(_07054_ ), .ZN(_07638_ ) );
OAI21_X1 _15676_ ( .A(_07052_ ), .B1(_06656_ ), .B2(_06662_ ), .ZN(_07639_ ) );
AOI21_X1 _15677_ ( .A(_06755_ ), .B1(_07638_ ), .B2(_07639_ ), .ZN(_07640_ ) );
AOI21_X1 _15678_ ( .A(_06547_ ), .B1(_07162_ ), .B2(_07163_ ), .ZN(_07641_ ) );
OAI21_X1 _15679_ ( .A(_05163_ ), .B1(_07640_ ), .B2(_07641_ ), .ZN(_07642_ ) );
NAND2_X1 _15680_ ( .A1(_04850_ ), .A2(_06687_ ), .ZN(_07643_ ) );
NOR3_X1 _15681_ ( .A1(_06539_ ), .A2(_06790_ ), .A3(_06710_ ), .ZN(_07644_ ) );
NAND2_X1 _15682_ ( .A1(_07644_ ), .A2(_06546_ ), .ZN(_07645_ ) );
OAI221_X1 _15683_ ( .A(_07643_ ), .B1(_05077_ ), .B2(_06797_ ), .C1(_07645_ ), .C2(_07166_ ), .ZN(_07646_ ) );
NAND3_X1 _15684_ ( .A1(_06497_ ), .A2(_06619_ ), .A3(_06495_ ), .ZN(_07647_ ) );
NAND4_X1 _15685_ ( .A1(_06467_ ), .A2(_06478_ ), .A3(_06480_ ), .A4(_07647_ ), .ZN(_07648_ ) );
AOI21_X1 _15686_ ( .A(_07002_ ), .B1(_07648_ ), .B2(_07645_ ), .ZN(_07649_ ) );
AOI211_X1 _15687_ ( .A(_07646_ ), .B(_07649_ ), .C1(_05076_ ), .C2(_06979_ ), .ZN(_07650_ ) );
NAND3_X1 _15688_ ( .A1(_07630_ ), .A2(_07642_ ), .A3(_07650_ ), .ZN(_07651_ ) );
AOI21_X1 _15689_ ( .A(_07624_ ), .B1(_07651_ ), .B2(_07498_ ), .ZN(_07652_ ) );
OAI21_X1 _15690_ ( .A(_07207_ ), .B1(_05199_ ), .B2(_07091_ ), .ZN(_07653_ ) );
OAI21_X1 _15691_ ( .A(_07619_ ), .B1(_07652_ ), .B2(_07653_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
NAND2_X1 _15692_ ( .A1(_05688_ ), .A2(_06094_ ), .ZN(_07654_ ) );
OAI21_X1 _15693_ ( .A(_06421_ ), .B1(_04462_ ), .B2(_05102_ ), .ZN(_07655_ ) );
AOI21_X1 _15694_ ( .A(_07655_ ), .B1(_04462_ ), .B2(_05102_ ), .ZN(_07656_ ) );
AND2_X1 _15695_ ( .A1(_05678_ ), .A2(_06404_ ), .ZN(_07657_ ) );
AND3_X1 _15696_ ( .A1(_06407_ ), .A2(\ID_EX_imm [1] ), .A3(_06997_ ), .ZN(_07658_ ) );
NOR3_X1 _15697_ ( .A1(_07656_ ), .A2(_07657_ ), .A3(_07658_ ), .ZN(_07659_ ) );
OAI21_X1 _15698_ ( .A(_05498_ ), .B1(_07659_ ), .B2(_06428_ ), .ZN(_07660_ ) );
AND3_X1 _15699_ ( .A1(_06952_ ), .A2(_06491_ ), .A3(_07277_ ), .ZN(_07661_ ) );
OR2_X1 _15700_ ( .A1(_06964_ ), .A2(_06546_ ), .ZN(_07662_ ) );
OAI21_X1 _15701_ ( .A(_07249_ ), .B1(_06633_ ), .B2(_06638_ ), .ZN(_07663_ ) );
OAI211_X1 _15702_ ( .A(_07663_ ), .B(_07377_ ), .C1(_07575_ ), .C2(_07249_ ), .ZN(_07664_ ) );
OAI211_X1 _15703_ ( .A(_07664_ ), .B(_06933_ ), .C1(_07377_ ), .C2(_07516_ ), .ZN(_07665_ ) );
OAI211_X1 _15704_ ( .A(_07258_ ), .B(_07665_ ), .C1(_07368_ ), .C2(_07054_ ), .ZN(_07666_ ) );
NAND2_X1 _15705_ ( .A1(_07662_ ), .A2(_07666_ ), .ZN(_07667_ ) );
OAI21_X1 _15706_ ( .A(_06432_ ), .B1(_07661_ ), .B2(_07667_ ), .ZN(_07668_ ) );
OAI21_X1 _15707_ ( .A(_07074_ ), .B1(_04949_ ), .B2(_06564_ ), .ZN(_07669_ ) );
OR2_X1 _15708_ ( .A1(_07669_ ), .A2(_06566_ ), .ZN(_07670_ ) );
AOI21_X1 _15709_ ( .A(_07166_ ), .B1(_07662_ ), .B2(_07666_ ), .ZN(_07671_ ) );
AND3_X1 _15710_ ( .A1(_06967_ ), .A2(_07054_ ), .A3(_07059_ ), .ZN(_07672_ ) );
NOR3_X1 _15711_ ( .A1(_04947_ ), .A2(_04948_ ), .A3(_05167_ ), .ZN(_07673_ ) );
OAI22_X1 _15712_ ( .A1(_06568_ ), .A2(_06795_ ), .B1(_04948_ ), .B2(_06797_ ), .ZN(_07674_ ) );
NOR4_X1 _15713_ ( .A1(_07671_ ), .A2(_07672_ ), .A3(_07673_ ), .A4(_07674_ ), .ZN(_07675_ ) );
NAND3_X1 _15714_ ( .A1(_07668_ ), .A2(_07670_ ), .A3(_07675_ ), .ZN(_07676_ ) );
AOI21_X1 _15715_ ( .A(_07660_ ), .B1(_07676_ ), .B2(_07498_ ), .ZN(_07677_ ) );
OAI21_X1 _15716_ ( .A(_07207_ ), .B1(_05182_ ), .B2(\ID_EX_pc [1] ), .ZN(_07678_ ) );
OAI21_X1 _15717_ ( .A(_07654_ ), .B1(_07677_ ), .B2(_07678_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
AND3_X1 _15718_ ( .A1(_05071_ ), .A2(_05083_ ), .A3(_06693_ ), .ZN(_07679_ ) );
NAND2_X1 _15719_ ( .A1(_04487_ ), .A2(_06421_ ), .ZN(_07680_ ) );
NAND3_X1 _15720_ ( .A1(_05725_ ), .A2(_06997_ ), .A3(_06401_ ), .ZN(_07681_ ) );
NAND3_X1 _15721_ ( .A1(_06407_ ), .A2(\ID_EX_imm [0] ), .A3(_06997_ ), .ZN(_07682_ ) );
NAND3_X1 _15722_ ( .A1(_07680_ ), .A2(_07681_ ), .A3(_07682_ ), .ZN(_07683_ ) );
OAI21_X1 _15723_ ( .A(_06425_ ), .B1(_07679_ ), .B2(_07683_ ), .ZN(_07684_ ) );
NAND4_X1 _15724_ ( .A1(_06708_ ), .A2(_04977_ ), .A3(_06430_ ), .A4(_06439_ ), .ZN(_07685_ ) );
OR3_X1 _15725_ ( .A1(_05074_ ), .A2(_05081_ ), .A3(_04830_ ), .ZN(_07686_ ) );
AOI21_X1 _15726_ ( .A(_07686_ ), .B1(_05082_ ), .B2(_05079_ ), .ZN(_07687_ ) );
NAND2_X1 _15727_ ( .A1(_05071_ ), .A2(_07687_ ), .ZN(_07688_ ) );
AOI21_X1 _15728_ ( .A(_06744_ ), .B1(_04950_ ), .B2(_06433_ ), .ZN(_07689_ ) );
MUX2_X1 _15729_ ( .A(_07599_ ), .B(_07689_ ), .S(_06487_ ), .Z(_07690_ ) );
MUX2_X1 _15730_ ( .A(_07544_ ), .B(_07690_ ), .S(_06435_ ), .Z(_07691_ ) );
AND2_X1 _15731_ ( .A1(_07691_ ), .A2(_06437_ ), .ZN(_07692_ ) );
AND3_X1 _15732_ ( .A1(_07402_ ), .A2(_04939_ ), .A3(_07406_ ), .ZN(_07693_ ) );
OR3_X1 _15733_ ( .A1(_07692_ ), .A2(_06645_ ), .A3(_07693_ ), .ZN(_07694_ ) );
OAI211_X1 _15734_ ( .A(_07694_ ), .B(_07037_ ), .C1(_06544_ ), .C2(_07012_ ), .ZN(_07695_ ) );
NAND3_X1 _15735_ ( .A1(_07025_ ), .A2(_06820_ ), .A3(_07058_ ), .ZN(_07696_ ) );
NAND3_X1 _15736_ ( .A1(_06892_ ), .A2(_04486_ ), .A3(_06686_ ), .ZN(_07697_ ) );
AOI22_X1 _15737_ ( .A1(_06892_ ), .A2(_04486_ ), .B1(_05167_ ), .B2(_06553_ ), .ZN(_07698_ ) );
OAI22_X1 _15738_ ( .A1(_07698_ ), .A2(_04827_ ), .B1(_04486_ ), .B2(_06892_ ), .ZN(_07699_ ) );
AND4_X1 _15739_ ( .A1(_07695_ ), .A2(_07696_ ), .A3(_07697_ ), .A4(_07699_ ), .ZN(_07700_ ) );
AND3_X1 _15740_ ( .A1(_07685_ ), .A2(_07688_ ), .A3(_07700_ ), .ZN(_07701_ ) );
OAI21_X1 _15741_ ( .A(_07684_ ), .B1(_07701_ ), .B2(_06695_ ), .ZN(_07702_ ) );
MUX2_X1 _15742_ ( .A(\ID_EX_pc [0] ), .B(_07702_ ), .S(_05180_ ), .Z(_07703_ ) );
MUX2_X1 _15743_ ( .A(_05724_ ), .B(_07703_ ), .S(_06099_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
NAND3_X1 _15744_ ( .A1(_06344_ ), .A2(_06345_ ), .A3(_06152_ ), .ZN(_07704_ ) );
OR2_X1 _15745_ ( .A1(_07269_ ), .A2(_04269_ ), .ZN(_07705_ ) );
AOI21_X1 _15746_ ( .A(_06886_ ), .B1(_07269_ ), .B2(_04269_ ), .ZN(_07706_ ) );
AND2_X1 _15747_ ( .A1(_07705_ ), .A2(_07706_ ), .ZN(_07707_ ) );
NOR2_X1 _15748_ ( .A1(_05483_ ), .A2(_06406_ ), .ZN(_07708_ ) );
AND3_X1 _15749_ ( .A1(_06407_ ), .A2(\ID_EX_imm [28] ), .A3(_06997_ ), .ZN(_07709_ ) );
NOR3_X1 _15750_ ( .A1(_07707_ ), .A2(_07708_ ), .A3(_07709_ ), .ZN(_07710_ ) );
OAI21_X1 _15751_ ( .A(_05498_ ), .B1(_07710_ ), .B2(_06427_ ), .ZN(_07711_ ) );
NOR3_X1 _15752_ ( .A1(_07225_ ), .A2(_04855_ ), .A3(_07228_ ), .ZN(_07712_ ) );
OR3_X1 _15753_ ( .A1(_07627_ ), .A2(_06554_ ), .A3(_07712_ ), .ZN(_07713_ ) );
NAND2_X1 _15754_ ( .A1(_04855_ ), .A2(_06879_ ), .ZN(_07714_ ) );
NAND3_X1 _15755_ ( .A1(_04853_ ), .A2(_02125_ ), .A3(_06979_ ), .ZN(_07715_ ) );
OAI21_X1 _15756_ ( .A(_07197_ ), .B1(_04853_ ), .B2(_02125_ ), .ZN(_07716_ ) );
AND3_X1 _15757_ ( .A1(_07714_ ), .A2(_07715_ ), .A3(_07716_ ), .ZN(_07717_ ) );
AND3_X1 _15758_ ( .A1(_06732_ ), .A2(_06844_ ), .A3(_07377_ ), .ZN(_07718_ ) );
NAND2_X1 _15759_ ( .A1(_07718_ ), .A2(_06546_ ), .ZN(_07719_ ) );
OR2_X1 _15760_ ( .A1(_07237_ ), .A2(_07185_ ), .ZN(_07720_ ) );
OAI211_X1 _15761_ ( .A(_07719_ ), .B(_07720_ ), .C1(_06482_ ), .C2(_06486_ ), .ZN(_07721_ ) );
NAND2_X1 _15762_ ( .A1(_07721_ ), .A2(_06432_ ), .ZN(_07722_ ) );
OAI211_X1 _15763_ ( .A(_06627_ ), .B(_06713_ ), .C1(_02815_ ), .C2(_06490_ ), .ZN(_07723_ ) );
OAI211_X1 _15764_ ( .A(_07723_ ), .B(_06770_ ), .C1(_06627_ ), .C2(_07248_ ), .ZN(_07724_ ) );
NOR2_X1 _15765_ ( .A1(_06723_ ), .A2(_06721_ ), .ZN(_07725_ ) );
MUX2_X1 _15766_ ( .A(_07725_ ), .B(_07251_ ), .S(_07249_ ), .Z(_07726_ ) );
OAI211_X1 _15767_ ( .A(_07724_ ), .B(_06844_ ), .C1(_07726_ ), .C2(_07377_ ), .ZN(_07727_ ) );
NAND3_X1 _15768_ ( .A1(_06763_ ), .A2(_06975_ ), .A3(_06771_ ), .ZN(_07728_ ) );
NAND3_X1 _15769_ ( .A1(_07727_ ), .A2(_06619_ ), .A3(_07728_ ), .ZN(_07729_ ) );
AND2_X1 _15770_ ( .A1(_07729_ ), .A2(_05163_ ), .ZN(_07730_ ) );
OAI21_X1 _15771_ ( .A(_07730_ ), .B1(_07191_ ), .B2(_06547_ ), .ZN(_07731_ ) );
NAND3_X1 _15772_ ( .A1(_07718_ ), .A2(_06547_ ), .A3(_06742_ ), .ZN(_07732_ ) );
AND3_X1 _15773_ ( .A1(_07722_ ), .A2(_07731_ ), .A3(_07732_ ), .ZN(_07733_ ) );
NAND3_X1 _15774_ ( .A1(_07713_ ), .A2(_07717_ ), .A3(_07733_ ), .ZN(_07734_ ) );
AOI21_X1 _15775_ ( .A(_07711_ ), .B1(_07734_ ), .B2(_07498_ ), .ZN(_07735_ ) );
OAI21_X1 _15776_ ( .A(_07207_ ), .B1(_05481_ ), .B2(_07091_ ), .ZN(_07736_ ) );
OAI21_X1 _15777_ ( .A(_07704_ ), .B1(_07735_ ), .B2(_07736_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND3_X1 _15778_ ( .A1(_06351_ ), .A2(_06352_ ), .A3(_06152_ ), .ZN(_07737_ ) );
NAND2_X1 _15779_ ( .A1(_07267_ ), .A2(_04434_ ), .ZN(_07738_ ) );
NAND2_X1 _15780_ ( .A1(_07738_ ), .A2(_05148_ ), .ZN(_07739_ ) );
AND2_X1 _15781_ ( .A1(_07739_ ), .A2(_04387_ ), .ZN(_07740_ ) );
OR3_X1 _15782_ ( .A1(_07740_ ), .A2(_04365_ ), .A3(_05143_ ), .ZN(_07741_ ) );
OAI21_X1 _15783_ ( .A(_04365_ ), .B1(_07740_ ), .B2(_05143_ ), .ZN(_07742_ ) );
AND3_X1 _15784_ ( .A1(_07741_ ), .A2(_06421_ ), .A3(_07742_ ), .ZN(_07743_ ) );
OAI22_X1 _15785_ ( .A1(_05709_ ), .A2(_06406_ ), .B1(_02819_ ), .B2(_06410_ ), .ZN(_07744_ ) );
OAI21_X1 _15786_ ( .A(_06425_ ), .B1(_07743_ ), .B2(_07744_ ), .ZN(_07745_ ) );
NAND2_X1 _15787_ ( .A1(_07745_ ), .A2(_05245_ ), .ZN(_07746_ ) );
AOI21_X1 _15788_ ( .A(_07210_ ), .B1(_07222_ ), .B2(_07224_ ), .ZN(_07747_ ) );
OR3_X1 _15789_ ( .A1(_07747_ ), .A2(_05040_ ), .A3(_05045_ ), .ZN(_07748_ ) );
OAI21_X1 _15790_ ( .A(_05040_ ), .B1(_07747_ ), .B2(_05045_ ), .ZN(_07749_ ) );
NAND3_X1 _15791_ ( .A1(_07748_ ), .A2(_07074_ ), .A3(_07749_ ), .ZN(_07750_ ) );
NOR2_X1 _15792_ ( .A1(_06545_ ), .A2(_06622_ ), .ZN(_07751_ ) );
AND2_X1 _15793_ ( .A1(_07299_ ), .A2(_07751_ ), .ZN(_07752_ ) );
OAI211_X1 _15794_ ( .A(_06664_ ), .B(_06665_ ), .C1(_06509_ ), .C2(_06530_ ), .ZN(_07753_ ) );
OAI21_X1 _15795_ ( .A(_06489_ ), .B1(_06529_ ), .B2(_06527_ ), .ZN(_07754_ ) );
AND2_X1 _15796_ ( .A1(_07753_ ), .A2(_07754_ ), .ZN(_07755_ ) );
NOR3_X1 _15797_ ( .A1(_06627_ ), .A2(_06514_ ), .A3(_06510_ ), .ZN(_07756_ ) );
NOR3_X1 _15798_ ( .A1(_06660_ ), .A2(_06489_ ), .A3(_06515_ ), .ZN(_07757_ ) );
OR2_X1 _15799_ ( .A1(_07756_ ), .A2(_07757_ ), .ZN(_07758_ ) );
MUX2_X1 _15800_ ( .A(_07755_ ), .B(_07758_ ), .S(_06494_ ), .Z(_07759_ ) );
MUX2_X1 _15801_ ( .A(_06843_ ), .B(_07759_ ), .S(_06933_ ), .Z(_07760_ ) );
AOI221_X4 _15802_ ( .A(_07752_ ), .B1(_07226_ ), .B2(_07197_ ), .C1(_07760_ ), .C2(_07059_ ), .ZN(_07761_ ) );
AOI22_X1 _15803_ ( .A1(_06481_ ), .A2(_06483_ ), .B1(_07258_ ), .B2(_07286_ ), .ZN(_07762_ ) );
OAI211_X1 _15804_ ( .A(_06708_ ), .B(_06484_ ), .C1(_06499_ ), .C2(_06863_ ), .ZN(_07763_ ) );
AOI21_X1 _15805_ ( .A(_07002_ ), .B1(_07762_ ), .B2(_07763_ ), .ZN(_07764_ ) );
NOR3_X1 _15806_ ( .A1(_05038_ ), .A2(_05039_ ), .A3(_05167_ ), .ZN(_07765_ ) );
NOR3_X1 _15807_ ( .A1(_05036_ ), .A2(_05037_ ), .A3(_06795_ ), .ZN(_07766_ ) );
AND3_X1 _15808_ ( .A1(_07286_ ), .A2(_07258_ ), .A3(_06741_ ), .ZN(_07767_ ) );
NOR4_X1 _15809_ ( .A1(_07764_ ), .A2(_07765_ ), .A3(_07766_ ), .A4(_07767_ ), .ZN(_07768_ ) );
NAND3_X1 _15810_ ( .A1(_07750_ ), .A2(_07761_ ), .A3(_07768_ ), .ZN(_07769_ ) );
AOI21_X1 _15811_ ( .A(_07746_ ), .B1(_07769_ ), .B2(_07498_ ), .ZN(_07770_ ) );
OAI21_X1 _15812_ ( .A(_07207_ ), .B1(_05693_ ), .B2(_07091_ ), .ZN(_07771_ ) );
OAI21_X1 _15813_ ( .A(_07737_ ), .B1(_07770_ ), .B2(_07771_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
NAND2_X1 _15814_ ( .A1(_05741_ ), .A2(_06111_ ), .ZN(_07772_ ) );
NOR2_X1 _15815_ ( .A1(_07739_ ), .A2(_04387_ ), .ZN(_07773_ ) );
NOR3_X1 _15816_ ( .A1(_07740_ ), .A2(_07773_ ), .A3(_06886_ ), .ZN(_07774_ ) );
OAI22_X1 _15817_ ( .A1(_05733_ ), .A2(_06406_ ), .B1(_02865_ ), .B2(_06410_ ), .ZN(_07775_ ) );
OAI21_X1 _15818_ ( .A(_06425_ ), .B1(_07774_ ), .B2(_07775_ ), .ZN(_07776_ ) );
NAND2_X1 _15819_ ( .A1(_07776_ ), .A2(_05245_ ), .ZN(_07777_ ) );
AND3_X1 _15820_ ( .A1(_07222_ ), .A2(_07210_ ), .A3(_07224_ ), .ZN(_07778_ ) );
OR3_X1 _15821_ ( .A1(_07778_ ), .A2(_07747_ ), .A3(_06554_ ), .ZN(_07779_ ) );
NOR2_X1 _15822_ ( .A1(_06901_ ), .A2(_07052_ ), .ZN(_07780_ ) );
NAND2_X1 _15823_ ( .A1(_07780_ ), .A2(_06547_ ), .ZN(_07781_ ) );
OAI21_X1 _15824_ ( .A(_07781_ ), .B1(_06482_ ), .B2(_06486_ ), .ZN(_07782_ ) );
AOI21_X1 _15825_ ( .A(_07322_ ), .B1(_06499_ ), .B2(_06708_ ), .ZN(_07783_ ) );
NOR2_X1 _15826_ ( .A1(_07783_ ), .A2(_06485_ ), .ZN(_07784_ ) );
OAI21_X1 _15827_ ( .A(_06432_ ), .B1(_07782_ ), .B2(_07784_ ), .ZN(_07785_ ) );
NAND3_X1 _15828_ ( .A1(_07780_ ), .A2(_06547_ ), .A3(_06742_ ), .ZN(_07786_ ) );
AND3_X1 _15829_ ( .A1(_07252_ ), .A2(_06776_ ), .A3(_07253_ ), .ZN(_07787_ ) );
AOI21_X1 _15830_ ( .A(_07787_ ), .B1(_06710_ ), .B2(_07244_ ), .ZN(_07788_ ) );
OAI21_X1 _15831_ ( .A(_07058_ ), .B1(_07788_ ), .B2(_06790_ ), .ZN(_07789_ ) );
AOI21_X1 _15832_ ( .A(_07789_ ), .B1(_07052_ ), .B2(_06932_ ), .ZN(_07790_ ) );
AND3_X1 _15833_ ( .A1(_07338_ ), .A2(_07339_ ), .A3(_07751_ ), .ZN(_07791_ ) );
NOR2_X1 _15834_ ( .A1(_07790_ ), .A2(_07791_ ), .ZN(_07792_ ) );
OR2_X1 _15835_ ( .A1(_05046_ ), .A2(_06797_ ), .ZN(_07793_ ) );
AOI22_X1 _15836_ ( .A1(_05047_ ), .A2(_06687_ ), .B1(_05045_ ), .B2(_06979_ ), .ZN(_07794_ ) );
AND4_X1 _15837_ ( .A1(_07786_ ), .A2(_07792_ ), .A3(_07793_ ), .A4(_07794_ ), .ZN(_07795_ ) );
NAND3_X1 _15838_ ( .A1(_07779_ ), .A2(_07785_ ), .A3(_07795_ ), .ZN(_07796_ ) );
AOI21_X1 _15839_ ( .A(_07777_ ), .B1(_07796_ ), .B2(_07498_ ), .ZN(_07797_ ) );
OAI21_X1 _15840_ ( .A(_06099_ ), .B1(_05730_ ), .B2(_07091_ ), .ZN(_07798_ ) );
OAI21_X1 _15841_ ( .A(_07772_ ), .B1(_07797_ ), .B2(_07798_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _15842_ ( .A1(_05750_ ), .A2(_06111_ ), .ZN(_07799_ ) );
AND2_X1 _15843_ ( .A1(_07267_ ), .A2(_04410_ ), .ZN(_07800_ ) );
OR3_X1 _15844_ ( .A1(_07800_ ), .A2(_04433_ ), .A3(_05147_ ), .ZN(_07801_ ) );
OAI21_X1 _15845_ ( .A(_04433_ ), .B1(_07800_ ), .B2(_05147_ ), .ZN(_07802_ ) );
AND3_X1 _15846_ ( .A1(_07801_ ), .A2(_06421_ ), .A3(_07802_ ), .ZN(_07803_ ) );
OAI22_X1 _15847_ ( .A1(_05760_ ), .A2(_06406_ ), .B1(_02867_ ), .B2(_06410_ ), .ZN(_07804_ ) );
OAI21_X1 _15848_ ( .A(_06425_ ), .B1(_07803_ ), .B2(_07804_ ), .ZN(_07805_ ) );
NAND2_X1 _15849_ ( .A1(_07805_ ), .A2(_05245_ ), .ZN(_07806_ ) );
AND3_X1 _15850_ ( .A1(_06960_ ), .A2(_06643_ ), .A3(_06962_ ), .ZN(_07807_ ) );
AND2_X1 _15851_ ( .A1(_07807_ ), .A2(_06545_ ), .ZN(_07808_ ) );
OR2_X1 _15852_ ( .A1(_06862_ ), .A2(_07808_ ), .ZN(_07809_ ) );
AOI21_X1 _15853_ ( .A(_07372_ ), .B1(_06499_ ), .B2(_06708_ ), .ZN(_07810_ ) );
NOR2_X1 _15854_ ( .A1(_07810_ ), .A2(_06485_ ), .ZN(_07811_ ) );
OAI21_X1 _15855_ ( .A(_06431_ ), .B1(_07809_ ), .B2(_07811_ ), .ZN(_07812_ ) );
NAND2_X1 _15856_ ( .A1(_07379_ ), .A2(_07751_ ), .ZN(_07813_ ) );
NAND3_X1 _15857_ ( .A1(_06659_ ), .A2(_06661_ ), .A3(_06710_ ), .ZN(_07814_ ) );
NAND3_X1 _15858_ ( .A1(_07631_ ), .A2(_07377_ ), .A3(_07632_ ), .ZN(_07815_ ) );
NAND3_X1 _15859_ ( .A1(_07814_ ), .A2(_07815_ ), .A3(_06933_ ), .ZN(_07816_ ) );
AND2_X1 _15860_ ( .A1(_07816_ ), .A2(_07059_ ), .ZN(_07817_ ) );
OAI21_X1 _15861_ ( .A(_07817_ ), .B1(_06972_ ), .B2(_07054_ ), .ZN(_07818_ ) );
NAND3_X1 _15862_ ( .A1(_07807_ ), .A2(_07258_ ), .A3(_06742_ ), .ZN(_07819_ ) );
AND4_X1 _15863_ ( .A1(_07812_ ), .A2(_07813_ ), .A3(_07818_ ), .A4(_07819_ ), .ZN(_07820_ ) );
AOI21_X1 _15864_ ( .A(_05056_ ), .B1(_07212_ ), .B2(_07219_ ), .ZN(_07821_ ) );
NOR3_X1 _15865_ ( .A1(_07821_ ), .A2(_05053_ ), .A3(_05060_ ), .ZN(_07822_ ) );
NOR2_X1 _15866_ ( .A1(_07822_ ), .A2(_06554_ ), .ZN(_07823_ ) );
OAI21_X1 _15867_ ( .A(_05060_ ), .B1(_07821_ ), .B2(_05053_ ), .ZN(_07824_ ) );
NAND2_X1 _15868_ ( .A1(_07823_ ), .A2(_07824_ ), .ZN(_07825_ ) );
NAND2_X1 _15869_ ( .A1(_05060_ ), .A2(_06879_ ), .ZN(_07826_ ) );
NAND3_X1 _15870_ ( .A1(_06463_ ), .A2(_02815_ ), .A3(_06979_ ), .ZN(_07827_ ) );
OAI21_X1 _15871_ ( .A(_07197_ ), .B1(_06463_ ), .B2(_02815_ ), .ZN(_07828_ ) );
AND3_X1 _15872_ ( .A1(_07826_ ), .A2(_07827_ ), .A3(_07828_ ), .ZN(_07829_ ) );
NAND3_X1 _15873_ ( .A1(_07820_ ), .A2(_07825_ ), .A3(_07829_ ), .ZN(_07830_ ) );
AOI21_X1 _15874_ ( .A(_07806_ ), .B1(_07830_ ), .B2(_07498_ ), .ZN(_07831_ ) );
OAI21_X1 _15875_ ( .A(_06099_ ), .B1(_05755_ ), .B2(_07091_ ), .ZN(_07832_ ) );
OAI21_X1 _15876_ ( .A(_07799_ ), .B1(_07831_ ), .B2(_07832_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND3_X1 _15877_ ( .A1(_05772_ ), .A2(_05780_ ), .A3(_06152_ ), .ZN(_07833_ ) );
NOR2_X1 _15878_ ( .A1(_07267_ ), .A2(_04410_ ), .ZN(_07834_ ) );
NOR3_X1 _15879_ ( .A1(_07800_ ), .A2(_07834_ ), .A3(_06886_ ), .ZN(_07835_ ) );
OAI22_X1 _15880_ ( .A1(_05770_ ), .A2(_06406_ ), .B1(_02788_ ), .B2(_06410_ ), .ZN(_07836_ ) );
OAI21_X1 _15881_ ( .A(_06425_ ), .B1(_07835_ ), .B2(_07836_ ), .ZN(_07837_ ) );
NAND2_X1 _15882_ ( .A1(_07837_ ), .A2(_05245_ ), .ZN(_07838_ ) );
INV_X1 _15883_ ( .A(_06436_ ), .ZN(_07839_ ) );
AOI21_X1 _15884_ ( .A(_07237_ ), .B1(_06844_ ), .B2(_07839_ ), .ZN(_07840_ ) );
NOR2_X1 _15885_ ( .A1(_07011_ ), .A2(_06542_ ), .ZN(_07841_ ) );
AND2_X1 _15886_ ( .A1(_07841_ ), .A2(_06545_ ), .ZN(_07842_ ) );
OR3_X1 _15887_ ( .A1(_06862_ ), .A2(_07840_ ), .A3(_07842_ ), .ZN(_07843_ ) );
NAND2_X1 _15888_ ( .A1(_07843_ ), .A2(_06431_ ), .ZN(_07844_ ) );
OAI21_X1 _15889_ ( .A(_07751_ ), .B1(_07415_ ), .B2(_07416_ ), .ZN(_07845_ ) );
OAI21_X1 _15890_ ( .A(_06844_ ), .B1(_06769_ ), .B2(_07377_ ), .ZN(_07846_ ) );
AOI21_X1 _15891_ ( .A(_07846_ ), .B1(_07377_ ), .B2(_07726_ ), .ZN(_07847_ ) );
NOR2_X1 _15892_ ( .A1(_07847_ ), .A2(_07161_ ), .ZN(_07848_ ) );
OAI21_X1 _15893_ ( .A(_07848_ ), .B1(_07054_ ), .B2(_07022_ ), .ZN(_07849_ ) );
NAND3_X1 _15894_ ( .A1(_07841_ ), .A2(_07258_ ), .A3(_06742_ ), .ZN(_07850_ ) );
AND4_X1 _15895_ ( .A1(_07844_ ), .A2(_07845_ ), .A3(_07849_ ), .A4(_07850_ ), .ZN(_07851_ ) );
AOI21_X1 _15896_ ( .A(_06554_ ), .B1(_07220_ ), .B2(_05056_ ), .ZN(_07852_ ) );
OAI21_X1 _15897_ ( .A(_07852_ ), .B1(_05056_ ), .B2(_07220_ ), .ZN(_07853_ ) );
NOR3_X1 _15898_ ( .A1(_05053_ ), .A2(_05054_ ), .A3(_05167_ ), .ZN(_07854_ ) );
NOR3_X1 _15899_ ( .A1(_05051_ ), .A2(_05052_ ), .A3(_06795_ ), .ZN(_07855_ ) );
AOI21_X1 _15900_ ( .A(_06797_ ), .B1(_05051_ ), .B2(_05052_ ), .ZN(_07856_ ) );
NOR3_X1 _15901_ ( .A1(_07854_ ), .A2(_07855_ ), .A3(_07856_ ), .ZN(_07857_ ) );
NAND3_X1 _15902_ ( .A1(_07851_ ), .A2(_07853_ ), .A3(_07857_ ), .ZN(_07858_ ) );
AOI21_X1 _15903_ ( .A(_07838_ ), .B1(_07858_ ), .B2(_07498_ ), .ZN(_07859_ ) );
OAI21_X1 _15904_ ( .A(_06099_ ), .B1(_05767_ ), .B2(_07091_ ), .ZN(_07860_ ) );
OAI21_X1 _15905_ ( .A(_07833_ ), .B1(_07859_ ), .B2(_07860_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _15906_ ( .A1(_05799_ ), .A2(_06111_ ), .ZN(_07861_ ) );
OAI22_X1 _15907_ ( .A1(_05791_ ), .A2(_06406_ ), .B1(_02177_ ), .B2(_06410_ ), .ZN(_07862_ ) );
OAI21_X1 _15908_ ( .A(_05123_ ), .B1(_06417_ ), .B2(_05121_ ), .ZN(_07863_ ) );
NAND2_X1 _15909_ ( .A1(_07863_ ), .A2(_04089_ ), .ZN(_07864_ ) );
OAI21_X1 _15910_ ( .A(_07864_ ), .B1(_04088_ ), .B2(_06392_ ), .ZN(_07865_ ) );
XOR2_X1 _15911_ ( .A(_07865_ ), .B(_04052_ ), .Z(_07866_ ) );
AOI21_X1 _15912_ ( .A(_07862_ ), .B1(_07866_ ), .B2(_06422_ ), .ZN(_07867_ ) );
OAI21_X1 _15913_ ( .A(_05245_ ), .B1(_07867_ ), .B2(_06428_ ), .ZN(_07868_ ) );
AOI211_X1 _15914_ ( .A(_07099_ ), .B(_07098_ ), .C1(_06486_ ), .C2(_06497_ ), .ZN(_07869_ ) );
AND2_X1 _15915_ ( .A1(_07447_ ), .A2(_06545_ ), .ZN(_07870_ ) );
OAI21_X1 _15916_ ( .A(_06431_ ), .B1(_07869_ ), .B2(_07870_ ), .ZN(_07871_ ) );
NAND3_X1 _15917_ ( .A1(_07447_ ), .A2(_06546_ ), .A3(_06741_ ), .ZN(_07872_ ) );
NAND2_X1 _15918_ ( .A1(_07871_ ), .A2(_07872_ ), .ZN(_07873_ ) );
OR3_X1 _15919_ ( .A1(_07051_ ), .A2(_06544_ ), .A3(_06789_ ), .ZN(_07874_ ) );
OAI21_X1 _15920_ ( .A(_06789_ ), .B1(_07055_ ), .B2(_07056_ ), .ZN(_07875_ ) );
NAND2_X1 _15921_ ( .A1(_06837_ ), .A2(_06494_ ), .ZN(_07876_ ) );
OAI21_X1 _15922_ ( .A(_06770_ ), .B1(_07756_ ), .B2(_07757_ ), .ZN(_07877_ ) );
NAND2_X1 _15923_ ( .A1(_07876_ ), .A2(_07877_ ), .ZN(_07878_ ) );
OAI211_X1 _15924_ ( .A(_07875_ ), .B(_06619_ ), .C1(_07878_ ), .C2(_06975_ ), .ZN(_07879_ ) );
AOI21_X1 _15925_ ( .A(_06622_ ), .B1(_07874_ ), .B2(_07879_ ), .ZN(_07880_ ) );
OR2_X1 _15926_ ( .A1(_07873_ ), .A2(_07880_ ), .ZN(_07881_ ) );
AND2_X1 _15927_ ( .A1(_04860_ ), .A2(_06687_ ), .ZN(_07882_ ) );
NOR3_X1 _15928_ ( .A1(_04859_ ), .A2(_04051_ ), .A3(_06795_ ), .ZN(_07883_ ) );
AOI21_X1 _15929_ ( .A(_06797_ ), .B1(_04859_ ), .B2(_04051_ ), .ZN(_00304_ ) );
NOR4_X1 _15930_ ( .A1(_07881_ ), .A2(_07882_ ), .A3(_07883_ ), .A4(_00304_ ), .ZN(_00305_ ) );
NAND2_X1 _15931_ ( .A1(_06739_ ), .A2(_07211_ ), .ZN(_00306_ ) );
AOI21_X1 _15932_ ( .A(_07213_ ), .B1(_00306_ ), .B2(_07214_ ), .ZN(_00307_ ) );
NOR3_X1 _15933_ ( .A1(_00307_ ), .A2(_04860_ ), .A3(_07217_ ), .ZN(_00308_ ) );
NOR2_X1 _15934_ ( .A1(_00308_ ), .A2(_06554_ ), .ZN(_00309_ ) );
OAI21_X1 _15935_ ( .A(_04860_ ), .B1(_00307_ ), .B2(_07217_ ), .ZN(_00310_ ) );
NAND2_X1 _15936_ ( .A1(_00309_ ), .A2(_00310_ ), .ZN(_00311_ ) );
AOI21_X1 _15937_ ( .A(_06696_ ), .B1(_00305_ ), .B2(_00311_ ), .ZN(_00312_ ) );
OAI22_X1 _15938_ ( .A1(_07868_ ), .A2(_00312_ ), .B1(_07091_ ), .B2(_05785_ ), .ZN(_00313_ ) );
OAI21_X1 _15939_ ( .A(_07861_ ), .B1(_00313_ ), .B2(_06211_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _15940_ ( .A1(_05815_ ), .A2(_05817_ ), .A3(_06152_ ), .ZN(_00314_ ) );
AOI21_X1 _15941_ ( .A(_06886_ ), .B1(_07863_ ), .B2(_04089_ ), .ZN(_00315_ ) );
OAI21_X1 _15942_ ( .A(_00315_ ), .B1(_04089_ ), .B2(_07863_ ), .ZN(_00316_ ) );
AOI22_X1 _15943_ ( .A1(_05806_ ), .A2(_06404_ ), .B1(\ID_EX_imm [22] ), .B2(_06408_ ), .ZN(_00317_ ) );
AOI21_X1 _15944_ ( .A(_06426_ ), .B1(_00316_ ), .B2(_00317_ ), .ZN(_00318_ ) );
OR2_X1 _15945_ ( .A1(_00318_ ), .A2(_03778_ ), .ZN(_00319_ ) );
AND2_X1 _15946_ ( .A1(_07477_ ), .A2(_06545_ ), .ZN(_00320_ ) );
OR2_X1 _15947_ ( .A1(_06862_ ), .A2(_00320_ ), .ZN(_00321_ ) );
NOR4_X1 _15948_ ( .A1(_07098_ ), .A2(_06497_ ), .A3(_06485_ ), .A4(_07100_ ), .ZN(_00322_ ) );
OAI21_X1 _15949_ ( .A(_06431_ ), .B1(_00321_ ), .B2(_00322_ ), .ZN(_00323_ ) );
OR3_X1 _15950_ ( .A1(_04867_ ), .A2(_04088_ ), .A3(_06795_ ), .ZN(_00324_ ) );
AOI21_X1 _15951_ ( .A(_04828_ ), .B1(_04867_ ), .B2(_04088_ ), .ZN(_00325_ ) );
AOI21_X1 _15952_ ( .A(_00325_ ), .B1(_04868_ ), .B2(_06687_ ), .ZN(_00326_ ) );
NAND3_X1 _15953_ ( .A1(_07477_ ), .A2(_07258_ ), .A3(_06741_ ), .ZN(_00327_ ) );
NAND4_X1 _15954_ ( .A1(_00323_ ), .A2(_00324_ ), .A3(_00326_ ), .A4(_00327_ ), .ZN(_00328_ ) );
AND3_X1 _15955_ ( .A1(_00306_ ), .A2(_07213_ ), .A3(_07214_ ), .ZN(_00329_ ) );
NOR3_X1 _15956_ ( .A1(_00329_ ), .A2(_00307_ ), .A3(_06553_ ), .ZN(_00330_ ) );
OR3_X1 _15957_ ( .A1(_07124_ ), .A2(_06546_ ), .A3(_06790_ ), .ZN(_00331_ ) );
NOR3_X1 _15958_ ( .A1(_07120_ ), .A2(_07054_ ), .A3(_07121_ ), .ZN(_00332_ ) );
AND3_X1 _15959_ ( .A1(_07241_ ), .A2(_06844_ ), .A3(_07245_ ), .ZN(_00333_ ) );
OAI21_X1 _15960_ ( .A(_07258_ ), .B1(_00332_ ), .B2(_00333_ ), .ZN(_00334_ ) );
AOI21_X1 _15961_ ( .A(_06622_ ), .B1(_00331_ ), .B2(_00334_ ), .ZN(_00335_ ) );
OR3_X1 _15962_ ( .A1(_00328_ ), .A2(_00330_ ), .A3(_00335_ ), .ZN(_00336_ ) );
AOI21_X1 _15963_ ( .A(_00319_ ), .B1(_06698_ ), .B2(_00336_ ), .ZN(_00337_ ) );
OAI21_X1 _15964_ ( .A(_06099_ ), .B1(_05804_ ), .B2(_07091_ ), .ZN(_00338_ ) );
OAI21_X1 _15965_ ( .A(_00314_ ), .B1(_00337_ ), .B2(_00338_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NAND3_X1 _15966_ ( .A1(_05308_ ), .A2(_05309_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_00339_ ) );
AND4_X1 _15967_ ( .A1(_05853_ ), .A2(_05854_ ), .A3(_05855_ ), .A4(_05856_ ), .ZN(_00340_ ) );
OAI21_X1 _15968_ ( .A(_00339_ ), .B1(_00340_ ), .B2(_03871_ ), .ZN(_00341_ ) );
NAND2_X1 _15969_ ( .A1(_00341_ ), .A2(_06111_ ), .ZN(_00342_ ) );
NOR2_X1 _15970_ ( .A1(_07234_ ), .A2(_04844_ ), .ZN(_00343_ ) );
AOI21_X1 _15971_ ( .A(_06554_ ), .B1(_00343_ ), .B2(_04841_ ), .ZN(_00344_ ) );
OAI21_X1 _15972_ ( .A(_00344_ ), .B1(_04841_ ), .B2(_00343_ ), .ZN(_00345_ ) );
AND2_X1 _15973_ ( .A1(_06439_ ), .A2(_02928_ ), .ZN(_00346_ ) );
OAI21_X1 _15974_ ( .A(_06431_ ), .B1(_06481_ ), .B2(_00346_ ), .ZN(_00347_ ) );
NAND3_X1 _15975_ ( .A1(_07053_ ), .A2(_07057_ ), .A3(_07751_ ), .ZN(_00348_ ) );
AOI21_X1 _15976_ ( .A(_06536_ ), .B1(_04838_ ), .B2(_06490_ ), .ZN(_00349_ ) );
MUX2_X1 _15977_ ( .A(_07635_ ), .B(_00349_ ), .S(_06489_ ), .Z(_00350_ ) );
MUX2_X1 _15978_ ( .A(_07755_ ), .B(_00350_ ), .S(_06776_ ), .Z(_00351_ ) );
MUX2_X1 _15979_ ( .A(_07878_ ), .B(_00351_ ), .S(_06933_ ), .Z(_00352_ ) );
NAND2_X1 _15980_ ( .A1(_00352_ ), .A2(_07059_ ), .ZN(_00353_ ) );
NAND3_X1 _15981_ ( .A1(_06439_ ), .A2(_02928_ ), .A3(_06741_ ), .ZN(_00354_ ) );
OR2_X1 _15982_ ( .A1(_04840_ ), .A2(_06795_ ), .ZN(_00355_ ) );
AND3_X1 _15983_ ( .A1(_04839_ ), .A2(_04840_ ), .A3(_05166_ ), .ZN(_00356_ ) );
AOI21_X1 _15984_ ( .A(_00356_ ), .B1(_04839_ ), .B2(_04827_ ), .ZN(_00357_ ) );
AND3_X1 _15985_ ( .A1(_00354_ ), .A2(_00355_ ), .A3(_00357_ ), .ZN(_00358_ ) );
AND4_X1 _15986_ ( .A1(_00347_ ), .A2(_00348_ ), .A3(_00353_ ), .A4(_00358_ ), .ZN(_00359_ ) );
AOI21_X1 _15987_ ( .A(_06696_ ), .B1(_00345_ ), .B2(_00359_ ), .ZN(_00360_ ) );
OR2_X1 _15988_ ( .A1(_05849_ ), .A2(_06406_ ), .ZN(_00361_ ) );
AOI21_X1 _15989_ ( .A(_05159_ ), .B1(_07271_ ), .B2(_04341_ ), .ZN(_00362_ ) );
XNOR2_X1 _15990_ ( .A(_00362_ ), .B(_04317_ ), .ZN(_00363_ ) );
AOI22_X1 _15991_ ( .A1(_00363_ ), .A2(_06422_ ), .B1(\ID_EX_imm [31] ), .B2(_06704_ ), .ZN(_00364_ ) );
AOI21_X1 _15992_ ( .A(_06427_ ), .B1(_00361_ ), .B2(_00364_ ), .ZN(_00365_ ) );
NOR3_X1 _15993_ ( .A1(_00360_ ), .A2(_05852_ ), .A3(_00365_ ), .ZN(_00366_ ) );
NAND2_X1 _15994_ ( .A1(_05862_ ), .A2(_05184_ ), .ZN(_00367_ ) );
NAND2_X1 _15995_ ( .A1(_00367_ ), .A2(_06234_ ), .ZN(_00368_ ) );
OAI21_X1 _15996_ ( .A(_00342_ ), .B1(_00366_ ), .B2(_00368_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
AND3_X1 _15997_ ( .A1(\myexu.state_$_ANDNOT__B_Y ), .A2(_03796_ ), .A3(_03798_ ), .ZN(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ) );
NOR2_X1 _15998_ ( .A1(_06024_ ), .A2(reset ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _15999_ ( .A1(_03282_ ), .A2(IDU_valid_EXU ), .ZN(_00369_ ) );
OAI21_X1 _16000_ ( .A(_00369_ ), .B1(_03220_ ), .B2(_03150_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16001_ ( .A1(_03217_ ), .A2(_03150_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16002_ ( .A1(_03217_ ), .A2(_03150_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16003_ ( .A1(_03527_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_02990_ ), .A4(_03146_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AND2_X1 _16004_ ( .A1(_03220_ ), .A2(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
AOI21_X1 _16005_ ( .A(_03729_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16006_ ( .A(_03147_ ), .ZN(_00370_ ) );
OAI21_X1 _16007_ ( .A(_00369_ ), .B1(_00370_ ), .B2(_03282_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16008_ ( .A1(_03147_ ), .A2(_03282_ ), .B1(_03792_ ), .B2(_03248_ ), .ZN(_00371_ ) );
INV_X1 _16009_ ( .A(loaduse_clear ), .ZN(_00372_ ) );
AOI221_X4 _16010_ ( .A(_00371_ ), .B1(\myidu.state [2] ), .B2(_00372_ ), .C1(_03217_ ), .C2(_03729_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
NAND3_X1 _16011_ ( .A1(_03060_ ), .A2(IDU_valid_EXU ), .A3(_05893_ ), .ZN(_00373_ ) );
NAND2_X1 _16012_ ( .A1(_00208_ ), .A2(loaduse_clear ), .ZN(_00374_ ) );
NAND4_X1 _16013_ ( .A1(_03191_ ), .A2(_03193_ ), .A3(_03213_ ), .A4(_03210_ ), .ZN(_00375_ ) );
NOR3_X1 _16014_ ( .A1(_03178_ ), .A2(_03182_ ), .A3(_00375_ ), .ZN(_00376_ ) );
AND2_X1 _16015_ ( .A1(_03071_ ), .A2(_03291_ ), .ZN(_00377_ ) );
BUF_X2 _16016_ ( .A(_00377_ ), .Z(_00378_ ) );
AOI21_X1 _16017_ ( .A(_03269_ ), .B1(_00376_ ), .B2(_00378_ ), .ZN(_00379_ ) );
INV_X1 _16018_ ( .A(_00379_ ), .ZN(_00380_ ) );
OAI21_X1 _16019_ ( .A(_03261_ ), .B1(_03279_ ), .B2(_03010_ ), .ZN(_00381_ ) );
NAND2_X1 _16020_ ( .A1(_00380_ ), .A2(_00381_ ), .ZN(_00382_ ) );
NAND3_X1 _16021_ ( .A1(_03147_ ), .A2(IDU_ready_IFU ), .A3(_02989_ ), .ZN(_00383_ ) );
OAI211_X1 _16022_ ( .A(_00373_ ), .B(_00374_ ), .C1(_00382_ ), .C2(_00383_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16023_ ( .A(_03060_ ), .B(_03775_ ), .C1(_03147_ ), .C2(_03282_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
OAI221_X1 _16024_ ( .A(_03145_ ), .B1(_03261_ ), .B2(_03268_ ), .C1(_03141_ ), .C2(_03142_ ), .ZN(_00384_ ) );
AOI21_X1 _16025_ ( .A(_00384_ ), .B1(_00376_ ), .B2(_00378_ ), .ZN(_00385_ ) );
OAI211_X1 _16026_ ( .A(_03145_ ), .B(_03261_ ), .C1(_03141_ ), .C2(_03142_ ), .ZN(_00386_ ) );
AOI21_X1 _16027_ ( .A(_00386_ ), .B1(_03278_ ), .B2(_03187_ ), .ZN(_00387_ ) );
OAI211_X1 _16028_ ( .A(IDU_ready_IFU ), .B(_03060_ ), .C1(_00385_ ), .C2(_00387_ ), .ZN(_00388_ ) );
NAND3_X1 _16029_ ( .A1(_03060_ ), .A2(\myidu.state [2] ), .A3(_00372_ ), .ZN(_00389_ ) );
NAND2_X1 _16030_ ( .A1(_00388_ ), .A2(_00389_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16031_ ( .A1(_03144_ ), .A2(IDU_ready_IFU ), .ZN(_00390_ ) );
NOR2_X1 _16032_ ( .A1(_03144_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00391_ ) );
NOR2_X1 _16033_ ( .A1(\myifu.state [0] ), .A2(\myifu.state [1] ), .ZN(_00392_ ) );
NOR4_X1 _16034_ ( .A1(_00390_ ), .A2(_00391_ ), .A3(reset ), .A4(_00392_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
CLKBUF_X2 _16035_ ( .A(_05954_ ), .Z(_00393_ ) );
OR3_X1 _16036_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00394_ ) );
OAI21_X1 _16037_ ( .A(_00394_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_05956_ ), .ZN(_00395_ ) );
MUX2_X1 _16038_ ( .A(\io_master_rdata [31] ), .B(_00395_ ), .S(_03707_ ), .Z(_00396_ ) );
AND2_X1 _16039_ ( .A1(_00396_ ), .A2(_01918_ ), .ZN(\myifu.data_in [31] ) );
CLKBUF_X2 _16040_ ( .A(_00393_ ), .Z(_00397_ ) );
OR3_X1 _16041_ ( .A1(_01916_ ), .A2(_01454_ ), .A3(_00397_ ), .ZN(_00398_ ) );
OAI211_X1 _16042_ ( .A(_03714_ ), .B(_00398_ ), .C1(_01575_ ), .C2(_05957_ ), .ZN(_00399_ ) );
OAI21_X1 _16043_ ( .A(\io_master_rdata [30] ), .B1(_01914_ ), .B2(_01988_ ), .ZN(_00400_ ) );
AOI21_X1 _16044_ ( .A(_05925_ ), .B1(_00399_ ), .B2(_00400_ ), .ZN(\myifu.data_in [30] ) );
AND2_X4 _16045_ ( .A1(_03719_ ), .A2(_03722_ ), .ZN(_00401_ ) );
BUF_X8 _16046_ ( .A(_00401_ ), .Z(_00402_ ) );
BUF_X4 _16047_ ( .A(_00402_ ), .Z(_00403_ ) );
BUF_X2 _16048_ ( .A(_00403_ ), .Z(_00404_ ) );
BUF_X2 _16049_ ( .A(_00404_ ), .Z(_00405_ ) );
OR2_X1 _16050_ ( .A1(_00405_ ), .A2(\io_master_rdata [21] ), .ZN(_00406_ ) );
CLKBUF_X2 _16051_ ( .A(_00397_ ), .Z(_00407_ ) );
OR3_X1 _16052_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00408_ ) );
OAI211_X1 _16053_ ( .A(_00405_ ), .B(_00408_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00409_ ) );
AND3_X1 _16054_ ( .A1(_00406_ ), .A2(_00409_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [21] ) );
OR3_X1 _16055_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00410_ ) );
OAI211_X1 _16056_ ( .A(_00403_ ), .B(_00410_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05956_ ), .ZN(_00411_ ) );
OAI21_X1 _16057_ ( .A(_00411_ ), .B1(_00403_ ), .B2(\io_master_rdata [20] ), .ZN(_00412_ ) );
NOR2_X1 _16058_ ( .A1(_00412_ ), .A2(_01993_ ), .ZN(\myifu.data_in [20] ) );
OR3_X1 _16059_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00413_ ) );
OAI211_X1 _16060_ ( .A(_00403_ ), .B(_00413_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05956_ ), .ZN(_00414_ ) );
OAI21_X1 _16061_ ( .A(_00414_ ), .B1(\io_master_rdata [19] ), .B2(_00403_ ), .ZN(_00415_ ) );
BUF_X4 _16062_ ( .A(_05932_ ), .Z(_00416_ ) );
NOR2_X1 _16063_ ( .A1(_00415_ ), .A2(_00416_ ), .ZN(\myifu.data_in [19] ) );
OR3_X1 _16064_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00417_ ) );
OAI211_X1 _16065_ ( .A(_00402_ ), .B(_00417_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05955_ ), .ZN(_00418_ ) );
OAI21_X1 _16066_ ( .A(_00418_ ), .B1(\io_master_rdata [18] ), .B2(_00402_ ), .ZN(_00419_ ) );
NOR2_X1 _16067_ ( .A1(_00419_ ), .A2(_05924_ ), .ZN(\myifu.data_in [18] ) );
OR3_X1 _16068_ ( .A1(_01869_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05954_ ), .ZN(_00420_ ) );
OAI211_X1 _16069_ ( .A(_00402_ ), .B(_00420_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05955_ ), .ZN(_00421_ ) );
OAI21_X2 _16070_ ( .A(_00421_ ), .B1(_00402_ ), .B2(\io_master_rdata [17] ), .ZN(_00422_ ) );
NOR2_X1 _16071_ ( .A1(_00422_ ), .A2(_00416_ ), .ZN(\myifu.data_in [17] ) );
OR2_X1 _16072_ ( .A1(_00405_ ), .A2(\io_master_rdata [16] ), .ZN(_00423_ ) );
OR3_X1 _16073_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00424_ ) );
OAI211_X1 _16074_ ( .A(_00405_ ), .B(_00424_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00425_ ) );
AND3_X1 _16075_ ( .A1(_00423_ ), .A2(_00425_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16076_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00426_ ) );
OAI211_X1 _16077_ ( .A(_00403_ ), .B(_00426_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05955_ ), .ZN(_00427_ ) );
OAI21_X1 _16078_ ( .A(_00427_ ), .B1(_00403_ ), .B2(\io_master_rdata [15] ), .ZN(_00428_ ) );
NOR2_X1 _16079_ ( .A1(_00428_ ), .A2(_00416_ ), .ZN(\myifu.data_in [15] ) );
BUF_X2 _16080_ ( .A(_00404_ ), .Z(_00429_ ) );
OR2_X1 _16081_ ( .A1(_00429_ ), .A2(\io_master_rdata [14] ), .ZN(_00430_ ) );
OR3_X1 _16082_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00431_ ) );
OAI211_X1 _16083_ ( .A(_00429_ ), .B(_00431_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00432_ ) );
AND3_X1 _16084_ ( .A1(_00430_ ), .A2(_00432_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16085_ ( .A1(_00405_ ), .A2(\io_master_rdata [13] ), .ZN(_00433_ ) );
OR3_X1 _16086_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00434_ ) );
OAI211_X1 _16087_ ( .A(_00429_ ), .B(_00434_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00435_ ) );
AND3_X1 _16088_ ( .A1(_00433_ ), .A2(_00435_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _16089_ ( .A1(_00404_ ), .A2(\io_master_rdata [12] ), .ZN(_00436_ ) );
OR3_X1 _16090_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00437_ ) );
OAI211_X1 _16091_ ( .A(_00404_ ), .B(_00437_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05957_ ), .ZN(_00438_ ) );
AND3_X1 _16092_ ( .A1(_00436_ ), .A2(_00438_ ), .A3(_01918_ ), .ZN(\myifu.data_in [12] ) );
MUX2_X1 _16093_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_05957_ ), .Z(_00439_ ) );
OR3_X1 _16094_ ( .A1(_01914_ ), .A2(_01988_ ), .A3(_00439_ ), .ZN(_00440_ ) );
OAI21_X1 _16095_ ( .A(\io_master_rdata [29] ), .B1(_01914_ ), .B2(_01988_ ), .ZN(_00441_ ) );
AOI21_X1 _16096_ ( .A(_05925_ ), .B1(_00440_ ), .B2(_00441_ ), .ZN(\myifu.data_in [29] ) );
OR3_X1 _16097_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00442_ ) );
OAI21_X1 _16098_ ( .A(_00442_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_05957_ ), .ZN(_00443_ ) );
MUX2_X1 _16099_ ( .A(\io_master_rdata [11] ), .B(_00443_ ), .S(_03707_ ), .Z(_00444_ ) );
AND2_X1 _16100_ ( .A1(_00444_ ), .A2(_01918_ ), .ZN(\myifu.data_in [11] ) );
OR3_X1 _16101_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00445_ ) );
OAI21_X1 _16102_ ( .A(_00445_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_05956_ ), .ZN(_00446_ ) );
MUX2_X1 _16103_ ( .A(\io_master_rdata [10] ), .B(_00446_ ), .S(_03714_ ), .Z(_00447_ ) );
AND2_X1 _16104_ ( .A1(_00447_ ), .A2(_01918_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16105_ ( .A1(_00404_ ), .A2(\io_master_rdata [9] ), .ZN(_00448_ ) );
OR3_X1 _16106_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00449_ ) );
OAI211_X1 _16107_ ( .A(_00404_ ), .B(_00449_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05957_ ), .ZN(_00450_ ) );
AND3_X1 _16108_ ( .A1(_00448_ ), .A2(_00450_ ), .A3(_01918_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16109_ ( .A1(_00429_ ), .A2(\io_master_rdata [8] ), .ZN(_00451_ ) );
OR3_X1 _16110_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00452_ ) );
OAI211_X1 _16111_ ( .A(_00429_ ), .B(_00452_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00453_ ) );
AND3_X1 _16112_ ( .A1(_00451_ ), .A2(_00453_ ), .A3(_01918_ ), .ZN(\myifu.data_in [8] ) );
OR3_X1 _16113_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00454_ ) );
OAI211_X1 _16114_ ( .A(_00404_ ), .B(_00454_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05957_ ), .ZN(_00455_ ) );
OAI21_X1 _16115_ ( .A(_00455_ ), .B1(\io_master_rdata [7] ), .B2(_00404_ ), .ZN(_00456_ ) );
NOR2_X1 _16116_ ( .A1(_00456_ ), .A2(_00416_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16117_ ( .A1(_01918_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00457_ ) );
OAI211_X1 _16118_ ( .A(_00429_ ), .B(_00457_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00458_ ) );
OAI21_X1 _16119_ ( .A(_00458_ ), .B1(\io_master_rdata [6] ), .B2(_00429_ ), .ZN(_00459_ ) );
NOR2_X1 _16120_ ( .A1(_00459_ ), .A2(_00416_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16121_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00460_ ) );
OAI211_X1 _16122_ ( .A(_00429_ ), .B(_00460_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00461_ ) );
OAI21_X1 _16123_ ( .A(_00461_ ), .B1(\io_master_rdata [5] ), .B2(_00429_ ), .ZN(_00462_ ) );
NOR2_X1 _16124_ ( .A1(_00462_ ), .A2(_00416_ ), .ZN(\myifu.data_in [5] ) );
BUF_X4 _16125_ ( .A(_00403_ ), .Z(_00463_ ) );
OR3_X1 _16126_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00464_ ) );
OAI211_X1 _16127_ ( .A(_00463_ ), .B(_00464_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05956_ ), .ZN(_00465_ ) );
OAI21_X1 _16128_ ( .A(_00465_ ), .B1(\io_master_rdata [4] ), .B2(_00463_ ), .ZN(_00466_ ) );
NOR2_X1 _16129_ ( .A1(_00466_ ), .A2(_01993_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16130_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00467_ ) );
OAI211_X1 _16131_ ( .A(_00463_ ), .B(_00467_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05956_ ), .ZN(_00468_ ) );
OAI21_X1 _16132_ ( .A(_00468_ ), .B1(\io_master_rdata [3] ), .B2(_00463_ ), .ZN(_00469_ ) );
NOR2_X1 _16133_ ( .A1(_00469_ ), .A2(_00416_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16134_ ( .A1(_01869_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05954_ ), .ZN(_00470_ ) );
OAI211_X1 _16135_ ( .A(_00402_ ), .B(_00470_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05955_ ), .ZN(_00471_ ) );
OAI21_X2 _16136_ ( .A(_00471_ ), .B1(\io_master_rdata [2] ), .B2(_00402_ ), .ZN(_00472_ ) );
NOR2_X1 _16137_ ( .A1(_00472_ ), .A2(_00416_ ), .ZN(\myifu.data_in [2] ) );
OR3_X1 _16138_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00473_ ) );
OAI211_X1 _16139_ ( .A(_00463_ ), .B(_00473_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05956_ ), .ZN(_00474_ ) );
OAI21_X1 _16140_ ( .A(_00474_ ), .B1(_00463_ ), .B2(\io_master_rdata [28] ), .ZN(_00475_ ) );
NOR2_X1 _16141_ ( .A1(_00475_ ), .A2(_00416_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16142_ ( .A1(_01869_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_05954_ ), .ZN(_00476_ ) );
OAI211_X1 _16143_ ( .A(_00402_ ), .B(_00476_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05955_ ), .ZN(_00477_ ) );
OAI21_X2 _16144_ ( .A(_00477_ ), .B1(\io_master_rdata [1] ), .B2(_00402_ ), .ZN(_00478_ ) );
NOR2_X1 _16145_ ( .A1(_00478_ ), .A2(_00416_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16146_ ( .A1(_01917_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00407_ ), .ZN(_00479_ ) );
OAI211_X1 _16147_ ( .A(_00405_ ), .B(_00479_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00480_ ) );
OAI21_X1 _16148_ ( .A(_00480_ ), .B1(\io_master_rdata [0] ), .B2(_00429_ ), .ZN(_00481_ ) );
NOR2_X1 _16149_ ( .A1(_00481_ ), .A2(_05925_ ), .ZN(\myifu.data_in [0] ) );
OR3_X1 _16150_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00482_ ) );
OAI211_X1 _16151_ ( .A(_00463_ ), .B(_00482_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05957_ ), .ZN(_00483_ ) );
OAI21_X1 _16152_ ( .A(_00483_ ), .B1(_00463_ ), .B2(\io_master_rdata [27] ), .ZN(_00484_ ) );
NOR2_X1 _16153_ ( .A1(_00484_ ), .A2(_05925_ ), .ZN(\myifu.data_in [27] ) );
OR3_X1 _16154_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00485_ ) );
OAI211_X1 _16155_ ( .A(_00403_ ), .B(_00485_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05956_ ), .ZN(_00486_ ) );
OAI21_X1 _16156_ ( .A(_00486_ ), .B1(_00463_ ), .B2(\io_master_rdata [26] ), .ZN(_00487_ ) );
NOR2_X1 _16157_ ( .A1(_00487_ ), .A2(_05925_ ), .ZN(\myifu.data_in [26] ) );
OR3_X1 _16158_ ( .A1(_01915_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00393_ ), .ZN(_00488_ ) );
OAI211_X1 _16159_ ( .A(_00403_ ), .B(_00488_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05956_ ), .ZN(_00489_ ) );
OAI21_X1 _16160_ ( .A(_00489_ ), .B1(_00463_ ), .B2(\io_master_rdata [25] ), .ZN(_00490_ ) );
NOR2_X1 _16161_ ( .A1(_00490_ ), .A2(_05925_ ), .ZN(\myifu.data_in [25] ) );
OR2_X1 _16162_ ( .A1(_00405_ ), .A2(\io_master_rdata [24] ), .ZN(_00491_ ) );
OR3_X1 _16163_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00492_ ) );
OAI211_X1 _16164_ ( .A(_00405_ ), .B(_00492_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05957_ ), .ZN(_00493_ ) );
AND3_X1 _16165_ ( .A1(_00491_ ), .A2(_00493_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16166_ ( .A1(_01916_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00397_ ), .ZN(_00494_ ) );
OAI211_X1 _16167_ ( .A(_00404_ ), .B(_00494_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_05957_ ), .ZN(_00495_ ) );
OAI21_X1 _16168_ ( .A(_00495_ ), .B1(\io_master_rdata [23] ), .B2(_00404_ ), .ZN(_00496_ ) );
NOR2_X1 _16169_ ( .A1(_00496_ ), .A2(_05925_ ), .ZN(\myifu.data_in [23] ) );
OR2_X1 _16170_ ( .A1(_00405_ ), .A2(\io_master_rdata [22] ), .ZN(_00497_ ) );
OR3_X1 _16171_ ( .A1(_01917_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00407_ ), .ZN(_00498_ ) );
OAI211_X1 _16172_ ( .A(_00405_ ), .B(_00498_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00499_ ) );
AND3_X1 _16173_ ( .A1(_00497_ ), .A2(_00499_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16174_ ( .A(_00242_ ), .ZN(_00500_ ) );
NAND2_X1 _16175_ ( .A1(_00500_ ), .A2(_01989_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16176_ ( .A1(_05892_ ), .A2(fanout_net_8 ), .ZN(_00501_ ) );
INV_X1 _16177_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00502_ ) );
OAI21_X1 _16178_ ( .A(_01989_ ), .B1(_00501_ ), .B2(_00502_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16179_ ( .A1(_03655_ ), .A2(fanout_net_12 ), .ZN(_00503_ ) );
OAI21_X1 _16180_ ( .A(_01989_ ), .B1(_00503_ ), .B2(_00502_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16181_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .ZN(_00504_ ) );
OAI21_X1 _16182_ ( .A(_01989_ ), .B1(_00504_ ), .B2(_00502_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
INV_X1 _16183_ ( .A(\IF_ID_inst [16] ), .ZN(_00505_ ) );
OR2_X1 _16184_ ( .A1(_03187_ ), .A2(_00505_ ), .ZN(_00506_ ) );
AND2_X1 _16185_ ( .A1(_00378_ ), .A2(_03235_ ), .ZN(_00507_ ) );
AOI211_X1 _16186_ ( .A(_03046_ ), .B(_03089_ ), .C1(_03048_ ), .C2(_03054_ ), .ZN(_00508_ ) );
AND4_X1 _16187_ ( .A1(_03187_ ), .A2(_00508_ ), .A3(_03315_ ), .A4(_03295_ ), .ZN(_00509_ ) );
NAND3_X1 _16188_ ( .A1(_00507_ ), .A2(_03183_ ), .A3(_00509_ ), .ZN(_00510_ ) );
AND2_X1 _16189_ ( .A1(_00510_ ), .A2(_03286_ ), .ZN(_00511_ ) );
OAI221_X1 _16190_ ( .A(_00506_ ), .B1(_03028_ ), .B2(_00378_ ), .C1(_00511_ ), .C2(_03006_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
NOR2_X1 _16191_ ( .A1(_03278_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00512_ ) );
INV_X1 _16192_ ( .A(_00512_ ), .ZN(_00513_ ) );
INV_X1 _16193_ ( .A(_03496_ ), .ZN(_00514_ ) );
BUF_X4 _16194_ ( .A(_00514_ ), .Z(_00515_ ) );
OAI211_X1 _16195_ ( .A(_00513_ ), .B(_00515_ ), .C1(_02988_ ), .C2(_00507_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
INV_X1 _16196_ ( .A(_03291_ ), .ZN(_00516_ ) );
OAI21_X1 _16197_ ( .A(\IF_ID_inst [31] ), .B1(_03072_ ), .B2(_00516_ ), .ZN(_00517_ ) );
AND2_X1 _16198_ ( .A1(_00513_ ), .A2(_00517_ ), .ZN(_00518_ ) );
BUF_X4 _16199_ ( .A(_00518_ ), .Z(_00519_ ) );
BUF_X4 _16200_ ( .A(_03235_ ), .Z(_00520_ ) );
OAI211_X1 _16201_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03005_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16202_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03006_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16203_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03011_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
INV_X1 _16204_ ( .A(\IF_ID_inst [19] ), .ZN(_00521_ ) );
NOR2_X1 _16205_ ( .A1(_03089_ ), .A2(_03094_ ), .ZN(_00522_ ) );
BUF_X4 _16206_ ( .A(_03278_ ), .Z(_00523_ ) );
OAI221_X1 _16207_ ( .A(_00517_ ), .B1(_00521_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
INV_X1 _16208_ ( .A(\IF_ID_inst [18] ), .ZN(_00524_ ) );
OAI221_X1 _16209_ ( .A(_00517_ ), .B1(_00524_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
INV_X1 _16210_ ( .A(\IF_ID_inst [17] ), .ZN(_00525_ ) );
OAI221_X1 _16211_ ( .A(_00517_ ), .B1(_00525_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16212_ ( .A(_00517_ ), .B1(_00505_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
INV_X1 _16213_ ( .A(\IF_ID_inst [15] ), .ZN(_00526_ ) );
OAI221_X1 _16214_ ( .A(_00517_ ), .B1(_00526_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16215_ ( .A(_00517_ ), .B1(_03167_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16216_ ( .A(_00517_ ), .B1(_03063_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16217_ ( .A(_00517_ ), .B1(_03067_ ), .B2(_00522_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16218_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03012_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
INV_X1 _16219_ ( .A(\IF_ID_inst [7] ), .ZN(_00527_ ) );
OR2_X1 _16220_ ( .A1(_03291_ ), .A2(_00527_ ), .ZN(_00528_ ) );
OR2_X1 _16221_ ( .A1(_03071_ ), .A2(_02988_ ), .ZN(_00529_ ) );
NAND4_X1 _16222_ ( .A1(_00513_ ), .A2(_03428_ ), .A3(_00528_ ), .A4(_00529_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16223_ ( .A(_03437_ ), .ZN(_00530_ ) );
OAI221_X1 _16224_ ( .A(_00530_ ), .B1(_00378_ ), .B2(_03005_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
INV_X1 _16225_ ( .A(_03433_ ), .ZN(_00531_ ) );
OAI221_X1 _16226_ ( .A(_00531_ ), .B1(_00378_ ), .B2(_03012_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00523_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16227_ ( .A(_03408_ ), .ZN(_00532_ ) );
OAI221_X1 _16228_ ( .A(_00532_ ), .B1(_00378_ ), .B2(_03013_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .C2(_03278_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
INV_X1 _16229_ ( .A(_03398_ ), .ZN(_00533_ ) );
OAI221_X1 _16230_ ( .A(_00533_ ), .B1(_00378_ ), .B2(_03014_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_03278_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16231_ ( .A(_03394_ ), .ZN(_00534_ ) );
OAI221_X1 _16232_ ( .A(_00534_ ), .B1(_00378_ ), .B2(_03015_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .C2(_03278_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16233_ ( .A(_03386_ ), .ZN(_00535_ ) );
OAI221_X1 _16234_ ( .A(_00535_ ), .B1(_00378_ ), .B2(_03016_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .C2(_03278_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16235_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03013_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16236_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03014_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16237_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03015_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16238_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03016_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16239_ ( .A(_00519_ ), .B(_00515_ ), .C1(_03017_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16240_ ( .A(_00519_ ), .B(_00514_ ), .C1(_03018_ ), .C2(_00520_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16241_ ( .A(_00518_ ), .B(_00514_ ), .C1(_03019_ ), .C2(_03235_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16242_ ( .A(\IF_ID_inst [11] ), .B1(_03072_ ), .B2(_00516_ ), .ZN(_00536_ ) );
OAI221_X1 _16243_ ( .A(_00536_ ), .B1(_00521_ ), .B2(_03187_ ), .C1(_00511_ ), .C2(_03017_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16244_ ( .A(\IF_ID_inst [10] ), .B1(_03072_ ), .B2(_00516_ ), .ZN(_00537_ ) );
OAI221_X1 _16245_ ( .A(_00537_ ), .B1(_00524_ ), .B2(_03187_ ), .C1(_00511_ ), .C2(_03018_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16246_ ( .A(\IF_ID_inst [9] ), .B1(_03072_ ), .B2(_00516_ ), .ZN(_00538_ ) );
OAI221_X1 _16247_ ( .A(_00538_ ), .B1(_00525_ ), .B2(_03187_ ), .C1(_00511_ ), .C2(_03019_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16248_ ( .A1(_03071_ ), .A2(_00527_ ), .ZN(_00539_ ) );
OAI221_X1 _16249_ ( .A(_00539_ ), .B1(_00526_ ), .B2(_03187_ ), .C1(_00510_ ), .C2(_03011_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
INV_X1 _16250_ ( .A(\myifu.state [2] ), .ZN(_00540_ ) );
BUF_X4 _16251_ ( .A(_00540_ ), .Z(_00541_ ) );
AND2_X2 _16252_ ( .A1(_03713_ ), .A2(_03725_ ), .ZN(_00542_ ) );
AOI21_X1 _16253_ ( .A(\IF_ID_pc [1] ), .B1(_03727_ ), .B2(\IF_ID_pc [2] ), .ZN(_00543_ ) );
INV_X1 _16254_ ( .A(_00543_ ), .ZN(_00544_ ) );
OAI21_X1 _16255_ ( .A(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .B1(_03727_ ), .B2(\IF_ID_pc [2] ), .ZN(_00545_ ) );
NOR2_X1 _16256_ ( .A1(_00544_ ), .A2(_00545_ ), .ZN(_00546_ ) );
AND2_X2 _16257_ ( .A1(_00542_ ), .A2(_00546_ ), .ZN(_00547_ ) );
INV_X1 _16258_ ( .A(_00547_ ), .ZN(_00548_ ) );
BUF_X4 _16259_ ( .A(_00548_ ), .Z(_00549_ ) );
AOI21_X1 _16260_ ( .A(_00541_ ), .B1(_00549_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_00550_ ) );
BUF_X2 _16261_ ( .A(_00548_ ), .Z(_00551_ ) );
OAI21_X1 _16262_ ( .A(_00550_ ), .B1(\myifu.data_in [8] ), .B2(_00551_ ), .ZN(_00552_ ) );
AND3_X1 _16263_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00553_ ) );
AND3_X1 _16264_ ( .A1(_05891_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00554_ ) );
AOI211_X1 _16265_ ( .A(_00553_ ), .B(_00554_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_05890_ ), .ZN(_00555_ ) );
NAND2_X1 _16266_ ( .A1(_00502_ ), .A2(\IF_ID_pc [2] ), .ZN(_00556_ ) );
BUF_X2 _16267_ ( .A(_00556_ ), .Z(_00557_ ) );
NAND2_X1 _16268_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00558_ ) );
BUF_X4 _16269_ ( .A(_00558_ ), .Z(_00559_ ) );
BUF_X4 _16270_ ( .A(_00559_ ), .Z(_00560_ ) );
NAND3_X1 _16271_ ( .A1(_03655_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00561_ ) );
NAND4_X1 _16272_ ( .A1(_00555_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00561_ ), .ZN(_00562_ ) );
NOR2_X1 _16273_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00563_ ) );
BUF_X4 _16274_ ( .A(_00563_ ), .Z(_00564_ ) );
BUF_X4 _16275_ ( .A(_00564_ ), .Z(_00565_ ) );
BUF_X4 _16276_ ( .A(_03636_ ), .Z(_00566_ ) );
BUF_X4 _16277_ ( .A(_00566_ ), .Z(_00567_ ) );
NAND3_X1 _16278_ ( .A1(_00567_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00568_ ) );
NAND3_X1 _16279_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00569_ ) );
AND2_X1 _16280_ ( .A1(_00568_ ), .A2(_00569_ ), .ZN(_00570_ ) );
NAND2_X1 _16281_ ( .A1(_00556_ ), .A2(_00558_ ), .ZN(_00571_ ) );
BUF_X2 _16282_ ( .A(_00571_ ), .Z(_00572_ ) );
BUF_X4 _16283_ ( .A(_03653_ ), .Z(_00573_ ) );
BUF_X4 _16284_ ( .A(_00573_ ), .Z(_00574_ ) );
BUF_X4 _16285_ ( .A(_00574_ ), .Z(_00575_ ) );
NAND3_X1 _16286_ ( .A1(_00575_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00576_ ) );
BUF_X4 _16287_ ( .A(_03654_ ), .Z(_00577_ ) );
NAND3_X1 _16288_ ( .A1(_05892_ ), .A2(_00577_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00578_ ) );
NAND4_X1 _16289_ ( .A1(_00570_ ), .A2(_00572_ ), .A3(_00576_ ), .A4(_00578_ ), .ZN(_00579_ ) );
NAND3_X1 _16290_ ( .A1(_00562_ ), .A2(_00565_ ), .A3(_00579_ ), .ZN(_00580_ ) );
NAND2_X1 _16291_ ( .A1(_00552_ ), .A2(_00580_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16292_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00581_ ) );
CLKBUF_X2 _16293_ ( .A(_03635_ ), .Z(_00582_ ) );
AND3_X1 _16294_ ( .A1(_00582_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00583_ ) );
BUF_X4 _16295_ ( .A(_05889_ ), .Z(_00584_ ) );
AOI211_X1 _16296_ ( .A(_00581_ ), .B(_00583_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00584_ ), .ZN(_00585_ ) );
BUF_X4 _16297_ ( .A(_00556_ ), .Z(_00586_ ) );
BUF_X4 _16298_ ( .A(_00586_ ), .Z(_00587_ ) );
BUF_X4 _16299_ ( .A(_00559_ ), .Z(_00588_ ) );
NAND3_X1 _16300_ ( .A1(_00577_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00589_ ) );
NAND4_X1 _16301_ ( .A1(_00585_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_00589_ ), .ZN(_00590_ ) );
BUF_X4 _16302_ ( .A(_00564_ ), .Z(_00591_ ) );
BUF_X4 _16303_ ( .A(_00566_ ), .Z(_00592_ ) );
NAND3_X1 _16304_ ( .A1(_00592_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00593_ ) );
NAND3_X1 _16305_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00594_ ) );
AND2_X1 _16306_ ( .A1(_00593_ ), .A2(_00594_ ), .ZN(_00595_ ) );
BUF_X4 _16307_ ( .A(_00571_ ), .Z(_00596_ ) );
BUF_X4 _16308_ ( .A(_00596_ ), .Z(_00597_ ) );
BUF_X4 _16309_ ( .A(_03653_ ), .Z(_00598_ ) );
BUF_X4 _16310_ ( .A(_00598_ ), .Z(_00599_ ) );
NAND3_X1 _16311_ ( .A1(_00599_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00600_ ) );
NAND3_X1 _16312_ ( .A1(_00567_ ), .A2(_00599_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00601_ ) );
NAND4_X1 _16313_ ( .A1(_00595_ ), .A2(_00597_ ), .A3(_00600_ ), .A4(_00601_ ), .ZN(_00602_ ) );
NAND3_X1 _16314_ ( .A1(_00590_ ), .A2(_00591_ ), .A3(_00602_ ), .ZN(_00603_ ) );
BUF_X4 _16315_ ( .A(_00542_ ), .Z(_00604_ ) );
INV_X1 _16316_ ( .A(_00604_ ), .ZN(_00605_ ) );
NOR4_X1 _16317_ ( .A1(\myifu.data_in [31] ), .A2(_00605_ ), .A3(_00545_ ), .A4(_00544_ ), .ZN(_00606_ ) );
OAI21_X1 _16318_ ( .A(\myifu.state [2] ), .B1(_00547_ ), .B2(_03419_ ), .ZN(_00607_ ) );
OAI21_X1 _16319_ ( .A(_00603_ ), .B1(_00606_ ), .B2(_00607_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
BUF_X4 _16320_ ( .A(_00604_ ), .Z(_00608_ ) );
BUF_X4 _16321_ ( .A(_00546_ ), .Z(_00609_ ) );
BUF_X4 _16322_ ( .A(_00609_ ), .Z(_00610_ ) );
AND2_X1 _16323_ ( .A1(_00399_ ), .A2(_00400_ ), .ZN(_00611_ ) );
OAI211_X1 _16324_ ( .A(_00608_ ), .B(_00610_ ), .C1(_00611_ ), .C2(_01993_ ), .ZN(_00612_ ) );
OAI211_X1 _16325_ ( .A(_00612_ ), .B(\myifu.state [2] ), .C1(_00547_ ), .C2(_03438_ ), .ZN(_00613_ ) );
AND3_X1 _16326_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00614_ ) );
AND3_X1 _16327_ ( .A1(_05891_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00615_ ) );
AOI211_X1 _16328_ ( .A(_00614_ ), .B(_00615_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_05890_ ), .ZN(_00616_ ) );
NAND3_X1 _16329_ ( .A1(_03655_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00617_ ) );
NAND4_X1 _16330_ ( .A1(_00616_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00617_ ), .ZN(_00618_ ) );
NAND3_X1 _16331_ ( .A1(_00567_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00619_ ) );
NAND3_X1 _16332_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00620_ ) );
AND2_X1 _16333_ ( .A1(_00619_ ), .A2(_00620_ ), .ZN(_00621_ ) );
NAND3_X1 _16334_ ( .A1(_00575_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00622_ ) );
NAND3_X1 _16335_ ( .A1(_05892_ ), .A2(_00577_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00623_ ) );
NAND4_X1 _16336_ ( .A1(_00621_ ), .A2(_00572_ ), .A3(_00622_ ), .A4(_00623_ ), .ZN(_00624_ ) );
NAND3_X1 _16337_ ( .A1(_00618_ ), .A2(_00565_ ), .A3(_00624_ ), .ZN(_00625_ ) );
NAND2_X1 _16338_ ( .A1(_00613_ ), .A2(_00625_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
NAND2_X1 _16339_ ( .A1(_00406_ ), .A2(_00409_ ), .ZN(_00626_ ) );
OAI211_X1 _16340_ ( .A(_00604_ ), .B(_00609_ ), .C1(_00626_ ), .C2(_05923_ ), .ZN(_00627_ ) );
NAND2_X1 _16341_ ( .A1(_00627_ ), .A2(\myifu.state [2] ), .ZN(_00628_ ) );
BUF_X4 _16342_ ( .A(_00548_ ), .Z(_00629_ ) );
AOI21_X1 _16343_ ( .A(_00628_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00629_ ), .ZN(_00630_ ) );
AND3_X1 _16344_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00631_ ) );
BUF_X4 _16345_ ( .A(_03635_ ), .Z(_00632_ ) );
AND3_X1 _16346_ ( .A1(_00632_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00633_ ) );
AOI211_X1 _16347_ ( .A(_00631_ ), .B(_00633_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_00584_ ), .ZN(_00634_ ) );
NAND3_X1 _16348_ ( .A1(_00574_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00635_ ) );
NAND4_X1 _16349_ ( .A1(_00634_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00635_ ), .ZN(_00636_ ) );
NAND3_X1 _16350_ ( .A1(_00566_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00637_ ) );
NAND3_X1 _16351_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00638_ ) );
AND2_X1 _16352_ ( .A1(_00637_ ), .A2(_00638_ ), .ZN(_00639_ ) );
NAND3_X1 _16353_ ( .A1(_00598_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00640_ ) );
BUF_X4 _16354_ ( .A(_00632_ ), .Z(_00641_ ) );
NAND3_X1 _16355_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00642_ ) );
NAND4_X1 _16356_ ( .A1(_00639_ ), .A2(_00596_ ), .A3(_00640_ ), .A4(_00642_ ), .ZN(_00643_ ) );
AND3_X1 _16357_ ( .A1(_00636_ ), .A2(_00564_ ), .A3(_00643_ ), .ZN(_00644_ ) );
OR2_X1 _16358_ ( .A1(_00630_ ), .A2(_00644_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
AND3_X1 _16359_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00645_ ) );
AND3_X1 _16360_ ( .A1(_00566_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00646_ ) );
AOI211_X1 _16361_ ( .A(_00645_ ), .B(_00646_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_00584_ ), .ZN(_00647_ ) );
NAND3_X1 _16362_ ( .A1(_00577_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00648_ ) );
NAND4_X1 _16363_ ( .A1(_00647_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_00648_ ), .ZN(_00649_ ) );
NAND3_X1 _16364_ ( .A1(_00592_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00650_ ) );
NAND3_X1 _16365_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00651_ ) );
AND2_X1 _16366_ ( .A1(_00650_ ), .A2(_00651_ ), .ZN(_00652_ ) );
NAND3_X1 _16367_ ( .A1(_00599_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00653_ ) );
NAND3_X1 _16368_ ( .A1(_00567_ ), .A2(_00574_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00654_ ) );
NAND4_X1 _16369_ ( .A1(_00652_ ), .A2(_00597_ ), .A3(_00653_ ), .A4(_00654_ ), .ZN(_00655_ ) );
NAND3_X1 _16370_ ( .A1(_00649_ ), .A2(_00591_ ), .A3(_00655_ ), .ZN(_00656_ ) );
AND2_X1 _16371_ ( .A1(_00551_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00657_ ) );
OAI21_X1 _16372_ ( .A(\myifu.state [2] ), .B1(_00551_ ), .B2(\myifu.data_in [20] ), .ZN(_00658_ ) );
OAI21_X1 _16373_ ( .A(_00656_ ), .B1(_00657_ ), .B2(_00658_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
AOI21_X1 _16374_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00659_ ) );
OAI211_X1 _16375_ ( .A(_00608_ ), .B(_00610_ ), .C1(_00415_ ), .C2(_05924_ ), .ZN(_00660_ ) );
NAND2_X1 _16376_ ( .A1(_00659_ ), .A2(_00660_ ), .ZN(_00661_ ) );
AND3_X1 _16377_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00662_ ) );
AND3_X1 _16378_ ( .A1(_05891_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00663_ ) );
AOI211_X1 _16379_ ( .A(_00662_ ), .B(_00663_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_05890_ ), .ZN(_00664_ ) );
NAND3_X1 _16380_ ( .A1(_03655_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00665_ ) );
NAND4_X1 _16381_ ( .A1(_00664_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00665_ ), .ZN(_00666_ ) );
BUF_X4 _16382_ ( .A(_00566_ ), .Z(_00667_ ) );
NAND3_X1 _16383_ ( .A1(_00667_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00668_ ) );
NAND3_X1 _16384_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00669_ ) );
AND2_X1 _16385_ ( .A1(_00668_ ), .A2(_00669_ ), .ZN(_00670_ ) );
NAND3_X1 _16386_ ( .A1(_00575_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00671_ ) );
NAND3_X1 _16387_ ( .A1(_05892_ ), .A2(_00577_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00672_ ) );
NAND4_X1 _16388_ ( .A1(_00670_ ), .A2(_00572_ ), .A3(_00671_ ), .A4(_00672_ ), .ZN(_00673_ ) );
NAND3_X1 _16389_ ( .A1(_00666_ ), .A2(_00565_ ), .A3(_00673_ ), .ZN(_00674_ ) );
NAND2_X1 _16390_ ( .A1(_00661_ ), .A2(_00674_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
AOI21_X1 _16391_ ( .A(_00540_ ), .B1(_00549_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00675_ ) );
OAI21_X1 _16392_ ( .A(_00675_ ), .B1(\myifu.data_in [18] ), .B2(_00551_ ), .ZN(_00676_ ) );
AND3_X1 _16393_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00677_ ) );
AND3_X1 _16394_ ( .A1(_05891_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00678_ ) );
AOI211_X1 _16395_ ( .A(_00677_ ), .B(_00678_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_05890_ ), .ZN(_00679_ ) );
NAND3_X1 _16396_ ( .A1(_03655_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00680_ ) );
NAND4_X1 _16397_ ( .A1(_00679_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00680_ ), .ZN(_00681_ ) );
NAND3_X1 _16398_ ( .A1(_00667_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00682_ ) );
NAND3_X1 _16399_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00683_ ) );
AND2_X1 _16400_ ( .A1(_00682_ ), .A2(_00683_ ), .ZN(_00684_ ) );
BUF_X4 _16401_ ( .A(_00596_ ), .Z(_00685_ ) );
NAND3_X1 _16402_ ( .A1(_00575_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00686_ ) );
NAND3_X1 _16403_ ( .A1(_05892_ ), .A2(_00577_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00687_ ) );
NAND4_X1 _16404_ ( .A1(_00684_ ), .A2(_00685_ ), .A3(_00686_ ), .A4(_00687_ ), .ZN(_00688_ ) );
NAND3_X1 _16405_ ( .A1(_00681_ ), .A2(_00565_ ), .A3(_00688_ ), .ZN(_00689_ ) );
NAND2_X1 _16406_ ( .A1(_00676_ ), .A2(_00689_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
OAI211_X1 _16407_ ( .A(_00604_ ), .B(_00609_ ), .C1(_05923_ ), .C2(_00422_ ), .ZN(_00690_ ) );
NAND2_X1 _16408_ ( .A1(_00690_ ), .A2(\myifu.state [2] ), .ZN(_00691_ ) );
AOI21_X1 _16409_ ( .A(_00691_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00549_ ), .ZN(_00692_ ) );
AND3_X1 _16410_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00693_ ) );
AND3_X1 _16411_ ( .A1(_00632_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00694_ ) );
AOI211_X1 _16412_ ( .A(_00693_ ), .B(_00694_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_00584_ ), .ZN(_00695_ ) );
NAND3_X1 _16413_ ( .A1(_00574_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00696_ ) );
NAND4_X1 _16414_ ( .A1(_00695_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00696_ ), .ZN(_00697_ ) );
NAND3_X1 _16415_ ( .A1(_00566_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00698_ ) );
NAND3_X1 _16416_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00699_ ) );
AND2_X1 _16417_ ( .A1(_00698_ ), .A2(_00699_ ), .ZN(_00700_ ) );
NAND3_X1 _16418_ ( .A1(_00598_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00701_ ) );
NAND3_X1 _16419_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00702_ ) );
NAND4_X1 _16420_ ( .A1(_00700_ ), .A2(_00596_ ), .A3(_00701_ ), .A4(_00702_ ), .ZN(_00703_ ) );
AND3_X1 _16421_ ( .A1(_00697_ ), .A2(_00564_ ), .A3(_00703_ ), .ZN(_00704_ ) );
OR2_X1 _16422_ ( .A1(_00692_ ), .A2(_00704_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NAND2_X1 _16423_ ( .A1(_00423_ ), .A2(_00425_ ), .ZN(_00705_ ) );
OAI211_X1 _16424_ ( .A(_00604_ ), .B(_00609_ ), .C1(_00705_ ), .C2(_05923_ ), .ZN(_00706_ ) );
NAND2_X1 _16425_ ( .A1(_00706_ ), .A2(\myifu.state [2] ), .ZN(_00707_ ) );
AOI21_X1 _16426_ ( .A(_00707_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00549_ ), .ZN(_00708_ ) );
AND3_X1 _16427_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00709_ ) );
AND3_X1 _16428_ ( .A1(_03636_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00710_ ) );
AOI211_X1 _16429_ ( .A(_00709_ ), .B(_00710_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_05889_ ), .ZN(_00711_ ) );
NAND3_X1 _16430_ ( .A1(_03654_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00712_ ) );
NAND4_X1 _16431_ ( .A1(_00711_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00712_ ), .ZN(_00713_ ) );
NAND3_X1 _16432_ ( .A1(_00632_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00714_ ) );
NAND3_X1 _16433_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00715_ ) );
AND2_X1 _16434_ ( .A1(_00714_ ), .A2(_00715_ ), .ZN(_00716_ ) );
NAND3_X1 _16435_ ( .A1(_00598_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00717_ ) );
NAND3_X1 _16436_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00718_ ) );
NAND4_X1 _16437_ ( .A1(_00716_ ), .A2(_00596_ ), .A3(_00717_ ), .A4(_00718_ ), .ZN(_00719_ ) );
AND3_X1 _16438_ ( .A1(_00713_ ), .A2(_00564_ ), .A3(_00719_ ), .ZN(_00720_ ) );
OR2_X1 _16439_ ( .A1(_00708_ ), .A2(_00720_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
OAI211_X1 _16440_ ( .A(_00604_ ), .B(_00609_ ), .C1(_05923_ ), .C2(_00428_ ), .ZN(_00721_ ) );
NAND2_X1 _16441_ ( .A1(_00721_ ), .A2(\myifu.state [2] ), .ZN(_00722_ ) );
AOI21_X1 _16442_ ( .A(_00722_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00549_ ), .ZN(_00723_ ) );
AND3_X1 _16443_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00724_ ) );
AND3_X1 _16444_ ( .A1(_03636_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00725_ ) );
AOI211_X1 _16445_ ( .A(_00724_ ), .B(_00725_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_05889_ ), .ZN(_00726_ ) );
NAND3_X1 _16446_ ( .A1(_03654_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00727_ ) );
NAND4_X1 _16447_ ( .A1(_00726_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00727_ ), .ZN(_00728_ ) );
NAND3_X1 _16448_ ( .A1(_00632_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00729_ ) );
NAND3_X1 _16449_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00730_ ) );
AND2_X1 _16450_ ( .A1(_00729_ ), .A2(_00730_ ), .ZN(_00731_ ) );
NAND3_X1 _16451_ ( .A1(_00598_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00732_ ) );
NAND3_X1 _16452_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00733_ ) );
NAND4_X1 _16453_ ( .A1(_00731_ ), .A2(_00596_ ), .A3(_00732_ ), .A4(_00733_ ), .ZN(_00734_ ) );
AND3_X1 _16454_ ( .A1(_00728_ ), .A2(_00564_ ), .A3(_00734_ ), .ZN(_00735_ ) );
OR2_X1 _16455_ ( .A1(_00723_ ), .A2(_00735_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
AOI21_X1 _16456_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00736_ ) );
NAND2_X1 _16457_ ( .A1(_00430_ ), .A2(_00432_ ), .ZN(_00737_ ) );
OAI211_X1 _16458_ ( .A(_00608_ ), .B(_00610_ ), .C1(_00737_ ), .C2(_05924_ ), .ZN(_00738_ ) );
NAND2_X1 _16459_ ( .A1(_00736_ ), .A2(_00738_ ), .ZN(_00739_ ) );
AND3_X1 _16460_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00740_ ) );
AND3_X1 _16461_ ( .A1(_05891_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00741_ ) );
AOI211_X1 _16462_ ( .A(_00740_ ), .B(_00741_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_05890_ ), .ZN(_00742_ ) );
BUF_X4 _16463_ ( .A(_00574_ ), .Z(_00743_ ) );
NAND3_X1 _16464_ ( .A1(_00743_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00744_ ) );
NAND4_X1 _16465_ ( .A1(_00742_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00744_ ), .ZN(_00745_ ) );
NAND3_X1 _16466_ ( .A1(_00667_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00746_ ) );
NAND3_X1 _16467_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00747_ ) );
AND2_X1 _16468_ ( .A1(_00746_ ), .A2(_00747_ ), .ZN(_00748_ ) );
NAND3_X1 _16469_ ( .A1(_00575_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00749_ ) );
BUF_X4 _16470_ ( .A(_03654_ ), .Z(_00750_ ) );
NAND3_X1 _16471_ ( .A1(_05892_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00751_ ) );
NAND4_X1 _16472_ ( .A1(_00748_ ), .A2(_00685_ ), .A3(_00749_ ), .A4(_00751_ ), .ZN(_00752_ ) );
NAND3_X1 _16473_ ( .A1(_00745_ ), .A2(_00565_ ), .A3(_00752_ ), .ZN(_00753_ ) );
NAND2_X1 _16474_ ( .A1(_00739_ ), .A2(_00753_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
NAND2_X1 _16475_ ( .A1(_00433_ ), .A2(_00435_ ), .ZN(_00754_ ) );
OAI211_X1 _16476_ ( .A(_00542_ ), .B(_00609_ ), .C1(_00754_ ), .C2(_05923_ ), .ZN(_00755_ ) );
NAND2_X1 _16477_ ( .A1(_00755_ ), .A2(\myifu.state [2] ), .ZN(_00756_ ) );
AOI21_X1 _16478_ ( .A(_00756_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00549_ ), .ZN(_00757_ ) );
AND3_X1 _16479_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00758_ ) );
AND3_X1 _16480_ ( .A1(_03636_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00759_ ) );
AOI211_X1 _16481_ ( .A(_00758_ ), .B(_00759_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_05889_ ), .ZN(_00760_ ) );
NAND3_X1 _16482_ ( .A1(_03654_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00761_ ) );
NAND4_X1 _16483_ ( .A1(_00760_ ), .A2(_00586_ ), .A3(_00558_ ), .A4(_00761_ ), .ZN(_00762_ ) );
NAND3_X1 _16484_ ( .A1(_00632_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00763_ ) );
NAND3_X1 _16485_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00764_ ) );
AND2_X1 _16486_ ( .A1(_00763_ ), .A2(_00764_ ), .ZN(_00765_ ) );
NAND3_X1 _16487_ ( .A1(_00598_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_00766_ ) );
NAND3_X1 _16488_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_00767_ ) );
NAND4_X1 _16489_ ( .A1(_00765_ ), .A2(_00596_ ), .A3(_00766_ ), .A4(_00767_ ), .ZN(_00768_ ) );
AND3_X1 _16490_ ( .A1(_00762_ ), .A2(_00564_ ), .A3(_00768_ ), .ZN(_00769_ ) );
OR2_X1 _16491_ ( .A1(_00757_ ), .A2(_00769_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
AND3_X1 _16492_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_00770_ ) );
AND3_X1 _16493_ ( .A1(_00566_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_00771_ ) );
AOI211_X1 _16494_ ( .A(_00770_ ), .B(_00771_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_00584_ ), .ZN(_00772_ ) );
NAND3_X1 _16495_ ( .A1(_00577_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_00773_ ) );
NAND4_X1 _16496_ ( .A1(_00772_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00773_ ), .ZN(_00774_ ) );
NAND3_X1 _16497_ ( .A1(_00592_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_00775_ ) );
NAND3_X1 _16498_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_00776_ ) );
AND2_X1 _16499_ ( .A1(_00775_ ), .A2(_00776_ ), .ZN(_00777_ ) );
NAND3_X1 _16500_ ( .A1(_00599_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_00778_ ) );
NAND3_X1 _16501_ ( .A1(_00567_ ), .A2(_00574_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_00779_ ) );
NAND4_X1 _16502_ ( .A1(_00777_ ), .A2(_00597_ ), .A3(_00778_ ), .A4(_00779_ ), .ZN(_00780_ ) );
NAND3_X1 _16503_ ( .A1(_00774_ ), .A2(_00591_ ), .A3(_00780_ ), .ZN(_00781_ ) );
AND2_X1 _16504_ ( .A1(_00551_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00782_ ) );
OAI21_X1 _16505_ ( .A(\myifu.state [2] ), .B1(_00551_ ), .B2(\myifu.data_in [12] ), .ZN(_00783_ ) );
OAI21_X1 _16506_ ( .A(_00781_ ), .B1(_00782_ ), .B2(_00783_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
AND2_X1 _16507_ ( .A1(_00440_ ), .A2(_00441_ ), .ZN(_00784_ ) );
OAI211_X1 _16508_ ( .A(_00608_ ), .B(_00610_ ), .C1(_00784_ ), .C2(_01993_ ), .ZN(_00785_ ) );
OAI211_X1 _16509_ ( .A(_00785_ ), .B(\myifu.state [2] ), .C1(_00547_ ), .C2(_03434_ ), .ZN(_00786_ ) );
AND3_X1 _16510_ ( .A1(fanout_net_14 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_00787_ ) );
AND3_X1 _16511_ ( .A1(_05891_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_00788_ ) );
AOI211_X1 _16512_ ( .A(_00787_ ), .B(_00788_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_05890_ ), .ZN(_00789_ ) );
NAND3_X1 _16513_ ( .A1(_00743_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_00790_ ) );
NAND4_X1 _16514_ ( .A1(_00789_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00790_ ), .ZN(_00791_ ) );
NAND3_X1 _16515_ ( .A1(_00667_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_00792_ ) );
NAND3_X1 _16516_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_00793_ ) );
AND2_X1 _16517_ ( .A1(_00792_ ), .A2(_00793_ ), .ZN(_00794_ ) );
NAND3_X1 _16518_ ( .A1(_00575_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_00795_ ) );
BUF_X4 _16519_ ( .A(_00641_ ), .Z(_00796_ ) );
NAND3_X1 _16520_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_00797_ ) );
NAND4_X1 _16521_ ( .A1(_00794_ ), .A2(_00685_ ), .A3(_00795_ ), .A4(_00797_ ), .ZN(_00798_ ) );
NAND3_X1 _16522_ ( .A1(_00791_ ), .A2(_00565_ ), .A3(_00798_ ), .ZN(_00799_ ) );
NAND2_X1 _16523_ ( .A1(_00786_ ), .A2(_00799_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
OR2_X1 _16524_ ( .A1(_00548_ ), .A2(\myifu.data_in [11] ), .ZN(_00800_ ) );
AOI21_X1 _16525_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_00801_ ) );
NAND2_X1 _16526_ ( .A1(_00800_ ), .A2(_00801_ ), .ZN(_00802_ ) );
AND3_X1 _16527_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_00803_ ) );
AND3_X1 _16528_ ( .A1(_05891_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_00804_ ) );
BUF_X4 _16529_ ( .A(_00584_ ), .Z(_00805_ ) );
AOI211_X1 _16530_ ( .A(_00803_ ), .B(_00804_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_00805_ ), .ZN(_00806_ ) );
NAND3_X1 _16531_ ( .A1(_00743_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_00807_ ) );
NAND4_X1 _16532_ ( .A1(_00806_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00807_ ), .ZN(_00808_ ) );
NAND3_X1 _16533_ ( .A1(_00667_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_00809_ ) );
NAND3_X1 _16534_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_00810_ ) );
AND2_X1 _16535_ ( .A1(_00809_ ), .A2(_00810_ ), .ZN(_00811_ ) );
NAND3_X1 _16536_ ( .A1(_00575_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_00812_ ) );
NAND3_X1 _16537_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_00813_ ) );
NAND4_X1 _16538_ ( .A1(_00811_ ), .A2(_00685_ ), .A3(_00812_ ), .A4(_00813_ ), .ZN(_00814_ ) );
NAND3_X1 _16539_ ( .A1(_00808_ ), .A2(_00565_ ), .A3(_00814_ ), .ZN(_00815_ ) );
NAND2_X1 _16540_ ( .A1(_00802_ ), .A2(_00815_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
AND3_X1 _16541_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_00816_ ) );
AND3_X1 _16542_ ( .A1(_00566_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_00817_ ) );
AOI211_X1 _16543_ ( .A(_00816_ ), .B(_00817_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_00584_ ), .ZN(_00818_ ) );
NAND3_X1 _16544_ ( .A1(_00577_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_00819_ ) );
NAND4_X1 _16545_ ( .A1(_00818_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00819_ ), .ZN(_00820_ ) );
NAND3_X1 _16546_ ( .A1(_00592_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_00821_ ) );
NAND3_X1 _16547_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_00822_ ) );
AND2_X1 _16548_ ( .A1(_00821_ ), .A2(_00822_ ), .ZN(_00823_ ) );
NAND3_X1 _16549_ ( .A1(_00599_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_00824_ ) );
NAND3_X1 _16550_ ( .A1(_00567_ ), .A2(_00574_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_00825_ ) );
NAND4_X1 _16551_ ( .A1(_00823_ ), .A2(_00597_ ), .A3(_00824_ ), .A4(_00825_ ), .ZN(_00826_ ) );
NAND3_X1 _16552_ ( .A1(_00820_ ), .A2(_00564_ ), .A3(_00826_ ), .ZN(_00827_ ) );
NOR4_X1 _16553_ ( .A1(_00605_ ), .A2(\myifu.data_in [10] ), .A3(_00545_ ), .A4(_00544_ ), .ZN(_00828_ ) );
OAI21_X1 _16554_ ( .A(\myifu.state [2] ), .B1(_00547_ ), .B2(_03377_ ), .ZN(_00829_ ) );
OAI21_X1 _16555_ ( .A(_00827_ ), .B1(_00828_ ), .B2(_00829_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
AND3_X1 _16556_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_00830_ ) );
AND3_X1 _16557_ ( .A1(_00566_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_00831_ ) );
AOI211_X1 _16558_ ( .A(_00830_ ), .B(_00831_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_00584_ ), .ZN(_00832_ ) );
NAND3_X1 _16559_ ( .A1(_00577_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_00833_ ) );
NAND4_X1 _16560_ ( .A1(_00832_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00833_ ), .ZN(_00834_ ) );
NAND3_X1 _16561_ ( .A1(_00592_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_00835_ ) );
NAND3_X1 _16562_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_00836_ ) );
AND2_X1 _16563_ ( .A1(_00835_ ), .A2(_00836_ ), .ZN(_00837_ ) );
NAND3_X1 _16564_ ( .A1(_00599_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_00838_ ) );
NAND3_X1 _16565_ ( .A1(_00567_ ), .A2(_00574_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_00839_ ) );
NAND4_X1 _16566_ ( .A1(_00837_ ), .A2(_00597_ ), .A3(_00838_ ), .A4(_00839_ ), .ZN(_00840_ ) );
NAND3_X1 _16567_ ( .A1(_00834_ ), .A2(_00564_ ), .A3(_00840_ ), .ZN(_00841_ ) );
AND2_X1 _16568_ ( .A1(_00551_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_00842_ ) );
OAI21_X1 _16569_ ( .A(\myifu.state [2] ), .B1(_00551_ ), .B2(\myifu.data_in [9] ), .ZN(_00843_ ) );
OAI21_X1 _16570_ ( .A(_00841_ ), .B1(_00842_ ), .B2(_00843_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
OAI211_X1 _16571_ ( .A(_00542_ ), .B(_00546_ ), .C1(_00456_ ), .C2(_05923_ ), .ZN(_00844_ ) );
NAND2_X1 _16572_ ( .A1(_00844_ ), .A2(\myifu.state [2] ), .ZN(_00845_ ) );
AOI21_X1 _16573_ ( .A(_00845_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_00549_ ), .ZN(_00846_ ) );
AND3_X1 _16574_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_00847_ ) );
AND3_X1 _16575_ ( .A1(_03636_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_00848_ ) );
AOI211_X1 _16576_ ( .A(_00847_ ), .B(_00848_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_05889_ ), .ZN(_00849_ ) );
NAND3_X1 _16577_ ( .A1(_03654_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_00850_ ) );
NAND4_X1 _16578_ ( .A1(_00849_ ), .A2(_00556_ ), .A3(_00558_ ), .A4(_00850_ ), .ZN(_00851_ ) );
NAND3_X1 _16579_ ( .A1(_00632_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_00852_ ) );
NAND3_X1 _16580_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_00853_ ) );
AND2_X1 _16581_ ( .A1(_00852_ ), .A2(_00853_ ), .ZN(_00854_ ) );
NAND3_X1 _16582_ ( .A1(_00598_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_00855_ ) );
NAND3_X1 _16583_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_00856_ ) );
NAND4_X1 _16584_ ( .A1(_00854_ ), .A2(_00596_ ), .A3(_00855_ ), .A4(_00856_ ), .ZN(_00857_ ) );
AND3_X1 _16585_ ( .A1(_00851_ ), .A2(_00563_ ), .A3(_00857_ ), .ZN(_00858_ ) );
OR2_X1 _16586_ ( .A1(_00846_ ), .A2(_00858_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AOI21_X1 _16587_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00859_ ) );
OAI211_X1 _16588_ ( .A(_00608_ ), .B(_00610_ ), .C1(_05924_ ), .C2(_00459_ ), .ZN(_00860_ ) );
NAND2_X1 _16589_ ( .A1(_00859_ ), .A2(_00860_ ), .ZN(_00861_ ) );
AND3_X1 _16590_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_00862_ ) );
AND3_X1 _16591_ ( .A1(_05891_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_00863_ ) );
AOI211_X1 _16592_ ( .A(_00862_ ), .B(_00863_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00805_ ), .ZN(_00864_ ) );
NAND3_X1 _16593_ ( .A1(_00743_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_00865_ ) );
NAND4_X1 _16594_ ( .A1(_00864_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00865_ ), .ZN(_00866_ ) );
NAND3_X1 _16595_ ( .A1(_00667_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_00867_ ) );
NAND3_X1 _16596_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_00868_ ) );
AND2_X1 _16597_ ( .A1(_00867_ ), .A2(_00868_ ), .ZN(_00869_ ) );
BUF_X4 _16598_ ( .A(_00574_ ), .Z(_00870_ ) );
NAND3_X1 _16599_ ( .A1(_00870_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_00871_ ) );
NAND3_X1 _16600_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_00872_ ) );
NAND4_X1 _16601_ ( .A1(_00869_ ), .A2(_00685_ ), .A3(_00871_ ), .A4(_00872_ ), .ZN(_00873_ ) );
NAND3_X1 _16602_ ( .A1(_00866_ ), .A2(_00565_ ), .A3(_00873_ ), .ZN(_00874_ ) );
NAND2_X1 _16603_ ( .A1(_00861_ ), .A2(_00874_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
AOI21_X1 _16604_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00875_ ) );
OAI211_X1 _16605_ ( .A(_00608_ ), .B(_00610_ ), .C1(_00462_ ), .C2(_05924_ ), .ZN(_00876_ ) );
NAND2_X1 _16606_ ( .A1(_00875_ ), .A2(_00876_ ), .ZN(_00877_ ) );
AND3_X1 _16607_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_00878_ ) );
AND3_X1 _16608_ ( .A1(_00582_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_00879_ ) );
AOI211_X1 _16609_ ( .A(_00878_ ), .B(_00879_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00805_ ), .ZN(_00880_ ) );
NAND3_X1 _16610_ ( .A1(_00743_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_00881_ ) );
NAND4_X1 _16611_ ( .A1(_00880_ ), .A2(_00557_ ), .A3(_00560_ ), .A4(_00881_ ), .ZN(_00882_ ) );
NAND3_X1 _16612_ ( .A1(_00667_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_00883_ ) );
NAND3_X1 _16613_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_00884_ ) );
AND2_X1 _16614_ ( .A1(_00883_ ), .A2(_00884_ ), .ZN(_00885_ ) );
NAND3_X1 _16615_ ( .A1(_00870_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_00886_ ) );
NAND3_X1 _16616_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_00887_ ) );
NAND4_X1 _16617_ ( .A1(_00885_ ), .A2(_00685_ ), .A3(_00886_ ), .A4(_00887_ ), .ZN(_00888_ ) );
NAND3_X1 _16618_ ( .A1(_00882_ ), .A2(_00565_ ), .A3(_00888_ ), .ZN(_00889_ ) );
NAND2_X1 _16619_ ( .A1(_00877_ ), .A2(_00889_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
AND3_X1 _16620_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_00890_ ) );
AND3_X1 _16621_ ( .A1(_00566_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_00891_ ) );
AOI211_X1 _16622_ ( .A(_00890_ ), .B(_00891_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00584_ ), .ZN(_00892_ ) );
NAND3_X1 _16623_ ( .A1(_00577_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_00893_ ) );
NAND4_X1 _16624_ ( .A1(_00892_ ), .A2(_00586_ ), .A3(_00559_ ), .A4(_00893_ ), .ZN(_00894_ ) );
NAND3_X1 _16625_ ( .A1(_00641_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_00895_ ) );
NAND3_X1 _16626_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_00896_ ) );
AND2_X1 _16627_ ( .A1(_00895_ ), .A2(_00896_ ), .ZN(_00897_ ) );
NAND3_X1 _16628_ ( .A1(_00599_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_00898_ ) );
NAND3_X1 _16629_ ( .A1(_00567_ ), .A2(_00574_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_00899_ ) );
NAND4_X1 _16630_ ( .A1(_00897_ ), .A2(_00597_ ), .A3(_00898_ ), .A4(_00899_ ), .ZN(_00900_ ) );
NAND3_X1 _16631_ ( .A1(_00894_ ), .A2(_00564_ ), .A3(_00900_ ), .ZN(_00901_ ) );
AND2_X1 _16632_ ( .A1(_00551_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00902_ ) );
OAI21_X1 _16633_ ( .A(\myifu.state [2] ), .B1(_00551_ ), .B2(\myifu.data_in [4] ), .ZN(_00903_ ) );
OAI21_X1 _16634_ ( .A(_00901_ ), .B1(_00902_ ), .B2(_00903_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _16635_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00904_ ) );
OAI211_X1 _16636_ ( .A(_00608_ ), .B(_00610_ ), .C1(_00469_ ), .C2(_05924_ ), .ZN(_00905_ ) );
NAND2_X1 _16637_ ( .A1(_00904_ ), .A2(_00905_ ), .ZN(_00906_ ) );
AND3_X1 _16638_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_00907_ ) );
AND3_X1 _16639_ ( .A1(_00582_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_00908_ ) );
AOI211_X1 _16640_ ( .A(_00907_ ), .B(_00908_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00805_ ), .ZN(_00909_ ) );
NAND3_X1 _16641_ ( .A1(_00743_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_00910_ ) );
NAND4_X1 _16642_ ( .A1(_00909_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_00910_ ), .ZN(_00911_ ) );
NAND3_X1 _16643_ ( .A1(_00667_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_00912_ ) );
NAND3_X1 _16644_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_00913_ ) );
AND2_X1 _16645_ ( .A1(_00912_ ), .A2(_00913_ ), .ZN(_00914_ ) );
NAND3_X1 _16646_ ( .A1(_00870_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_00915_ ) );
NAND3_X1 _16647_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_00916_ ) );
NAND4_X1 _16648_ ( .A1(_00914_ ), .A2(_00685_ ), .A3(_00915_ ), .A4(_00916_ ), .ZN(_00917_ ) );
NAND3_X1 _16649_ ( .A1(_00911_ ), .A2(_00565_ ), .A3(_00917_ ), .ZN(_00918_ ) );
NAND2_X1 _16650_ ( .A1(_00906_ ), .A2(_00918_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
OAI211_X1 _16651_ ( .A(_00542_ ), .B(_00546_ ), .C1(_05923_ ), .C2(_00472_ ), .ZN(_00919_ ) );
NAND2_X1 _16652_ ( .A1(_00919_ ), .A2(\myifu.state [2] ), .ZN(_00920_ ) );
AOI21_X1 _16653_ ( .A(_00920_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00549_ ), .ZN(_00921_ ) );
AND3_X1 _16654_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_00922_ ) );
AND3_X1 _16655_ ( .A1(_03636_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_00923_ ) );
AOI211_X1 _16656_ ( .A(_00922_ ), .B(_00923_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_05889_ ), .ZN(_00924_ ) );
NAND3_X1 _16657_ ( .A1(_03654_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_00925_ ) );
NAND4_X1 _16658_ ( .A1(_00924_ ), .A2(_00556_ ), .A3(_00558_ ), .A4(_00925_ ), .ZN(_00926_ ) );
NAND3_X1 _16659_ ( .A1(_00632_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_00927_ ) );
NAND3_X1 _16660_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_00928_ ) );
AND2_X1 _16661_ ( .A1(_00927_ ), .A2(_00928_ ), .ZN(_00929_ ) );
NAND3_X1 _16662_ ( .A1(_00598_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_00930_ ) );
NAND3_X1 _16663_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_00931_ ) );
NAND4_X1 _16664_ ( .A1(_00929_ ), .A2(_00596_ ), .A3(_00930_ ), .A4(_00931_ ), .ZN(_00932_ ) );
AND3_X1 _16665_ ( .A1(_00926_ ), .A2(_00563_ ), .A3(_00932_ ), .ZN(_00933_ ) );
OR2_X1 _16666_ ( .A1(_00921_ ), .A2(_00933_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
OAI211_X1 _16667_ ( .A(_00542_ ), .B(_00546_ ), .C1(_00478_ ), .C2(_05923_ ), .ZN(_00934_ ) );
NAND2_X1 _16668_ ( .A1(_00934_ ), .A2(\myifu.state [2] ), .ZN(_00935_ ) );
AOI21_X1 _16669_ ( .A(_00935_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00549_ ), .ZN(_00936_ ) );
AND3_X1 _16670_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_00937_ ) );
AND3_X1 _16671_ ( .A1(_03636_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_00938_ ) );
AOI211_X1 _16672_ ( .A(_00937_ ), .B(_00938_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_05889_ ), .ZN(_00939_ ) );
NAND3_X1 _16673_ ( .A1(_03654_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_00940_ ) );
NAND4_X1 _16674_ ( .A1(_00939_ ), .A2(_00556_ ), .A3(_00558_ ), .A4(_00940_ ), .ZN(_00941_ ) );
NAND3_X1 _16675_ ( .A1(_00632_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_00942_ ) );
NAND3_X1 _16676_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_00943_ ) );
AND2_X1 _16677_ ( .A1(_00942_ ), .A2(_00943_ ), .ZN(_00944_ ) );
NAND3_X1 _16678_ ( .A1(_00598_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_00945_ ) );
NAND3_X1 _16679_ ( .A1(_00641_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_00946_ ) );
NAND4_X1 _16680_ ( .A1(_00944_ ), .A2(_00596_ ), .A3(_00945_ ), .A4(_00946_ ), .ZN(_00947_ ) );
AND3_X1 _16681_ ( .A1(_00941_ ), .A2(_00563_ ), .A3(_00947_ ), .ZN(_00948_ ) );
OR2_X1 _16682_ ( .A1(_00936_ ), .A2(_00948_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
OAI211_X1 _16683_ ( .A(_00604_ ), .B(_00609_ ), .C1(_01993_ ), .C2(_00475_ ), .ZN(_00949_ ) );
OAI211_X1 _16684_ ( .A(_00949_ ), .B(\myifu.state [2] ), .C1(_00547_ ), .C2(_03409_ ), .ZN(_00950_ ) );
AND3_X1 _16685_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_00951_ ) );
AND3_X1 _16686_ ( .A1(_00582_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_00952_ ) );
AOI211_X1 _16687_ ( .A(_00951_ ), .B(_00952_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00805_ ), .ZN(_00953_ ) );
NAND3_X1 _16688_ ( .A1(_00743_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_00954_ ) );
NAND4_X1 _16689_ ( .A1(_00953_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_00954_ ), .ZN(_00955_ ) );
NAND3_X1 _16690_ ( .A1(_00667_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_00956_ ) );
NAND3_X1 _16691_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_00957_ ) );
AND2_X1 _16692_ ( .A1(_00956_ ), .A2(_00957_ ), .ZN(_00958_ ) );
NAND3_X1 _16693_ ( .A1(_00870_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_00959_ ) );
NAND3_X1 _16694_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_00960_ ) );
NAND4_X1 _16695_ ( .A1(_00958_ ), .A2(_00685_ ), .A3(_00959_ ), .A4(_00960_ ), .ZN(_00961_ ) );
NAND3_X1 _16696_ ( .A1(_00955_ ), .A2(_00591_ ), .A3(_00961_ ), .ZN(_00962_ ) );
NAND2_X1 _16697_ ( .A1(_00950_ ), .A2(_00962_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
OAI211_X1 _16698_ ( .A(_00542_ ), .B(_00546_ ), .C1(_05923_ ), .C2(_00481_ ), .ZN(_00963_ ) );
NAND2_X1 _16699_ ( .A1(_00963_ ), .A2(\myifu.state [2] ), .ZN(_00964_ ) );
AOI21_X1 _16700_ ( .A(_00964_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00549_ ), .ZN(_00965_ ) );
AND3_X1 _16701_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_00966_ ) );
AND3_X1 _16702_ ( .A1(_03636_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_00967_ ) );
AOI211_X1 _16703_ ( .A(_00966_ ), .B(_00967_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_05889_ ), .ZN(_00968_ ) );
NAND3_X1 _16704_ ( .A1(_03654_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_00969_ ) );
NAND4_X1 _16705_ ( .A1(_00968_ ), .A2(_00556_ ), .A3(_00558_ ), .A4(_00969_ ), .ZN(_00970_ ) );
NAND3_X1 _16706_ ( .A1(_00632_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_00971_ ) );
NAND3_X1 _16707_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_00972_ ) );
AND2_X1 _16708_ ( .A1(_00971_ ), .A2(_00972_ ), .ZN(_00973_ ) );
NAND3_X1 _16709_ ( .A1(_00598_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_00974_ ) );
NAND3_X1 _16710_ ( .A1(_05891_ ), .A2(_00573_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_00975_ ) );
NAND4_X1 _16711_ ( .A1(_00973_ ), .A2(_00571_ ), .A3(_00974_ ), .A4(_00975_ ), .ZN(_00976_ ) );
AND3_X1 _16712_ ( .A1(_00970_ ), .A2(_00563_ ), .A3(_00976_ ), .ZN(_00977_ ) );
OR2_X1 _16713_ ( .A1(_00965_ ), .A2(_00977_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
OAI211_X1 _16714_ ( .A(_00604_ ), .B(_00609_ ), .C1(_01993_ ), .C2(_00484_ ), .ZN(_00978_ ) );
OAI211_X1 _16715_ ( .A(_00978_ ), .B(\myifu.state [2] ), .C1(_00547_ ), .C2(_03399_ ), .ZN(_00979_ ) );
AND3_X1 _16716_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_00980_ ) );
AND3_X1 _16717_ ( .A1(_00582_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_00981_ ) );
AOI211_X1 _16718_ ( .A(_00980_ ), .B(_00981_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00805_ ), .ZN(_00982_ ) );
NAND3_X1 _16719_ ( .A1(_00743_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_00983_ ) );
NAND4_X1 _16720_ ( .A1(_00982_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_00983_ ), .ZN(_00984_ ) );
NAND3_X1 _16721_ ( .A1(_00667_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_00985_ ) );
NAND3_X1 _16722_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_00986_ ) );
AND2_X1 _16723_ ( .A1(_00985_ ), .A2(_00986_ ), .ZN(_00987_ ) );
NAND3_X1 _16724_ ( .A1(_00870_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_00988_ ) );
NAND3_X1 _16725_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_00989_ ) );
NAND4_X1 _16726_ ( .A1(_00987_ ), .A2(_00685_ ), .A3(_00988_ ), .A4(_00989_ ), .ZN(_00990_ ) );
NAND3_X1 _16727_ ( .A1(_00984_ ), .A2(_00591_ ), .A3(_00990_ ), .ZN(_00991_ ) );
NAND2_X1 _16728_ ( .A1(_00979_ ), .A2(_00991_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
OAI211_X1 _16729_ ( .A(_00604_ ), .B(_00609_ ), .C1(_01993_ ), .C2(_00487_ ), .ZN(_00992_ ) );
OAI211_X1 _16730_ ( .A(_00992_ ), .B(\myifu.state [2] ), .C1(_00547_ ), .C2(_03395_ ), .ZN(_00993_ ) );
AND3_X1 _16731_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_00994_ ) );
AND3_X1 _16732_ ( .A1(_00582_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_00995_ ) );
AOI211_X1 _16733_ ( .A(_00994_ ), .B(_00995_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_00805_ ), .ZN(_00996_ ) );
NAND3_X1 _16734_ ( .A1(_00743_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_00997_ ) );
NAND4_X1 _16735_ ( .A1(_00996_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_00997_ ), .ZN(_00998_ ) );
NAND3_X1 _16736_ ( .A1(_00592_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_00999_ ) );
NAND3_X1 _16737_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01000_ ) );
AND2_X1 _16738_ ( .A1(_00999_ ), .A2(_01000_ ), .ZN(_01001_ ) );
NAND3_X1 _16739_ ( .A1(_00870_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01002_ ) );
NAND3_X1 _16740_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01003_ ) );
NAND4_X1 _16741_ ( .A1(_01001_ ), .A2(_00685_ ), .A3(_01002_ ), .A4(_01003_ ), .ZN(_01004_ ) );
NAND3_X1 _16742_ ( .A1(_00998_ ), .A2(_00591_ ), .A3(_01004_ ), .ZN(_01005_ ) );
NAND2_X1 _16743_ ( .A1(_00993_ ), .A2(_01005_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
OAI211_X1 _16744_ ( .A(_00604_ ), .B(_00609_ ), .C1(_01993_ ), .C2(_00490_ ), .ZN(_01006_ ) );
OAI211_X1 _16745_ ( .A(_01006_ ), .B(\myifu.state [2] ), .C1(_00547_ ), .C2(_03387_ ), .ZN(_01007_ ) );
AND3_X1 _16746_ ( .A1(\IF_ID_pc [4] ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01008_ ) );
AND3_X1 _16747_ ( .A1(_00582_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01009_ ) );
AOI211_X1 _16748_ ( .A(_01008_ ), .B(_01009_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00805_ ), .ZN(_01010_ ) );
NAND3_X1 _16749_ ( .A1(_00743_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01011_ ) );
NAND4_X1 _16750_ ( .A1(_01010_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_01011_ ), .ZN(_01012_ ) );
NAND3_X1 _16751_ ( .A1(_00592_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01013_ ) );
NAND3_X1 _16752_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01014_ ) );
AND2_X1 _16753_ ( .A1(_01013_ ), .A2(_01014_ ), .ZN(_01015_ ) );
NAND3_X1 _16754_ ( .A1(_00870_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01016_ ) );
NAND3_X1 _16755_ ( .A1(_00796_ ), .A2(_00750_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01017_ ) );
NAND4_X1 _16756_ ( .A1(_01015_ ), .A2(_00597_ ), .A3(_01016_ ), .A4(_01017_ ), .ZN(_01018_ ) );
NAND3_X1 _16757_ ( .A1(_01012_ ), .A2(_00591_ ), .A3(_01018_ ), .ZN(_01019_ ) );
NAND2_X1 _16758_ ( .A1(_01007_ ), .A2(_01019_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
AOI21_X1 _16759_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01020_ ) );
NAND2_X1 _16760_ ( .A1(_00491_ ), .A2(_00493_ ), .ZN(_01021_ ) );
OAI211_X1 _16761_ ( .A(_00608_ ), .B(_00610_ ), .C1(_01021_ ), .C2(_05924_ ), .ZN(_01022_ ) );
NAND2_X1 _16762_ ( .A1(_01020_ ), .A2(_01022_ ), .ZN(_01023_ ) );
AND3_X1 _16763_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01024_ ) );
AND3_X1 _16764_ ( .A1(_00582_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01025_ ) );
AOI211_X1 _16765_ ( .A(_01024_ ), .B(_01025_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_00805_ ), .ZN(_01026_ ) );
NAND3_X1 _16766_ ( .A1(_00575_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01027_ ) );
NAND4_X1 _16767_ ( .A1(_01026_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_01027_ ), .ZN(_01028_ ) );
NAND3_X1 _16768_ ( .A1(_00592_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01029_ ) );
NAND3_X1 _16769_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01030_ ) );
AND2_X1 _16770_ ( .A1(_01029_ ), .A2(_01030_ ), .ZN(_01031_ ) );
NAND3_X1 _16771_ ( .A1(_00870_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01032_ ) );
NAND3_X1 _16772_ ( .A1(_00796_ ), .A2(_00599_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01033_ ) );
NAND4_X1 _16773_ ( .A1(_01031_ ), .A2(_00597_ ), .A3(_01032_ ), .A4(_01033_ ), .ZN(_01034_ ) );
NAND3_X1 _16774_ ( .A1(_01028_ ), .A2(_00591_ ), .A3(_01034_ ), .ZN(_01035_ ) );
NAND2_X1 _16775_ ( .A1(_01023_ ), .A2(_01035_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
AOI21_X1 _16776_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01036_ ) );
OAI211_X1 _16777_ ( .A(_00608_ ), .B(_00610_ ), .C1(_00496_ ), .C2(_05924_ ), .ZN(_01037_ ) );
NAND2_X1 _16778_ ( .A1(_01036_ ), .A2(_01037_ ), .ZN(_01038_ ) );
AND3_X1 _16779_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01039_ ) );
AND3_X1 _16780_ ( .A1(_00582_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01040_ ) );
AOI211_X1 _16781_ ( .A(_01039_ ), .B(_01040_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_00805_ ), .ZN(_01041_ ) );
NAND3_X1 _16782_ ( .A1(_00575_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01042_ ) );
NAND4_X1 _16783_ ( .A1(_01041_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_01042_ ), .ZN(_01043_ ) );
NAND3_X1 _16784_ ( .A1(_00592_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01044_ ) );
NAND3_X1 _16785_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01045_ ) );
AND2_X1 _16786_ ( .A1(_01044_ ), .A2(_01045_ ), .ZN(_01046_ ) );
NAND3_X1 _16787_ ( .A1(_00870_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01047_ ) );
NAND3_X1 _16788_ ( .A1(_00567_ ), .A2(_00599_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01048_ ) );
NAND4_X1 _16789_ ( .A1(_01046_ ), .A2(_00597_ ), .A3(_01047_ ), .A4(_01048_ ), .ZN(_01049_ ) );
NAND3_X1 _16790_ ( .A1(_01043_ ), .A2(_00591_ ), .A3(_01049_ ), .ZN(_01050_ ) );
NAND2_X1 _16791_ ( .A1(_01038_ ), .A2(_01050_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
AOI21_X1 _16792_ ( .A(_00541_ ), .B1(_00629_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_01051_ ) );
NAND2_X1 _16793_ ( .A1(_00497_ ), .A2(_00499_ ), .ZN(_01052_ ) );
OAI211_X1 _16794_ ( .A(_00608_ ), .B(_00610_ ), .C1(_01052_ ), .C2(_05924_ ), .ZN(_01053_ ) );
NAND2_X1 _16795_ ( .A1(_01051_ ), .A2(_01053_ ), .ZN(_01054_ ) );
AND3_X1 _16796_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01055_ ) );
AND3_X1 _16797_ ( .A1(_00582_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01056_ ) );
AOI211_X1 _16798_ ( .A(_01055_ ), .B(_01056_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_00584_ ), .ZN(_01057_ ) );
NAND3_X1 _16799_ ( .A1(_00575_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01058_ ) );
NAND4_X1 _16800_ ( .A1(_01057_ ), .A2(_00587_ ), .A3(_00588_ ), .A4(_01058_ ), .ZN(_01059_ ) );
NAND3_X1 _16801_ ( .A1(_00592_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01060_ ) );
NAND3_X1 _16802_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01061_ ) );
AND2_X1 _16803_ ( .A1(_01060_ ), .A2(_01061_ ), .ZN(_01062_ ) );
NAND3_X1 _16804_ ( .A1(_00870_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01063_ ) );
NAND3_X1 _16805_ ( .A1(_00567_ ), .A2(_00599_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01064_ ) );
NAND4_X1 _16806_ ( .A1(_01062_ ), .A2(_00597_ ), .A3(_01063_ ), .A4(_01064_ ), .ZN(_01065_ ) );
NAND3_X1 _16807_ ( .A1(_01059_ ), .A2(_00591_ ), .A3(_01065_ ), .ZN(_01066_ ) );
NAND2_X1 _16808_ ( .A1(_01054_ ), .A2(_01066_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI21_X1 _16809_ ( .A(_03656_ ), .B1(_03546_ ), .B2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _16810_ ( .A1(_03713_ ), .A2(_03716_ ), .A3(_03725_ ), .A4(\myifu.state [2] ), .ZN(_01067_ ) );
INV_X1 _16811_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01068_ ) );
AND4_X1 _16812_ ( .A1(_01068_ ), .A2(_01797_ ), .A3(\myifu.state [0] ), .A4(_01863_ ), .ZN(_01069_ ) );
NOR2_X1 _16813_ ( .A1(_01069_ ), .A2(_00390_ ), .ZN(_01070_ ) );
AOI21_X1 _16814_ ( .A(reset ), .B1(_01067_ ), .B2(_01070_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _16815_ ( .A1(_05873_ ), .A2(_01883_ ), .ZN(_01071_ ) );
INV_X1 _16816_ ( .A(_01071_ ), .ZN(_01072_ ) );
NAND3_X1 _16817_ ( .A1(_01072_ ), .A2(_01068_ ), .A3(_01890_ ), .ZN(_01073_ ) );
NAND2_X1 _16818_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01074_ ) );
NAND4_X1 _16819_ ( .A1(_01073_ ), .A2(_01545_ ), .A3(_03656_ ), .A4(_01074_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _16820_ ( .A1(_03726_ ), .A2(_01545_ ), .A3(\myifu.state [2] ), .ZN(_01075_ ) );
NAND3_X1 _16821_ ( .A1(_01071_ ), .A2(_01890_ ), .A3(_01989_ ), .ZN(_01076_ ) );
NAND2_X1 _16822_ ( .A1(_01075_ ), .A2(_01076_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _16823_ ( .A1(_03713_ ), .A2(\myifu.state [2] ), .A3(_03725_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16824_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01077_ ) );
NOR3_X1 _16825_ ( .A1(_01077_ ), .A2(_00503_ ), .A3(_00572_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NOR3_X1 _16826_ ( .A1(_01077_ ), .A2(_00504_ ), .A3(_00572_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _16827_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00572_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _16828_ ( .A1(\IF_ID_pc [4] ), .A2(_05888_ ), .A3(_03655_ ), .A4(_00572_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
NOR3_X1 _16829_ ( .A1(_01077_ ), .A2(_00501_ ), .A3(_00572_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _16830_ ( .A1(_05892_ ), .A2(_05888_ ), .A3(\IF_ID_pc [3] ), .A4(_00572_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
AND3_X1 _16831_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05890_ ), .A3(_00572_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _16832_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05890_ ), .A3(_00557_ ), .A4(_00560_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
AND3_X1 _16833_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_05892_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
AND3_X1 _16834_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_03655_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
AND3_X1 _16835_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
AND3_X1 _16836_ ( .A1(_01989_ ), .A2(_05890_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
AND2_X1 _16837_ ( .A1(_01797_ ), .A2(_01863_ ), .ZN(_01078_ ) );
NAND2_X1 _16838_ ( .A1(_01078_ ), .A2(\myifu.state [0] ), .ZN(_01079_ ) );
OAI21_X1 _16839_ ( .A(\myifu.state [1] ), .B1(_03282_ ), .B2(_03333_ ), .ZN(_01080_ ) );
NAND2_X1 _16840_ ( .A1(_00392_ ), .A2(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01081_ ) );
NAND4_X1 _16841_ ( .A1(_01079_ ), .A2(_01074_ ), .A3(_01080_ ), .A4(_01081_ ), .ZN(_01082_ ) );
AOI221_X4 _16842_ ( .A(_01082_ ), .B1(_01072_ ), .B2(\myifu.state [0] ), .C1(_01891_ ), .C2(_03726_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _16843_ ( .A1(_03527_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03146_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16844_ ( .A(_03223_ ), .ZN(_01083_ ) );
AOI211_X1 _16845_ ( .A(_03282_ ), .B(_00370_ ), .C1(_03187_ ), .C2(_01083_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
NAND4_X1 _16846_ ( .A1(_01080_ ), .A2(_01081_ ), .A3(_01459_ ), .A4(_01074_ ), .ZN(_01084_ ) );
AOI21_X1 _16847_ ( .A(_01084_ ), .B1(_01864_ ), .B2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _16848_ ( .A(_05969_ ), .B(_03793_ ), .S(\mylsu.state [0] ), .Z(_01085_ ) );
NOR2_X1 _16849_ ( .A1(_05973_ ), .A2(_01085_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ) );
NOR3_X1 _16850_ ( .A1(_05973_ ), .A2(_03801_ ), .A3(_01085_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
NOR4_X1 _16851_ ( .A1(_05873_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A3(_03763_ ), .A4(_05878_ ), .ZN(_01086_ ) );
NOR2_X1 _16852_ ( .A1(_03800_ ), .A2(_03740_ ), .ZN(_01087_ ) );
AND2_X1 _16853_ ( .A1(_01941_ ), .A2(_01087_ ), .ZN(_01088_ ) );
NAND3_X1 _16854_ ( .A1(_01086_ ), .A2(\mylsu.state [0] ), .A3(_01088_ ), .ZN(_01089_ ) );
AND2_X1 _16855_ ( .A1(_05972_ ), .A2(_03725_ ), .ZN(_01090_ ) );
OAI21_X1 _16856_ ( .A(_01089_ ), .B1(_05909_ ), .B2(_01090_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
INV_X1 _16857_ ( .A(io_master_wready ), .ZN(_01091_ ) );
NAND3_X1 _16858_ ( .A1(_03790_ ), .A2(\mylsu.state [2] ), .A3(_01091_ ), .ZN(_01092_ ) );
INV_X1 _16859_ ( .A(_01951_ ), .ZN(_01093_ ) );
BUF_X2 _16860_ ( .A(_01944_ ), .Z(_01094_ ) );
NAND4_X1 _16861_ ( .A1(_01094_ ), .A2(_03790_ ), .A3(io_master_awready ), .A4(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_01095_ ) );
AND2_X1 _16862_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01096_ ) );
OR3_X1 _16863_ ( .A1(_01095_ ), .A2(_03740_ ), .A3(_01096_ ), .ZN(_01097_ ) );
OAI21_X1 _16864_ ( .A(_01092_ ), .B1(_01093_ ), .B2(_01097_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
AND3_X1 _16865_ ( .A1(_03787_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .A3(_03788_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
INV_X1 _16866_ ( .A(_01950_ ), .ZN(_01098_ ) );
AND3_X1 _16867_ ( .A1(_01087_ ), .A2(_05960_ ), .A3(_01096_ ), .ZN(_01099_ ) );
NAND3_X1 _16868_ ( .A1(_05904_ ), .A2(_01098_ ), .A3(_01099_ ), .ZN(_01100_ ) );
NAND3_X1 _16869_ ( .A1(_03790_ ), .A2(\mylsu.state [4] ), .A3(io_master_awready ), .ZN(_01101_ ) );
NAND4_X1 _16870_ ( .A1(_03796_ ), .A2(\mylsu.state [2] ), .A3(_03798_ ), .A4(io_master_wready ), .ZN(_01102_ ) );
OAI211_X1 _16871_ ( .A(\mylsu.state [1] ), .B(_03790_ ), .C1(_05975_ ), .C2(_05977_ ), .ZN(_01103_ ) );
NAND4_X1 _16872_ ( .A1(_01100_ ), .A2(_01101_ ), .A3(_01102_ ), .A4(_01103_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
OAI211_X1 _16873_ ( .A(_05871_ ), .B(_01088_ ), .C1(_05873_ ), .C2(_05879_ ), .ZN(_01104_ ) );
OR2_X1 _16874_ ( .A1(_01104_ ), .A2(_05884_ ), .ZN(_01105_ ) );
NAND3_X1 _16875_ ( .A1(_05972_ ), .A2(_03725_ ), .A3(_00283_ ), .ZN(_01106_ ) );
NAND3_X1 _16876_ ( .A1(_05900_ ), .A2(_03744_ ), .A3(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .ZN(_01107_ ) );
AND4_X1 _16877_ ( .A1(_01922_ ), .A2(_01098_ ), .A3(_01087_ ), .A4(_05960_ ), .ZN(_01108_ ) );
AND2_X1 _16878_ ( .A1(_01951_ ), .A2(\mylsu.state [0] ), .ZN(_01109_ ) );
AND3_X1 _16879_ ( .A1(_01944_ ), .A2(_01091_ ), .A3(_05881_ ), .ZN(_01110_ ) );
NAND3_X1 _16880_ ( .A1(_01109_ ), .A2(_05886_ ), .A3(_01110_ ), .ZN(_01111_ ) );
NAND4_X1 _16881_ ( .A1(_01087_ ), .A2(_05960_ ), .A3(_01949_ ), .A4(_01947_ ), .ZN(_01112_ ) );
NAND2_X1 _16882_ ( .A1(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .A2(_03740_ ), .ZN(_01113_ ) );
AOI221_X4 _16883_ ( .A(_03800_ ), .B1(\mylsu.state [0] ), .B2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .C1(_05978_ ), .C2(\mylsu.state [1] ), .ZN(_01114_ ) );
NAND4_X1 _16884_ ( .A1(_01111_ ), .A2(_01112_ ), .A3(_01113_ ), .A4(_01114_ ), .ZN(_01115_ ) );
NOR4_X1 _16885_ ( .A1(_05887_ ), .A2(_03744_ ), .A3(_01944_ ), .A4(_03740_ ), .ZN(_01116_ ) );
AOI211_X1 _16886_ ( .A(_01108_ ), .B(_01115_ ), .C1(\mylsu.state [0] ), .C2(_01116_ ), .ZN(_01117_ ) );
NAND4_X1 _16887_ ( .A1(_01105_ ), .A2(_01106_ ), .A3(_01107_ ), .A4(_01117_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
AND2_X1 _16888_ ( .A1(_01094_ ), .A2(EXU_valid_LSU ), .ZN(_01118_ ) );
NAND4_X1 _16889_ ( .A1(_01109_ ), .A2(io_master_wready ), .A3(_01087_ ), .A4(_01118_ ), .ZN(_01119_ ) );
NAND3_X1 _16890_ ( .A1(_03796_ ), .A2(\mylsu.state [4] ), .A3(_03798_ ), .ZN(_01120_ ) );
AOI21_X1 _16891_ ( .A(io_master_awready ), .B1(_01119_ ), .B2(_01120_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
AOI211_X1 _16892_ ( .A(\mylsu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__A_B ), .B(_03800_ ), .C1(_01091_ ), .C2(_05881_ ), .ZN(_01121_ ) );
AND4_X1 _16893_ ( .A1(_05904_ ), .A2(_01121_ ), .A3(_01098_ ), .A4(_01118_ ), .ZN(\mylsu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ) );
MUX2_X1 _16894_ ( .A(\LS_WB_wdata_csreg [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_03735_ ), .Z(_01122_ ) );
INV_X1 _16895_ ( .A(_03741_ ), .ZN(_01123_ ) );
OR2_X1 _16896_ ( .A1(_03732_ ), .A2(_01123_ ), .ZN(_01124_ ) );
BUF_X4 _16897_ ( .A(_01124_ ), .Z(_01125_ ) );
BUF_X4 _16898_ ( .A(_01125_ ), .Z(_01126_ ) );
MUX2_X1 _16899_ ( .A(_01122_ ), .B(\EX_LS_pc [21] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
BUF_X4 _16900_ ( .A(_02039_ ), .Z(_01127_ ) );
MUX2_X1 _16901_ ( .A(\LS_WB_wdata_csreg [20] ), .B(\EX_LS_result_csreg_mem [20] ), .S(_01127_ ), .Z(_01128_ ) );
MUX2_X1 _16902_ ( .A(_01128_ ), .B(\EX_LS_pc [20] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
OAI22_X1 _16903_ ( .A1(_03735_ ), .A2(_02005_ ), .B1(_03749_ ), .B2(_05997_ ), .ZN(_01129_ ) );
MUX2_X1 _16904_ ( .A(_01129_ ), .B(\EX_LS_pc [19] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
AOI21_X1 _16905_ ( .A(\EX_LS_pc [18] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01130_ ) );
MUX2_X1 _16906_ ( .A(\LS_WB_wdata_csreg [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_02039_ ), .Z(_01131_ ) );
NOR3_X1 _16907_ ( .A1(_03732_ ), .A2(_01123_ ), .A3(_01131_ ), .ZN(_01132_ ) );
NOR2_X1 _16908_ ( .A1(_01130_ ), .A2(_01132_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
OAI22_X1 _16909_ ( .A1(_03735_ ), .A2(_02006_ ), .B1(_03748_ ), .B2(_05350_ ), .ZN(_01133_ ) );
MUX2_X1 _16910_ ( .A(_01133_ ), .B(\EX_LS_pc [17] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _16911_ ( .A(\EX_LS_pc [16] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01134_ ) );
INV_X2 _16912_ ( .A(_02039_ ), .ZN(_01135_ ) );
OAI21_X1 _16913_ ( .A(_03742_ ), .B1(_01135_ ), .B2(_05364_ ), .ZN(_01136_ ) );
BUF_X4 _16914_ ( .A(_01135_ ), .Z(_01137_ ) );
AOI221_X4 _16915_ ( .A(_01136_ ), .B1(\LS_WB_wdata_csreg [16] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01138_ ) );
NOR2_X1 _16916_ ( .A1(_01134_ ), .A2(_01138_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _16917_ ( .A(\LS_WB_wdata_csreg [15] ), .B(\EX_LS_result_csreg_mem [15] ), .S(_01127_ ), .Z(_01139_ ) );
MUX2_X1 _16918_ ( .A(_01139_ ), .B(\EX_LS_pc [15] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _16919_ ( .A(\EX_LS_pc [14] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01140_ ) );
OAI21_X1 _16920_ ( .A(_03742_ ), .B1(_01135_ ), .B2(_05404_ ), .ZN(_01141_ ) );
AOI221_X4 _16921_ ( .A(_01141_ ), .B1(\LS_WB_wdata_csreg [14] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01142_ ) );
NOR2_X1 _16922_ ( .A1(_01140_ ), .A2(_01142_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
OAI22_X1 _16923_ ( .A1(_03735_ ), .A2(_02007_ ), .B1(_03748_ ), .B2(_05428_ ), .ZN(_01143_ ) );
MUX2_X1 _16924_ ( .A(_01143_ ), .B(\EX_LS_pc [13] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _16925_ ( .A(\LS_WB_wdata_csreg [12] ), .B(\EX_LS_result_csreg_mem [12] ), .S(_01127_ ), .Z(_01144_ ) );
MUX2_X1 _16926_ ( .A(_01144_ ), .B(\EX_LS_pc [12] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _16927_ ( .A(\EX_LS_pc [30] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01145_ ) );
MUX2_X1 _16928_ ( .A(\LS_WB_wdata_csreg [30] ), .B(\EX_LS_result_csreg_mem [30] ), .S(_02039_ ), .Z(_01146_ ) );
NOR3_X1 _16929_ ( .A1(_03732_ ), .A2(_01123_ ), .A3(_01146_ ), .ZN(_01147_ ) );
NOR2_X1 _16930_ ( .A1(_01145_ ), .A2(_01147_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
AOI21_X1 _16931_ ( .A(\EX_LS_pc [11] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01148_ ) );
OAI21_X1 _16932_ ( .A(_03741_ ), .B1(_01135_ ), .B2(_05469_ ), .ZN(_01149_ ) );
AOI221_X4 _16933_ ( .A(_01149_ ), .B1(\LS_WB_wdata_csreg [11] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01150_ ) );
NOR2_X1 _16934_ ( .A1(_01148_ ), .A2(_01150_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _16935_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_01127_ ), .Z(_01151_ ) );
MUX2_X1 _16936_ ( .A(_01151_ ), .B(\EX_LS_pc [10] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
AOI21_X1 _16937_ ( .A(\EX_LS_pc [9] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01152_ ) );
OAI21_X1 _16938_ ( .A(_03741_ ), .B1(_01135_ ), .B2(_06001_ ), .ZN(_01153_ ) );
AOI221_X4 _16939_ ( .A(_01153_ ), .B1(\LS_WB_wdata_csreg [9] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01154_ ) );
NOR2_X1 _16940_ ( .A1(_01152_ ), .A2(_01154_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _16941_ ( .A(\EX_LS_pc [8] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01155_ ) );
OAI21_X1 _16942_ ( .A(_03741_ ), .B1(_01135_ ), .B2(_05544_ ), .ZN(_01156_ ) );
AOI221_X4 _16943_ ( .A(_01156_ ), .B1(\LS_WB_wdata_csreg [8] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01157_ ) );
NOR2_X1 _16944_ ( .A1(_01155_ ), .A2(_01157_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _16945_ ( .A(\LS_WB_wdata_csreg [7] ), .B(\EX_LS_result_csreg_mem [7] ), .S(_01127_ ), .Z(_01158_ ) );
MUX2_X1 _16946_ ( .A(_01158_ ), .B(\EX_LS_pc [7] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
AOI221_X4 _16947_ ( .A(_01125_ ), .B1(\LS_WB_wdata_csreg [6] ), .B2(_03748_ ), .C1(\EX_LS_result_csreg_mem [6] ), .C2(_03735_ ), .ZN(_01159_ ) );
AOI21_X1 _16948_ ( .A(\EX_LS_pc [6] ), .B1(_03733_ ), .B2(_03742_ ), .ZN(_01160_ ) );
NOR2_X1 _16949_ ( .A1(_01159_ ), .A2(_01160_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _16950_ ( .A(\LS_WB_wdata_csreg [5] ), .B(\EX_LS_result_csreg_mem [5] ), .S(_01127_ ), .Z(_01161_ ) );
MUX2_X1 _16951_ ( .A(_01161_ ), .B(\EX_LS_pc [5] ), .S(_01126_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _16952_ ( .A(\LS_WB_wdata_csreg [4] ), .B(\EX_LS_result_csreg_mem [4] ), .S(_01127_ ), .Z(_01162_ ) );
MUX2_X1 _16953_ ( .A(_01162_ ), .B(\EX_LS_pc [4] ), .S(_01125_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
AOI221_X4 _16954_ ( .A(_01125_ ), .B1(_03748_ ), .B2(\LS_WB_wdata_csreg [3] ), .C1(\EX_LS_result_csreg_mem [3] ), .C2(_03735_ ), .ZN(_01163_ ) );
AOI21_X1 _16955_ ( .A(\EX_LS_pc [3] ), .B1(_03733_ ), .B2(_03742_ ), .ZN(_01164_ ) );
NOR2_X1 _16956_ ( .A1(_01163_ ), .A2(_01164_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
AOI21_X1 _16957_ ( .A(\EX_LS_pc [2] ), .B1(_03734_ ), .B2(_03743_ ), .ZN(_01165_ ) );
OAI21_X1 _16958_ ( .A(_03741_ ), .B1(_01135_ ), .B2(_05983_ ), .ZN(_01166_ ) );
AOI221_X4 _16959_ ( .A(_01166_ ), .B1(\LS_WB_wdata_csreg [2] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01167_ ) );
NOR2_X1 _16960_ ( .A1(_01165_ ), .A2(_01167_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
AOI21_X1 _16961_ ( .A(\EX_LS_pc [29] ), .B1(_03733_ ), .B2(_03743_ ), .ZN(_01168_ ) );
OAI21_X1 _16962_ ( .A(_03741_ ), .B1(_01135_ ), .B2(_05239_ ), .ZN(_01169_ ) );
AOI221_X4 _16963_ ( .A(_01169_ ), .B1(\LS_WB_wdata_csreg [29] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01170_ ) );
NOR2_X1 _16964_ ( .A1(_01168_ ), .A2(_01170_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _16965_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\EX_LS_result_csreg_mem [1] ), .S(_01127_ ), .Z(_01171_ ) );
MUX2_X1 _16966_ ( .A(_01171_ ), .B(\EX_LS_pc [1] ), .S(_01125_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI21_X1 _16967_ ( .A(\EX_LS_pc [0] ), .B1(_03733_ ), .B2(_03742_ ), .ZN(_01172_ ) );
OAI21_X1 _16968_ ( .A(_03741_ ), .B1(_01135_ ), .B2(_05722_ ), .ZN(_01173_ ) );
AOI221_X4 _16969_ ( .A(_01173_ ), .B1(\LS_WB_wdata_csreg [0] ), .B2(_01137_ ), .C1(_01093_ ), .C2(_01094_ ), .ZN(_01174_ ) );
NOR2_X1 _16970_ ( .A1(_01172_ ), .A2(_01174_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
AOI221_X4 _16971_ ( .A(_01125_ ), .B1(\LS_WB_wdata_csreg [28] ), .B2(_01137_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [28] ), .ZN(_01175_ ) );
AOI21_X1 _16972_ ( .A(\EX_LS_pc [28] ), .B1(_03733_ ), .B2(_03742_ ), .ZN(_01176_ ) );
NOR2_X1 _16973_ ( .A1(_01175_ ), .A2(_01176_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _16974_ ( .A(\LS_WB_wdata_csreg [27] ), .B(\EX_LS_result_csreg_mem [27] ), .S(_01127_ ), .Z(_01177_ ) );
MUX2_X1 _16975_ ( .A(_01177_ ), .B(\EX_LS_pc [27] ), .S(_01125_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI221_X4 _16976_ ( .A(_01124_ ), .B1(\LS_WB_wdata_csreg [26] ), .B2(_03748_ ), .C1(\EX_LS_result_csreg_mem [26] ), .C2(_03735_ ), .ZN(_01178_ ) );
AOI21_X1 _16977_ ( .A(\EX_LS_pc [26] ), .B1(_03733_ ), .B2(_03742_ ), .ZN(_01179_ ) );
NOR2_X1 _16978_ ( .A1(_01178_ ), .A2(_01179_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _16979_ ( .A(\LS_WB_wdata_csreg [25] ), .B(\EX_LS_result_csreg_mem [25] ), .S(_01127_ ), .Z(_01180_ ) );
MUX2_X1 _16980_ ( .A(_01180_ ), .B(\EX_LS_pc [25] ), .S(_01125_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _16981_ ( .A(\LS_WB_wdata_csreg [24] ), .B(\EX_LS_result_csreg_mem [24] ), .S(_02039_ ), .Z(_01181_ ) );
MUX2_X1 _16982_ ( .A(_01181_ ), .B(\EX_LS_pc [24] ), .S(_01125_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
AOI221_X4 _16983_ ( .A(_01124_ ), .B1(\LS_WB_wdata_csreg [23] ), .B2(_03748_ ), .C1(\EX_LS_result_csreg_mem [23] ), .C2(_03735_ ), .ZN(_01182_ ) );
AOI21_X1 _16984_ ( .A(\EX_LS_pc [23] ), .B1(_03733_ ), .B2(_03742_ ), .ZN(_01183_ ) );
NOR2_X1 _16985_ ( .A1(_01182_ ), .A2(_01183_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _16986_ ( .A(\LS_WB_wdata_csreg [22] ), .B(\EX_LS_result_csreg_mem [22] ), .S(_02039_ ), .Z(_01184_ ) );
MUX2_X1 _16987_ ( .A(_01184_ ), .B(\EX_LS_pc [22] ), .S(_01125_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
AOI221_X4 _16988_ ( .A(_01124_ ), .B1(\LS_WB_wdata_csreg [31] ), .B2(_01137_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [31] ), .ZN(_01185_ ) );
AOI21_X1 _16989_ ( .A(\EX_LS_pc [31] ), .B1(_03733_ ), .B2(_03742_ ), .ZN(_01186_ ) );
NOR2_X1 _16990_ ( .A1(_01185_ ), .A2(_01186_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X2 _16991_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01187_ ) );
INV_X1 _16992_ ( .A(_01187_ ), .ZN(_01188_ ) );
OR3_X1 _16993_ ( .A1(_00428_ ), .A2(_05875_ ), .A3(_01188_ ), .ZN(_01189_ ) );
NAND3_X1 _16994_ ( .A1(_00396_ ), .A2(_01884_ ), .A3(_01188_ ), .ZN(_01190_ ) );
AND2_X1 _16995_ ( .A1(_01189_ ), .A2(_01190_ ), .ZN(_01191_ ) );
AND2_X2 _16996_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01192_ ) );
INV_X1 _16997_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01193_ ) );
AND2_X1 _16998_ ( .A1(_01192_ ), .A2(_01193_ ), .ZN(_01194_ ) );
BUF_X4 _16999_ ( .A(_01194_ ), .Z(_01195_ ) );
AND2_X1 _17000_ ( .A1(_01191_ ), .A2(_01195_ ), .ZN(_01196_ ) );
AND2_X1 _17001_ ( .A1(_01193_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01197_ ) );
INV_X1 _17002_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_01198_ ) );
AND2_X1 _17003_ ( .A1(_01197_ ), .A2(_01198_ ), .ZN(_01199_ ) );
NAND2_X1 _17004_ ( .A1(_01198_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01200_ ) );
NOR2_X1 _17005_ ( .A1(_01200_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01201_ ) );
OR2_X1 _17006_ ( .A1(_01199_ ), .A2(_01201_ ), .ZN(_01202_ ) );
NOR2_X4 _17007_ ( .A1(_01196_ ), .A2(_01202_ ), .ZN(_01203_ ) );
BUF_X4 _17008_ ( .A(_01203_ ), .Z(_01204_ ) );
AND2_X1 _17009_ ( .A1(_01192_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01205_ ) );
BUF_X4 _17010_ ( .A(_01205_ ), .Z(_01206_ ) );
INV_X1 _17011_ ( .A(_01206_ ), .ZN(_01207_ ) );
AND4_X1 _17012_ ( .A1(\io_master_arid [1] ), .A2(_00406_ ), .A3(_00409_ ), .A4(_01207_ ), .ZN(_01208_ ) );
OAI21_X1 _17013_ ( .A(_01204_ ), .B1(_01208_ ), .B2(_01195_ ), .ZN(_01209_ ) );
INV_X2 _17014_ ( .A(_01199_ ), .ZN(_01210_ ) );
BUF_X4 _17015_ ( .A(_01210_ ), .Z(_01211_ ) );
NOR2_X1 _17016_ ( .A1(_00496_ ), .A2(_05877_ ), .ZN(_01212_ ) );
NOR2_X1 _17017_ ( .A1(_05915_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01213_ ) );
NOR2_X1 _17018_ ( .A1(_00428_ ), .A2(_05877_ ), .ZN(_01214_ ) );
NOR2_X1 _17019_ ( .A1(_05918_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01215_ ) );
AOI22_X1 _17020_ ( .A1(_01212_ ), .A2(_01213_ ), .B1(_01214_ ), .B2(_01215_ ), .ZN(_01216_ ) );
OR3_X1 _17021_ ( .A1(_00456_ ), .A2(_05877_ ), .A3(_01188_ ), .ZN(_01217_ ) );
NAND4_X1 _17022_ ( .A1(_00396_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_01884_ ), .ZN(_01218_ ) );
AND3_X1 _17023_ ( .A1(_01216_ ), .A2(_01217_ ), .A3(_01218_ ), .ZN(_01219_ ) );
BUF_X4 _17024_ ( .A(_01219_ ), .Z(_01220_ ) );
OAI21_X1 _17025_ ( .A(_01209_ ), .B1(_01211_ ), .B2(_01220_ ), .ZN(_01221_ ) );
MUX2_X1 _17026_ ( .A(\EX_LS_result_reg [21] ), .B(_01221_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
BUF_X4 _17027_ ( .A(_01195_ ), .Z(_01222_ ) );
NOR3_X1 _17028_ ( .A1(_00412_ ), .A2(_05878_ ), .A3(_01206_ ), .ZN(_01223_ ) );
OAI21_X1 _17029_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01223_ ), .ZN(_01224_ ) );
OAI21_X1 _17030_ ( .A(_01224_ ), .B1(_01211_ ), .B2(_01220_ ), .ZN(_01225_ ) );
MUX2_X1 _17031_ ( .A(\EX_LS_result_reg [20] ), .B(_01225_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NOR3_X1 _17032_ ( .A1(_00415_ ), .A2(_05878_ ), .A3(_01206_ ), .ZN(_01226_ ) );
OAI21_X1 _17033_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01226_ ), .ZN(_01227_ ) );
OAI21_X1 _17034_ ( .A(_01227_ ), .B1(_01211_ ), .B2(_01220_ ), .ZN(_01228_ ) );
MUX2_X1 _17035_ ( .A(\EX_LS_result_reg [19] ), .B(_01228_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
AND2_X1 _17036_ ( .A1(_01203_ ), .A2(_01207_ ), .ZN(_01229_ ) );
NOR2_X2 _17037_ ( .A1(_00419_ ), .A2(_05874_ ), .ZN(_01230_ ) );
OAI21_X1 _17038_ ( .A(_01229_ ), .B1(_01192_ ), .B2(_01230_ ), .ZN(_01231_ ) );
OAI21_X1 _17039_ ( .A(_01231_ ), .B1(_01211_ ), .B2(_01220_ ), .ZN(_01232_ ) );
MUX2_X1 _17040_ ( .A(\EX_LS_result_reg [18] ), .B(_01232_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NOR3_X1 _17041_ ( .A1(_00422_ ), .A2(_05878_ ), .A3(_01206_ ), .ZN(_01233_ ) );
OAI21_X1 _17042_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01233_ ), .ZN(_01234_ ) );
OAI21_X1 _17043_ ( .A(_01234_ ), .B1(_01211_ ), .B2(_01220_ ), .ZN(_01235_ ) );
MUX2_X1 _17044_ ( .A(\EX_LS_result_reg [17] ), .B(_01235_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
AND4_X1 _17045_ ( .A1(\io_master_arid [1] ), .A2(_00423_ ), .A3(_00425_ ), .A4(_01207_ ), .ZN(_01236_ ) );
OAI21_X1 _17046_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01236_ ), .ZN(_01237_ ) );
BUF_X4 _17047_ ( .A(_01219_ ), .Z(_01238_ ) );
OAI21_X1 _17048_ ( .A(_01237_ ), .B1(_01211_ ), .B2(_01238_ ), .ZN(_01239_ ) );
MUX2_X1 _17049_ ( .A(\EX_LS_result_reg [16] ), .B(_01239_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
NOR2_X1 _17050_ ( .A1(_01219_ ), .A2(_01210_ ), .ZN(_01240_ ) );
NOR2_X1 _17051_ ( .A1(_01240_ ), .A2(_05969_ ), .ZN(_01241_ ) );
INV_X1 _17052_ ( .A(_01192_ ), .ZN(_01242_ ) );
AOI21_X1 _17053_ ( .A(_01242_ ), .B1(_01189_ ), .B2(_01190_ ), .ZN(_01243_ ) );
NOR3_X1 _17054_ ( .A1(_01199_ ), .A2(_01192_ ), .A3(_01201_ ), .ZN(_01244_ ) );
AOI21_X1 _17055_ ( .A(_01243_ ), .B1(_01214_ ), .B2(_01244_ ), .ZN(_01245_ ) );
AOI22_X1 _17056_ ( .A1(_01241_ ), .A2(_01245_ ), .B1(_05969_ ), .B2(_04583_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
NOR2_X1 _17057_ ( .A1(_01242_ ), .A2(_01187_ ), .ZN(_01246_ ) );
INV_X1 _17058_ ( .A(_01246_ ), .ZN(_01247_ ) );
OR3_X1 _17059_ ( .A1(_00611_ ), .A2(_05878_ ), .A3(_01247_ ), .ZN(_01248_ ) );
NOR2_X1 _17060_ ( .A1(_01202_ ), .A2(_01246_ ), .ZN(_01249_ ) );
AND2_X1 _17061_ ( .A1(\io_master_arid [1] ), .A2(_01249_ ), .ZN(_01250_ ) );
NAND3_X1 _17062_ ( .A1(_00430_ ), .A2(_00432_ ), .A3(_01250_ ), .ZN(_01251_ ) );
BUF_X4 _17063_ ( .A(_01210_ ), .Z(_01252_ ) );
OAI211_X1 _17064_ ( .A(_01248_ ), .B(_01251_ ), .C1(_01220_ ), .C2(_01252_ ), .ZN(_01253_ ) );
MUX2_X1 _17065_ ( .A(\EX_LS_result_reg [14] ), .B(_01253_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
OR3_X1 _17066_ ( .A1(_00784_ ), .A2(_05877_ ), .A3(_01247_ ), .ZN(_01254_ ) );
NAND3_X1 _17067_ ( .A1(_00433_ ), .A2(_00435_ ), .A3(_01250_ ), .ZN(_01255_ ) );
OAI211_X1 _17068_ ( .A(_01254_ ), .B(_01255_ ), .C1(_01220_ ), .C2(_01252_ ), .ZN(_01256_ ) );
MUX2_X1 _17069_ ( .A(\EX_LS_result_reg [13] ), .B(_01256_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _17070_ ( .A1(_00436_ ), .A2(_00438_ ), .A3(_01250_ ), .ZN(_01257_ ) );
NOR2_X1 _17071_ ( .A1(_00475_ ), .A2(_05876_ ), .ZN(_01258_ ) );
INV_X1 _17072_ ( .A(_01258_ ), .ZN(_01259_ ) );
OAI221_X1 _17073_ ( .A(_01257_ ), .B1(_01247_ ), .B2(_01259_ ), .C1(_01238_ ), .C2(_01252_ ), .ZN(_01260_ ) );
MUX2_X1 _17074_ ( .A(\EX_LS_result_reg [12] ), .B(_01260_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
AOI211_X1 _17075_ ( .A(_05877_ ), .B(_01192_ ), .C1(_00399_ ), .C2(_00400_ ), .ZN(_01261_ ) );
OAI21_X1 _17076_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01261_ ), .ZN(_01262_ ) );
OAI21_X1 _17077_ ( .A(_01262_ ), .B1(_01211_ ), .B2(_01238_ ), .ZN(_01263_ ) );
MUX2_X1 _17078_ ( .A(\EX_LS_result_reg [30] ), .B(_01263_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _17079_ ( .A1(_00444_ ), .A2(\io_master_arid [1] ), .A3(_01249_ ), .ZN(_01264_ ) );
NOR2_X1 _17080_ ( .A1(_00484_ ), .A2(_05876_ ), .ZN(_01265_ ) );
INV_X1 _17081_ ( .A(_01265_ ), .ZN(_01266_ ) );
OAI221_X1 _17082_ ( .A(_01264_ ), .B1(_01247_ ), .B2(_01266_ ), .C1(_01238_ ), .C2(_01252_ ), .ZN(_01267_ ) );
MUX2_X1 _17083_ ( .A(\EX_LS_result_reg [11] ), .B(_01267_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
OR3_X1 _17084_ ( .A1(_00487_ ), .A2(_05877_ ), .A3(_01247_ ), .ZN(_01268_ ) );
NAND3_X1 _17085_ ( .A1(_00447_ ), .A2(\io_master_arid [1] ), .A3(_01249_ ), .ZN(_01269_ ) );
OAI211_X1 _17086_ ( .A(_01268_ ), .B(_01269_ ), .C1(_01220_ ), .C2(_01252_ ), .ZN(_01270_ ) );
MUX2_X1 _17087_ ( .A(\EX_LS_result_reg [10] ), .B(_01270_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
OR3_X1 _17088_ ( .A1(_00490_ ), .A2(_05877_ ), .A3(_01247_ ), .ZN(_01271_ ) );
NAND3_X1 _17089_ ( .A1(_00448_ ), .A2(_00450_ ), .A3(_01250_ ), .ZN(_01272_ ) );
OAI211_X1 _17090_ ( .A(_01271_ ), .B(_01272_ ), .C1(_01220_ ), .C2(_01252_ ), .ZN(_01273_ ) );
MUX2_X1 _17091_ ( .A(\EX_LS_result_reg [9] ), .B(_01273_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _17092_ ( .A1(_00451_ ), .A2(_00453_ ), .A3(_01250_ ), .ZN(_01274_ ) );
NAND4_X1 _17093_ ( .A1(_00491_ ), .A2(_00493_ ), .A3(\io_master_arid [1] ), .A4(_01246_ ), .ZN(_01275_ ) );
OAI211_X1 _17094_ ( .A(_01274_ ), .B(_01275_ ), .C1(_01220_ ), .C2(_01252_ ), .ZN(_01276_ ) );
MUX2_X1 _17095_ ( .A(\EX_LS_result_reg [8] ), .B(_01276_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
AND4_X1 _17096_ ( .A1(_01202_ ), .A2(_01216_ ), .A3(_01217_ ), .A4(_01218_ ), .ZN(_01277_ ) );
OAI21_X1 _17097_ ( .A(_01249_ ), .B1(_00456_ ), .B2(_05879_ ), .ZN(_01278_ ) );
OAI211_X1 _17098_ ( .A(_01278_ ), .B(fanout_net_44 ), .C1(_01212_ ), .C2(_01247_ ), .ZN(_01279_ ) );
OAI22_X1 _17099_ ( .A1(_01277_ ), .A2(_01279_ ), .B1(fanout_net_44 ), .B2(_04726_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _17100_ ( .A1(_05969_ ), .A2(\EX_LS_result_reg [6] ), .ZN(_01280_ ) );
MUX2_X1 _17101_ ( .A(_00611_ ), .B(_00737_ ), .S(_05915_ ), .Z(_01281_ ) );
AND2_X1 _17102_ ( .A1(_01202_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01282_ ) );
AND2_X1 _17103_ ( .A1(_01281_ ), .A2(_01282_ ), .ZN(_01283_ ) );
NOR2_X1 _17104_ ( .A1(_01244_ ), .A2(_01187_ ), .ZN(_01284_ ) );
INV_X1 _17105_ ( .A(_01284_ ), .ZN(_01285_ ) );
AOI211_X1 _17106_ ( .A(_05969_ ), .B(_05879_ ), .C1(_00459_ ), .C2(_01285_ ), .ZN(_01286_ ) );
NOR2_X1 _17107_ ( .A1(_01285_ ), .A2(_01282_ ), .ZN(_01287_ ) );
NAND2_X1 _17108_ ( .A1(_01052_ ), .A2(_01287_ ), .ZN(_01288_ ) );
NAND2_X1 _17109_ ( .A1(_01286_ ), .A2(_01288_ ), .ZN(_01289_ ) );
OAI21_X1 _17110_ ( .A(_01280_ ), .B1(_01283_ ), .B2(_01289_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
AOI211_X1 _17111_ ( .A(_05968_ ), .B(_05878_ ), .C1(_00626_ ), .C2(_01287_ ), .ZN(_01290_ ) );
NAND2_X1 _17112_ ( .A1(_00462_ ), .A2(_01285_ ), .ZN(_01291_ ) );
NAND2_X1 _17113_ ( .A1(_01290_ ), .A2(_01291_ ), .ZN(_01292_ ) );
MUX2_X1 _17114_ ( .A(_00784_ ), .B(_00754_ ), .S(_05915_ ), .Z(_01293_ ) );
AOI21_X1 _17115_ ( .A(_01292_ ), .B1(_01282_ ), .B2(_01293_ ), .ZN(_01294_ ) );
AND2_X1 _17116_ ( .A1(_05969_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01295_ ) );
OR2_X1 _17117_ ( .A1(_01294_ ), .A2(_01295_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
NOR3_X1 _17118_ ( .A1(_00466_ ), .A2(_05875_ ), .A3(_01188_ ), .ZN(_01296_ ) );
INV_X1 _17119_ ( .A(_01296_ ), .ZN(_01297_ ) );
AND4_X1 _17120_ ( .A1(_01884_ ), .A2(_00436_ ), .A3(_00438_ ), .A4(_01215_ ), .ZN(_01298_ ) );
OR4_X1 _17121_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(_00412_ ), .A3(_05915_ ), .A4(_05875_ ), .ZN(_01299_ ) );
OAI21_X1 _17122_ ( .A(_01299_ ), .B1(_01213_ ), .B2(_01259_ ), .ZN(_01300_ ) );
INV_X1 _17123_ ( .A(_01215_ ), .ZN(_01301_ ) );
AOI21_X1 _17124_ ( .A(_01298_ ), .B1(_01300_ ), .B2(_01301_ ), .ZN(_01302_ ) );
OAI21_X1 _17125_ ( .A(_01297_ ), .B1(_01302_ ), .B2(_01187_ ), .ZN(_01303_ ) );
NOR3_X1 _17126_ ( .A1(_00412_ ), .A2(_05876_ ), .A3(_01187_ ), .ZN(_01304_ ) );
OAI21_X1 _17127_ ( .A(_01195_ ), .B1(_01296_ ), .B2(_01304_ ), .ZN(_01305_ ) );
OAI21_X1 _17128_ ( .A(_01206_ ), .B1(_01296_ ), .B2(_01304_ ), .ZN(_01306_ ) );
OR3_X1 _17129_ ( .A1(_00466_ ), .A2(_05876_ ), .A3(_01205_ ), .ZN(_01307_ ) );
AND2_X1 _17130_ ( .A1(_01306_ ), .A2(_01307_ ), .ZN(_01308_ ) );
OAI21_X1 _17131_ ( .A(_01305_ ), .B1(_01308_ ), .B2(_01195_ ), .ZN(_01309_ ) );
MUX2_X1 _17132_ ( .A(_01309_ ), .B(_01303_ ), .S(_01201_ ), .Z(_01310_ ) );
MUX2_X1 _17133_ ( .A(_01303_ ), .B(_01310_ ), .S(_01210_ ), .Z(_01311_ ) );
MUX2_X1 _17134_ ( .A(\EX_LS_result_reg [4] ), .B(_01311_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
NOR3_X1 _17135_ ( .A1(_00469_ ), .A2(_05875_ ), .A3(_01188_ ), .ZN(_01312_ ) );
INV_X1 _17136_ ( .A(_01312_ ), .ZN(_01313_ ) );
AND3_X1 _17137_ ( .A1(_00444_ ), .A2(_01884_ ), .A3(_01215_ ), .ZN(_01314_ ) );
OR4_X1 _17138_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(_00415_ ), .A3(_05915_ ), .A4(_05875_ ), .ZN(_01315_ ) );
OAI21_X1 _17139_ ( .A(_01315_ ), .B1(_01213_ ), .B2(_01266_ ), .ZN(_01316_ ) );
AOI21_X1 _17140_ ( .A(_01314_ ), .B1(_01316_ ), .B2(_01301_ ), .ZN(_01317_ ) );
OAI21_X1 _17141_ ( .A(_01313_ ), .B1(_01317_ ), .B2(_01187_ ), .ZN(_01318_ ) );
NOR3_X1 _17142_ ( .A1(_00415_ ), .A2(_05876_ ), .A3(_01187_ ), .ZN(_01319_ ) );
OAI21_X1 _17143_ ( .A(_01195_ ), .B1(_01312_ ), .B2(_01319_ ), .ZN(_01320_ ) );
OAI21_X1 _17144_ ( .A(_01206_ ), .B1(_01312_ ), .B2(_01319_ ), .ZN(_01321_ ) );
OR3_X1 _17145_ ( .A1(_00469_ ), .A2(_05876_ ), .A3(_01205_ ), .ZN(_01322_ ) );
AND2_X1 _17146_ ( .A1(_01321_ ), .A2(_01322_ ), .ZN(_01323_ ) );
OAI21_X1 _17147_ ( .A(_01320_ ), .B1(_01323_ ), .B2(_01195_ ), .ZN(_01324_ ) );
MUX2_X1 _17148_ ( .A(_01324_ ), .B(_01318_ ), .S(_01201_ ), .Z(_01325_ ) );
MUX2_X1 _17149_ ( .A(_01318_ ), .B(_01325_ ), .S(_01210_ ), .Z(_01326_ ) );
MUX2_X1 _17150_ ( .A(\EX_LS_result_reg [3] ), .B(_01326_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
OR3_X1 _17151_ ( .A1(_00472_ ), .A2(_05876_ ), .A3(_01188_ ), .ZN(_01327_ ) );
AND3_X1 _17152_ ( .A1(_00447_ ), .A2(_01884_ ), .A3(_01215_ ), .ZN(_01328_ ) );
NOR2_X1 _17153_ ( .A1(_00487_ ), .A2(_05876_ ), .ZN(_01329_ ) );
MUX2_X1 _17154_ ( .A(_01329_ ), .B(_01230_ ), .S(_01213_ ), .Z(_01330_ ) );
AOI21_X1 _17155_ ( .A(_01328_ ), .B1(_01330_ ), .B2(_01301_ ), .ZN(_01331_ ) );
OAI21_X1 _17156_ ( .A(_01327_ ), .B1(_01331_ ), .B2(_01187_ ), .ZN(_01332_ ) );
NOR2_X2 _17157_ ( .A1(_00472_ ), .A2(_05875_ ), .ZN(_01333_ ) );
MUX2_X2 _17158_ ( .A(_01333_ ), .B(_01230_ ), .S(_01188_ ), .Z(_01334_ ) );
MUX2_X2 _17159_ ( .A(_01333_ ), .B(_01334_ ), .S(_01206_ ), .Z(_01335_ ) );
INV_X1 _17160_ ( .A(_01195_ ), .ZN(_01336_ ) );
MUX2_X1 _17161_ ( .A(_01334_ ), .B(_01335_ ), .S(_01336_ ), .Z(_01337_ ) );
INV_X1 _17162_ ( .A(_01201_ ), .ZN(_01338_ ) );
MUX2_X1 _17163_ ( .A(_01332_ ), .B(_01337_ ), .S(_01338_ ), .Z(_01339_ ) );
MUX2_X1 _17164_ ( .A(_01332_ ), .B(_01339_ ), .S(_01210_ ), .Z(_01340_ ) );
MUX2_X1 _17165_ ( .A(\EX_LS_result_reg [2] ), .B(_01340_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
AOI211_X1 _17166_ ( .A(_05877_ ), .B(_01192_ ), .C1(_00440_ ), .C2(_00441_ ), .ZN(_01341_ ) );
OAI21_X1 _17167_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01341_ ), .ZN(_01342_ ) );
OAI21_X1 _17168_ ( .A(_01342_ ), .B1(_01211_ ), .B2(_01238_ ), .ZN(_01343_ ) );
MUX2_X1 _17169_ ( .A(\EX_LS_result_reg [29] ), .B(_01343_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
OR3_X1 _17170_ ( .A1(_00478_ ), .A2(_05876_ ), .A3(_01188_ ), .ZN(_01344_ ) );
AND4_X1 _17171_ ( .A1(_01884_ ), .A2(_00448_ ), .A3(_00450_ ), .A4(_01215_ ), .ZN(_01345_ ) );
NOR2_X1 _17172_ ( .A1(_00490_ ), .A2(_05875_ ), .ZN(_01346_ ) );
NOR2_X1 _17173_ ( .A1(_00422_ ), .A2(_05875_ ), .ZN(_01347_ ) );
MUX2_X1 _17174_ ( .A(_01346_ ), .B(_01347_ ), .S(_01213_ ), .Z(_01348_ ) );
AOI21_X1 _17175_ ( .A(_01345_ ), .B1(_01348_ ), .B2(_01301_ ), .ZN(_01349_ ) );
OAI21_X1 _17176_ ( .A(_01344_ ), .B1(_01349_ ), .B2(_01187_ ), .ZN(_01350_ ) );
NOR2_X1 _17177_ ( .A1(_00478_ ), .A2(_05875_ ), .ZN(_01351_ ) );
MUX2_X2 _17178_ ( .A(_01347_ ), .B(_01351_ ), .S(_01187_ ), .Z(_01352_ ) );
MUX2_X2 _17179_ ( .A(_01351_ ), .B(_01352_ ), .S(_01205_ ), .Z(_01353_ ) );
MUX2_X1 _17180_ ( .A(_01352_ ), .B(_01353_ ), .S(_01336_ ), .Z(_01354_ ) );
MUX2_X1 _17181_ ( .A(_01350_ ), .B(_01354_ ), .S(_01338_ ), .Z(_01355_ ) );
MUX2_X1 _17182_ ( .A(_01350_ ), .B(_01355_ ), .S(_01210_ ), .Z(_01356_ ) );
MUX2_X1 _17183_ ( .A(\EX_LS_result_reg [1] ), .B(_01356_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
AOI211_X1 _17184_ ( .A(_05969_ ), .B(_05879_ ), .C1(_00705_ ), .C2(_01287_ ), .ZN(_01357_ ) );
NAND2_X1 _17185_ ( .A1(_00481_ ), .A2(_01285_ ), .ZN(_01358_ ) );
NAND2_X1 _17186_ ( .A1(_01357_ ), .A2(_01358_ ), .ZN(_01359_ ) );
NAND3_X1 _17187_ ( .A1(_00491_ ), .A2(\mylsu.araddr_tmp [1] ), .A3(_00493_ ), .ZN(_01360_ ) );
NAND3_X1 _17188_ ( .A1(_00451_ ), .A2(_05915_ ), .A3(_00453_ ), .ZN(_01361_ ) );
AND3_X1 _17189_ ( .A1(_01360_ ), .A2(_01361_ ), .A3(_01282_ ), .ZN(_01362_ ) );
OAI22_X1 _17190_ ( .A1(_01359_ ), .A2(_01362_ ), .B1(fanout_net_44 ), .B2(_04463_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
NOR3_X1 _17191_ ( .A1(_00475_ ), .A2(_05878_ ), .A3(_01206_ ), .ZN(_01363_ ) );
OAI21_X1 _17192_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01363_ ), .ZN(_01364_ ) );
OAI21_X1 _17193_ ( .A(_01364_ ), .B1(_01211_ ), .B2(_01238_ ), .ZN(_01365_ ) );
MUX2_X1 _17194_ ( .A(\EX_LS_result_reg [28] ), .B(_01365_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
OR3_X1 _17195_ ( .A1(_00484_ ), .A2(_05877_ ), .A3(_01206_ ), .ZN(_01366_ ) );
AOI211_X1 _17196_ ( .A(_01202_ ), .B(_01196_ ), .C1(_01336_ ), .C2(_01366_ ), .ZN(_01367_ ) );
OAI21_X1 _17197_ ( .A(fanout_net_44 ), .B1(_01367_ ), .B2(_01240_ ), .ZN(_01368_ ) );
OAI21_X1 _17198_ ( .A(_01368_ ), .B1(fanout_net_44 ), .B2(_04361_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
NOR3_X1 _17199_ ( .A1(_00487_ ), .A2(_05878_ ), .A3(_01206_ ), .ZN(_01369_ ) );
OAI21_X1 _17200_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01369_ ), .ZN(_01370_ ) );
OAI21_X1 _17201_ ( .A(_01370_ ), .B1(_01211_ ), .B2(_01238_ ), .ZN(_01371_ ) );
MUX2_X1 _17202_ ( .A(\EX_LS_result_reg [26] ), .B(_01371_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
OAI21_X1 _17203_ ( .A(_01229_ ), .B1(_01192_ ), .B2(_01346_ ), .ZN(_01372_ ) );
AOI22_X1 _17204_ ( .A1(_01372_ ), .A2(_01241_ ), .B1(_05969_ ), .B2(_04411_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
AND4_X1 _17205_ ( .A1(\io_master_arid [1] ), .A2(_00491_ ), .A3(_00493_ ), .A4(_01242_ ), .ZN(_01373_ ) );
OAI21_X1 _17206_ ( .A(_01204_ ), .B1(_01222_ ), .B2(_01373_ ), .ZN(_01374_ ) );
OAI21_X1 _17207_ ( .A(_01374_ ), .B1(_01252_ ), .B2(_01238_ ), .ZN(_01375_ ) );
MUX2_X1 _17208_ ( .A(\EX_LS_result_reg [24] ), .B(_01375_ ), .S(fanout_net_44 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
OAI21_X1 _17209_ ( .A(_01229_ ), .B1(_01192_ ), .B2(_01212_ ), .ZN(_01376_ ) );
AOI22_X1 _17210_ ( .A1(_01376_ ), .A2(_01241_ ), .B1(_05969_ ), .B2(_04015_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
AND4_X1 _17211_ ( .A1(\io_master_arid [1] ), .A2(_00497_ ), .A3(_00499_ ), .A4(_01207_ ), .ZN(_01377_ ) );
OAI21_X1 _17212_ ( .A(_01203_ ), .B1(_01222_ ), .B2(_01377_ ), .ZN(_01378_ ) );
OAI21_X1 _17213_ ( .A(_01378_ ), .B1(_01252_ ), .B2(_01238_ ), .ZN(_01379_ ) );
MUX2_X1 _17214_ ( .A(\EX_LS_result_reg [22] ), .B(_01379_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17215_ ( .A1(_00396_ ), .A2(\io_master_arid [1] ), .A3(_01242_ ), .ZN(_01380_ ) );
OAI21_X1 _17216_ ( .A(_01203_ ), .B1(_01195_ ), .B2(_01380_ ), .ZN(_01381_ ) );
OAI21_X1 _17217_ ( .A(_01381_ ), .B1(_01252_ ), .B2(_01238_ ), .ZN(_01382_ ) );
MUX2_X1 _17218_ ( .A(\EX_LS_result_reg [31] ), .B(_01382_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
INV_X1 _17219_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01383_ ) );
NOR2_X1 _17220_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(\LS_WB_waddr_reg [2] ), .ZN(_01384_ ) );
INV_X1 _17221_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01385_ ) );
INV_X1 _17222_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01386_ ) );
NAND3_X1 _17223_ ( .A1(_01384_ ), .A2(_01385_ ), .A3(_01386_ ), .ZN(_01387_ ) );
AND2_X1 _17224_ ( .A1(_01459_ ), .A2(LS_WB_wen_reg ), .ZN(_01388_ ) );
NAND2_X1 _17225_ ( .A1(_01387_ ), .A2(_01388_ ), .ZN(_01389_ ) );
BUF_X4 _17226_ ( .A(_01389_ ), .Z(_01390_ ) );
NOR2_X1 _17227_ ( .A1(_01390_ ), .A2(_01386_ ), .ZN(_01391_ ) );
INV_X1 _17228_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01392_ ) );
NOR2_X1 _17229_ ( .A1(_01390_ ), .A2(_01392_ ), .ZN(_01393_ ) );
AND4_X1 _17230_ ( .A1(_01383_ ), .A2(_01391_ ), .A3(_01393_ ), .A4(_01385_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _17231_ ( .A1(_01389_ ), .A2(_01385_ ), .ZN(_01394_ ) );
AND4_X1 _17232_ ( .A1(_01383_ ), .A2(_01394_ ), .A3(_01393_ ), .A4(_01386_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
AOI21_X1 _17233_ ( .A(_01390_ ), .B1(_01385_ ), .B2(_01386_ ), .ZN(_01395_ ) );
NOR4_X1 _17234_ ( .A1(_01395_ ), .A2(_01383_ ), .A3(_01392_ ), .A4(_01390_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
CLKBUF_X1 _17235_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
AOI21_X1 _17236_ ( .A(_01390_ ), .B1(_01383_ ), .B2(_01392_ ), .ZN(_01396_ ) );
NOR4_X1 _17237_ ( .A1(_01396_ ), .A2(_01394_ ), .A3(_01386_ ), .A4(_01390_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
NOR4_X1 _17238_ ( .A1(_01396_ ), .A2(_01391_ ), .A3(_01385_ ), .A4(_01390_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17239_ ( .A1(_01396_ ), .A2(_01385_ ), .A3(_01386_ ), .A4(_01390_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17240_ ( .A1(_01383_ ), .A2(_01394_ ), .A3(_01393_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
NOR4_X1 _17241_ ( .A1(_01395_ ), .A2(_01393_ ), .A3(_01383_ ), .A4(_01390_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR2_X1 _17242_ ( .A1(_01389_ ), .A2(_01383_ ), .ZN(_01397_ ) );
AND4_X1 _17243_ ( .A1(_01392_ ), .A2(_01391_ ), .A3(_01397_ ), .A4(_01385_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17244_ ( .A1(_01392_ ), .A2(_01394_ ), .A3(_01397_ ), .A4(_01386_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17245_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01391_ ), .A3(_01397_ ), .A4(_01385_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17246_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01394_ ), .A3(_01397_ ), .A4(_01386_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17247_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(_01394_ ), .A3(_01393_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17248_ ( .A1(_01392_ ), .A2(_01394_ ), .A3(_01397_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17249_ ( .A1(_01395_ ), .A2(_01397_ ), .A3(_01392_ ), .A4(_01390_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17250_ ( .A1(_01867_ ), .A2(_01545_ ), .A3(_01876_ ), .ZN(_01398_ ) );
NAND2_X1 _17251_ ( .A1(_01398_ ), .A2(_01545_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17252_ ( .A(reset ), .B(_01867_ ), .C1(_01868_ ), .C2(_05938_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17253_ ( .A(_01387_ ), .Z(_01399_ ) );
CLKBUF_X2 _17254_ ( .A(_01388_ ), .Z(_01400_ ) );
AND3_X1 _17255_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17256_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17257_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17258_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17259_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17260_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17261_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17262_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17263_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17264_ ( .A1(_01399_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01400_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17265_ ( .A(_01387_ ), .Z(_01401_ ) );
CLKBUF_X2 _17266_ ( .A(_01388_ ), .Z(_01402_ ) );
AND3_X1 _17267_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17268_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17269_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17270_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17271_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17272_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17273_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17274_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17275_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17276_ ( .A1(_01401_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01402_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17277_ ( .A(_01387_ ), .Z(_01403_ ) );
CLKBUF_X2 _17278_ ( .A(_01388_ ), .Z(_01404_ ) );
AND3_X1 _17279_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17280_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17281_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17282_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17283_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17284_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17285_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17286_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17287_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17288_ ( .A1(_01403_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01404_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17289_ ( .A1(_01387_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01388_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17290_ ( .A1(_01387_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01388_ ), .ZN(\myreg.Reg[6]_$_DFFE_PP__Q_D ) );
AND3_X1 _17291_ ( .A1(_01545_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17292_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01405_ ) );
AND2_X1 _17293_ ( .A1(_01405_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01406_ ) );
INV_X1 _17294_ ( .A(_01406_ ), .ZN(_01407_ ) );
NOR2_X1 _17295_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01408_ ) );
OAI211_X1 _17296_ ( .A(_01459_ ), .B(\mysc.state [0] ), .C1(_01407_ ), .C2(_01408_ ), .ZN(_01409_ ) );
INV_X1 _17297_ ( .A(_01409_ ), .ZN(_01410_ ) );
OR3_X1 _17298_ ( .A1(_01410_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17299_ ( .A1(_01407_ ), .A2(reset ), .A3(_01408_ ), .ZN(_01411_ ) );
NAND2_X1 _17300_ ( .A1(_01411_ ), .A2(\mysc.state [0] ), .ZN(_01412_ ) );
OR3_X1 _17301_ ( .A1(_03774_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01413_ ) );
NAND2_X1 _17302_ ( .A1(_01412_ ), .A2(_01413_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17303_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07884_ ) );
CLKGATE_X1 _17304_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07885_ ) );
CLKGATE_X1 _17305_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07886_ ) );
CLKGATE_X1 _17306_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07887_ ) );
CLKGATE_X1 _17307_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07888_ ) );
CLKGATE_X1 _17308_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_07889_ ) );
CLKGATE_X1 _17309_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_07890_ ) );
CLKGATE_X1 _17310_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_07891_ ) );
CLKGATE_X1 _17311_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_07892_ ) );
CLKGATE_X1 _17312_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_07893_ ) );
CLKGATE_X1 _17313_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_07894_ ) );
CLKGATE_X1 _17314_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07895_ ) );
CLKGATE_X1 _17315_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07896_ ) );
CLKGATE_X1 _17316_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_07897_ ) );
CLKGATE_X1 _17317_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_07898_ ) );
CLKGATE_X1 _17318_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07899_ ) );
CLKGATE_X1 _17319_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07900_ ) );
CLKGATE_X1 _17320_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_07901_ ) );
CLKGATE_X1 _17321_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_07902_ ) );
CLKGATE_X1 _17322_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ), .GCK(_07903_ ) );
CLKGATE_X1 _17323_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .GCK(_07904_ ) );
CLKGATE_X1 _17324_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07905_ ) );
CLKGATE_X1 _17325_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_07906_ ) );
CLKGATE_X1 _17326_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_07907_ ) );
CLKGATE_X1 _17327_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_07908_ ) );
CLKGATE_X1 _17328_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_07909_ ) );
CLKGATE_X1 _17329_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_07910_ ) );
CLKGATE_X1 _17330_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_07911_ ) );
CLKGATE_X1 _17331_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_07912_ ) );
CLKGATE_X1 _17332_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_07913_ ) );
CLKGATE_X1 _17333_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_07914_ ) );
CLKGATE_X1 _17334_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_07915_ ) );
CLKGATE_X1 _17335_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_07916_ ) );
CLKGATE_X1 _17336_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_07917_ ) );
CLKGATE_X1 _17337_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_07918_ ) );
CLKGATE_X1 _17338_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07919_ ) );
CLKGATE_X1 _17339_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07920_ ) );
CLKGATE_X1 _17340_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07921_ ) );
CLKGATE_X1 _17341_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07922_ ) );
CLKGATE_X1 _17342_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07923_ ) );
CLKGATE_X1 _17343_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07924_ ) );
CLKGATE_X1 _17344_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07925_ ) );
CLKGATE_X1 _17345_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07926_ ) );
CLKGATE_X1 _17346_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07927_ ) );
CLKGATE_X1 _17347_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_07928_ ) );
CLKGATE_X1 _17348_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_07929_ ) );
CLKGATE_X1 _17349_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_07930_ ) );
CLKGATE_X1 _17350_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_07931_ ) );
CLKGATE_X1 _17351_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07932_ ) );
CLKGATE_X1 _17352_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07933_ ) );
CLKGATE_X1 _17353_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07934_ ) );
CLKGATE_X1 _17354_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_07935_ ) );
CLKGATE_X1 _17355_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07936_ ) );
CLKGATE_X1 _17356_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_07937_ ) );
CLKGATE_X1 _17357_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_07938_ ) );
CLKGATE_X1 _17358_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_07939_ ) );
CLKGATE_X1 _17359_ ( .CK(clock ), .E(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07940_ ) );
CLKGATE_X1 _17360_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_07941_ ) );
CLKGATE_X1 _17361_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ), .GCK(_07942_ ) );
CLKGATE_X1 _17362_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_07943_ ) );
CLKGATE_X1 _17363_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07944_ ) );
CLKGATE_X1 _17364_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07945_ ) );
CLKGATE_X1 _17365_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07946_ ) );
CLKGATE_X1 _17366_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07947_ ) );
CLKGATE_X1 _17367_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07948_ ) );
LOGIC1_X1 _17368_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17369_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08178_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08179_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08180_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08181_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08182_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08183_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08184_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08185_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08186_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08187_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08188_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08189_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08190_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08191_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08192_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08193_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08194_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08195_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08196_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08197_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08198_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08199_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08200_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08201_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08202_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08203_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08204_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08205_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08206_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08207_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08208_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07948_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08209_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07947_ ), .Q(\mtvec [31] ), .QN(_08210_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07947_ ), .Q(\mtvec [30] ), .QN(_08211_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07947_ ), .Q(\mtvec [21] ), .QN(_08212_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07947_ ), .Q(\mtvec [20] ), .QN(_08213_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07947_ ), .Q(\mtvec [19] ), .QN(_08214_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07947_ ), .Q(\mtvec [18] ), .QN(_08215_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07947_ ), .Q(\mtvec [17] ), .QN(_08216_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07947_ ), .Q(\mtvec [16] ), .QN(_08217_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07947_ ), .Q(\mtvec [15] ), .QN(_08218_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07947_ ), .Q(\mtvec [14] ), .QN(_08219_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07947_ ), .Q(\mtvec [13] ), .QN(_08220_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07947_ ), .Q(\mtvec [12] ), .QN(_08221_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07947_ ), .Q(\mtvec [29] ), .QN(_08222_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07947_ ), .Q(\mtvec [11] ), .QN(_08223_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07947_ ), .Q(\mtvec [10] ), .QN(_08224_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07947_ ), .Q(\mtvec [9] ), .QN(_08225_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07947_ ), .Q(\mtvec [8] ), .QN(_08226_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07947_ ), .Q(\mtvec [7] ), .QN(_08227_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07947_ ), .Q(\mtvec [6] ), .QN(_08228_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07947_ ), .Q(\mtvec [5] ), .QN(_08229_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07947_ ), .Q(\mtvec [4] ), .QN(_08230_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07947_ ), .Q(\mtvec [3] ), .QN(_08231_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07947_ ), .Q(\mtvec [2] ), .QN(_08232_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07947_ ), .Q(\mtvec [28] ), .QN(_08233_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07947_ ), .Q(\mtvec [1] ), .QN(_08234_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07947_ ), .Q(\mtvec [0] ), .QN(_08235_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07947_ ), .Q(\mtvec [27] ), .QN(_08236_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07947_ ), .Q(\mtvec [26] ), .QN(_08237_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07947_ ), .Q(\mtvec [25] ), .QN(_08238_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07947_ ), .Q(\mtvec [24] ), .QN(_08239_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07947_ ), .Q(\mtvec [23] ), .QN(_08240_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07947_ ), .Q(\mtvec [22] ), .QN(_08241_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07946_ ), .Q(\mepc [31] ), .QN(_08242_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07946_ ), .Q(\mepc [30] ), .QN(_08243_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07946_ ), .Q(\mepc [21] ), .QN(_08244_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07946_ ), .Q(\mepc [20] ), .QN(_08245_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07946_ ), .Q(\mepc [19] ), .QN(_08246_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07946_ ), .Q(\mepc [18] ), .QN(_08247_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07946_ ), .Q(\mepc [17] ), .QN(_08248_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07946_ ), .Q(\mepc [16] ), .QN(_08249_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07946_ ), .Q(\mepc [15] ), .QN(_08250_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07946_ ), .Q(\mepc [14] ), .QN(_08251_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07946_ ), .Q(\mepc [13] ), .QN(_08252_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07946_ ), .Q(\mepc [12] ), .QN(_08253_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07946_ ), .Q(\mepc [29] ), .QN(_08254_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07946_ ), .Q(\mepc [11] ), .QN(_08255_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07946_ ), .Q(\mepc [10] ), .QN(_08256_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07946_ ), .Q(\mepc [9] ), .QN(_08257_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07946_ ), .Q(\mepc [8] ), .QN(_08258_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07946_ ), .Q(\mepc [7] ), .QN(_08259_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07946_ ), .Q(\mepc [6] ), .QN(_08260_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07946_ ), .Q(\mepc [5] ), .QN(_08261_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07946_ ), .Q(\mepc [4] ), .QN(_08262_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07946_ ), .Q(\mepc [3] ), .QN(_08263_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07946_ ), .Q(\mepc [2] ), .QN(_08264_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07946_ ), .Q(\mepc [28] ), .QN(_08265_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07946_ ), .Q(\mepc [1] ), .QN(_08266_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07946_ ), .Q(\mepc [0] ), .QN(_08267_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07946_ ), .Q(\mepc [27] ), .QN(_08268_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07946_ ), .Q(\mepc [26] ), .QN(_08269_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07946_ ), .Q(\mepc [25] ), .QN(_08270_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07946_ ), .Q(\mepc [24] ), .QN(_08271_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07946_ ), .Q(\mepc [23] ), .QN(_08272_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07946_ ), .Q(\mepc [22] ), .QN(_08273_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08274_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08275_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08276_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08177_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08176_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08175_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08174_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08173_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08172_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08171_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08170_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08169_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08168_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08167_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08166_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08165_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08164_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08163_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08162_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08161_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08160_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08159_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08158_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08157_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08156_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00086_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08155_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00087_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08154_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00088_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08153_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00089_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08152_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00090_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08151_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00091_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08150_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00092_ ), .CK(_07945_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08277_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PP0__Q ( .D(_00093_ ), .CK(clock ), .Q(excp_written ), .QN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08149_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08278_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08279_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08280_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08281_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08282_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08283_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08284_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08285_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08286_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08287_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08288_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08289_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08290_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08291_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08292_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08293_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08294_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08295_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08296_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08297_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08298_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08299_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08300_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08301_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08302_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08303_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08304_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08305_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08306_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08307_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_07944_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08148_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00094_ ), .CK(_07943_ ), .Q(\myec.state [1] ), .QN(_08147_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00095_ ), .CK(_07943_ ), .Q(\myec.state [0] ), .QN(_08308_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PN0__Q ( .D(_00096_ ), .CK(clock ), .Q(check_quest ), .QN(_08309_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08146_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08310_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08311_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08312_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08313_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08314_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08315_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08316_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08317_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08318_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08319_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08145_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00097_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08144_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00098_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08143_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00099_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08142_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00100_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08141_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00101_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08140_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00102_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08139_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00103_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08138_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00104_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08137_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00105_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08136_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00106_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08135_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00107_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08134_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00108_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08133_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00109_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08132_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00110_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08131_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00111_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08130_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00112_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08129_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00113_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08128_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00114_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08127_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00115_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08126_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00116_ ), .CK(_07942_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08125_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q ( .D(_00117_ ), .CK(_07941_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08124_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_1 ( .D(_00118_ ), .CK(_07941_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08123_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_2 ( .D(_00119_ ), .CK(_07941_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08122_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_3 ( .D(_00120_ ), .CK(_07941_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08121_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_4 ( .D(_00121_ ), .CK(_07941_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08120_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q ( .D(_00122_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [30] ), .QN(_08119_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_1 ( .D(_00123_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [29] ), .QN(_08118_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_10 ( .D(_00124_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [20] ), .QN(_08117_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_11 ( .D(_00125_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [19] ), .QN(_08116_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_12 ( .D(_00126_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [18] ), .QN(_08115_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_13 ( .D(_00127_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [17] ), .QN(_08114_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_14 ( .D(_00128_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [16] ), .QN(_08113_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_15 ( .D(_00129_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [15] ), .QN(_08112_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_16 ( .D(_00130_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [14] ), .QN(_08111_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_17 ( .D(_00131_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [13] ), .QN(_08110_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_18 ( .D(_00132_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [12] ), .QN(_08109_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_19 ( .D(_00133_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [11] ), .QN(_08108_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_2 ( .D(_00134_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [28] ), .QN(_08107_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_20 ( .D(_00135_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [10] ), .QN(_08106_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_21 ( .D(_00136_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [9] ), .QN(_08105_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_22 ( .D(_00137_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [8] ), .QN(_08104_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_23 ( .D(_00138_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [7] ), .QN(_08103_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_24 ( .D(_00139_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [6] ), .QN(_08102_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_25 ( .D(_00140_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [5] ), .QN(_08101_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_26 ( .D(_00141_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [4] ), .QN(_08100_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_27 ( .D(_00142_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [3] ), .QN(_08099_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_28 ( .D(_00143_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [2] ), .QN(_08098_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_29 ( .D(_00144_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [1] ), .QN(_08097_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_3 ( .D(_00145_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [27] ), .QN(_08096_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_30 ( .D(_00146_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [0] ), .QN(_08095_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_4 ( .D(_00147_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [26] ), .QN(_08094_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_5 ( .D(_00148_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [25] ), .QN(_08093_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_6 ( .D(_00149_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [24] ), .QN(_08092_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_7 ( .D(_00150_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [23] ), .QN(_08091_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_8 ( .D(_00151_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [22] ), .QN(_08090_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_9 ( .D(_00152_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [21] ), .QN(_08089_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN1P__Q ( .D(_00153_ ), .CK(_07940_ ), .Q(\myexu.pc_jump [31] ), .QN(_08088_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q ( .D(_00154_ ), .CK(_07941_ ), .Q(\EX_LS_pc [31] ), .QN(_08087_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_1 ( .D(_00155_ ), .CK(_07941_ ), .Q(\EX_LS_pc [30] ), .QN(_08086_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_10 ( .D(_00156_ ), .CK(_07941_ ), .Q(\EX_LS_pc [21] ), .QN(_08085_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_11 ( .D(_00157_ ), .CK(_07941_ ), .Q(\EX_LS_pc [20] ), .QN(_08084_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_12 ( .D(_00158_ ), .CK(_07941_ ), .Q(\EX_LS_pc [19] ), .QN(_08083_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_13 ( .D(_00159_ ), .CK(_07941_ ), .Q(\EX_LS_pc [18] ), .QN(_08082_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_14 ( .D(_00160_ ), .CK(_07941_ ), .Q(\EX_LS_pc [17] ), .QN(_08081_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_15 ( .D(_00161_ ), .CK(_07941_ ), .Q(\EX_LS_pc [16] ), .QN(_08080_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_16 ( .D(_00162_ ), .CK(_07941_ ), .Q(\EX_LS_pc [15] ), .QN(_08079_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_17 ( .D(_00163_ ), .CK(_07941_ ), .Q(\EX_LS_pc [14] ), .QN(_08078_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_18 ( .D(_00164_ ), .CK(_07941_ ), .Q(\EX_LS_pc [13] ), .QN(_08077_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_19 ( .D(_00165_ ), .CK(_07941_ ), .Q(\EX_LS_pc [12] ), .QN(_08076_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_2 ( .D(_00166_ ), .CK(_07941_ ), .Q(\EX_LS_pc [29] ), .QN(_08075_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_20 ( .D(_00167_ ), .CK(_07941_ ), .Q(\EX_LS_pc [11] ), .QN(_08074_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_21 ( .D(_00168_ ), .CK(_07941_ ), .Q(\EX_LS_pc [10] ), .QN(_08073_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_22 ( .D(_00169_ ), .CK(_07941_ ), .Q(\EX_LS_pc [9] ), .QN(_08072_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_23 ( .D(_00170_ ), .CK(_07941_ ), .Q(\EX_LS_pc [8] ), .QN(_08071_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_24 ( .D(_00171_ ), .CK(_07941_ ), .Q(\EX_LS_pc [7] ), .QN(_08070_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_25 ( .D(_00172_ ), .CK(_07941_ ), .Q(\EX_LS_pc [6] ), .QN(_08069_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_26 ( .D(_00173_ ), .CK(_07941_ ), .Q(\EX_LS_pc [5] ), .QN(_08068_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_27 ( .D(_00174_ ), .CK(_07941_ ), .Q(\EX_LS_pc [4] ), .QN(_08067_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_28 ( .D(_00175_ ), .CK(_07941_ ), .Q(\EX_LS_pc [3] ), .QN(_08066_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_29 ( .D(_00176_ ), .CK(_07941_ ), .Q(\EX_LS_pc [2] ), .QN(_08065_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_3 ( .D(_00177_ ), .CK(_07941_ ), .Q(\EX_LS_pc [28] ), .QN(_08064_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_30 ( .D(_00178_ ), .CK(_07941_ ), .Q(\EX_LS_pc [1] ), .QN(_08063_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_31 ( .D(_00179_ ), .CK(_07941_ ), .Q(\EX_LS_pc [0] ), .QN(_08062_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_4 ( .D(_00180_ ), .CK(_07941_ ), .Q(\EX_LS_pc [27] ), .QN(_08061_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_5 ( .D(_00181_ ), .CK(_07941_ ), .Q(\EX_LS_pc [26] ), .QN(_08060_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_6 ( .D(_00182_ ), .CK(_07941_ ), .Q(\EX_LS_pc [25] ), .QN(_08059_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_7 ( .D(_00183_ ), .CK(_07941_ ), .Q(\EX_LS_pc [24] ), .QN(_08058_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_8 ( .D(_00184_ ), .CK(_07941_ ), .Q(\EX_LS_pc [23] ), .QN(_08057_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_9 ( .D(_00185_ ), .CK(_07941_ ), .Q(\EX_LS_pc [22] ), .QN(_08320_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08321_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08322_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08323_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08324_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08325_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08326_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08327_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08328_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08329_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08330_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08331_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08332_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08333_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08334_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08335_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08336_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08337_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08338_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08339_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08340_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08341_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08342_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08343_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08344_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08345_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08346_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08347_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08348_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08349_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08350_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08351_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07942_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08352_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_07942_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PN0__Q ( .D(_00187_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q ( .D(_00186_ ), .CK(_07941_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_1 ( .D(_00188_ ), .CK(_07941_ ), .Q(\EX_LS_flag [1] ), .QN(_08056_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_2 ( .D(_00189_ ), .CK(_07941_ ), .Q(\EX_LS_flag [0] ), .QN(_08055_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_3 ( .D(_00190_ ), .CK(_07941_ ), .Q(\EX_LS_typ [4] ), .QN(_08054_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_4 ( .D(_00191_ ), .CK(_07941_ ), .Q(\EX_LS_typ [3] ), .QN(_08053_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_5 ( .D(_00192_ ), .CK(_07941_ ), .Q(\EX_LS_typ [2] ), .QN(_08052_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_6 ( .D(_00193_ ), .CK(_07941_ ), .Q(\EX_LS_typ [1] ), .QN(_08051_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_7 ( .D(_00194_ ), .CK(_07941_ ), .Q(\EX_LS_typ [0] ), .QN(_08050_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00195_ ), .CK(_07939_ ), .Q(\ID_EX_csr [11] ), .QN(_08049_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00196_ ), .CK(_07939_ ), .Q(\ID_EX_csr [10] ), .QN(_08048_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00197_ ), .CK(_07939_ ), .Q(\ID_EX_csr [1] ), .QN(_08047_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00198_ ), .CK(_07939_ ), .Q(\ID_EX_csr [0] ), .QN(_08046_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00199_ ), .CK(_07939_ ), .Q(\ID_EX_csr [9] ), .QN(_08045_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00200_ ), .CK(_07939_ ), .Q(\ID_EX_csr [8] ), .QN(_08044_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00201_ ), .CK(_07939_ ), .Q(\ID_EX_csr [7] ), .QN(_08043_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00202_ ), .CK(_07939_ ), .Q(\ID_EX_csr [6] ), .QN(_08042_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00203_ ), .CK(_07939_ ), .Q(\ID_EX_csr [5] ), .QN(_08041_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00204_ ), .CK(_07939_ ), .Q(\ID_EX_csr [4] ), .QN(_08040_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00205_ ), .CK(_07939_ ), .Q(\ID_EX_csr [3] ), .QN(_08039_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00206_ ), .CK(_07939_ ), .Q(\ID_EX_csr [2] ), .QN(_08038_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00207_ ), .CK(_07938_ ), .Q(exception_quest_IDU ), .QN(_08037_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00208_ ), .CK(_07937_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_07936_ ), .Q(\ID_EX_imm [31] ), .QN(_08353_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_07936_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_07936_ ), .Q(\ID_EX_imm [21] ), .QN(_08354_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_07936_ ), .Q(\ID_EX_imm [20] ), .QN(_08355_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_07936_ ), .Q(\ID_EX_imm [19] ), .QN(_08356_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_07936_ ), .Q(\ID_EX_imm [18] ), .QN(_08357_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_07936_ ), .Q(\ID_EX_imm [17] ), .QN(_08358_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_07936_ ), .Q(\ID_EX_imm [16] ), .QN(_08359_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_07936_ ), .Q(\ID_EX_imm [15] ), .QN(_08360_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_07936_ ), .Q(\ID_EX_imm [14] ), .QN(_08361_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_07936_ ), .Q(\ID_EX_imm [13] ), .QN(_08362_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_07936_ ), .Q(\ID_EX_imm [12] ), .QN(_08363_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_07936_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_07936_ ), .Q(\ID_EX_imm [11] ), .QN(_08364_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_07936_ ), .Q(\ID_EX_imm [10] ), .QN(_08365_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_07936_ ), .Q(\ID_EX_imm [9] ), .QN(_08366_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_07936_ ), .Q(\ID_EX_imm [8] ), .QN(_08367_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_07936_ ), .Q(\ID_EX_imm [7] ), .QN(_08368_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_07936_ ), .Q(\ID_EX_imm [6] ), .QN(_08369_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_07936_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_07936_ ), .Q(\ID_EX_imm [4] ), .QN(_08370_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_07936_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_07936_ ), .Q(\ID_EX_imm [2] ), .QN(_08371_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_07936_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_07936_ ), .Q(\ID_EX_imm [1] ), .QN(_08372_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_07936_ ), .Q(\ID_EX_imm [0] ), .QN(_08373_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_07936_ ), .Q(\ID_EX_imm [27] ), .QN(_08374_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_07936_ ), .Q(\ID_EX_imm [26] ), .QN(_08375_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_07936_ ), .Q(\ID_EX_imm [25] ), .QN(_08376_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_07936_ ), .Q(\ID_EX_imm [24] ), .QN(_08377_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_07936_ ), .Q(\ID_EX_imm [23] ), .QN(_08378_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_07936_ ), .Q(\ID_EX_imm [22] ), .QN(_08379_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07935_ ), .Q(\ID_EX_pc [31] ), .QN(_08380_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07935_ ), .Q(\ID_EX_pc [30] ), .QN(_08381_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07935_ ), .Q(\ID_EX_pc [21] ), .QN(_08382_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07935_ ), .Q(\ID_EX_pc [20] ), .QN(_08383_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07935_ ), .Q(\ID_EX_pc [19] ), .QN(_08384_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07935_ ), .Q(\ID_EX_pc [18] ), .QN(_08385_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07935_ ), .Q(\ID_EX_pc [17] ), .QN(_08386_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07935_ ), .Q(\ID_EX_pc [16] ), .QN(_08387_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07935_ ), .Q(\ID_EX_pc [15] ), .QN(_08388_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07935_ ), .Q(\ID_EX_pc [14] ), .QN(_08389_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07935_ ), .Q(\ID_EX_pc [13] ), .QN(_08390_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07935_ ), .Q(\ID_EX_pc [12] ), .QN(_08391_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07935_ ), .Q(\ID_EX_pc [29] ), .QN(_08392_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07935_ ), .Q(\ID_EX_pc [11] ), .QN(_08393_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07935_ ), .Q(\ID_EX_pc [10] ), .QN(_08394_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07935_ ), .Q(\ID_EX_pc [9] ), .QN(_08395_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07935_ ), .Q(\ID_EX_pc [8] ), .QN(_08396_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07935_ ), .Q(\ID_EX_pc [7] ), .QN(_08397_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07935_ ), .Q(\ID_EX_pc [6] ), .QN(_08398_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07935_ ), .Q(\ID_EX_pc [5] ), .QN(_08399_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07935_ ), .Q(\ID_EX_pc [4] ), .QN(_08400_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_07935_ ), .Q(\ID_EX_pc [3] ), .QN(_08401_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_07935_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07935_ ), .Q(\ID_EX_pc [28] ), .QN(_08402_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_07935_ ), .Q(\ID_EX_pc [1] ), .QN(_08403_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_07935_ ), .Q(\ID_EX_pc [0] ), .QN(_08404_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07935_ ), .Q(\ID_EX_pc [27] ), .QN(_08405_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07935_ ), .Q(\ID_EX_pc [26] ), .QN(_08406_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07935_ ), .Q(\ID_EX_pc [25] ), .QN(_08407_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07935_ ), .Q(\ID_EX_pc [24] ), .QN(_08408_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07935_ ), .Q(\ID_EX_pc [23] ), .QN(_08409_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07935_ ), .Q(\ID_EX_pc [22] ), .QN(_08036_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00209_ ), .CK(_07934_ ), .Q(\ID_EX_rd [4] ), .QN(_08035_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00210_ ), .CK(_07934_ ), .Q(\ID_EX_rd [3] ), .QN(_08034_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00211_ ), .CK(_07934_ ), .Q(\ID_EX_rd [2] ), .QN(_08033_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00212_ ), .CK(_07934_ ), .Q(\ID_EX_rd [1] ), .QN(_08032_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00213_ ), .CK(_07934_ ), .Q(\ID_EX_rd [0] ), .QN(_08031_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00214_ ), .CK(_07933_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08030_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00215_ ), .CK(_07933_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08029_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00217_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08027_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00216_ ), .CK(_07933_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08028_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00219_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08025_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00218_ ), .CK(_07933_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08026_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00221_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08023_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00220_ ), .CK(_07933_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08024_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00223_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08021_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00222_ ), .CK(_07932_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08022_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00224_ ), .CK(_07932_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08020_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00226_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08018_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00225_ ), .CK(_07932_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08019_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00228_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08016_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00227_ ), .CK(_07932_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08017_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00230_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08014_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00229_ ), .CK(_07932_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08015_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00232_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08012_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_07931_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08013_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00233_ ), .CK(_07930_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08011_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08411_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00234_ ), .CK(_07929_ ), .Q(\ID_EX_typ [7] ), .QN(_08410_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00235_ ), .CK(_07929_ ), .Q(\ID_EX_typ [6] ), .QN(_08010_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00236_ ), .CK(_07929_ ), .Q(\ID_EX_typ [5] ), .QN(_08009_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00237_ ), .CK(_07929_ ), .Q(\ID_EX_typ [4] ), .QN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00238_ ), .CK(_07929_ ), .Q(\ID_EX_typ [3] ), .QN(_08008_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00239_ ), .CK(_07929_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00240_ ), .CK(_07929_ ), .Q(\ID_EX_typ [1] ), .QN(_08007_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00241_ ), .CK(_07929_ ), .Q(\ID_EX_typ [0] ), .QN(_08412_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_07928_ ), .Q(check_assert ), .QN(_08413_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_07927_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_07927_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_07927_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_07927_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_07927_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_07927_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_07927_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_07927_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_07927_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_07927_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_07927_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_07927_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_07927_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_07927_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_07927_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_07927_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_07927_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_07927_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_07927_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_07927_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_07927_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_07927_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_07927_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_07927_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_07927_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_07927_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_07927_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_07927_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_07927_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_07927_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_07927_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_07927_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08414_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08415_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08416_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08417_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08418_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08419_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08420_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08421_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08422_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08423_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08424_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08425_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08426_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08427_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08428_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08429_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08430_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08431_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08432_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08433_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08434_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08435_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08436_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08437_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08438_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08439_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08440_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08441_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08442_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08443_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08444_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07926_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08445_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08446_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08447_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08448_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08449_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08450_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08451_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08452_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08453_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08454_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08455_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08456_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08457_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08458_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08459_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08460_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08461_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08462_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08463_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08464_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08465_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08466_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08467_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08468_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08469_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08470_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08471_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08472_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08473_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08474_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08475_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08476_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07925_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08477_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08478_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08479_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08480_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08481_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08482_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08483_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08484_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08485_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08486_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08487_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08488_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08489_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08490_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08491_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08492_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08493_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08494_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08495_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08496_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08497_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08498_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08499_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08500_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08501_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08502_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08503_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08504_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08505_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08506_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08507_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08508_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07924_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08509_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08510_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08511_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08512_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08513_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08514_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08515_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08516_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08517_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08518_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08519_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08520_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08521_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08522_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08523_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08524_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08525_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08526_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08527_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08528_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08529_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08530_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08531_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08532_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08533_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08534_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08535_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08536_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08537_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08538_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08539_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08540_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07923_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08541_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08542_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08543_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08544_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08545_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08546_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08547_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08548_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08549_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08550_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08551_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08552_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08553_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08554_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08555_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08556_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08557_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08558_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08559_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08560_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08561_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08562_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08563_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08564_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08565_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08566_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08567_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07922_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07921_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07920_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07919_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07918_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07917_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07916_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07915_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08006_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00242_ ), .CK(_07914_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08005_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00243_ ), .CK(_07913_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08004_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00244_ ), .CK(_07912_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_07911_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08003_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_07910_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_07909_ ), .Q(\IF_ID_pc [30] ), .QN(_08002_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00247_ ), .CK(_07909_ ), .Q(\IF_ID_pc [21] ), .QN(_08001_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00248_ ), .CK(_07909_ ), .Q(\IF_ID_pc [20] ), .QN(_08000_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00249_ ), .CK(_07909_ ), .Q(\IF_ID_pc [19] ), .QN(_07999_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00250_ ), .CK(_07909_ ), .Q(\IF_ID_pc [18] ), .QN(_07998_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00251_ ), .CK(_07909_ ), .Q(\IF_ID_pc [17] ), .QN(_07997_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00252_ ), .CK(_07909_ ), .Q(\IF_ID_pc [16] ), .QN(_07996_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00253_ ), .CK(_07909_ ), .Q(\IF_ID_pc [15] ), .QN(_07995_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00254_ ), .CK(_07909_ ), .Q(\IF_ID_pc [14] ), .QN(_07994_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00255_ ), .CK(_07909_ ), .Q(\IF_ID_pc [13] ), .QN(_07993_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00256_ ), .CK(_07909_ ), .Q(\IF_ID_pc [12] ), .QN(_07992_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00257_ ), .CK(_07909_ ), .Q(\IF_ID_pc [29] ), .QN(_07991_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00258_ ), .CK(_07909_ ), .Q(\IF_ID_pc [11] ), .QN(_07990_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00259_ ), .CK(_07909_ ), .Q(\IF_ID_pc [10] ), .QN(_07989_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00260_ ), .CK(_07909_ ), .Q(\IF_ID_pc [9] ), .QN(_07988_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00261_ ), .CK(_07909_ ), .Q(\IF_ID_pc [8] ), .QN(_07987_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00262_ ), .CK(_07909_ ), .Q(\IF_ID_pc [7] ), .QN(_07986_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00263_ ), .CK(_07909_ ), .Q(\IF_ID_pc [6] ), .QN(_07985_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00264_ ), .CK(_07909_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00265_ ), .CK(_07909_ ), .Q(\IF_ID_pc [4] ), .QN(_07984_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00267_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_07983_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00266_ ), .CK(_07909_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00269_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_07981_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00268_ ), .CK(_07909_ ), .Q(\IF_ID_pc [2] ), .QN(_07982_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00270_ ), .CK(_07909_ ), .Q(\IF_ID_pc [28] ), .QN(_07980_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00271_ ), .CK(_07909_ ), .Q(\IF_ID_pc [1] ), .QN(_07979_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00272_ ), .CK(_07909_ ), .Q(\IF_ID_pc [27] ), .QN(_07978_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00273_ ), .CK(_07909_ ), .Q(\IF_ID_pc [26] ), .QN(_07977_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00274_ ), .CK(_07909_ ), .Q(\IF_ID_pc [25] ), .QN(_07976_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00275_ ), .CK(_07909_ ), .Q(\IF_ID_pc [24] ), .QN(_07975_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00276_ ), .CK(_07909_ ), .Q(\IF_ID_pc [23] ), .QN(_07974_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00277_ ), .CK(_07909_ ), .Q(\IF_ID_pc [22] ), .QN(_07973_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00278_ ), .CK(_07909_ ), .Q(\IF_ID_pc [31] ), .QN(_07972_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08779_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_07971_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00279_ ), .CK(_07908_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08778_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00281_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00280_ ), .CK(_07907_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_07970_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08780_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08781_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08782_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08783_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08784_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08785_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08786_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08787_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08788_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08789_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08790_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08791_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08792_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08793_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08794_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08795_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08796_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08797_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08798_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08799_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08800_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08801_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08802_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08803_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08804_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08805_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08806_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08807_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08808_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08809_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08810_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07906_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08811_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08812_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08813_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08814_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08815_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08816_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08817_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08818_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08819_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08820_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08821_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08822_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08823_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08824_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08825_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08826_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08827_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08828_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08829_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08830_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08831_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08832_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08833_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08834_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08835_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08836_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08837_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08838_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08839_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08840_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08841_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08842_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07905_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_07969_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PN0P__Q ( .D(_00282_ ), .CK(_07904_ ), .Q(LS_WB_pc ), .QN(_07968_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PN0P__Q ( .D(_00283_ ), .CK(_07903_ ), .Q(\mylsu.previous_load_done ), .QN(_08843_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08844_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08845_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08846_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(\mylsu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__A_B ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_07906_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_07906_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08847_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_07906_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_07967_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00284_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_07966_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00285_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_07965_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00286_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_07964_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00287_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_07963_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00288_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_07962_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00289_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_07961_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00290_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_07960_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00291_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_07959_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00292_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_07958_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00293_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_07957_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00294_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_07956_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00295_ ), .CK(_07906_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08848_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_07906_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08849_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_07906_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08850_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_07906_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08851_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_07906_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08852_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08853_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08854_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08855_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08856_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08857_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08858_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08859_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08860_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08861_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08862_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08863_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08864_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08865_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08866_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08867_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08868_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08869_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08870_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08871_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08872_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08873_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08874_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08875_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08876_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08877_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08878_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08879_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08880_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08881_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08882_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08883_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_07906_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08884_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08885_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_08886_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_08887_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_08888_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_08889_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_08890_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_08891_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_08892_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_08893_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_08894_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_08895_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_08896_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_08897_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_08898_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_08899_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_08900_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_08901_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_08902_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_08903_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_08904_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_08905_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_08906_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_08907_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_08908_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_08909_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_08910_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_08911_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_08912_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_08913_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_08914_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_08915_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_07902_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_07955_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q ( .D(_00296_ ), .CK(_07901_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(\myec.state_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A_$_OR__Y_B_$_ANDNOT__A_B_$_ANDNOT__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_B_$_OR__B_Y_$_OR__A_Y_$_OR__A_B ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_1 ( .D(_00297_ ), .CK(_07901_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_07954_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_2 ( .D(_00298_ ), .CK(_07901_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_07953_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_3 ( .D(_00299_ ), .CK(_07901_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_07952_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_4 ( .D(_00300_ ), .CK(_07901_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_07951_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_5 ( .D(_00301_ ), .CK(_07901_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_07950_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PN0P__Q ( .D(_00302_ ), .CK(_07901_ ), .Q(LS_WB_wen_reg ), .QN(_08916_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_08917_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_08918_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07900_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07899_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07898_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07897_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07896_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07895_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07894_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07893_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07892_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07891_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07890_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07889_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07888_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07887_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07886_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_1_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_10_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_11_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_12_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_13_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_14_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_15_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_16_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_17_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_18_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_19_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_2_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_20_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_21_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_22_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_23_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_24_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_25_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_26_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_27_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_28_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_29_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_3_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_30_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_31_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_4_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_5_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_6_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_7_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_8_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[6]_$_DFFE_PP__Q_9_D ), .CK(_07885_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00303_ ), .CK(_07884_ ), .Q(loaduse_clear ), .QN(_08919_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_08920_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_08921_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_07949_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\ID_EX_typ [2] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(fanout_net_24 ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(fanout_net_24 ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(fanout_net_37 ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(fanout_net_37 ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\myifu.to_reset ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(\mylsu.state [3] ), .Z(fanout_net_44 ) );

endmodule
