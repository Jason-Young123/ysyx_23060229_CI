//Generate the verilog at 2025-09-29T16:37:28 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire _09036_ ;
wire _09037_ ;
wire _09038_ ;
wire _09039_ ;
wire _09040_ ;
wire _09041_ ;
wire _09042_ ;
wire _09043_ ;
wire _09044_ ;
wire _09045_ ;
wire _09046_ ;
wire _09047_ ;
wire _09048_ ;
wire _09049_ ;
wire _09050_ ;
wire _09051_ ;
wire _09052_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[2]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire fanout_net_45 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

AND3_X4 _09053_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [1] ), .A3(\myclint.mtime [0] ), .ZN(_01535_ ) );
AND3_X1 _09054_ ( .A1(_01535_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01536_ ) );
AND3_X4 _09055_ ( .A1(_01536_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01537_ ) );
AND2_X2 _09056_ ( .A1(_01537_ ), .A2(\myclint.mtime [7] ), .ZN(_01538_ ) );
AND4_X1 _09057_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01539_ ) );
AND2_X1 _09058_ ( .A1(\myclint.mtime [8] ), .A2(\myclint.mtime [9] ), .ZN(_01540_ ) );
AND4_X1 _09059_ ( .A1(\myclint.mtime [10] ), .A2(_01539_ ), .A3(\myclint.mtime [11] ), .A4(_01540_ ), .ZN(_01541_ ) );
AND2_X1 _09060_ ( .A1(_01538_ ), .A2(_01541_ ), .ZN(_01542_ ) );
AND2_X1 _09061_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01543_ ) );
AND2_X1 _09062_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_01544_ ) );
NAND3_X1 _09063_ ( .A1(_01544_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01545_ ) );
NAND4_X1 _09064_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01546_ ) );
NOR2_X1 _09065_ ( .A1(_01545_ ), .A2(_01546_ ), .ZN(_01547_ ) );
AND2_X1 _09066_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01548_ ) );
AND2_X1 _09067_ ( .A1(\myclint.mtime [24] ), .A2(\myclint.mtime [25] ), .ZN(_01549_ ) );
AND3_X1 _09068_ ( .A1(_01549_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [27] ), .ZN(_01550_ ) );
AND4_X1 _09069_ ( .A1(_01543_ ), .A2(_01547_ ), .A3(_01548_ ), .A4(_01550_ ), .ZN(_01551_ ) );
NAND2_X1 _09070_ ( .A1(_01542_ ), .A2(_01551_ ), .ZN(_01552_ ) );
AND2_X1 _09071_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01553_ ) );
AND3_X1 _09072_ ( .A1(_01553_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01554_ ) );
AND2_X1 _09073_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01555_ ) );
AND3_X1 _09074_ ( .A1(_01555_ ), .A2(\myclint.mtime [42] ), .A3(\myclint.mtime [43] ), .ZN(_01556_ ) );
AND4_X1 _09075_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01557_ ) );
NAND2_X1 _09076_ ( .A1(\myclint.mtime [34] ), .A2(\myclint.mtime [35] ), .ZN(_01558_ ) );
INV_X1 _09077_ ( .A(\myclint.mtime [33] ), .ZN(_01559_ ) );
INV_X1 _09078_ ( .A(\myclint.mtime [32] ), .ZN(_01560_ ) );
NOR3_X1 _09079_ ( .A1(_01558_ ), .A2(_01559_ ), .A3(_01560_ ), .ZN(_01561_ ) );
AND4_X1 _09080_ ( .A1(_01554_ ), .A2(_01556_ ), .A3(_01557_ ), .A4(_01561_ ), .ZN(_01562_ ) );
INV_X1 _09081_ ( .A(_01562_ ), .ZN(_01563_ ) );
NOR2_X1 _09082_ ( .A1(_01552_ ), .A2(_01563_ ), .ZN(_01564_ ) );
AND2_X1 _09083_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01565_ ) );
AND2_X1 _09084_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01566_ ) );
AND2_X1 _09085_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01567_ ) );
AND2_X1 _09086_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01568_ ) );
AND4_X1 _09087_ ( .A1(_01565_ ), .A2(_01566_ ), .A3(_01567_ ), .A4(_01568_ ), .ZN(_01569_ ) );
AND2_X1 _09088_ ( .A1(_01564_ ), .A2(_01569_ ), .ZN(_01570_ ) );
AND2_X1 _09089_ ( .A1(\myclint.mtime [60] ), .A2(\myclint.mtime [61] ), .ZN(_01571_ ) );
AND4_X1 _09090_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01572_ ) );
NAND3_X1 _09091_ ( .A1(_01570_ ), .A2(_01571_ ), .A3(_01572_ ), .ZN(_01573_ ) );
OR3_X1 _09092_ ( .A1(_01573_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [63] ), .ZN(_01574_ ) );
OAI21_X1 _09093_ ( .A(\myclint.mtime [63] ), .B1(_01573_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01575_ ) );
AOI21_X1 _09094_ ( .A(fanout_net_1 ), .B1(_01574_ ), .B2(_01575_ ), .ZN(_00000_ ) );
OR2_X1 _09095_ ( .A1(_01573_ ), .A2(\myclint.mtime [62] ), .ZN(_01576_ ) );
NAND2_X1 _09096_ ( .A1(_01573_ ), .A2(\myclint.mtime [62] ), .ZN(_01577_ ) );
AOI21_X1 _09097_ ( .A(fanout_net_1 ), .B1(_01576_ ), .B2(_01577_ ), .ZN(_00001_ ) );
AND2_X1 _09098_ ( .A1(_01567_ ), .A2(_01568_ ), .ZN(_01578_ ) );
NAND2_X1 _09099_ ( .A1(_01564_ ), .A2(_01578_ ), .ZN(_01579_ ) );
OR3_X1 _09100_ ( .A1(_01579_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [53] ), .ZN(_01580_ ) );
OAI21_X1 _09101_ ( .A(\myclint.mtime [53] ), .B1(_01579_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01581_ ) );
AOI21_X1 _09102_ ( .A(fanout_net_1 ), .B1(_01580_ ), .B2(_01581_ ), .ZN(_00002_ ) );
XNOR2_X1 _09103_ ( .A(_01579_ ), .B(\myclint.mtime [52] ), .ZN(_01582_ ) );
INV_X1 _09104_ ( .A(fanout_net_1 ), .ZN(_01583_ ) );
BUF_X4 _09105_ ( .A(_01583_ ), .Z(_01584_ ) );
BUF_X2 _09106_ ( .A(_01584_ ), .Z(_01585_ ) );
AND2_X1 _09107_ ( .A1(_01582_ ), .A2(_01585_ ), .ZN(_00003_ ) );
INV_X1 _09108_ ( .A(_01552_ ), .ZN(_01586_ ) );
NAND3_X1 _09109_ ( .A1(_01586_ ), .A2(_01568_ ), .A3(_01562_ ), .ZN(_01587_ ) );
OR3_X1 _09110_ ( .A1(_01587_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [51] ), .ZN(_01588_ ) );
OAI21_X1 _09111_ ( .A(\myclint.mtime [51] ), .B1(_01587_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01589_ ) );
AOI21_X1 _09112_ ( .A(fanout_net_1 ), .B1(_01588_ ), .B2(_01589_ ), .ZN(_00004_ ) );
OR2_X1 _09113_ ( .A1(_01587_ ), .A2(\myclint.mtime [50] ), .ZN(_01590_ ) );
NAND2_X1 _09114_ ( .A1(_01587_ ), .A2(\myclint.mtime [50] ), .ZN(_01591_ ) );
AOI21_X1 _09115_ ( .A(fanout_net_1 ), .B1(_01590_ ), .B2(_01591_ ), .ZN(_00005_ ) );
AND3_X4 _09116_ ( .A1(_01537_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01592_ ) );
AND3_X4 _09117_ ( .A1(_01592_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01593_ ) );
AND3_X1 _09118_ ( .A1(_01593_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01594_ ) );
AND3_X2 _09119_ ( .A1(_01594_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01595_ ) );
AND3_X4 _09120_ ( .A1(_01595_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01596_ ) );
AND3_X1 _09121_ ( .A1(_01596_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01597_ ) );
AND3_X4 _09122_ ( .A1(_01597_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01598_ ) );
AND3_X4 _09123_ ( .A1(_01598_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01599_ ) );
AND3_X4 _09124_ ( .A1(_01599_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01600_ ) );
AND3_X2 _09125_ ( .A1(_01600_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01601_ ) );
AND2_X4 _09126_ ( .A1(_01601_ ), .A2(\myclint.mtime [27] ), .ZN(_01602_ ) );
AND4_X1 _09127_ ( .A1(\myclint.mtime [33] ), .A2(_01602_ ), .A3(_01543_ ), .A4(_01548_ ), .ZN(_01603_ ) );
AND3_X2 _09128_ ( .A1(_01603_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01604_ ) );
AND2_X1 _09129_ ( .A1(_01604_ ), .A2(\myclint.mtime [35] ), .ZN(_01605_ ) );
AND2_X1 _09130_ ( .A1(\myclint.mtime [36] ), .A2(\myclint.mtime [37] ), .ZN(_01606_ ) );
AND2_X1 _09131_ ( .A1(_01605_ ), .A2(_01606_ ), .ZN(_01607_ ) );
AND3_X1 _09132_ ( .A1(_01607_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [39] ), .ZN(_01608_ ) );
AND3_X4 _09133_ ( .A1(_01608_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01609_ ) );
AND2_X4 _09134_ ( .A1(_01609_ ), .A2(\myclint.mtime [42] ), .ZN(_01610_ ) );
AND2_X4 _09135_ ( .A1(_01610_ ), .A2(\myclint.mtime [43] ), .ZN(_01611_ ) );
INV_X1 _09136_ ( .A(_01611_ ), .ZN(_01612_ ) );
INV_X1 _09137_ ( .A(_01554_ ), .ZN(_01613_ ) );
NOR3_X4 _09138_ ( .A1(_01612_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01613_ ), .ZN(_01614_ ) );
AND2_X1 _09139_ ( .A1(_01614_ ), .A2(\myclint.mtime [49] ), .ZN(_01615_ ) );
BUF_X4 _09140_ ( .A(_01584_ ), .Z(_01616_ ) );
OAI21_X1 _09141_ ( .A(_01616_ ), .B1(_01614_ ), .B2(\myclint.mtime [49] ), .ZN(_01617_ ) );
NOR2_X1 _09142_ ( .A1(_01615_ ), .A2(_01617_ ), .ZN(_00006_ ) );
NAND2_X1 _09143_ ( .A1(_01538_ ), .A2(_01541_ ), .ZN(_01618_ ) );
NAND4_X1 _09144_ ( .A1(_01547_ ), .A2(_01543_ ), .A3(_01548_ ), .A4(_01550_ ), .ZN(_01619_ ) );
OR4_X1 _09145_ ( .A1(\myclint.mtime [48] ), .A2(_01618_ ), .A3(_01619_ ), .A4(_01563_ ), .ZN(_01620_ ) );
OAI21_X1 _09146_ ( .A(\myclint.mtime [48] ), .B1(_01552_ ), .B2(_01563_ ), .ZN(_01621_ ) );
AOI21_X1 _09147_ ( .A(fanout_net_1 ), .B1(_01620_ ), .B2(_01621_ ), .ZN(_00007_ ) );
NAND3_X1 _09148_ ( .A1(_01610_ ), .A2(\myclint.mtime [43] ), .A3(_01553_ ), .ZN(_01622_ ) );
NOR2_X1 _09149_ ( .A1(_01622_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01623_ ) );
OAI21_X1 _09150_ ( .A(_01584_ ), .B1(_01623_ ), .B2(\myclint.mtime [47] ), .ZN(_01624_ ) );
NAND3_X1 _09151_ ( .A1(_01610_ ), .A2(\myclint.mtime [44] ), .A3(\myclint.mtime [43] ), .ZN(_01625_ ) );
INV_X1 _09152_ ( .A(\myclint.mtime [45] ), .ZN(_01626_ ) );
NOR3_X1 _09153_ ( .A1(_01625_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01626_ ), .ZN(_01627_ ) );
AOI21_X1 _09154_ ( .A(_01624_ ), .B1(\myclint.mtime [47] ), .B2(_01627_ ), .ZN(_00008_ ) );
AND2_X1 _09155_ ( .A1(_01561_ ), .A2(_01557_ ), .ZN(_01628_ ) );
AND2_X1 _09156_ ( .A1(_01586_ ), .A2(_01628_ ), .ZN(_01629_ ) );
AND3_X1 _09157_ ( .A1(_01629_ ), .A2(_01553_ ), .A3(_01556_ ), .ZN(_01630_ ) );
XNOR2_X1 _09158_ ( .A(_01630_ ), .B(\myclint.mtime [46] ), .ZN(_01631_ ) );
NOR2_X1 _09159_ ( .A1(_01631_ ), .A2(fanout_net_1 ), .ZN(_00009_ ) );
INV_X1 _09160_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01632_ ) );
AND3_X1 _09161_ ( .A1(_01610_ ), .A2(_01632_ ), .A3(\myclint.mtime [43] ), .ZN(_01633_ ) );
AND2_X1 _09162_ ( .A1(_01633_ ), .A2(\myclint.mtime [45] ), .ZN(_01634_ ) );
OAI21_X1 _09163_ ( .A(_01616_ ), .B1(_01633_ ), .B2(\myclint.mtime [45] ), .ZN(_01635_ ) );
NOR2_X1 _09164_ ( .A1(_01634_ ), .A2(_01635_ ), .ZN(_00010_ ) );
AND2_X1 _09165_ ( .A1(_01629_ ), .A2(_01556_ ), .ZN(_01636_ ) );
XNOR2_X1 _09166_ ( .A(_01636_ ), .B(\myclint.mtime [44] ), .ZN(_01637_ ) );
NOR2_X1 _09167_ ( .A1(_01637_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
INV_X1 _09168_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01638_ ) );
NAND3_X1 _09169_ ( .A1(_01570_ ), .A2(_01638_ ), .A3(_01572_ ), .ZN(_01639_ ) );
OR2_X1 _09170_ ( .A1(_01639_ ), .A2(\myclint.mtime [61] ), .ZN(_01640_ ) );
NAND2_X1 _09171_ ( .A1(_01639_ ), .A2(\myclint.mtime [61] ), .ZN(_01641_ ) );
AOI21_X1 _09172_ ( .A(fanout_net_1 ), .B1(_01640_ ), .B2(_01641_ ), .ZN(_00012_ ) );
INV_X1 _09173_ ( .A(_01609_ ), .ZN(_01642_ ) );
NOR2_X1 _09174_ ( .A1(_01642_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01643_ ) );
AND2_X1 _09175_ ( .A1(_01643_ ), .A2(\myclint.mtime [43] ), .ZN(_01644_ ) );
OAI21_X1 _09176_ ( .A(_01616_ ), .B1(_01643_ ), .B2(\myclint.mtime [43] ), .ZN(_01645_ ) );
NOR2_X1 _09177_ ( .A1(_01644_ ), .A2(_01645_ ), .ZN(_00013_ ) );
OAI21_X1 _09178_ ( .A(_01616_ ), .B1(_01609_ ), .B2(\myclint.mtime [42] ), .ZN(_01646_ ) );
NOR2_X1 _09179_ ( .A1(_01610_ ), .A2(_01646_ ), .ZN(_00014_ ) );
INV_X1 _09180_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01647_ ) );
AND2_X1 _09181_ ( .A1(_01608_ ), .A2(_01647_ ), .ZN(_01648_ ) );
OAI21_X1 _09182_ ( .A(_01585_ ), .B1(_01648_ ), .B2(\myclint.mtime [41] ), .ZN(_01649_ ) );
AND3_X1 _09183_ ( .A1(_01608_ ), .A2(\myclint.mtime [41] ), .A3(_01647_ ), .ZN(_01650_ ) );
NOR2_X1 _09184_ ( .A1(_01649_ ), .A2(_01650_ ), .ZN(_00015_ ) );
XNOR2_X1 _09185_ ( .A(_01629_ ), .B(\myclint.mtime [40] ), .ZN(_01651_ ) );
NOR2_X1 _09186_ ( .A1(_01651_ ), .A2(fanout_net_1 ), .ZN(_00016_ ) );
NAND3_X1 _09187_ ( .A1(_01586_ ), .A2(_01606_ ), .A3(_01561_ ), .ZN(_01652_ ) );
OR3_X1 _09188_ ( .A1(_01652_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [39] ), .ZN(_01653_ ) );
OAI21_X1 _09189_ ( .A(\myclint.mtime [39] ), .B1(_01652_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01654_ ) );
AOI21_X1 _09190_ ( .A(fanout_net_1 ), .B1(_01653_ ), .B2(_01654_ ), .ZN(_00017_ ) );
OR2_X1 _09191_ ( .A1(_01652_ ), .A2(\myclint.mtime [38] ), .ZN(_01655_ ) );
NAND2_X1 _09192_ ( .A1(_01652_ ), .A2(\myclint.mtime [38] ), .ZN(_01656_ ) );
AOI21_X1 _09193_ ( .A(fanout_net_1 ), .B1(_01655_ ), .B2(_01656_ ), .ZN(_00018_ ) );
INV_X1 _09194_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01657_ ) );
AND3_X1 _09195_ ( .A1(_01604_ ), .A2(_01657_ ), .A3(\myclint.mtime [35] ), .ZN(_01658_ ) );
AND2_X1 _09196_ ( .A1(_01658_ ), .A2(\myclint.mtime [37] ), .ZN(_01659_ ) );
OAI21_X1 _09197_ ( .A(_01616_ ), .B1(_01658_ ), .B2(\myclint.mtime [37] ), .ZN(_01660_ ) );
NOR2_X1 _09198_ ( .A1(_01659_ ), .A2(_01660_ ), .ZN(_00019_ ) );
NAND2_X1 _09199_ ( .A1(_01586_ ), .A2(_01561_ ), .ZN(_01661_ ) );
OR2_X1 _09200_ ( .A1(_01661_ ), .A2(\myclint.mtime [36] ), .ZN(_01662_ ) );
NAND2_X1 _09201_ ( .A1(_01661_ ), .A2(\myclint.mtime [36] ), .ZN(_01663_ ) );
AOI21_X1 _09202_ ( .A(fanout_net_1 ), .B1(_01662_ ), .B2(_01663_ ), .ZN(_00020_ ) );
NAND4_X1 _09203_ ( .A1(_01602_ ), .A2(\myclint.mtime [33] ), .A3(_01543_ ), .A4(_01548_ ), .ZN(_01664_ ) );
NOR3_X1 _09204_ ( .A1(_01664_ ), .A2(_01560_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01665_ ) );
AND2_X1 _09205_ ( .A1(_01665_ ), .A2(\myclint.mtime [35] ), .ZN(_01666_ ) );
OAI21_X1 _09206_ ( .A(_01616_ ), .B1(_01665_ ), .B2(\myclint.mtime [35] ), .ZN(_01667_ ) );
NOR2_X1 _09207_ ( .A1(_01666_ ), .A2(_01667_ ), .ZN(_00021_ ) );
NOR2_X1 _09208_ ( .A1(_01664_ ), .A2(_01560_ ), .ZN(_01668_ ) );
OAI21_X1 _09209_ ( .A(_01585_ ), .B1(_01668_ ), .B2(\myclint.mtime [34] ), .ZN(_01669_ ) );
NOR2_X1 _09210_ ( .A1(_01669_ ), .A2(_01604_ ), .ZN(_00022_ ) );
AND2_X1 _09211_ ( .A1(_01570_ ), .A2(_01572_ ), .ZN(_01670_ ) );
XNOR2_X1 _09212_ ( .A(_01670_ ), .B(\myclint.mtime [60] ), .ZN(_01671_ ) );
NOR2_X1 _09213_ ( .A1(_01671_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
NOR3_X1 _09214_ ( .A1(_01618_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_01619_ ), .ZN(_01672_ ) );
XNOR2_X1 _09215_ ( .A(_01672_ ), .B(\myclint.mtime [33] ), .ZN(_01673_ ) );
NOR2_X1 _09216_ ( .A1(_01673_ ), .A2(fanout_net_1 ), .ZN(_00024_ ) );
OAI21_X1 _09217_ ( .A(\myclint.mtime [32] ), .B1(_01618_ ), .B2(_01619_ ), .ZN(_01674_ ) );
NAND4_X1 _09218_ ( .A1(_01538_ ), .A2(_01560_ ), .A3(_01541_ ), .A4(_01551_ ), .ZN(_01675_ ) );
AOI21_X1 _09219_ ( .A(fanout_net_1 ), .B1(_01674_ ), .B2(_01675_ ), .ZN(_00025_ ) );
AND2_X1 _09220_ ( .A1(_01542_ ), .A2(_01547_ ), .ZN(_01676_ ) );
NAND3_X1 _09221_ ( .A1(_01676_ ), .A2(_01548_ ), .A3(_01550_ ), .ZN(_01677_ ) );
OR3_X1 _09222_ ( .A1(_01677_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [31] ), .ZN(_01678_ ) );
OAI21_X1 _09223_ ( .A(\myclint.mtime [31] ), .B1(_01677_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01679_ ) );
AOI21_X1 _09224_ ( .A(fanout_net_1 ), .B1(_01678_ ), .B2(_01679_ ), .ZN(_00026_ ) );
OR2_X1 _09225_ ( .A1(_01677_ ), .A2(\myclint.mtime [30] ), .ZN(_01680_ ) );
NAND2_X1 _09226_ ( .A1(_01677_ ), .A2(\myclint.mtime [30] ), .ZN(_01681_ ) );
AOI21_X1 _09227_ ( .A(fanout_net_1 ), .B1(_01680_ ), .B2(_01681_ ), .ZN(_00027_ ) );
INV_X1 _09228_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01682_ ) );
AND3_X1 _09229_ ( .A1(_01601_ ), .A2(_01682_ ), .A3(\myclint.mtime [27] ), .ZN(_01683_ ) );
AND2_X1 _09230_ ( .A1(_01683_ ), .A2(\myclint.mtime [29] ), .ZN(_01684_ ) );
OAI21_X1 _09231_ ( .A(_01616_ ), .B1(_01683_ ), .B2(\myclint.mtime [29] ), .ZN(_01685_ ) );
NOR2_X1 _09232_ ( .A1(_01684_ ), .A2(_01685_ ), .ZN(_00028_ ) );
NAND2_X1 _09233_ ( .A1(_01676_ ), .A2(_01550_ ), .ZN(_01686_ ) );
OR2_X1 _09234_ ( .A1(_01686_ ), .A2(\myclint.mtime [28] ), .ZN(_01687_ ) );
NAND2_X1 _09235_ ( .A1(_01686_ ), .A2(\myclint.mtime [28] ), .ZN(_01688_ ) );
AOI21_X1 _09236_ ( .A(fanout_net_1 ), .B1(_01687_ ), .B2(_01688_ ), .ZN(_00029_ ) );
NAND3_X1 _09237_ ( .A1(_01542_ ), .A2(_01549_ ), .A3(_01547_ ), .ZN(_01689_ ) );
OR3_X1 _09238_ ( .A1(_01689_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01690_ ) );
OAI21_X1 _09239_ ( .A(\myclint.mtime [27] ), .B1(_01689_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01691_ ) );
AOI21_X1 _09240_ ( .A(fanout_net_1 ), .B1(_01690_ ), .B2(_01691_ ), .ZN(_00030_ ) );
AND2_X1 _09241_ ( .A1(_01600_ ), .A2(\myclint.mtime [25] ), .ZN(_01692_ ) );
OAI21_X1 _09242_ ( .A(_01585_ ), .B1(_01692_ ), .B2(\myclint.mtime [26] ), .ZN(_01693_ ) );
NOR2_X1 _09243_ ( .A1(_01693_ ), .A2(_01601_ ), .ZN(_00031_ ) );
INV_X1 _09244_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01694_ ) );
AND3_X1 _09245_ ( .A1(_01599_ ), .A2(_01694_ ), .A3(\myclint.mtime [23] ), .ZN(_01695_ ) );
AND2_X1 _09246_ ( .A1(_01695_ ), .A2(\myclint.mtime [25] ), .ZN(_01696_ ) );
OAI21_X1 _09247_ ( .A(_01616_ ), .B1(_01695_ ), .B2(\myclint.mtime [25] ), .ZN(_01697_ ) );
NOR2_X1 _09248_ ( .A1(_01696_ ), .A2(_01697_ ), .ZN(_00032_ ) );
BUF_X4 _09249_ ( .A(_01584_ ), .Z(_01698_ ) );
AND2_X1 _09250_ ( .A1(_01599_ ), .A2(\myclint.mtime [23] ), .ZN(_01699_ ) );
OAI21_X1 _09251_ ( .A(_01698_ ), .B1(_01699_ ), .B2(\myclint.mtime [24] ), .ZN(_01700_ ) );
NOR2_X1 _09252_ ( .A1(_01700_ ), .A2(_01600_ ), .ZN(_00033_ ) );
NAND3_X1 _09253_ ( .A1(_01570_ ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .ZN(_01701_ ) );
OR3_X1 _09254_ ( .A1(_01701_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [59] ), .ZN(_01702_ ) );
OAI21_X1 _09255_ ( .A(\myclint.mtime [59] ), .B1(_01701_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01703_ ) );
AOI21_X1 _09256_ ( .A(fanout_net_1 ), .B1(_01702_ ), .B2(_01703_ ), .ZN(_00034_ ) );
NOR2_X1 _09257_ ( .A1(_01618_ ), .A2(_01545_ ), .ZN(_01704_ ) );
NAND3_X1 _09258_ ( .A1(_01704_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01705_ ) );
OR3_X1 _09259_ ( .A1(_01705_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01706_ ) );
OAI21_X1 _09260_ ( .A(\myclint.mtime [23] ), .B1(_01705_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01707_ ) );
AOI21_X1 _09261_ ( .A(fanout_net_1 ), .B1(_01706_ ), .B2(_01707_ ), .ZN(_00035_ ) );
AND2_X1 _09262_ ( .A1(_01598_ ), .A2(\myclint.mtime [21] ), .ZN(_01708_ ) );
OAI21_X1 _09263_ ( .A(_01698_ ), .B1(_01708_ ), .B2(\myclint.mtime [22] ), .ZN(_01709_ ) );
NOR2_X1 _09264_ ( .A1(_01709_ ), .A2(_01599_ ), .ZN(_00036_ ) );
OR3_X1 _09265_ ( .A1(_01618_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01545_ ), .ZN(_01710_ ) );
NAND2_X1 _09266_ ( .A1(_01710_ ), .A2(\myclint.mtime [21] ), .ZN(_01711_ ) );
OR4_X1 _09267_ ( .A1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01618_ ), .A3(\myclint.mtime [21] ), .A4(_01545_ ), .ZN(_01712_ ) );
AOI21_X1 _09268_ ( .A(fanout_net_1 ), .B1(_01711_ ), .B2(_01712_ ), .ZN(_00037_ ) );
AND2_X1 _09269_ ( .A1(_01597_ ), .A2(\myclint.mtime [19] ), .ZN(_01713_ ) );
OAI21_X1 _09270_ ( .A(_01698_ ), .B1(_01713_ ), .B2(\myclint.mtime [20] ), .ZN(_01714_ ) );
NOR2_X1 _09271_ ( .A1(_01714_ ), .A2(_01598_ ), .ZN(_00038_ ) );
NAND3_X1 _09272_ ( .A1(_01542_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01715_ ) );
OR3_X1 _09273_ ( .A1(_01715_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01716_ ) );
OAI21_X1 _09274_ ( .A(\myclint.mtime [19] ), .B1(_01715_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01717_ ) );
AOI21_X1 _09275_ ( .A(fanout_net_1 ), .B1(_01716_ ), .B2(_01717_ ), .ZN(_00039_ ) );
AND2_X1 _09276_ ( .A1(_01596_ ), .A2(\myclint.mtime [17] ), .ZN(_01718_ ) );
OAI21_X1 _09277_ ( .A(_01698_ ), .B1(_01718_ ), .B2(\myclint.mtime [18] ), .ZN(_01719_ ) );
NOR2_X1 _09278_ ( .A1(_01719_ ), .A2(_01597_ ), .ZN(_00040_ ) );
INV_X1 _09279_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01720_ ) );
AND3_X1 _09280_ ( .A1(_01595_ ), .A2(_01720_ ), .A3(\myclint.mtime [15] ), .ZN(_01721_ ) );
AND2_X1 _09281_ ( .A1(_01721_ ), .A2(\myclint.mtime [17] ), .ZN(_01722_ ) );
OAI21_X1 _09282_ ( .A(_01616_ ), .B1(_01721_ ), .B2(\myclint.mtime [17] ), .ZN(_01723_ ) );
NOR2_X1 _09283_ ( .A1(_01722_ ), .A2(_01723_ ), .ZN(_00041_ ) );
AND2_X1 _09284_ ( .A1(_01595_ ), .A2(\myclint.mtime [15] ), .ZN(_01724_ ) );
OAI21_X1 _09285_ ( .A(_01698_ ), .B1(_01724_ ), .B2(\myclint.mtime [16] ), .ZN(_01725_ ) );
NOR2_X1 _09286_ ( .A1(_01725_ ), .A2(_01596_ ), .ZN(_00042_ ) );
AND3_X1 _09287_ ( .A1(_01540_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [11] ), .ZN(_01726_ ) );
AND2_X1 _09288_ ( .A1(_01538_ ), .A2(_01726_ ), .ZN(_01727_ ) );
NAND3_X1 _09289_ ( .A1(_01727_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01728_ ) );
OR3_X1 _09290_ ( .A1(_01728_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01729_ ) );
OAI21_X1 _09291_ ( .A(\myclint.mtime [15] ), .B1(_01728_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01730_ ) );
AOI21_X1 _09292_ ( .A(fanout_net_1 ), .B1(_01729_ ), .B2(_01730_ ), .ZN(_00043_ ) );
AND2_X1 _09293_ ( .A1(_01594_ ), .A2(\myclint.mtime [13] ), .ZN(_01731_ ) );
OAI21_X1 _09294_ ( .A(_01698_ ), .B1(_01731_ ), .B2(\myclint.mtime [14] ), .ZN(_01732_ ) );
NOR2_X1 _09295_ ( .A1(_01732_ ), .A2(_01595_ ), .ZN(_00044_ ) );
OR2_X1 _09296_ ( .A1(_01701_ ), .A2(\myclint.mtime [58] ), .ZN(_01733_ ) );
NAND2_X1 _09297_ ( .A1(_01701_ ), .A2(\myclint.mtime [58] ), .ZN(_01734_ ) );
AOI21_X1 _09298_ ( .A(fanout_net_1 ), .B1(_01733_ ), .B2(_01734_ ), .ZN(_00045_ ) );
INV_X1 _09299_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01735_ ) );
AND3_X1 _09300_ ( .A1(_01593_ ), .A2(_01735_ ), .A3(\myclint.mtime [11] ), .ZN(_01736_ ) );
AND2_X1 _09301_ ( .A1(_01736_ ), .A2(\myclint.mtime [13] ), .ZN(_01737_ ) );
OAI21_X1 _09302_ ( .A(_01616_ ), .B1(_01736_ ), .B2(\myclint.mtime [13] ), .ZN(_01738_ ) );
NOR2_X1 _09303_ ( .A1(_01737_ ), .A2(_01738_ ), .ZN(_00046_ ) );
XNOR2_X1 _09304_ ( .A(_01727_ ), .B(\myclint.mtime [12] ), .ZN(_01739_ ) );
NOR2_X1 _09305_ ( .A1(_01739_ ), .A2(fanout_net_1 ), .ZN(_00047_ ) );
INV_X1 _09306_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01740_ ) );
AND3_X1 _09307_ ( .A1(_01592_ ), .A2(_01740_ ), .A3(\myclint.mtime [9] ), .ZN(_01741_ ) );
OAI21_X1 _09308_ ( .A(_01584_ ), .B1(_01741_ ), .B2(\myclint.mtime [11] ), .ZN(_01742_ ) );
AOI21_X1 _09309_ ( .A(_01742_ ), .B1(\myclint.mtime [11] ), .B2(_01741_ ), .ZN(_00048_ ) );
AOI21_X1 _09310_ ( .A(\myclint.mtime [10] ), .B1(_01592_ ), .B2(\myclint.mtime [9] ), .ZN(_01743_ ) );
NOR3_X1 _09311_ ( .A1(_01593_ ), .A2(_01743_ ), .A3(fanout_net_1 ), .ZN(_00049_ ) );
INV_X1 _09312_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01744_ ) );
AND3_X1 _09313_ ( .A1(_01538_ ), .A2(\myclint.mtime [9] ), .A3(_01744_ ), .ZN(_01745_ ) );
AOI21_X1 _09314_ ( .A(\myclint.mtime [9] ), .B1(_01538_ ), .B2(_01744_ ), .ZN(_01746_ ) );
NOR3_X1 _09315_ ( .A1(_01745_ ), .A2(_01746_ ), .A3(fanout_net_1 ), .ZN(_00050_ ) );
OAI21_X1 _09316_ ( .A(_01698_ ), .B1(_01538_ ), .B2(\myclint.mtime [8] ), .ZN(_01747_ ) );
NOR2_X1 _09317_ ( .A1(_01747_ ), .A2(_01592_ ), .ZN(_00051_ ) );
AND2_X1 _09318_ ( .A1(_01536_ ), .A2(\myclint.mtime [5] ), .ZN(_01748_ ) );
INV_X1 _09319_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01749_ ) );
AND3_X1 _09320_ ( .A1(_01748_ ), .A2(_01749_ ), .A3(\myclint.mtime [7] ), .ZN(_01750_ ) );
AOI21_X1 _09321_ ( .A(\myclint.mtime [7] ), .B1(_01748_ ), .B2(_01749_ ), .ZN(_01751_ ) );
NOR3_X1 _09322_ ( .A1(_01750_ ), .A2(_01751_ ), .A3(fanout_net_2 ), .ZN(_00052_ ) );
OAI21_X1 _09323_ ( .A(_01698_ ), .B1(_01748_ ), .B2(\myclint.mtime [6] ), .ZN(_01752_ ) );
NOR2_X1 _09324_ ( .A1(_01752_ ), .A2(_01537_ ), .ZN(_00053_ ) );
AND2_X1 _09325_ ( .A1(_01535_ ), .A2(\myclint.mtime [3] ), .ZN(_01753_ ) );
INV_X1 _09326_ ( .A(_01753_ ), .ZN(_01754_ ) );
OR3_X1 _09327_ ( .A1(_01754_ ), .A2(\myclint.mtime [5] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01755_ ) );
OAI21_X1 _09328_ ( .A(\myclint.mtime [5] ), .B1(_01754_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01756_ ) );
AOI21_X1 _09329_ ( .A(fanout_net_2 ), .B1(_01755_ ), .B2(_01756_ ), .ZN(_00054_ ) );
OAI21_X1 _09330_ ( .A(_01698_ ), .B1(_01753_ ), .B2(\myclint.mtime [4] ), .ZN(_01757_ ) );
NOR2_X1 _09331_ ( .A1(_01757_ ), .A2(_01536_ ), .ZN(_00055_ ) );
INV_X1 _09332_ ( .A(_01570_ ), .ZN(_01758_ ) );
OR3_X1 _09333_ ( .A1(_01758_ ), .A2(\myclint.mtime [57] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01759_ ) );
OAI21_X1 _09334_ ( .A(\myclint.mtime [57] ), .B1(_01758_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01760_ ) );
AOI21_X1 _09335_ ( .A(fanout_net_2 ), .B1(_01759_ ), .B2(_01760_ ), .ZN(_00056_ ) );
AND2_X1 _09336_ ( .A1(\myclint.mtime [1] ), .A2(\myclint.mtime [0] ), .ZN(_01761_ ) );
INV_X1 _09337_ ( .A(_01761_ ), .ZN(_01762_ ) );
OR3_X1 _09338_ ( .A1(_01762_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01763_ ) );
OAI21_X1 _09339_ ( .A(\myclint.mtime [3] ), .B1(_01762_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01764_ ) );
AOI21_X1 _09340_ ( .A(fanout_net_2 ), .B1(_01763_ ), .B2(_01764_ ), .ZN(_00057_ ) );
AOI21_X1 _09341_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [1] ), .B2(\myclint.mtime [0] ), .ZN(_01765_ ) );
NOR3_X1 _09342_ ( .A1(_01535_ ), .A2(_01765_ ), .A3(fanout_net_2 ), .ZN(_00058_ ) );
NOR2_X1 _09343_ ( .A1(\myclint.mtime [1] ), .A2(\myclint.mtime [0] ), .ZN(_01766_ ) );
NOR3_X1 _09344_ ( .A1(_01761_ ), .A2(_01766_ ), .A3(fanout_net_2 ), .ZN(_00059_ ) );
AND2_X1 _09345_ ( .A1(_01585_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_00060_ ) );
OR2_X1 _09346_ ( .A1(_01758_ ), .A2(\myclint.mtime [56] ), .ZN(_01767_ ) );
NAND2_X1 _09347_ ( .A1(_01758_ ), .A2(\myclint.mtime [56] ), .ZN(_01768_ ) );
AOI21_X1 _09348_ ( .A(fanout_net_2 ), .B1(_01767_ ), .B2(_01768_ ), .ZN(_00061_ ) );
NAND3_X1 _09349_ ( .A1(_01564_ ), .A2(_01566_ ), .A3(_01578_ ), .ZN(_01769_ ) );
OR3_X1 _09350_ ( .A1(_01769_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01770_ ) );
OAI21_X1 _09351_ ( .A(\myclint.mtime [55] ), .B1(_01769_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01771_ ) );
AOI21_X1 _09352_ ( .A(fanout_net_2 ), .B1(_01770_ ), .B2(_01771_ ), .ZN(_00062_ ) );
OR2_X1 _09353_ ( .A1(_01769_ ), .A2(\myclint.mtime [54] ), .ZN(_01772_ ) );
NAND2_X1 _09354_ ( .A1(_01769_ ), .A2(\myclint.mtime [54] ), .ZN(_01773_ ) );
AOI21_X1 _09355_ ( .A(fanout_net_2 ), .B1(_01772_ ), .B2(_01773_ ), .ZN(_00063_ ) );
OR2_X1 _09356_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[0][26] ), .ZN(_01774_ ) );
INV_X8 _09357_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01775_ ) );
BUF_X4 _09358_ ( .A(_01775_ ), .Z(_01776_ ) );
INV_X32 _09359_ ( .A(fanout_net_43 ), .ZN(_01777_ ) );
BUF_X32 _09360_ ( .A(_01777_ ), .Z(_01778_ ) );
BUF_X16 _09361_ ( .A(_01778_ ), .Z(_01779_ ) );
OAI211_X1 _09362_ ( .A(_01774_ ), .B(_01776_ ), .C1(_01779_ ), .C2(\myifu.myicache.tag[1][26] ), .ZN(_01780_ ) );
OR2_X1 _09363_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[2][26] ), .ZN(_01781_ ) );
BUF_X16 _09364_ ( .A(_01777_ ), .Z(_01782_ ) );
OAI211_X1 _09365_ ( .A(_01781_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01782_ ), .C2(\myifu.myicache.tag[3][26] ), .ZN(_01783_ ) );
AND3_X1 _09366_ ( .A1(_01780_ ), .A2(_01783_ ), .A3(\IF_ID_pc [31] ), .ZN(_01784_ ) );
OR2_X4 _09367_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[3][0] ), .ZN(_01785_ ) );
OAI211_X2 _09368_ ( .A(_01785_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[2][0] ), .ZN(_01786_ ) );
OR2_X1 _09369_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[0][0] ), .ZN(_01787_ ) );
OAI211_X1 _09370_ ( .A(_01787_ ), .B(_01775_ ), .C1(_01782_ ), .C2(\myifu.myicache.tag[1][0] ), .ZN(_01788_ ) );
NAND2_X2 _09371_ ( .A1(_01786_ ), .A2(_01788_ ), .ZN(_01789_ ) );
XNOR2_X2 _09372_ ( .A(_01789_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01790_ ) );
OR2_X1 _09373_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.valid [2] ), .ZN(_01791_ ) );
BUF_X4 _09374_ ( .A(_01779_ ), .Z(_01792_ ) );
OAI211_X1 _09375_ ( .A(_01791_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01792_ ), .C2(\myifu.myicache.valid [3] ), .ZN(_01793_ ) );
OR2_X1 _09376_ ( .A1(\myifu.myicache.valid [0] ), .A2(fanout_net_43 ), .ZN(_01794_ ) );
BUF_X4 _09377_ ( .A(_01776_ ), .Z(_01795_ ) );
OAI211_X1 _09378_ ( .A(_01794_ ), .B(_01795_ ), .C1(\myifu.myicache.valid [1] ), .C2(_01792_ ), .ZN(_01796_ ) );
AOI211_X1 _09379_ ( .A(_01784_ ), .B(_01790_ ), .C1(_01793_ ), .C2(_01796_ ), .ZN(_01797_ ) );
AOI21_X1 _09380_ ( .A(\IF_ID_pc [31] ), .B1(_01780_ ), .B2(_01783_ ), .ZN(_01798_ ) );
OR2_X4 _09381_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[3][25] ), .ZN(_01799_ ) );
OAI211_X2 _09382_ ( .A(_01799_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[2][25] ), .ZN(_01800_ ) );
OR2_X1 _09383_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[0][25] ), .ZN(_01801_ ) );
OAI211_X1 _09384_ ( .A(_01801_ ), .B(_01775_ ), .C1(_01782_ ), .C2(\myifu.myicache.tag[1][25] ), .ZN(_01802_ ) );
NAND2_X2 _09385_ ( .A1(_01800_ ), .A2(_01802_ ), .ZN(_01803_ ) );
INV_X1 _09386_ ( .A(\IF_ID_pc [30] ), .ZN(_01804_ ) );
XNOR2_X1 _09387_ ( .A(_01803_ ), .B(_01804_ ), .ZN(_01805_ ) );
MUX2_X1 _09388_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(fanout_net_43 ), .Z(_01806_ ) );
OR2_X1 _09389_ ( .A1(_01806_ ), .A2(_01776_ ), .ZN(_01807_ ) );
MUX2_X1 _09390_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(fanout_net_43 ), .Z(_01808_ ) );
OAI21_X1 _09391_ ( .A(_01807_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01808_ ), .ZN(_01809_ ) );
AOI211_X1 _09392_ ( .A(_01798_ ), .B(_01805_ ), .C1(\IF_ID_pc [29] ), .C2(_01809_ ), .ZN(_01810_ ) );
AND2_X1 _09393_ ( .A1(_01797_ ), .A2(_01810_ ), .ZN(_01811_ ) );
OR2_X1 _09394_ ( .A1(_01779_ ), .A2(\myifu.myicache.tag[1][21] ), .ZN(_01812_ ) );
OAI211_X1 _09395_ ( .A(_01812_ ), .B(_01795_ ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[0][21] ), .ZN(_01813_ ) );
OR2_X1 _09396_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[2][21] ), .ZN(_01814_ ) );
OAI211_X1 _09397_ ( .A(_01814_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01792_ ), .C2(\myifu.myicache.tag[3][21] ), .ZN(_01815_ ) );
NAND2_X1 _09398_ ( .A1(_01813_ ), .A2(_01815_ ), .ZN(_01816_ ) );
XNOR2_X1 _09399_ ( .A(_01816_ ), .B(\IF_ID_pc [26] ), .ZN(_01817_ ) );
AND2_X1 _09400_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[3][23] ), .ZN(_01818_ ) );
AOI211_X1 _09401_ ( .A(_01795_ ), .B(_01818_ ), .C1(_01792_ ), .C2(\myifu.myicache.tag[2][23] ), .ZN(_01819_ ) );
AND2_X1 _09402_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[1][23] ), .ZN(_01820_ ) );
AOI211_X1 _09403_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B(_01820_ ), .C1(_01792_ ), .C2(\myifu.myicache.tag[0][23] ), .ZN(_01821_ ) );
NOR2_X1 _09404_ ( .A1(_01819_ ), .A2(_01821_ ), .ZN(_01822_ ) );
XNOR2_X1 _09405_ ( .A(_01822_ ), .B(\IF_ID_pc [28] ), .ZN(_01823_ ) );
OR2_X2 _09406_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[1][20] ), .ZN(_01824_ ) );
OAI211_X2 _09407_ ( .A(_01824_ ), .B(_01775_ ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[0][20] ), .ZN(_01825_ ) );
OR2_X4 _09408_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[3][20] ), .ZN(_01826_ ) );
OAI211_X2 _09409_ ( .A(_01826_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[2][20] ), .ZN(_01827_ ) );
NAND2_X1 _09410_ ( .A1(_01825_ ), .A2(_01827_ ), .ZN(_01828_ ) );
INV_X1 _09411_ ( .A(\IF_ID_pc [25] ), .ZN(_01829_ ) );
NAND2_X1 _09412_ ( .A1(_01828_ ), .A2(_01829_ ), .ZN(_01830_ ) );
INV_X1 _09413_ ( .A(\IF_ID_pc [23] ), .ZN(_01831_ ) );
MUX2_X1 _09414_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(fanout_net_43 ), .Z(_01832_ ) );
MUX2_X1 _09415_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(fanout_net_43 ), .Z(_01833_ ) );
MUX2_X1 _09416_ ( .A(_01832_ ), .B(_01833_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01834_ ) );
OAI21_X2 _09417_ ( .A(_01830_ ), .B1(_01831_ ), .B2(_01834_ ), .ZN(_01835_ ) );
MUX2_X1 _09418_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(fanout_net_43 ), .Z(_01836_ ) );
AND2_X2 _09419_ ( .A1(_01836_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01837_ ) );
MUX2_X1 _09420_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(fanout_net_43 ), .Z(_01838_ ) );
AOI21_X4 _09421_ ( .A(_01837_ ), .B1(_01795_ ), .B2(_01838_ ), .ZN(_01839_ ) );
AOI221_X1 _09422_ ( .A(_01835_ ), .B1(_01831_ ), .B2(_01834_ ), .C1(\IF_ID_pc [21] ), .C2(_01839_ ), .ZN(_01840_ ) );
NAND4_X1 _09423_ ( .A1(_01811_ ), .A2(_01817_ ), .A3(_01823_ ), .A4(_01840_ ), .ZN(_01841_ ) );
MUX2_X1 _09424_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_43 ), .Z(_01842_ ) );
AND2_X2 _09425_ ( .A1(_01842_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01843_ ) );
MUX2_X1 _09426_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_43 ), .Z(_01844_ ) );
AOI21_X2 _09427_ ( .A(_01843_ ), .B1(_01795_ ), .B2(_01844_ ), .ZN(_01845_ ) );
NOR2_X1 _09428_ ( .A1(_01845_ ), .A2(\IF_ID_pc [16] ), .ZN(_01846_ ) );
OR2_X4 _09429_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[1][8] ), .ZN(_01847_ ) );
OAI211_X1 _09430_ ( .A(_01847_ ), .B(_01776_ ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[0][8] ), .ZN(_01848_ ) );
OR2_X1 _09431_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[2][8] ), .ZN(_01849_ ) );
OAI211_X1 _09432_ ( .A(_01849_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01782_ ), .C2(\myifu.myicache.tag[3][8] ), .ZN(_01850_ ) );
AND3_X1 _09433_ ( .A1(_01848_ ), .A2(_01850_ ), .A3(\IF_ID_pc [13] ), .ZN(_01851_ ) );
AOI21_X1 _09434_ ( .A(\IF_ID_pc [13] ), .B1(_01848_ ), .B2(_01850_ ), .ZN(_01852_ ) );
OR2_X4 _09435_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[3][9] ), .ZN(_01853_ ) );
OAI211_X2 _09436_ ( .A(_01853_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[2][9] ), .ZN(_01854_ ) );
OR2_X1 _09437_ ( .A1(fanout_net_43 ), .A2(\myifu.myicache.tag[0][9] ), .ZN(_01855_ ) );
OAI211_X1 _09438_ ( .A(_01855_ ), .B(_01775_ ), .C1(_01782_ ), .C2(\myifu.myicache.tag[1][9] ), .ZN(_01856_ ) );
AND3_X1 _09439_ ( .A1(_01854_ ), .A2(\IF_ID_pc [14] ), .A3(_01856_ ), .ZN(_01857_ ) );
NOR4_X1 _09440_ ( .A1(_01846_ ), .A2(_01851_ ), .A3(_01852_ ), .A4(_01857_ ), .ZN(_01858_ ) );
OR2_X4 _09441_ ( .A1(_01782_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01859_ ) );
OAI211_X1 _09442_ ( .A(_01859_ ), .B(_01776_ ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01860_ ) );
OR2_X4 _09443_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[3][12] ), .ZN(_01861_ ) );
OAI211_X1 _09444_ ( .A(_01861_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[2][12] ), .ZN(_01862_ ) );
AND3_X1 _09445_ ( .A1(_01860_ ), .A2(_01862_ ), .A3(\IF_ID_pc [17] ), .ZN(_01863_ ) );
OR2_X4 _09446_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[1][14] ), .ZN(_01864_ ) );
OAI211_X1 _09447_ ( .A(_01864_ ), .B(_01776_ ), .C1(fanout_net_43 ), .C2(\myifu.myicache.tag[0][14] ), .ZN(_01865_ ) );
OR2_X4 _09448_ ( .A1(_01778_ ), .A2(\myifu.myicache.tag[3][14] ), .ZN(_01866_ ) );
OAI211_X2 _09449_ ( .A(_01866_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][14] ), .ZN(_01867_ ) );
AND3_X1 _09450_ ( .A1(_01865_ ), .A2(_01867_ ), .A3(\IF_ID_pc [19] ), .ZN(_01868_ ) );
AOI21_X1 _09451_ ( .A(\IF_ID_pc [17] ), .B1(_01860_ ), .B2(_01862_ ), .ZN(_01869_ ) );
AOI21_X1 _09452_ ( .A(\IF_ID_pc [19] ), .B1(_01865_ ), .B2(_01867_ ), .ZN(_01870_ ) );
NOR4_X1 _09453_ ( .A1(_01863_ ), .A2(_01868_ ), .A3(_01869_ ), .A4(_01870_ ), .ZN(_01871_ ) );
AND2_X1 _09454_ ( .A1(_01858_ ), .A2(_01871_ ), .ZN(_01872_ ) );
OR2_X1 _09455_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][4] ), .ZN(_01873_ ) );
OAI211_X1 _09456_ ( .A(_01873_ ), .B(_01795_ ), .C1(_01792_ ), .C2(\myifu.myicache.tag[1][4] ), .ZN(_01874_ ) );
OR2_X1 _09457_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][4] ), .ZN(_01875_ ) );
OAI211_X1 _09458_ ( .A(_01875_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01792_ ), .C2(\myifu.myicache.tag[3][4] ), .ZN(_01876_ ) );
NAND2_X1 _09459_ ( .A1(_01874_ ), .A2(_01876_ ), .ZN(_01877_ ) );
XNOR2_X1 _09460_ ( .A(_01877_ ), .B(\IF_ID_pc [9] ), .ZN(_01878_ ) );
OR2_X1 _09461_ ( .A1(_01782_ ), .A2(\myifu.myicache.tag[3][3] ), .ZN(_01879_ ) );
OAI211_X1 _09462_ ( .A(_01879_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][3] ), .ZN(_01880_ ) );
OR2_X1 _09463_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][3] ), .ZN(_01881_ ) );
OAI211_X1 _09464_ ( .A(_01881_ ), .B(_01776_ ), .C1(_01779_ ), .C2(\myifu.myicache.tag[1][3] ), .ZN(_01882_ ) );
AOI21_X1 _09465_ ( .A(\IF_ID_pc [8] ), .B1(_01880_ ), .B2(_01882_ ), .ZN(_01883_ ) );
NAND3_X1 _09466_ ( .A1(_01880_ ), .A2(\IF_ID_pc [8] ), .A3(_01882_ ), .ZN(_01884_ ) );
OAI21_X1 _09467_ ( .A(_01884_ ), .B1(_01839_ ), .B2(\IF_ID_pc [21] ), .ZN(_01885_ ) );
MUX2_X1 _09468_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01886_ ) );
OR2_X2 _09469_ ( .A1(_01886_ ), .A2(_01775_ ), .ZN(_01887_ ) );
MUX2_X1 _09470_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01888_ ) );
OAI21_X1 _09471_ ( .A(_01887_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01888_ ), .ZN(_01889_ ) );
AOI211_X1 _09472_ ( .A(_01883_ ), .B(_01885_ ), .C1(\IF_ID_pc [12] ), .C2(_01889_ ), .ZN(_01890_ ) );
AND2_X1 _09473_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[3][6] ), .ZN(_01891_ ) );
AOI211_X1 _09474_ ( .A(_01795_ ), .B(_01891_ ), .C1(_01792_ ), .C2(\myifu.myicache.tag[2][6] ), .ZN(_01892_ ) );
AND2_X1 _09475_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_01893_ ) );
AOI211_X1 _09476_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B(_01893_ ), .C1(_01792_ ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_01894_ ) );
NOR2_X2 _09477_ ( .A1(_01892_ ), .A2(_01894_ ), .ZN(_01895_ ) );
XNOR2_X1 _09478_ ( .A(_01895_ ), .B(\IF_ID_pc [11] ), .ZN(_01896_ ) );
NAND4_X1 _09479_ ( .A1(_01872_ ), .A2(_01878_ ), .A3(_01890_ ), .A4(_01896_ ), .ZN(_01897_ ) );
NOR2_X2 _09480_ ( .A1(_01841_ ), .A2(_01897_ ), .ZN(_01898_ ) );
AND3_X1 _09481_ ( .A1(_01825_ ), .A2(_01827_ ), .A3(\IF_ID_pc [25] ), .ZN(_01899_ ) );
INV_X1 _09482_ ( .A(\IF_ID_pc [27] ), .ZN(_01900_ ) );
MUX2_X1 _09483_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01901_ ) );
MUX2_X1 _09484_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01902_ ) );
MUX2_X1 _09485_ ( .A(_01901_ ), .B(_01902_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01903_ ) );
AOI21_X1 _09486_ ( .A(_01899_ ), .B1(_01900_ ), .B2(_01903_ ), .ZN(_01904_ ) );
OAI221_X1 _09487_ ( .A(_01904_ ), .B1(\IF_ID_pc [29] ), .B2(_01809_ ), .C1(_01900_ ), .C2(_01903_ ), .ZN(_01905_ ) );
OR2_X1 _09488_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][17] ), .ZN(_01906_ ) );
OAI211_X1 _09489_ ( .A(_01906_ ), .B(_01776_ ), .C1(_01779_ ), .C2(\myifu.myicache.tag[1][17] ), .ZN(_01907_ ) );
OR2_X1 _09490_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][17] ), .ZN(_01908_ ) );
OAI211_X1 _09491_ ( .A(_01908_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01779_ ), .C2(\myifu.myicache.tag[3][17] ), .ZN(_01909_ ) );
NAND2_X1 _09492_ ( .A1(_01907_ ), .A2(_01909_ ), .ZN(_01910_ ) );
INV_X1 _09493_ ( .A(\IF_ID_pc [22] ), .ZN(_01911_ ) );
XNOR2_X1 _09494_ ( .A(_01910_ ), .B(_01911_ ), .ZN(_01912_ ) );
OR2_X1 _09495_ ( .A1(_01782_ ), .A2(\myifu.myicache.tag[3][19] ), .ZN(_01913_ ) );
OAI211_X1 _09496_ ( .A(_01913_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][19] ), .ZN(_01914_ ) );
OR2_X1 _09497_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][19] ), .ZN(_01915_ ) );
OAI211_X1 _09498_ ( .A(_01915_ ), .B(_01795_ ), .C1(_01792_ ), .C2(\myifu.myicache.tag[1][19] ), .ZN(_01916_ ) );
AND3_X1 _09499_ ( .A1(_01914_ ), .A2(\IF_ID_pc [24] ), .A3(_01916_ ), .ZN(_01917_ ) );
AOI21_X1 _09500_ ( .A(\IF_ID_pc [24] ), .B1(_01914_ ), .B2(_01916_ ), .ZN(_01918_ ) );
NOR4_X1 _09501_ ( .A1(_01905_ ), .A2(_01912_ ), .A3(_01917_ ), .A4(_01918_ ), .ZN(_01919_ ) );
MUX2_X1 _09502_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01920_ ) );
OR2_X2 _09503_ ( .A1(_01920_ ), .A2(_01776_ ), .ZN(_01921_ ) );
MUX2_X1 _09504_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01922_ ) );
OAI21_X1 _09505_ ( .A(_01921_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01922_ ), .ZN(_01923_ ) );
OR2_X2 _09506_ ( .A1(_01923_ ), .A2(\IF_ID_pc [20] ), .ZN(_01924_ ) );
MUX2_X1 _09507_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01925_ ) );
OR2_X2 _09508_ ( .A1(_01925_ ), .A2(_01775_ ), .ZN(_01926_ ) );
MUX2_X1 _09509_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01927_ ) );
OAI21_X1 _09510_ ( .A(_01926_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01927_ ), .ZN(_01928_ ) );
OR2_X1 _09511_ ( .A1(_01928_ ), .A2(\IF_ID_pc [18] ), .ZN(_01929_ ) );
NAND2_X1 _09512_ ( .A1(_01928_ ), .A2(\IF_ID_pc [18] ), .ZN(_01930_ ) );
NAND2_X1 _09513_ ( .A1(_01845_ ), .A2(\IF_ID_pc [16] ), .ZN(_01931_ ) );
NAND4_X1 _09514_ ( .A1(_01924_ ), .A2(_01929_ ), .A3(_01930_ ), .A4(_01931_ ), .ZN(_01932_ ) );
OR2_X4 _09515_ ( .A1(_01779_ ), .A2(\myifu.myicache.tag[1][10] ), .ZN(_01933_ ) );
OAI211_X1 _09516_ ( .A(_01933_ ), .B(_01795_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][10] ), .ZN(_01934_ ) );
OR2_X1 _09517_ ( .A1(_01782_ ), .A2(\myifu.myicache.tag[3][10] ), .ZN(_01935_ ) );
OAI211_X1 _09518_ ( .A(_01935_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][10] ), .ZN(_01936_ ) );
AND3_X1 _09519_ ( .A1(_01934_ ), .A2(_01936_ ), .A3(\IF_ID_pc [15] ), .ZN(_01937_ ) );
AOI21_X1 _09520_ ( .A(\IF_ID_pc [15] ), .B1(_01934_ ), .B2(_01936_ ), .ZN(_01938_ ) );
AOI21_X1 _09521_ ( .A(\IF_ID_pc [14] ), .B1(_01854_ ), .B2(_01856_ ), .ZN(_01939_ ) );
NOR4_X1 _09522_ ( .A1(_01932_ ), .A2(_01937_ ), .A3(_01938_ ), .A4(_01939_ ), .ZN(_01940_ ) );
MUX2_X1 _09523_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01941_ ) );
OR2_X2 _09524_ ( .A1(_01941_ ), .A2(_01775_ ), .ZN(_01942_ ) );
MUX2_X1 _09525_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01943_ ) );
OAI21_X1 _09526_ ( .A(_01942_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01943_ ), .ZN(_01944_ ) );
OR2_X1 _09527_ ( .A1(_01944_ ), .A2(\IF_ID_pc [10] ), .ZN(_01945_ ) );
OR2_X1 _09528_ ( .A1(_01889_ ), .A2(\IF_ID_pc [12] ), .ZN(_01946_ ) );
NAND2_X1 _09529_ ( .A1(_01923_ ), .A2(\IF_ID_pc [20] ), .ZN(_01947_ ) );
NAND2_X1 _09530_ ( .A1(_01944_ ), .A2(\IF_ID_pc [10] ), .ZN(_01948_ ) );
NAND4_X1 _09531_ ( .A1(_01945_ ), .A2(_01946_ ), .A3(_01947_ ), .A4(_01948_ ), .ZN(_01949_ ) );
OR2_X1 _09532_ ( .A1(_01782_ ), .A2(\myifu.myicache.tag[3][1] ), .ZN(_01950_ ) );
OAI211_X1 _09533_ ( .A(_01950_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][1] ), .ZN(_01951_ ) );
OR2_X1 _09534_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_01952_ ) );
OAI211_X1 _09535_ ( .A(_01952_ ), .B(_01776_ ), .C1(_01779_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_01953_ ) );
NAND2_X1 _09536_ ( .A1(_01951_ ), .A2(_01953_ ), .ZN(_01954_ ) );
INV_X1 _09537_ ( .A(\IF_ID_pc [6] ), .ZN(_01955_ ) );
XNOR2_X1 _09538_ ( .A(_01954_ ), .B(_01955_ ), .ZN(_01956_ ) );
OR2_X1 _09539_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][2] ), .ZN(_01957_ ) );
OAI211_X1 _09540_ ( .A(_01957_ ), .B(_01795_ ), .C1(_01779_ ), .C2(\myifu.myicache.tag[1][2] ), .ZN(_01958_ ) );
OR2_X1 _09541_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][2] ), .ZN(_01959_ ) );
OAI211_X1 _09542_ ( .A(_01959_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01779_ ), .C2(\myifu.myicache.tag[3][2] ), .ZN(_01960_ ) );
AOI21_X1 _09543_ ( .A(\IF_ID_pc [7] ), .B1(_01958_ ), .B2(_01960_ ), .ZN(_01961_ ) );
AND3_X1 _09544_ ( .A1(_01958_ ), .A2(_01960_ ), .A3(\IF_ID_pc [7] ), .ZN(_01962_ ) );
NOR4_X1 _09545_ ( .A1(_01949_ ), .A2(_01956_ ), .A3(_01961_ ), .A4(_01962_ ), .ZN(_01963_ ) );
AND3_X2 _09546_ ( .A1(_01919_ ), .A2(_01940_ ), .A3(_01963_ ), .ZN(_01964_ ) );
AND2_X4 _09547_ ( .A1(_01898_ ), .A2(_01964_ ), .ZN(_01965_ ) );
INV_X1 _09548_ ( .A(\myifu.state [0] ), .ZN(_01966_ ) );
NOR2_X4 _09549_ ( .A1(_01965_ ), .A2(_01966_ ), .ZN(_01967_ ) );
INV_X1 _09550_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01968_ ) );
NOR2_X4 _09551_ ( .A1(_01967_ ), .A2(_01968_ ), .ZN(_01969_ ) );
NOR2_X1 _09552_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01970_ ) );
NOR2_X4 _09553_ ( .A1(_01969_ ), .A2(_01970_ ), .ZN(_01971_ ) );
INV_X32 _09554_ ( .A(\EX_LS_flag [2] ), .ZN(_01972_ ) );
NAND4_X1 _09555_ ( .A1(_01972_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(\mylsu.state [0] ), .ZN(_01973_ ) );
INV_X1 _09556_ ( .A(EXU_valid_LSU ), .ZN(_01974_ ) );
NOR2_X1 _09557_ ( .A1(_01973_ ), .A2(_01974_ ), .ZN(_01975_ ) );
INV_X1 _09558_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01976_ ) );
NOR2_X1 _09559_ ( .A1(_01975_ ), .A2(_01976_ ), .ZN(_01977_ ) );
NOR2_X4 _09560_ ( .A1(_01971_ ), .A2(_01977_ ), .ZN(_01978_ ) );
BUF_X8 _09561_ ( .A(_01978_ ), .Z(_01979_ ) );
CLKBUF_X2 _09562_ ( .A(_01974_ ), .Z(_01980_ ) );
OR3_X1 _09563_ ( .A1(_01973_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(_01980_ ), .ZN(_01981_ ) );
BUF_X4 _09564_ ( .A(_01975_ ), .Z(_01982_ ) );
OAI211_X1 _09565_ ( .A(_01979_ ), .B(_01981_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01982_ ), .ZN(_01983_ ) );
INV_X4 _09566_ ( .A(_01971_ ), .ZN(_01984_ ) );
OAI21_X1 _09567_ ( .A(_01983_ ), .B1(_01804_ ), .B2(_01984_ ), .ZN(\io_master_araddr [30] ) );
CLKBUF_X2 _09568_ ( .A(_01973_ ), .Z(_01985_ ) );
OR3_X1 _09569_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(_01980_ ), .ZN(_01986_ ) );
OAI211_X1 _09570_ ( .A(_01979_ ), .B(_01986_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01982_ ), .ZN(_01987_ ) );
BUF_X4 _09571_ ( .A(_01967_ ), .Z(_01988_ ) );
OAI221_X1 _09572_ ( .A(\IF_ID_pc [27] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01988_ ), .C2(_01968_ ), .ZN(_01989_ ) );
AND2_X1 _09573_ ( .A1(_01987_ ), .A2(_01989_ ), .ZN(_01990_ ) );
INV_X1 _09574_ ( .A(_01990_ ), .ZN(\io_master_araddr [27] ) );
OR3_X1 _09575_ ( .A1(_01973_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(_01974_ ), .ZN(_01991_ ) );
OAI211_X1 _09576_ ( .A(_01978_ ), .B(_01991_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01982_ ), .ZN(_01992_ ) );
INV_X1 _09577_ ( .A(\IF_ID_pc [28] ), .ZN(_01993_ ) );
OAI21_X1 _09578_ ( .A(_01992_ ), .B1(_01993_ ), .B2(_01984_ ), .ZN(\io_master_araddr [28] ) );
OR3_X1 _09579_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(_01980_ ), .ZN(_01994_ ) );
BUF_X4 _09580_ ( .A(_01982_ ), .Z(_01995_ ) );
OAI211_X1 _09581_ ( .A(_01979_ ), .B(_01994_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01995_ ), .ZN(_01996_ ) );
INV_X1 _09582_ ( .A(\IF_ID_pc [24] ), .ZN(_01997_ ) );
BUF_X4 _09583_ ( .A(_01984_ ), .Z(_01998_ ) );
OAI21_X1 _09584_ ( .A(_01996_ ), .B1(_01997_ ), .B2(_01998_ ), .ZN(\io_master_araddr [24] ) );
OR4_X1 _09585_ ( .A1(\io_master_araddr [30] ), .A2(\io_master_araddr [27] ), .A3(\io_master_araddr [28] ), .A4(\io_master_araddr [24] ), .ZN(_01999_ ) );
BUF_X8 _09586_ ( .A(_01979_ ), .Z(_02000_ ) );
OR3_X1 _09587_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(_01980_ ), .ZN(_02001_ ) );
OAI211_X1 _09588_ ( .A(_02000_ ), .B(_02001_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01995_ ), .ZN(_02002_ ) );
OAI221_X1 _09589_ ( .A(\IF_ID_pc [26] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01988_ ), .C2(_01968_ ), .ZN(_02003_ ) );
AND2_X1 _09590_ ( .A1(_02002_ ), .A2(_02003_ ), .ZN(_02004_ ) );
CLKBUF_X2 _09591_ ( .A(_01974_ ), .Z(_02005_ ) );
OR3_X1 _09592_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [25] ), .A3(_02005_ ), .ZN(_02006_ ) );
OAI211_X4 _09593_ ( .A(_02000_ ), .B(_02006_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_01995_ ), .ZN(_02007_ ) );
OAI21_X1 _09594_ ( .A(_02007_ ), .B1(_01829_ ), .B2(_01998_ ), .ZN(\io_master_araddr [25] ) );
NAND2_X1 _09595_ ( .A1(_02004_ ), .A2(\io_master_araddr [25] ), .ZN(_02008_ ) );
OR3_X1 _09596_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(_02005_ ), .ZN(_02009_ ) );
OAI211_X1 _09597_ ( .A(_02000_ ), .B(_02009_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01995_ ), .ZN(_02010_ ) );
INV_X1 _09598_ ( .A(\IF_ID_pc [17] ), .ZN(_02011_ ) );
OAI21_X1 _09599_ ( .A(_02010_ ), .B1(_02011_ ), .B2(_01998_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09600_ ( .A1(_01973_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(_01974_ ), .ZN(_02012_ ) );
OAI211_X1 _09601_ ( .A(_01978_ ), .B(_02012_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01982_ ), .ZN(_02013_ ) );
OAI21_X2 _09602_ ( .A(_02013_ ), .B1(_01911_ ), .B2(_01984_ ), .ZN(\io_master_araddr [22] ) );
NOR4_X4 _09603_ ( .A1(_01999_ ), .A2(_02008_ ), .A3(\io_master_araddr [17] ), .A4(\io_master_araddr [22] ), .ZN(_02014_ ) );
INV_X1 _09604_ ( .A(_01995_ ), .ZN(_02015_ ) );
OR2_X1 _09605_ ( .A1(\EX_LS_dest_csreg_mem [27] ), .A2(\EX_LS_dest_csreg_mem [26] ), .ZN(_02016_ ) );
OR3_X1 _09606_ ( .A1(_02016_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(\EX_LS_dest_csreg_mem [25] ), .ZN(_02017_ ) );
OR4_X1 _09607_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(_02017_ ), .A3(\EX_LS_dest_csreg_mem [30] ), .A4(\EX_LS_dest_csreg_mem [29] ), .ZN(_02018_ ) );
NOR2_X1 _09608_ ( .A1(_02018_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .ZN(_02019_ ) );
AND2_X4 _09609_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02020_ ) );
AND2_X4 _09610_ ( .A1(_02020_ ), .A2(_01972_ ), .ZN(_02021_ ) );
AND2_X1 _09611_ ( .A1(_02019_ ), .A2(_02021_ ), .ZN(_02022_ ) );
INV_X1 _09612_ ( .A(_02022_ ), .ZN(_02023_ ) );
NOR2_X1 _09613_ ( .A1(fanout_net_5 ), .A2(fanout_net_6 ), .ZN(_02024_ ) );
INV_X1 _09614_ ( .A(_02024_ ), .ZN(_02025_ ) );
INV_X1 _09615_ ( .A(\EX_LS_typ [3] ), .ZN(_02026_ ) );
NOR2_X1 _09616_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [0] ), .ZN(_02027_ ) );
NAND4_X1 _09617_ ( .A1(_02025_ ), .A2(_02026_ ), .A3(\EX_LS_typ [2] ), .A4(_02027_ ), .ZN(_02028_ ) );
NOR2_X1 _09618_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02029_ ) );
INV_X1 _09619_ ( .A(_02029_ ), .ZN(_02030_ ) );
AND2_X1 _09620_ ( .A1(fanout_net_5 ), .A2(\EX_LS_typ [1] ), .ZN(_02031_ ) );
INV_X1 _09621_ ( .A(_02031_ ), .ZN(_02032_ ) );
OAI21_X1 _09622_ ( .A(_02028_ ), .B1(_02030_ ), .B2(_02032_ ), .ZN(_02033_ ) );
INV_X1 _09623_ ( .A(\EX_LS_typ [4] ), .ZN(_02034_ ) );
AND2_X1 _09624_ ( .A1(_02021_ ), .A2(_02034_ ), .ZN(_02035_ ) );
NAND2_X1 _09625_ ( .A1(_02033_ ), .A2(_02035_ ), .ZN(_02036_ ) );
AND2_X2 _09626_ ( .A1(_02023_ ), .A2(_02036_ ), .ZN(_02037_ ) );
INV_X32 _09627_ ( .A(\EX_LS_flag [1] ), .ZN(_02038_ ) );
NOR2_X4 _09628_ ( .A1(_02038_ ), .A2(\EX_LS_flag [0] ), .ZN(_02039_ ) );
AND2_X2 _09629_ ( .A1(_02039_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02040_ ) );
AND2_X1 _09630_ ( .A1(_02019_ ), .A2(_02040_ ), .ZN(_02041_ ) );
NAND3_X1 _09631_ ( .A1(_01972_ ), .A2(_02034_ ), .A3(\EX_LS_typ [0] ), .ZN(_02042_ ) );
NOR3_X1 _09632_ ( .A1(_02042_ ), .A2(_02038_ ), .A3(\EX_LS_flag [0] ), .ZN(_02043_ ) );
INV_X1 _09633_ ( .A(_02043_ ), .ZN(_02044_ ) );
AND3_X1 _09634_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02045_ ) );
AOI22_X1 _09635_ ( .A1(_02025_ ), .A2(_02045_ ), .B1(_02031_ ), .B2(_02029_ ), .ZN(_02046_ ) );
NOR2_X1 _09636_ ( .A1(_02044_ ), .A2(_02046_ ), .ZN(_02047_ ) );
NOR2_X1 _09637_ ( .A1(_02041_ ), .A2(_02047_ ), .ZN(_02048_ ) );
AND2_X1 _09638_ ( .A1(_02037_ ), .A2(_02048_ ), .ZN(_02049_ ) );
INV_X1 _09639_ ( .A(_02049_ ), .ZN(_02050_ ) );
OAI21_X1 _09640_ ( .A(_01998_ ), .B1(_02015_ ), .B2(_02050_ ), .ZN(_02051_ ) );
CLKBUF_X2 _09641_ ( .A(_01971_ ), .Z(_02052_ ) );
CLKBUF_X2 _09642_ ( .A(_02052_ ), .Z(_02053_ ) );
CLKBUF_X2 _09643_ ( .A(_02053_ ), .Z(_02054_ ) );
CLKBUF_X2 _09644_ ( .A(_02054_ ), .Z(_02055_ ) );
NOR2_X1 _09645_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02056_ ) );
INV_X2 _09646_ ( .A(_02056_ ), .ZN(_02057_ ) );
OAI21_X1 _09647_ ( .A(_02055_ ), .B1(_01966_ ), .B2(_02057_ ), .ZN(_02058_ ) );
OR3_X1 _09648_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(_01980_ ), .ZN(_02059_ ) );
OAI211_X1 _09649_ ( .A(_01979_ ), .B(_02059_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01995_ ), .ZN(_02060_ ) );
INV_X1 _09650_ ( .A(\IF_ID_pc [19] ), .ZN(_02061_ ) );
OAI21_X1 _09651_ ( .A(_02060_ ), .B1(_02061_ ), .B2(_01998_ ), .ZN(\io_master_araddr [19] ) );
OR3_X1 _09652_ ( .A1(_01973_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(_01980_ ), .ZN(_02062_ ) );
OAI211_X1 _09653_ ( .A(_01979_ ), .B(_02062_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01982_ ), .ZN(_02063_ ) );
INV_X1 _09654_ ( .A(\IF_ID_pc [20] ), .ZN(_02064_ ) );
OAI21_X1 _09655_ ( .A(_02063_ ), .B1(_02064_ ), .B2(_01984_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09656_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(_01980_ ), .ZN(_02065_ ) );
OAI211_X1 _09657_ ( .A(_01979_ ), .B(_02065_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01982_ ), .ZN(_02066_ ) );
INV_X1 _09658_ ( .A(\IF_ID_pc [18] ), .ZN(_02067_ ) );
OAI21_X1 _09659_ ( .A(_02066_ ), .B1(_02067_ ), .B2(_01984_ ), .ZN(\io_master_araddr [18] ) );
OR3_X1 _09660_ ( .A1(_01973_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(_01974_ ), .ZN(_02068_ ) );
OAI211_X1 _09661_ ( .A(_01978_ ), .B(_02068_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01982_ ), .ZN(_02069_ ) );
INV_X1 _09662_ ( .A(\IF_ID_pc [21] ), .ZN(_02070_ ) );
OAI21_X1 _09663_ ( .A(_02069_ ), .B1(_02070_ ), .B2(_01984_ ), .ZN(\io_master_araddr [21] ) );
NOR4_X1 _09664_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [18] ), .A4(\io_master_araddr [21] ), .ZN(_02071_ ) );
OR3_X1 _09665_ ( .A1(_01973_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(_01980_ ), .ZN(_02072_ ) );
OAI211_X1 _09666_ ( .A(_01979_ ), .B(_02072_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01982_ ), .ZN(_02073_ ) );
INV_X1 _09667_ ( .A(\IF_ID_pc [29] ), .ZN(_02074_ ) );
OAI21_X1 _09668_ ( .A(_02073_ ), .B1(_02074_ ), .B2(_01984_ ), .ZN(\io_master_araddr [29] ) );
OR3_X1 _09669_ ( .A1(_01973_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(_01980_ ), .ZN(_02075_ ) );
OAI211_X1 _09670_ ( .A(_01979_ ), .B(_02075_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01982_ ), .ZN(_02076_ ) );
OAI21_X1 _09671_ ( .A(_02076_ ), .B1(_01831_ ), .B2(_01984_ ), .ZN(\io_master_araddr [23] ) );
OR3_X1 _09672_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(_01980_ ), .ZN(_02077_ ) );
OAI211_X1 _09673_ ( .A(_01979_ ), .B(_02077_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01995_ ), .ZN(_02078_ ) );
OAI221_X1 _09674_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01988_ ), .C2(_01968_ ), .ZN(_02079_ ) );
NAND2_X1 _09675_ ( .A1(_02078_ ), .A2(_02079_ ), .ZN(\io_master_araddr [31] ) );
OR3_X1 _09676_ ( .A1(_01985_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(_02005_ ), .ZN(_02080_ ) );
OAI211_X1 _09677_ ( .A(_02000_ ), .B(_02080_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01995_ ), .ZN(_02081_ ) );
OAI221_X1 _09678_ ( .A(\IF_ID_pc [16] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01988_ ), .C2(_01968_ ), .ZN(_02082_ ) );
NAND2_X1 _09679_ ( .A1(_02081_ ), .A2(_02082_ ), .ZN(\io_master_araddr [16] ) );
NOR4_X1 _09680_ ( .A1(\io_master_araddr [29] ), .A2(\io_master_araddr [23] ), .A3(\io_master_araddr [31] ), .A4(\io_master_araddr [16] ), .ZN(_02083_ ) );
AND2_X1 _09681_ ( .A1(_02071_ ), .A2(_02083_ ), .ZN(_02084_ ) );
NAND4_X1 _09682_ ( .A1(_02014_ ), .A2(_02051_ ), .A3(_02058_ ), .A4(_02084_ ), .ZN(_02085_ ) );
INV_X1 _09683_ ( .A(\myclint.rvalid ), .ZN(_02086_ ) );
AOI211_X1 _09684_ ( .A(_01968_ ), .B(_01998_ ), .C1(_01988_ ), .C2(_02056_ ), .ZN(_02087_ ) );
BUF_X4 _09685_ ( .A(_01995_ ), .Z(_02088_ ) );
AOI211_X1 _09686_ ( .A(_01976_ ), .B(_02055_ ), .C1(_02088_ ), .C2(_02049_ ), .ZN(_02089_ ) );
NOR2_X1 _09687_ ( .A1(_02087_ ), .A2(_02089_ ), .ZN(_02090_ ) );
AND3_X1 _09688_ ( .A1(_02014_ ), .A2(\myclint.rvalid ), .A3(_02084_ ), .ZN(_02091_ ) );
AOI221_X4 _09689_ ( .A(fanout_net_2 ), .B1(_02085_ ), .B2(_02086_ ), .C1(_02090_ ), .C2(_02091_ ), .ZN(_00064_ ) );
INV_X1 _09690_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02092_ ) );
CLKBUF_X2 _09691_ ( .A(_02092_ ), .Z(_02093_ ) );
AND2_X1 _09692_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00065_ ) );
AND2_X1 _09693_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [4] ), .ZN(_00066_ ) );
INV_X1 _09694_ ( .A(\LS_WB_wdata_csreg [23] ), .ZN(_02094_ ) );
NOR2_X1 _09695_ ( .A1(_02094_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00067_ ) );
AND2_X1 _09696_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00068_ ) );
AND2_X1 _09697_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00069_ ) );
AND2_X1 _09698_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [20] ), .ZN(_00070_ ) );
INV_X1 _09699_ ( .A(\LS_WB_wdata_csreg [19] ), .ZN(_02095_ ) );
NOR2_X1 _09700_ ( .A1(_02095_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00071_ ) );
INV_X1 _09701_ ( .A(\LS_WB_wdata_csreg [18] ), .ZN(_02096_ ) );
NOR2_X1 _09702_ ( .A1(_02096_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00072_ ) );
INV_X1 _09703_ ( .A(\LS_WB_wdata_csreg [17] ), .ZN(_02097_ ) );
NOR2_X1 _09704_ ( .A1(_02097_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00073_ ) );
AND2_X1 _09705_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00074_ ) );
AND2_X1 _09706_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00075_ ) );
AND2_X1 _09707_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00076_ ) );
AND2_X1 _09708_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00077_ ) );
AND2_X1 _09709_ ( .A1(_02093_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00078_ ) );
INV_X1 _09710_ ( .A(\LS_WB_wdata_csreg [12] ), .ZN(_02098_ ) );
NOR2_X1 _09711_ ( .A1(_02098_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00079_ ) );
CLKBUF_X2 _09712_ ( .A(_02092_ ), .Z(_02099_ ) );
AND2_X1 _09713_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00080_ ) );
AND2_X1 _09714_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00081_ ) );
AND2_X1 _09715_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00082_ ) );
INV_X1 _09716_ ( .A(\LS_WB_wdata_csreg [8] ), .ZN(_02100_ ) );
NOR2_X1 _09717_ ( .A1(_02100_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00083_ ) );
INV_X1 _09718_ ( .A(\LS_WB_wdata_csreg [7] ), .ZN(_02101_ ) );
NOR2_X1 _09719_ ( .A1(_02101_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00084_ ) );
INV_X1 _09720_ ( .A(\LS_WB_wdata_csreg [6] ), .ZN(_02102_ ) );
NOR2_X1 _09721_ ( .A1(_02102_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00085_ ) );
AND2_X1 _09722_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00086_ ) );
AND2_X1 _09723_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00087_ ) );
AND2_X1 _09724_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00088_ ) );
AND2_X1 _09725_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00089_ ) );
AND2_X1 _09726_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00090_ ) );
AND2_X1 _09727_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00091_ ) );
AND2_X1 _09728_ ( .A1(_02099_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00092_ ) );
INV_X1 _09729_ ( .A(_02037_ ), .ZN(_02103_ ) );
INV_X1 _09730_ ( .A(_02048_ ), .ZN(_02104_ ) );
BUF_X2 _09731_ ( .A(_02104_ ), .Z(_02105_ ) );
NOR2_X1 _09732_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02106_ ) );
NAND2_X1 _09733_ ( .A1(_02106_ ), .A2(_01584_ ), .ZN(_02107_ ) );
OR2_X1 _09734_ ( .A1(\myexu.pc_jump [27] ), .A2(\myexu.pc_jump [26] ), .ZN(_02108_ ) );
OR3_X1 _09735_ ( .A1(_02108_ ), .A2(\myexu.pc_jump [25] ), .A3(\myexu.pc_jump [24] ), .ZN(_02109_ ) );
OR4_X1 _09736_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02110_ ) );
NOR2_X1 _09737_ ( .A1(_02109_ ), .A2(_02110_ ), .ZN(_02111_ ) );
NOR2_X1 _09738_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02112_ ) );
INV_X1 _09739_ ( .A(_02112_ ), .ZN(_02113_ ) );
NOR3_X1 _09740_ ( .A1(_02111_ ), .A2(exception_quest_IDU ), .A3(_02113_ ), .ZN(_02114_ ) );
NOR4_X1 _09741_ ( .A1(_02103_ ), .A2(_02105_ ), .A3(_02107_ ), .A4(_02114_ ), .ZN(_00094_ ) );
AOI21_X1 _09742_ ( .A(_02107_ ), .B1(_02049_ ), .B2(exception_quest_IDU ), .ZN(_00095_ ) );
NOR2_X1 _09743_ ( .A1(fanout_net_2 ), .A2(fanout_net_17 ), .ZN(_02115_ ) );
INV_X1 _09744_ ( .A(IDU_valid_EXU ), .ZN(_02116_ ) );
NOR2_X1 _09745_ ( .A1(_02116_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _09746_ ( .A(check_quest ), .ZN(_02117_ ) );
NOR2_X1 _09747_ ( .A1(_02117_ ), .A2(check_assert ), .ZN(_02118_ ) );
OAI21_X1 _09748_ ( .A(_02115_ ), .B1(\myexu.state_$_ANDNOT__B_Y ), .B2(_02118_ ), .ZN(_02119_ ) );
INV_X1 _09749_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_02120_ ) );
INV_X1 _09750_ ( .A(\ID_EX_typ [6] ), .ZN(_02121_ ) );
NAND2_X1 _09751_ ( .A1(_02121_ ), .A2(\ID_EX_typ [7] ), .ZN(_02122_ ) );
INV_X1 _09752_ ( .A(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_02123_ ) );
NOR3_X1 _09753_ ( .A1(_02122_ ), .A2(\ID_EX_typ [5] ), .A3(_02123_ ), .ZN(_02124_ ) );
AOI211_X1 _09754_ ( .A(_02120_ ), .B(_02124_ ), .C1(_02118_ ), .C2(_02122_ ), .ZN(_02125_ ) );
INV_X1 _09755_ ( .A(\ID_EX_typ [5] ), .ZN(_02126_ ) );
NOR2_X1 _09756_ ( .A1(_02122_ ), .A2(_02126_ ), .ZN(_02127_ ) );
AND2_X2 _09757_ ( .A1(_02127_ ), .A2(fanout_net_7 ), .ZN(_02128_ ) );
INV_X1 _09758_ ( .A(_02128_ ), .ZN(_02129_ ) );
BUF_X4 _09759_ ( .A(_02129_ ), .Z(_02130_ ) );
AOI21_X1 _09760_ ( .A(_02119_ ), .B1(_02125_ ), .B2(_02130_ ), .ZN(_00096_ ) );
INV_X1 _09761_ ( .A(fanout_net_18 ), .ZN(_02131_ ) );
CLKBUF_X2 _09762_ ( .A(_02131_ ), .Z(_02132_ ) );
CLKBUF_X2 _09763_ ( .A(_02132_ ), .Z(_02133_ ) );
CLKBUF_X2 _09764_ ( .A(_02133_ ), .Z(_02134_ ) );
CLKBUF_X2 _09765_ ( .A(_02134_ ), .Z(_02135_ ) );
BUF_X2 _09766_ ( .A(_02135_ ), .Z(_02136_ ) );
NOR2_X1 _09767_ ( .A1(_02136_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02137_ ) );
OAI21_X1 _09768_ ( .A(fanout_net_26 ), .B1(fanout_net_18 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02138_ ) );
NOR2_X1 _09769_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02139_ ) );
INV_X2 _09770_ ( .A(fanout_net_26 ), .ZN(_02140_ ) );
BUF_X4 _09771_ ( .A(_02140_ ), .Z(_02141_ ) );
BUF_X4 _09772_ ( .A(_02141_ ), .Z(_02142_ ) );
BUF_X4 _09773_ ( .A(_02142_ ), .Z(_02143_ ) );
BUF_X4 _09774_ ( .A(_02143_ ), .Z(_02144_ ) );
BUF_X4 _09775_ ( .A(_02144_ ), .Z(_02145_ ) );
OAI21_X1 _09776_ ( .A(_02145_ ), .B1(_02136_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02146_ ) );
OAI221_X1 _09777_ ( .A(fanout_net_29 ), .B1(_02137_ ), .B2(_02138_ ), .C1(_02139_ ), .C2(_02146_ ), .ZN(_02147_ ) );
MUX2_X1 _09778_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02148_ ) );
MUX2_X1 _09779_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02149_ ) );
MUX2_X1 _09780_ ( .A(_02148_ ), .B(_02149_ ), .S(_02145_ ), .Z(_02150_ ) );
OAI211_X1 _09781_ ( .A(fanout_net_30 ), .B(_02147_ ), .C1(_02150_ ), .C2(fanout_net_29 ), .ZN(_02151_ ) );
MUX2_X1 _09782_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02152_ ) );
AND2_X1 _09783_ ( .A1(_02152_ ), .A2(fanout_net_26 ), .ZN(_02153_ ) );
MUX2_X1 _09784_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02154_ ) );
AOI211_X1 _09785_ ( .A(fanout_net_29 ), .B(_02153_ ), .C1(_02145_ ), .C2(_02154_ ), .ZN(_02155_ ) );
INV_X1 _09786_ ( .A(fanout_net_30 ), .ZN(_02156_ ) );
BUF_X4 _09787_ ( .A(_02156_ ), .Z(_02157_ ) );
BUF_X4 _09788_ ( .A(_02157_ ), .Z(_02158_ ) );
BUF_X4 _09789_ ( .A(_02158_ ), .Z(_02159_ ) );
MUX2_X1 _09790_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02160_ ) );
MUX2_X1 _09791_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02161_ ) );
MUX2_X1 _09792_ ( .A(_02160_ ), .B(_02161_ ), .S(fanout_net_26 ), .Z(_02162_ ) );
INV_X2 _09793_ ( .A(fanout_net_29 ), .ZN(_02163_ ) );
BUF_X4 _09794_ ( .A(_02163_ ), .Z(_02164_ ) );
BUF_X4 _09795_ ( .A(_02164_ ), .Z(_02165_ ) );
BUF_X4 _09796_ ( .A(_02165_ ), .Z(_02166_ ) );
BUF_X4 _09797_ ( .A(_02166_ ), .Z(_02167_ ) );
OAI21_X1 _09798_ ( .A(_02159_ ), .B1(_02162_ ), .B2(_02167_ ), .ZN(_02168_ ) );
INV_X1 _09799_ ( .A(\EX_LS_flag [0] ), .ZN(_02169_ ) );
NOR2_X2 _09800_ ( .A1(_02169_ ), .A2(\EX_LS_flag [1] ), .ZN(_02170_ ) );
AND2_X2 _09801_ ( .A1(_02170_ ), .A2(\EX_LS_flag [2] ), .ZN(_02171_ ) );
AOI211_X1 _09802_ ( .A(_02021_ ), .B(_02171_ ), .C1(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .C2(_02170_ ), .ZN(_02172_ ) );
AND2_X4 _09803_ ( .A1(_02039_ ), .A2(\EX_LS_flag [2] ), .ZN(_02173_ ) );
INV_X4 _09804_ ( .A(_02173_ ), .ZN(_02174_ ) );
NAND2_X2 _09805_ ( .A1(_02172_ ), .A2(_02174_ ), .ZN(_02175_ ) );
XNOR2_X1 _09806_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02176_ ) );
OR4_X1 _09807_ ( .A1(\EX_LS_dest_reg [3] ), .A2(\EX_LS_dest_reg [2] ), .A3(\EX_LS_dest_reg [1] ), .A4(\EX_LS_dest_reg [0] ), .ZN(_02177_ ) );
OR2_X4 _09808_ ( .A1(_02177_ ), .A2(\EX_LS_dest_reg [4] ), .ZN(_02178_ ) );
INV_X1 _09809_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02179_ ) );
NAND2_X1 _09810_ ( .A1(_02179_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02180_ ) );
NAND4_X4 _09811_ ( .A1(_02175_ ), .A2(_02176_ ), .A3(_02178_ ), .A4(_02180_ ), .ZN(_02181_ ) );
BUF_X16 _09812_ ( .A(_02181_ ), .Z(_02182_ ) );
BUF_X16 _09813_ ( .A(_02182_ ), .Z(_02183_ ) );
BUF_X2 _09814_ ( .A(_02183_ ), .Z(_02184_ ) );
BUF_X2 _09815_ ( .A(_02184_ ), .Z(_02185_ ) );
XNOR2_X1 _09816_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .ZN(_02186_ ) );
INV_X1 _09817_ ( .A(\ID_EX_rs1 [3] ), .ZN(_02187_ ) );
NAND2_X1 _09818_ ( .A1(_02187_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02188_ ) );
NAND3_X1 _09819_ ( .A1(_02186_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y ), .A3(_02188_ ), .ZN(_02189_ ) );
XOR2_X1 _09820_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .Z(_02190_ ) );
OAI22_X1 _09821_ ( .A1(_02187_ ), .A2(\EX_LS_dest_reg [3] ), .B1(_02179_ ), .B2(\ID_EX_rs1 [1] ), .ZN(_02191_ ) );
OR3_X2 _09822_ ( .A1(_02189_ ), .A2(_02190_ ), .A3(_02191_ ), .ZN(_02192_ ) );
BUF_X2 _09823_ ( .A(_02192_ ), .Z(_02193_ ) );
BUF_X2 _09824_ ( .A(_02193_ ), .Z(_02194_ ) );
BUF_X2 _09825_ ( .A(_02194_ ), .Z(_02195_ ) );
BUF_X2 _09826_ ( .A(_02195_ ), .Z(_02196_ ) );
OAI221_X1 _09827_ ( .A(_02151_ ), .B1(_02155_ ), .B2(_02168_ ), .C1(_02185_ ), .C2(_02196_ ), .ZN(_02197_ ) );
OR3_X1 _09828_ ( .A1(_02185_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02196_ ), .ZN(_02198_ ) );
AND2_X2 _09829_ ( .A1(_02197_ ), .A2(_02198_ ), .ZN(_02199_ ) );
XNOR2_X1 _09830_ ( .A(_02199_ ), .B(\ID_EX_imm [30] ), .ZN(_02200_ ) );
OR3_X1 _09831_ ( .A1(_02185_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02196_ ), .ZN(_02201_ ) );
OR2_X1 _09832_ ( .A1(_02136_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02202_ ) );
OAI211_X1 _09833_ ( .A(_02202_ ), .B(_02145_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02203_ ) );
INV_X1 _09834_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02204_ ) );
NAND2_X1 _09835_ ( .A1(_02204_ ), .A2(fanout_net_18 ), .ZN(_02205_ ) );
OAI211_X1 _09836_ ( .A(_02205_ ), .B(fanout_net_26 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02206_ ) );
NAND3_X1 _09837_ ( .A1(_02203_ ), .A2(_02206_ ), .A3(_02167_ ), .ZN(_02207_ ) );
MUX2_X1 _09838_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02208_ ) );
MUX2_X1 _09839_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02209_ ) );
BUF_X4 _09840_ ( .A(_02144_ ), .Z(_02210_ ) );
MUX2_X1 _09841_ ( .A(_02208_ ), .B(_02209_ ), .S(_02210_ ), .Z(_02211_ ) );
OAI211_X1 _09842_ ( .A(_02159_ ), .B(_02207_ ), .C1(_02211_ ), .C2(_02167_ ), .ZN(_02212_ ) );
CLKBUF_X2 _09843_ ( .A(_02135_ ), .Z(_02213_ ) );
OR2_X1 _09844_ ( .A1(_02213_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02214_ ) );
OAI211_X1 _09845_ ( .A(_02214_ ), .B(fanout_net_26 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02215_ ) );
OR2_X1 _09846_ ( .A1(_02213_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02216_ ) );
OAI211_X1 _09847_ ( .A(_02216_ ), .B(_02145_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02217_ ) );
NAND3_X1 _09848_ ( .A1(_02215_ ), .A2(_02217_ ), .A3(fanout_net_29 ), .ZN(_02218_ ) );
MUX2_X1 _09849_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02219_ ) );
MUX2_X1 _09850_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02220_ ) );
MUX2_X1 _09851_ ( .A(_02219_ ), .B(_02220_ ), .S(fanout_net_26 ), .Z(_02221_ ) );
OAI211_X1 _09852_ ( .A(fanout_net_30 ), .B(_02218_ ), .C1(_02221_ ), .C2(fanout_net_29 ), .ZN(_02222_ ) );
OAI211_X1 _09853_ ( .A(_02212_ ), .B(_02222_ ), .C1(_02185_ ), .C2(_02196_ ), .ZN(_02223_ ) );
NAND2_X1 _09854_ ( .A1(_02201_ ), .A2(_02223_ ), .ZN(_02224_ ) );
XNOR2_X1 _09855_ ( .A(_02224_ ), .B(\ID_EX_imm [28] ), .ZN(_02225_ ) );
OR3_X1 _09856_ ( .A1(_02185_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02195_ ), .ZN(_02226_ ) );
INV_X1 _09857_ ( .A(\ID_EX_imm [27] ), .ZN(_02227_ ) );
OR2_X1 _09858_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02228_ ) );
OAI211_X1 _09859_ ( .A(_02228_ ), .B(_02145_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02229_ ) );
OR2_X1 _09860_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02230_ ) );
OAI211_X1 _09861_ ( .A(_02230_ ), .B(fanout_net_26 ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02231_ ) );
NAND3_X1 _09862_ ( .A1(_02229_ ), .A2(_02231_ ), .A3(_02166_ ), .ZN(_02232_ ) );
MUX2_X1 _09863_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02233_ ) );
MUX2_X1 _09864_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02234_ ) );
MUX2_X1 _09865_ ( .A(_02233_ ), .B(_02234_ ), .S(_02210_ ), .Z(_02235_ ) );
OAI211_X1 _09866_ ( .A(_02159_ ), .B(_02232_ ), .C1(_02235_ ), .C2(_02167_ ), .ZN(_02236_ ) );
OR2_X1 _09867_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02237_ ) );
OAI211_X1 _09868_ ( .A(_02237_ ), .B(_02210_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02238_ ) );
NOR2_X1 _09869_ ( .A1(_02136_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02239_ ) );
OAI21_X1 _09870_ ( .A(fanout_net_26 ), .B1(fanout_net_18 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02240_ ) );
OAI211_X1 _09871_ ( .A(_02238_ ), .B(fanout_net_29 ), .C1(_02239_ ), .C2(_02240_ ), .ZN(_02241_ ) );
MUX2_X1 _09872_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02242_ ) );
MUX2_X1 _09873_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02243_ ) );
MUX2_X1 _09874_ ( .A(_02242_ ), .B(_02243_ ), .S(fanout_net_26 ), .Z(_02244_ ) );
OAI211_X1 _09875_ ( .A(_02241_ ), .B(fanout_net_30 ), .C1(_02244_ ), .C2(fanout_net_29 ), .ZN(_02245_ ) );
OAI211_X1 _09876_ ( .A(_02236_ ), .B(_02245_ ), .C1(_02185_ ), .C2(_02196_ ), .ZN(_02246_ ) );
AND3_X1 _09877_ ( .A1(_02226_ ), .A2(_02227_ ), .A3(_02246_ ), .ZN(_02247_ ) );
AOI21_X1 _09878_ ( .A(_02227_ ), .B1(_02226_ ), .B2(_02246_ ), .ZN(_02248_ ) );
NOR2_X1 _09879_ ( .A1(_02247_ ), .A2(_02248_ ), .ZN(_02249_ ) );
INV_X1 _09880_ ( .A(_02249_ ), .ZN(_02250_ ) );
OR3_X1 _09881_ ( .A1(_02184_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02195_ ), .ZN(_02251_ ) );
OR2_X1 _09882_ ( .A1(_02135_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02252_ ) );
OAI211_X1 _09883_ ( .A(_02252_ ), .B(_02210_ ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02253_ ) );
OR2_X1 _09884_ ( .A1(_02135_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02254_ ) );
OAI211_X1 _09885_ ( .A(_02254_ ), .B(fanout_net_26 ), .C1(fanout_net_18 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02255_ ) );
NAND3_X1 _09886_ ( .A1(_02253_ ), .A2(_02255_ ), .A3(_02166_ ), .ZN(_02256_ ) );
MUX2_X1 _09887_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02257_ ) );
MUX2_X1 _09888_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02258_ ) );
MUX2_X1 _09889_ ( .A(_02257_ ), .B(_02258_ ), .S(_02144_ ), .Z(_02259_ ) );
OAI211_X1 _09890_ ( .A(_02159_ ), .B(_02256_ ), .C1(_02259_ ), .C2(_02167_ ), .ZN(_02260_ ) );
OR2_X1 _09891_ ( .A1(_02135_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02261_ ) );
OAI211_X1 _09892_ ( .A(_02261_ ), .B(_02144_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02262_ ) );
NOR2_X1 _09893_ ( .A1(_02136_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02263_ ) );
OAI21_X1 _09894_ ( .A(fanout_net_26 ), .B1(fanout_net_19 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02264_ ) );
OAI211_X1 _09895_ ( .A(_02262_ ), .B(fanout_net_29 ), .C1(_02263_ ), .C2(_02264_ ), .ZN(_02265_ ) );
MUX2_X1 _09896_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02266_ ) );
MUX2_X1 _09897_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02267_ ) );
MUX2_X1 _09898_ ( .A(_02266_ ), .B(_02267_ ), .S(fanout_net_26 ), .Z(_02268_ ) );
OAI211_X1 _09899_ ( .A(_02265_ ), .B(fanout_net_30 ), .C1(_02268_ ), .C2(fanout_net_29 ), .ZN(_02269_ ) );
OAI211_X1 _09900_ ( .A(_02260_ ), .B(_02269_ ), .C1(_02184_ ), .C2(_02196_ ), .ZN(_02270_ ) );
NAND2_X2 _09901_ ( .A1(_02251_ ), .A2(_02270_ ), .ZN(_02271_ ) );
INV_X1 _09902_ ( .A(\ID_EX_imm [26] ), .ZN(_02272_ ) );
XNOR2_X1 _09903_ ( .A(_02271_ ), .B(_02272_ ), .ZN(_02273_ ) );
INV_X1 _09904_ ( .A(_02273_ ), .ZN(_02274_ ) );
OR3_X1 _09905_ ( .A1(_02184_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02195_ ), .ZN(_02275_ ) );
OR2_X1 _09906_ ( .A1(_02135_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02276_ ) );
OAI211_X1 _09907_ ( .A(_02276_ ), .B(_02210_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02277_ ) );
INV_X1 _09908_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02278_ ) );
NAND2_X1 _09909_ ( .A1(_02278_ ), .A2(fanout_net_19 ), .ZN(_02279_ ) );
OAI211_X1 _09910_ ( .A(_02279_ ), .B(fanout_net_26 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02280_ ) );
NAND3_X1 _09911_ ( .A1(_02277_ ), .A2(_02280_ ), .A3(_02166_ ), .ZN(_02281_ ) );
MUX2_X1 _09912_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02282_ ) );
MUX2_X1 _09913_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02283_ ) );
MUX2_X1 _09914_ ( .A(_02282_ ), .B(_02283_ ), .S(_02144_ ), .Z(_02284_ ) );
OAI211_X1 _09915_ ( .A(_02159_ ), .B(_02281_ ), .C1(_02284_ ), .C2(_02167_ ), .ZN(_02285_ ) );
OR2_X1 _09916_ ( .A1(_02135_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02286_ ) );
OAI211_X1 _09917_ ( .A(_02286_ ), .B(fanout_net_26 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02287_ ) );
OR2_X1 _09918_ ( .A1(_02135_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02288_ ) );
OAI211_X1 _09919_ ( .A(_02288_ ), .B(_02144_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02289_ ) );
NAND3_X1 _09920_ ( .A1(_02287_ ), .A2(_02289_ ), .A3(fanout_net_29 ), .ZN(_02290_ ) );
MUX2_X1 _09921_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02291_ ) );
MUX2_X1 _09922_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02292_ ) );
MUX2_X1 _09923_ ( .A(_02291_ ), .B(_02292_ ), .S(fanout_net_26 ), .Z(_02293_ ) );
OAI211_X1 _09924_ ( .A(fanout_net_30 ), .B(_02290_ ), .C1(_02293_ ), .C2(fanout_net_29 ), .ZN(_02294_ ) );
OAI211_X1 _09925_ ( .A(_02285_ ), .B(_02294_ ), .C1(_02184_ ), .C2(_02195_ ), .ZN(_02295_ ) );
NAND2_X1 _09926_ ( .A1(_02275_ ), .A2(_02295_ ), .ZN(_02296_ ) );
INV_X1 _09927_ ( .A(\ID_EX_imm [24] ), .ZN(_02297_ ) );
XNOR2_X1 _09928_ ( .A(_02296_ ), .B(_02297_ ), .ZN(_02298_ ) );
INV_X1 _09929_ ( .A(_02298_ ), .ZN(_02299_ ) );
OR3_X1 _09930_ ( .A1(_02184_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02195_ ), .ZN(_02300_ ) );
OR2_X1 _09931_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02301_ ) );
OAI211_X1 _09932_ ( .A(_02301_ ), .B(_02210_ ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02302_ ) );
OR2_X1 _09933_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02303_ ) );
OAI211_X1 _09934_ ( .A(_02303_ ), .B(fanout_net_26 ), .C1(fanout_net_19 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02304_ ) );
NAND3_X1 _09935_ ( .A1(_02302_ ), .A2(_02304_ ), .A3(fanout_net_29 ), .ZN(_02305_ ) );
MUX2_X1 _09936_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02306_ ) );
MUX2_X1 _09937_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02307_ ) );
MUX2_X1 _09938_ ( .A(_02306_ ), .B(_02307_ ), .S(_02210_ ), .Z(_02308_ ) );
OAI211_X1 _09939_ ( .A(_02159_ ), .B(_02305_ ), .C1(_02308_ ), .C2(fanout_net_29 ), .ZN(_02309_ ) );
NOR2_X1 _09940_ ( .A1(_02136_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02310_ ) );
OAI21_X1 _09941_ ( .A(fanout_net_26 ), .B1(fanout_net_19 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02311_ ) );
NOR2_X1 _09942_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02312_ ) );
OAI21_X1 _09943_ ( .A(_02210_ ), .B1(_02136_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02313_ ) );
OAI221_X1 _09944_ ( .A(_02166_ ), .B1(_02310_ ), .B2(_02311_ ), .C1(_02312_ ), .C2(_02313_ ), .ZN(_02314_ ) );
MUX2_X1 _09945_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02315_ ) );
MUX2_X1 _09946_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02316_ ) );
MUX2_X1 _09947_ ( .A(_02315_ ), .B(_02316_ ), .S(fanout_net_26 ), .Z(_02317_ ) );
OAI211_X1 _09948_ ( .A(fanout_net_30 ), .B(_02314_ ), .C1(_02317_ ), .C2(_02167_ ), .ZN(_02318_ ) );
OAI211_X1 _09949_ ( .A(_02309_ ), .B(_02318_ ), .C1(_02185_ ), .C2(_02196_ ), .ZN(_02319_ ) );
NAND2_X2 _09950_ ( .A1(_02300_ ), .A2(_02319_ ), .ZN(_02320_ ) );
INV_X1 _09951_ ( .A(\ID_EX_imm [25] ), .ZN(_02321_ ) );
XNOR2_X1 _09952_ ( .A(_02320_ ), .B(_02321_ ), .ZN(_02322_ ) );
INV_X1 _09953_ ( .A(_02322_ ), .ZN(_02323_ ) );
BUF_X8 _09954_ ( .A(_02181_ ), .Z(_02324_ ) );
CLKBUF_X3 _09955_ ( .A(_02324_ ), .Z(_02325_ ) );
BUF_X2 _09956_ ( .A(_02192_ ), .Z(_02326_ ) );
CLKBUF_X2 _09957_ ( .A(_02326_ ), .Z(_02327_ ) );
OR3_X1 _09958_ ( .A1(_02325_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02328_ ) );
CLKBUF_X2 _09959_ ( .A(_02134_ ), .Z(_02329_ ) );
OR2_X1 _09960_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02330_ ) );
OAI211_X1 _09961_ ( .A(_02330_ ), .B(_02144_ ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02331_ ) );
OR2_X1 _09962_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02332_ ) );
OAI211_X1 _09963_ ( .A(_02332_ ), .B(fanout_net_26 ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02333_ ) );
BUF_X4 _09964_ ( .A(_02165_ ), .Z(_02334_ ) );
NAND3_X1 _09965_ ( .A1(_02331_ ), .A2(_02333_ ), .A3(_02334_ ), .ZN(_02335_ ) );
MUX2_X1 _09966_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02336_ ) );
MUX2_X1 _09967_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02337_ ) );
BUF_X4 _09968_ ( .A(_02140_ ), .Z(_02338_ ) );
BUF_X4 _09969_ ( .A(_02338_ ), .Z(_02339_ ) );
BUF_X4 _09970_ ( .A(_02339_ ), .Z(_02340_ ) );
BUF_X4 _09971_ ( .A(_02340_ ), .Z(_02341_ ) );
MUX2_X1 _09972_ ( .A(_02336_ ), .B(_02337_ ), .S(_02341_ ), .Z(_02342_ ) );
OAI211_X1 _09973_ ( .A(_02159_ ), .B(_02335_ ), .C1(_02342_ ), .C2(_02166_ ), .ZN(_02343_ ) );
OR2_X1 _09974_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02344_ ) );
OAI211_X1 _09975_ ( .A(_02344_ ), .B(fanout_net_26 ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02345_ ) );
CLKBUF_X2 _09976_ ( .A(_02131_ ), .Z(_02346_ ) );
CLKBUF_X2 _09977_ ( .A(_02346_ ), .Z(_02347_ ) );
CLKBUF_X2 _09978_ ( .A(_02347_ ), .Z(_02348_ ) );
CLKBUF_X2 _09979_ ( .A(_02348_ ), .Z(_02349_ ) );
OR2_X1 _09980_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02350_ ) );
OAI211_X1 _09981_ ( .A(_02350_ ), .B(_02144_ ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02351_ ) );
NAND3_X1 _09982_ ( .A1(_02345_ ), .A2(_02351_ ), .A3(fanout_net_29 ), .ZN(_02352_ ) );
MUX2_X1 _09983_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02353_ ) );
MUX2_X1 _09984_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02354_ ) );
MUX2_X1 _09985_ ( .A(_02353_ ), .B(_02354_ ), .S(fanout_net_26 ), .Z(_02355_ ) );
OAI211_X1 _09986_ ( .A(fanout_net_30 ), .B(_02352_ ), .C1(_02355_ ), .C2(fanout_net_29 ), .ZN(_02356_ ) );
OAI211_X1 _09987_ ( .A(_02343_ ), .B(_02356_ ), .C1(_02184_ ), .C2(_02195_ ), .ZN(_02357_ ) );
NAND2_X2 _09988_ ( .A1(_02328_ ), .A2(_02357_ ), .ZN(_02358_ ) );
INV_X1 _09989_ ( .A(\ID_EX_imm [20] ), .ZN(_02359_ ) );
XNOR2_X1 _09990_ ( .A(_02358_ ), .B(_02359_ ), .ZN(_02360_ ) );
OR3_X1 _09991_ ( .A1(_02325_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02361_ ) );
INV_X1 _09992_ ( .A(\ID_EX_imm [21] ), .ZN(_02362_ ) );
OR2_X1 _09993_ ( .A1(_02134_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02363_ ) );
OAI211_X1 _09994_ ( .A(_02363_ ), .B(_02341_ ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02364_ ) );
OR2_X1 _09995_ ( .A1(_02134_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02365_ ) );
OAI211_X1 _09996_ ( .A(_02365_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02366_ ) );
NAND3_X1 _09997_ ( .A1(_02364_ ), .A2(_02366_ ), .A3(fanout_net_29 ), .ZN(_02367_ ) );
MUX2_X1 _09998_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02368_ ) );
MUX2_X1 _09999_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02369_ ) );
MUX2_X1 _10000_ ( .A(_02368_ ), .B(_02369_ ), .S(_02143_ ), .Z(_02370_ ) );
OAI211_X1 _10001_ ( .A(_02158_ ), .B(_02367_ ), .C1(_02370_ ), .C2(fanout_net_29 ), .ZN(_02371_ ) );
NOR2_X1 _10002_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02372_ ) );
OAI21_X1 _10003_ ( .A(fanout_net_26 ), .B1(fanout_net_20 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02373_ ) );
NOR2_X1 _10004_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02374_ ) );
OAI21_X1 _10005_ ( .A(_02143_ ), .B1(_02329_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02375_ ) );
OAI221_X1 _10006_ ( .A(_02334_ ), .B1(_02372_ ), .B2(_02373_ ), .C1(_02374_ ), .C2(_02375_ ), .ZN(_02376_ ) );
MUX2_X1 _10007_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02377_ ) );
MUX2_X1 _10008_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02378_ ) );
MUX2_X1 _10009_ ( .A(_02377_ ), .B(_02378_ ), .S(fanout_net_26 ), .Z(_02379_ ) );
OAI211_X1 _10010_ ( .A(fanout_net_30 ), .B(_02376_ ), .C1(_02379_ ), .C2(_02334_ ), .ZN(_02380_ ) );
OAI211_X1 _10011_ ( .A(_02371_ ), .B(_02380_ ), .C1(_02325_ ), .C2(_02327_ ), .ZN(_02381_ ) );
AND3_X1 _10012_ ( .A1(_02361_ ), .A2(_02362_ ), .A3(_02381_ ), .ZN(_02382_ ) );
AOI21_X1 _10013_ ( .A(_02362_ ), .B1(_02361_ ), .B2(_02381_ ), .ZN(_02383_ ) );
NOR2_X1 _10014_ ( .A1(_02382_ ), .A2(_02383_ ), .ZN(_02384_ ) );
AND2_X1 _10015_ ( .A1(_02360_ ), .A2(_02384_ ), .ZN(_02385_ ) );
OR3_X1 _10016_ ( .A1(_02183_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02194_ ), .ZN(_02386_ ) );
OR2_X1 _10017_ ( .A1(_02134_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02387_ ) );
OAI211_X1 _10018_ ( .A(_02387_ ), .B(_02143_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02388_ ) );
OR2_X1 _10019_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02389_ ) );
OAI211_X1 _10020_ ( .A(_02389_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02390_ ) );
NAND3_X1 _10021_ ( .A1(_02388_ ), .A2(_02390_ ), .A3(_02165_ ), .ZN(_02391_ ) );
MUX2_X1 _10022_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02392_ ) );
MUX2_X1 _10023_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02393_ ) );
MUX2_X1 _10024_ ( .A(_02392_ ), .B(_02393_ ), .S(_02340_ ), .Z(_02394_ ) );
OAI211_X1 _10025_ ( .A(_02158_ ), .B(_02391_ ), .C1(_02394_ ), .C2(_02165_ ), .ZN(_02395_ ) );
OR2_X1 _10026_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02396_ ) );
OAI211_X1 _10027_ ( .A(_02396_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02397_ ) );
OR2_X1 _10028_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02398_ ) );
OAI211_X1 _10029_ ( .A(_02398_ ), .B(_02143_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02399_ ) );
NAND3_X1 _10030_ ( .A1(_02397_ ), .A2(_02399_ ), .A3(fanout_net_29 ), .ZN(_02400_ ) );
MUX2_X1 _10031_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02401_ ) );
MUX2_X1 _10032_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02402_ ) );
MUX2_X1 _10033_ ( .A(_02401_ ), .B(_02402_ ), .S(fanout_net_26 ), .Z(_02403_ ) );
OAI211_X1 _10034_ ( .A(fanout_net_30 ), .B(_02400_ ), .C1(_02403_ ), .C2(fanout_net_29 ), .ZN(_02404_ ) );
OAI211_X1 _10035_ ( .A(_02395_ ), .B(_02404_ ), .C1(_02325_ ), .C2(_02327_ ), .ZN(_02405_ ) );
NAND2_X2 _10036_ ( .A1(_02386_ ), .A2(_02405_ ), .ZN(_02406_ ) );
INV_X1 _10037_ ( .A(\ID_EX_imm [23] ), .ZN(_02407_ ) );
XNOR2_X1 _10038_ ( .A(_02406_ ), .B(_02407_ ), .ZN(_02408_ ) );
OR3_X1 _10039_ ( .A1(_02325_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02409_ ) );
OR2_X1 _10040_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02410_ ) );
OAI211_X1 _10041_ ( .A(_02410_ ), .B(_02341_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02411_ ) );
OR2_X1 _10042_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02412_ ) );
OAI211_X1 _10043_ ( .A(_02412_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02413_ ) );
NAND3_X1 _10044_ ( .A1(_02411_ ), .A2(_02413_ ), .A3(_02334_ ), .ZN(_02414_ ) );
MUX2_X1 _10045_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02415_ ) );
MUX2_X1 _10046_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02416_ ) );
MUX2_X1 _10047_ ( .A(_02415_ ), .B(_02416_ ), .S(_02341_ ), .Z(_02417_ ) );
OAI211_X1 _10048_ ( .A(fanout_net_30 ), .B(_02414_ ), .C1(_02417_ ), .C2(_02166_ ), .ZN(_02418_ ) );
OR2_X1 _10049_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02419_ ) );
OAI211_X1 _10050_ ( .A(_02419_ ), .B(_02341_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02420_ ) );
OR2_X1 _10051_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02421_ ) );
OAI211_X1 _10052_ ( .A(_02421_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02422_ ) );
NAND3_X1 _10053_ ( .A1(_02420_ ), .A2(_02422_ ), .A3(_02334_ ), .ZN(_02423_ ) );
MUX2_X1 _10054_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02424_ ) );
MUX2_X1 _10055_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02425_ ) );
MUX2_X1 _10056_ ( .A(_02424_ ), .B(_02425_ ), .S(_02143_ ), .Z(_02426_ ) );
OAI211_X1 _10057_ ( .A(_02158_ ), .B(_02423_ ), .C1(_02426_ ), .C2(_02334_ ), .ZN(_02427_ ) );
OAI211_X1 _10058_ ( .A(_02418_ ), .B(_02427_ ), .C1(_02325_ ), .C2(_02327_ ), .ZN(_02428_ ) );
NAND2_X2 _10059_ ( .A1(_02409_ ), .A2(_02428_ ), .ZN(_02429_ ) );
INV_X1 _10060_ ( .A(\ID_EX_imm [22] ), .ZN(_02430_ ) );
XNOR2_X1 _10061_ ( .A(_02429_ ), .B(_02430_ ), .ZN(_02431_ ) );
AND3_X1 _10062_ ( .A1(_02385_ ), .A2(_02408_ ), .A3(_02431_ ), .ZN(_02432_ ) );
OR3_X1 _10063_ ( .A1(_02184_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02433_ ) );
OR2_X1 _10064_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02434_ ) );
OAI211_X1 _10065_ ( .A(_02434_ ), .B(_02144_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02435_ ) );
OR2_X1 _10066_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02436_ ) );
OAI211_X1 _10067_ ( .A(_02436_ ), .B(fanout_net_27 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02437_ ) );
NAND3_X1 _10068_ ( .A1(_02435_ ), .A2(_02437_ ), .A3(_02334_ ), .ZN(_02438_ ) );
MUX2_X1 _10069_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02439_ ) );
MUX2_X1 _10070_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02440_ ) );
MUX2_X1 _10071_ ( .A(_02439_ ), .B(_02440_ ), .S(_02341_ ), .Z(_02441_ ) );
OAI211_X1 _10072_ ( .A(_02159_ ), .B(_02438_ ), .C1(_02441_ ), .C2(_02166_ ), .ZN(_02442_ ) );
OR2_X1 _10073_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02443_ ) );
OAI211_X1 _10074_ ( .A(_02443_ ), .B(fanout_net_27 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02444_ ) );
OR2_X1 _10075_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02445_ ) );
OAI211_X1 _10076_ ( .A(_02445_ ), .B(_02144_ ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02446_ ) );
NAND3_X1 _10077_ ( .A1(_02444_ ), .A2(_02446_ ), .A3(fanout_net_29 ), .ZN(_02447_ ) );
MUX2_X1 _10078_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02448_ ) );
MUX2_X1 _10079_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02449_ ) );
MUX2_X1 _10080_ ( .A(_02448_ ), .B(_02449_ ), .S(fanout_net_27 ), .Z(_02450_ ) );
OAI211_X1 _10081_ ( .A(fanout_net_30 ), .B(_02447_ ), .C1(_02450_ ), .C2(fanout_net_29 ), .ZN(_02451_ ) );
OAI211_X1 _10082_ ( .A(_02442_ ), .B(_02451_ ), .C1(_02184_ ), .C2(_02195_ ), .ZN(_02452_ ) );
NAND2_X2 _10083_ ( .A1(_02433_ ), .A2(_02452_ ), .ZN(_02453_ ) );
INV_X1 _10084_ ( .A(\ID_EX_imm [16] ), .ZN(_02454_ ) );
XNOR2_X1 _10085_ ( .A(_02453_ ), .B(_02454_ ), .ZN(_02455_ ) );
OR3_X1 _10086_ ( .A1(_02325_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02456_ ) );
OR2_X1 _10087_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02457_ ) );
OAI211_X1 _10088_ ( .A(_02457_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02458_ ) );
OR2_X1 _10089_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02459_ ) );
OAI211_X1 _10090_ ( .A(_02459_ ), .B(_02341_ ), .C1(_02135_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02460_ ) );
NAND3_X1 _10091_ ( .A1(_02458_ ), .A2(fanout_net_29 ), .A3(_02460_ ), .ZN(_02461_ ) );
MUX2_X1 _10092_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02462_ ) );
MUX2_X1 _10093_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02463_ ) );
MUX2_X1 _10094_ ( .A(_02462_ ), .B(_02463_ ), .S(_02143_ ), .Z(_02464_ ) );
OAI211_X1 _10095_ ( .A(_02158_ ), .B(_02461_ ), .C1(_02464_ ), .C2(fanout_net_29 ), .ZN(_02465_ ) );
NOR2_X1 _10096_ ( .A1(_02329_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02466_ ) );
OAI21_X1 _10097_ ( .A(fanout_net_27 ), .B1(fanout_net_21 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02467_ ) );
NOR2_X1 _10098_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02468_ ) );
OAI21_X1 _10099_ ( .A(_02143_ ), .B1(_02135_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02469_ ) );
OAI221_X1 _10100_ ( .A(_02334_ ), .B1(_02466_ ), .B2(_02467_ ), .C1(_02468_ ), .C2(_02469_ ), .ZN(_02470_ ) );
MUX2_X1 _10101_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02471_ ) );
MUX2_X1 _10102_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02472_ ) );
MUX2_X1 _10103_ ( .A(_02471_ ), .B(_02472_ ), .S(fanout_net_27 ), .Z(_02473_ ) );
OAI211_X1 _10104_ ( .A(fanout_net_30 ), .B(_02470_ ), .C1(_02473_ ), .C2(_02334_ ), .ZN(_02474_ ) );
OAI211_X1 _10105_ ( .A(_02465_ ), .B(_02474_ ), .C1(_02325_ ), .C2(_02195_ ), .ZN(_02475_ ) );
NAND2_X1 _10106_ ( .A1(_02456_ ), .A2(_02475_ ), .ZN(_02476_ ) );
INV_X1 _10107_ ( .A(\ID_EX_imm [17] ), .ZN(_02477_ ) );
XNOR2_X1 _10108_ ( .A(_02476_ ), .B(_02477_ ), .ZN(_02478_ ) );
AND2_X1 _10109_ ( .A1(_02455_ ), .A2(_02478_ ), .ZN(_02479_ ) );
OR3_X1 _10110_ ( .A1(_02325_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02327_ ), .ZN(_02480_ ) );
OR2_X1 _10111_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02481_ ) );
OAI211_X1 _10112_ ( .A(_02481_ ), .B(_02341_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02482_ ) );
OR2_X1 _10113_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02483_ ) );
OAI211_X1 _10114_ ( .A(_02483_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02484_ ) );
NAND3_X1 _10115_ ( .A1(_02482_ ), .A2(_02484_ ), .A3(_02334_ ), .ZN(_02485_ ) );
MUX2_X1 _10116_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02486_ ) );
MUX2_X1 _10117_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02487_ ) );
MUX2_X1 _10118_ ( .A(_02486_ ), .B(_02487_ ), .S(_02341_ ), .Z(_02488_ ) );
OAI211_X1 _10119_ ( .A(_02158_ ), .B(_02485_ ), .C1(_02488_ ), .C2(_02166_ ), .ZN(_02489_ ) );
OR2_X1 _10120_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02490_ ) );
OAI211_X1 _10121_ ( .A(_02490_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02491_ ) );
OR2_X1 _10122_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02492_ ) );
OAI211_X1 _10123_ ( .A(_02492_ ), .B(_02341_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02493_ ) );
NAND3_X1 _10124_ ( .A1(_02491_ ), .A2(_02493_ ), .A3(fanout_net_29 ), .ZN(_02494_ ) );
MUX2_X1 _10125_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02495_ ) );
MUX2_X1 _10126_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02496_ ) );
MUX2_X1 _10127_ ( .A(_02495_ ), .B(_02496_ ), .S(fanout_net_27 ), .Z(_02497_ ) );
OAI211_X1 _10128_ ( .A(fanout_net_30 ), .B(_02494_ ), .C1(_02497_ ), .C2(fanout_net_29 ), .ZN(_02498_ ) );
OAI211_X1 _10129_ ( .A(_02489_ ), .B(_02498_ ), .C1(_02184_ ), .C2(_02195_ ), .ZN(_02499_ ) );
NAND2_X1 _10130_ ( .A1(_02480_ ), .A2(_02499_ ), .ZN(_02500_ ) );
BUF_X4 _10131_ ( .A(_02500_ ), .Z(_02501_ ) );
INV_X1 _10132_ ( .A(\ID_EX_imm [18] ), .ZN(_02502_ ) );
XNOR2_X1 _10133_ ( .A(_02501_ ), .B(_02502_ ), .ZN(_02503_ ) );
OR3_X1 _10134_ ( .A1(_02183_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02194_ ), .ZN(_02504_ ) );
OR2_X1 _10135_ ( .A1(_02134_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02505_ ) );
OAI211_X1 _10136_ ( .A(_02505_ ), .B(_02143_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02506_ ) );
OR2_X1 _10137_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02507_ ) );
OAI211_X1 _10138_ ( .A(_02507_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02508_ ) );
NAND3_X1 _10139_ ( .A1(_02506_ ), .A2(_02508_ ), .A3(_02165_ ), .ZN(_02509_ ) );
MUX2_X1 _10140_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02510_ ) );
MUX2_X1 _10141_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02511_ ) );
MUX2_X1 _10142_ ( .A(_02510_ ), .B(_02511_ ), .S(_02340_ ), .Z(_02512_ ) );
OAI211_X1 _10143_ ( .A(_02158_ ), .B(_02509_ ), .C1(_02512_ ), .C2(_02165_ ), .ZN(_02513_ ) );
OR2_X1 _10144_ ( .A1(_02134_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02514_ ) );
OAI211_X1 _10145_ ( .A(_02514_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02515_ ) );
OR2_X1 _10146_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02516_ ) );
OAI211_X1 _10147_ ( .A(_02516_ ), .B(_02143_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02517_ ) );
NAND3_X1 _10148_ ( .A1(_02515_ ), .A2(_02517_ ), .A3(fanout_net_29 ), .ZN(_02518_ ) );
MUX2_X1 _10149_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02519_ ) );
MUX2_X1 _10150_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02520_ ) );
MUX2_X1 _10151_ ( .A(_02519_ ), .B(_02520_ ), .S(fanout_net_27 ), .Z(_02521_ ) );
OAI211_X1 _10152_ ( .A(fanout_net_30 ), .B(_02518_ ), .C1(_02521_ ), .C2(fanout_net_29 ), .ZN(_02522_ ) );
OAI211_X1 _10153_ ( .A(_02513_ ), .B(_02522_ ), .C1(_02325_ ), .C2(_02327_ ), .ZN(_02523_ ) );
NAND2_X2 _10154_ ( .A1(_02504_ ), .A2(_02523_ ), .ZN(_02524_ ) );
INV_X1 _10155_ ( .A(\ID_EX_imm [19] ), .ZN(_02525_ ) );
XNOR2_X1 _10156_ ( .A(_02524_ ), .B(_02525_ ), .ZN(_02526_ ) );
AND2_X1 _10157_ ( .A1(_02503_ ), .A2(_02526_ ), .ZN(_02527_ ) );
AND2_X1 _10158_ ( .A1(_02479_ ), .A2(_02527_ ), .ZN(_02528_ ) );
OR3_X1 _10159_ ( .A1(_02324_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02326_ ), .ZN(_02529_ ) );
CLKBUF_X2 _10160_ ( .A(_02131_ ), .Z(_02530_ ) );
CLKBUF_X2 _10161_ ( .A(_02530_ ), .Z(_02531_ ) );
OR2_X1 _10162_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02532_ ) );
OAI211_X1 _10163_ ( .A(_02532_ ), .B(_02340_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02533_ ) );
OR2_X1 _10164_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02534_ ) );
OAI211_X1 _10165_ ( .A(_02534_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02535_ ) );
BUF_X4 _10166_ ( .A(_02163_ ), .Z(_02536_ ) );
BUF_X4 _10167_ ( .A(_02536_ ), .Z(_02537_ ) );
NAND3_X1 _10168_ ( .A1(_02533_ ), .A2(_02535_ ), .A3(_02537_ ), .ZN(_02538_ ) );
MUX2_X1 _10169_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02539_ ) );
MUX2_X1 _10170_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02540_ ) );
MUX2_X1 _10171_ ( .A(_02539_ ), .B(_02540_ ), .S(_02142_ ), .Z(_02541_ ) );
OAI211_X1 _10172_ ( .A(_02158_ ), .B(_02538_ ), .C1(_02541_ ), .C2(_02165_ ), .ZN(_02542_ ) );
OR2_X1 _10173_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02543_ ) );
OAI211_X1 _10174_ ( .A(_02543_ ), .B(fanout_net_27 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02544_ ) );
OR2_X1 _10175_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02545_ ) );
OAI211_X1 _10176_ ( .A(_02545_ ), .B(_02340_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02546_ ) );
NAND3_X1 _10177_ ( .A1(_02544_ ), .A2(_02546_ ), .A3(fanout_net_29 ), .ZN(_02547_ ) );
MUX2_X1 _10178_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02548_ ) );
MUX2_X1 _10179_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02549_ ) );
MUX2_X1 _10180_ ( .A(_02548_ ), .B(_02549_ ), .S(fanout_net_27 ), .Z(_02550_ ) );
OAI211_X1 _10181_ ( .A(fanout_net_30 ), .B(_02547_ ), .C1(_02550_ ), .C2(fanout_net_29 ), .ZN(_02551_ ) );
OAI211_X2 _10182_ ( .A(_02542_ ), .B(_02551_ ), .C1(_02183_ ), .C2(_02194_ ), .ZN(_02552_ ) );
NAND2_X2 _10183_ ( .A1(_02529_ ), .A2(_02552_ ), .ZN(_02553_ ) );
XOR2_X1 _10184_ ( .A(_02553_ ), .B(\ID_EX_imm [15] ), .Z(_02554_ ) );
OR3_X1 _10185_ ( .A1(_02324_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02326_ ), .ZN(_02555_ ) );
OR2_X1 _10186_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02556_ ) );
OAI211_X1 _10187_ ( .A(_02556_ ), .B(_02142_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02557_ ) );
OR2_X1 _10188_ ( .A1(_02133_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02558_ ) );
OAI211_X1 _10189_ ( .A(_02558_ ), .B(fanout_net_27 ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02559_ ) );
NAND3_X1 _10190_ ( .A1(_02557_ ), .A2(_02559_ ), .A3(_02537_ ), .ZN(_02560_ ) );
MUX2_X1 _10191_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02561_ ) );
MUX2_X1 _10192_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02562_ ) );
MUX2_X1 _10193_ ( .A(_02561_ ), .B(_02562_ ), .S(_02142_ ), .Z(_02563_ ) );
OAI211_X1 _10194_ ( .A(_02157_ ), .B(_02560_ ), .C1(_02563_ ), .C2(_02537_ ), .ZN(_02564_ ) );
OR2_X1 _10195_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02565_ ) );
OAI211_X1 _10196_ ( .A(_02565_ ), .B(_02142_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02566_ ) );
OR2_X1 _10197_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02567_ ) );
OAI211_X1 _10198_ ( .A(_02567_ ), .B(fanout_net_27 ), .C1(_02134_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02568_ ) );
NAND3_X1 _10199_ ( .A1(_02566_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02568_ ), .ZN(_02569_ ) );
MUX2_X1 _10200_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02570_ ) );
MUX2_X1 _10201_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02571_ ) );
MUX2_X1 _10202_ ( .A(_02570_ ), .B(_02571_ ), .S(fanout_net_27 ), .Z(_02572_ ) );
OAI211_X1 _10203_ ( .A(fanout_net_30 ), .B(_02569_ ), .C1(_02572_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02573_ ) );
OAI211_X4 _10204_ ( .A(_02564_ ), .B(_02573_ ), .C1(_02183_ ), .C2(_02194_ ), .ZN(_02574_ ) );
NAND2_X4 _10205_ ( .A1(_02555_ ), .A2(_02574_ ), .ZN(_02575_ ) );
INV_X1 _10206_ ( .A(\ID_EX_imm [14] ), .ZN(_02576_ ) );
XNOR2_X1 _10207_ ( .A(_02575_ ), .B(_02576_ ), .ZN(_02577_ ) );
NAND2_X1 _10208_ ( .A1(_02554_ ), .A2(_02577_ ), .ZN(_02578_ ) );
OR3_X1 _10209_ ( .A1(_02324_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02326_ ), .ZN(_02579_ ) );
OR2_X1 _10210_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02580_ ) );
OAI211_X1 _10211_ ( .A(_02580_ ), .B(_02340_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02581_ ) );
OR2_X1 _10212_ ( .A1(_02531_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02582_ ) );
OAI211_X1 _10213_ ( .A(_02582_ ), .B(fanout_net_27 ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02583_ ) );
NAND3_X1 _10214_ ( .A1(_02581_ ), .A2(_02583_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02584_ ) );
MUX2_X1 _10215_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02585_ ) );
MUX2_X1 _10216_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02586_ ) );
MUX2_X1 _10217_ ( .A(_02585_ ), .B(_02586_ ), .S(_02340_ ), .Z(_02587_ ) );
OAI211_X1 _10218_ ( .A(_02158_ ), .B(_02584_ ), .C1(_02587_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02588_ ) );
NOR2_X1 _10219_ ( .A1(_02134_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02589_ ) );
OAI21_X1 _10220_ ( .A(fanout_net_27 ), .B1(fanout_net_22 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02590_ ) );
NOR2_X1 _10221_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02591_ ) );
OAI21_X1 _10222_ ( .A(_02142_ ), .B1(_02134_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02592_ ) );
OAI221_X1 _10223_ ( .A(_02537_ ), .B1(_02589_ ), .B2(_02590_ ), .C1(_02591_ ), .C2(_02592_ ), .ZN(_02593_ ) );
MUX2_X1 _10224_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02594_ ) );
MUX2_X1 _10225_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02595_ ) );
MUX2_X1 _10226_ ( .A(_02594_ ), .B(_02595_ ), .S(fanout_net_27 ), .Z(_02596_ ) );
OAI211_X1 _10227_ ( .A(fanout_net_30 ), .B(_02593_ ), .C1(_02596_ ), .C2(_02165_ ), .ZN(_02597_ ) );
OAI211_X1 _10228_ ( .A(_02588_ ), .B(_02597_ ), .C1(_02183_ ), .C2(_02194_ ), .ZN(_02598_ ) );
NAND2_X1 _10229_ ( .A1(_02579_ ), .A2(_02598_ ), .ZN(_02599_ ) );
BUF_X2 _10230_ ( .A(_02599_ ), .Z(_02600_ ) );
XNOR2_X1 _10231_ ( .A(_02600_ ), .B(\ID_EX_imm [13] ), .ZN(_02601_ ) );
OR3_X1 _10232_ ( .A1(_02183_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02194_ ), .ZN(_02602_ ) );
OR2_X1 _10233_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02603_ ) );
OAI211_X1 _10234_ ( .A(_02603_ ), .B(_02340_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02604_ ) );
OR2_X1 _10235_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02605_ ) );
OAI211_X1 _10236_ ( .A(_02605_ ), .B(fanout_net_27 ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02606_ ) );
NAND3_X1 _10237_ ( .A1(_02604_ ), .A2(_02606_ ), .A3(_02165_ ), .ZN(_02607_ ) );
MUX2_X1 _10238_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02608_ ) );
MUX2_X1 _10239_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02609_ ) );
MUX2_X1 _10240_ ( .A(_02608_ ), .B(_02609_ ), .S(_02340_ ), .Z(_02610_ ) );
OAI211_X1 _10241_ ( .A(_02158_ ), .B(_02607_ ), .C1(_02610_ ), .C2(_02165_ ), .ZN(_02611_ ) );
OR2_X1 _10242_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02612_ ) );
OAI211_X1 _10243_ ( .A(_02612_ ), .B(fanout_net_27 ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02613_ ) );
OR2_X1 _10244_ ( .A1(_02348_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02614_ ) );
OAI211_X1 _10245_ ( .A(_02614_ ), .B(_02340_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02615_ ) );
NAND3_X1 _10246_ ( .A1(_02613_ ), .A2(_02615_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02616_ ) );
MUX2_X1 _10247_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02617_ ) );
MUX2_X1 _10248_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02618_ ) );
MUX2_X1 _10249_ ( .A(_02617_ ), .B(_02618_ ), .S(fanout_net_27 ), .Z(_02619_ ) );
OAI211_X1 _10250_ ( .A(fanout_net_30 ), .B(_02616_ ), .C1(_02619_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02620_ ) );
OAI211_X1 _10251_ ( .A(_02611_ ), .B(_02620_ ), .C1(_02183_ ), .C2(_02194_ ), .ZN(_02621_ ) );
NAND2_X2 _10252_ ( .A1(_02602_ ), .A2(_02621_ ), .ZN(_02622_ ) );
INV_X1 _10253_ ( .A(\ID_EX_imm [12] ), .ZN(_02623_ ) );
XNOR2_X1 _10254_ ( .A(_02622_ ), .B(_02623_ ), .ZN(_02624_ ) );
INV_X1 _10255_ ( .A(_02624_ ), .ZN(_02625_ ) );
OR3_X1 _10256_ ( .A1(_02578_ ), .A2(_02601_ ), .A3(_02625_ ), .ZN(_02626_ ) );
OR3_X1 _10257_ ( .A1(_02181_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02192_ ), .ZN(_02627_ ) );
OR2_X1 _10258_ ( .A1(_02132_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02628_ ) );
OAI211_X1 _10259_ ( .A(_02628_ ), .B(_02338_ ), .C1(fanout_net_22 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02629_ ) );
OR2_X1 _10260_ ( .A1(_02132_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02630_ ) );
OAI211_X1 _10261_ ( .A(_02630_ ), .B(fanout_net_27 ), .C1(fanout_net_22 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02631_ ) );
NAND3_X1 _10262_ ( .A1(_02629_ ), .A2(_02631_ ), .A3(_02536_ ), .ZN(_02632_ ) );
MUX2_X1 _10263_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02633_ ) );
MUX2_X1 _10264_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02634_ ) );
MUX2_X1 _10265_ ( .A(_02633_ ), .B(_02634_ ), .S(_02338_ ), .Z(_02635_ ) );
OAI211_X1 _10266_ ( .A(fanout_net_30 ), .B(_02632_ ), .C1(_02635_ ), .C2(_02536_ ), .ZN(_02636_ ) );
OR2_X1 _10267_ ( .A1(_02132_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02637_ ) );
OAI211_X1 _10268_ ( .A(_02637_ ), .B(_02338_ ), .C1(fanout_net_23 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02638_ ) );
OR2_X1 _10269_ ( .A1(_02132_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02639_ ) );
OAI211_X1 _10270_ ( .A(_02639_ ), .B(fanout_net_27 ), .C1(fanout_net_23 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02640_ ) );
NAND3_X1 _10271_ ( .A1(_02638_ ), .A2(_02640_ ), .A3(_02163_ ), .ZN(_02641_ ) );
MUX2_X1 _10272_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02642_ ) );
MUX2_X1 _10273_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02643_ ) );
MUX2_X1 _10274_ ( .A(_02642_ ), .B(_02643_ ), .S(_02338_ ), .Z(_02644_ ) );
OAI211_X1 _10275_ ( .A(_02157_ ), .B(_02641_ ), .C1(_02644_ ), .C2(_02536_ ), .ZN(_02645_ ) );
OAI211_X1 _10276_ ( .A(_02636_ ), .B(_02645_ ), .C1(_02182_ ), .C2(_02193_ ), .ZN(_02646_ ) );
NAND2_X1 _10277_ ( .A1(_02627_ ), .A2(_02646_ ), .ZN(_02647_ ) );
INV_X1 _10278_ ( .A(\ID_EX_imm [8] ), .ZN(_02648_ ) );
XNOR2_X1 _10279_ ( .A(_02647_ ), .B(_02648_ ), .ZN(_02649_ ) );
OR3_X1 _10280_ ( .A1(_02181_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02192_ ), .ZN(_02650_ ) );
OR2_X1 _10281_ ( .A1(_02132_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02651_ ) );
OAI211_X1 _10282_ ( .A(_02651_ ), .B(_02338_ ), .C1(fanout_net_23 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02652_ ) );
OR2_X1 _10283_ ( .A1(_02132_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02653_ ) );
OAI211_X1 _10284_ ( .A(_02653_ ), .B(fanout_net_27 ), .C1(fanout_net_23 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02654_ ) );
NAND3_X1 _10285_ ( .A1(_02652_ ), .A2(_02654_ ), .A3(_02163_ ), .ZN(_02655_ ) );
MUX2_X1 _10286_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02656_ ) );
MUX2_X1 _10287_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02657_ ) );
MUX2_X1 _10288_ ( .A(_02656_ ), .B(_02657_ ), .S(_02140_ ), .Z(_02658_ ) );
OAI211_X1 _10289_ ( .A(_02156_ ), .B(_02655_ ), .C1(_02658_ ), .C2(_02536_ ), .ZN(_02659_ ) );
OR2_X1 _10290_ ( .A1(_02132_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02660_ ) );
OAI211_X1 _10291_ ( .A(_02660_ ), .B(fanout_net_27 ), .C1(fanout_net_23 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02661_ ) );
OR2_X1 _10292_ ( .A1(_02346_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02662_ ) );
OAI211_X1 _10293_ ( .A(_02662_ ), .B(_02338_ ), .C1(fanout_net_23 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02663_ ) );
NAND3_X1 _10294_ ( .A1(_02661_ ), .A2(_02663_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02664_ ) );
MUX2_X1 _10295_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02665_ ) );
MUX2_X1 _10296_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02666_ ) );
MUX2_X1 _10297_ ( .A(_02665_ ), .B(_02666_ ), .S(fanout_net_27 ), .Z(_02667_ ) );
OAI211_X1 _10298_ ( .A(fanout_net_30 ), .B(_02664_ ), .C1(_02667_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02668_ ) );
OAI211_X1 _10299_ ( .A(_02659_ ), .B(_02668_ ), .C1(_02182_ ), .C2(_02193_ ), .ZN(_02669_ ) );
NAND2_X2 _10300_ ( .A1(_02650_ ), .A2(_02669_ ), .ZN(_02670_ ) );
INV_X1 _10301_ ( .A(\ID_EX_imm [9] ), .ZN(_02671_ ) );
XNOR2_X1 _10302_ ( .A(_02670_ ), .B(_02671_ ), .ZN(_02672_ ) );
AND2_X1 _10303_ ( .A1(_02649_ ), .A2(_02672_ ), .ZN(_02673_ ) );
OR3_X4 _10304_ ( .A1(_02182_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_02193_ ), .ZN(_02674_ ) );
OR2_X1 _10305_ ( .A1(_02530_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02675_ ) );
OAI211_X1 _10306_ ( .A(_02675_ ), .B(_02141_ ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02676_ ) );
OR2_X1 _10307_ ( .A1(_02132_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02677_ ) );
OAI211_X1 _10308_ ( .A(_02677_ ), .B(fanout_net_27 ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02678_ ) );
NAND3_X1 _10309_ ( .A1(_02676_ ), .A2(_02678_ ), .A3(_02536_ ), .ZN(_02679_ ) );
MUX2_X1 _10310_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02680_ ) );
MUX2_X1 _10311_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02681_ ) );
MUX2_X1 _10312_ ( .A(_02680_ ), .B(_02681_ ), .S(_02338_ ), .Z(_02682_ ) );
OAI211_X1 _10313_ ( .A(_02157_ ), .B(_02679_ ), .C1(_02682_ ), .C2(_02164_ ), .ZN(_02683_ ) );
OR2_X1 _10314_ ( .A1(_02530_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02684_ ) );
OAI211_X1 _10315_ ( .A(_02684_ ), .B(fanout_net_28 ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02685_ ) );
OR2_X1 _10316_ ( .A1(_02132_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02686_ ) );
OAI211_X1 _10317_ ( .A(_02686_ ), .B(_02141_ ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02687_ ) );
NAND3_X1 _10318_ ( .A1(_02685_ ), .A2(_02687_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02688_ ) );
MUX2_X1 _10319_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02689_ ) );
MUX2_X1 _10320_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02690_ ) );
MUX2_X1 _10321_ ( .A(_02689_ ), .B(_02690_ ), .S(fanout_net_28 ), .Z(_02691_ ) );
OAI211_X1 _10322_ ( .A(fanout_net_30 ), .B(_02688_ ), .C1(_02691_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02692_ ) );
OAI211_X1 _10323_ ( .A(_02683_ ), .B(_02692_ ), .C1(_02182_ ), .C2(_02326_ ), .ZN(_02693_ ) );
NAND2_X4 _10324_ ( .A1(_02674_ ), .A2(_02693_ ), .ZN(_02694_ ) );
INV_X1 _10325_ ( .A(\ID_EX_imm [11] ), .ZN(_02695_ ) );
XNOR2_X1 _10326_ ( .A(_02694_ ), .B(_02695_ ), .ZN(_02696_ ) );
OR3_X1 _10327_ ( .A1(_02324_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02326_ ), .ZN(_02697_ ) );
OR2_X1 _10328_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02698_ ) );
OAI211_X1 _10329_ ( .A(_02698_ ), .B(_02142_ ), .C1(fanout_net_23 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02699_ ) );
OR2_X1 _10330_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02700_ ) );
OAI211_X1 _10331_ ( .A(_02700_ ), .B(fanout_net_28 ), .C1(fanout_net_23 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02701_ ) );
NAND3_X1 _10332_ ( .A1(_02699_ ), .A2(_02701_ ), .A3(_02164_ ), .ZN(_02702_ ) );
MUX2_X1 _10333_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02703_ ) );
MUX2_X1 _10334_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02704_ ) );
MUX2_X1 _10335_ ( .A(_02703_ ), .B(_02704_ ), .S(_02339_ ), .Z(_02705_ ) );
OAI211_X1 _10336_ ( .A(_02157_ ), .B(_02702_ ), .C1(_02705_ ), .C2(_02537_ ), .ZN(_02706_ ) );
OR2_X1 _10337_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02707_ ) );
OAI211_X1 _10338_ ( .A(_02707_ ), .B(fanout_net_28 ), .C1(fanout_net_23 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02708_ ) );
OR2_X1 _10339_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02709_ ) );
OAI211_X1 _10340_ ( .A(_02709_ ), .B(_02142_ ), .C1(fanout_net_23 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02710_ ) );
NAND3_X1 _10341_ ( .A1(_02708_ ), .A2(_02710_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02711_ ) );
MUX2_X1 _10342_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02712_ ) );
MUX2_X1 _10343_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02713_ ) );
MUX2_X1 _10344_ ( .A(_02712_ ), .B(_02713_ ), .S(fanout_net_28 ), .Z(_02714_ ) );
OAI211_X1 _10345_ ( .A(fanout_net_30 ), .B(_02711_ ), .C1(_02714_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02715_ ) );
OAI211_X1 _10346_ ( .A(_02706_ ), .B(_02715_ ), .C1(_02183_ ), .C2(_02194_ ), .ZN(_02716_ ) );
NAND2_X1 _10347_ ( .A1(_02697_ ), .A2(_02716_ ), .ZN(_02717_ ) );
BUF_X4 _10348_ ( .A(_02717_ ), .Z(_02718_ ) );
XOR2_X1 _10349_ ( .A(_02718_ ), .B(\ID_EX_imm [10] ), .Z(_02719_ ) );
NAND3_X1 _10350_ ( .A1(_02673_ ), .A2(_02696_ ), .A3(_02719_ ), .ZN(_02720_ ) );
OR3_X1 _10351_ ( .A1(_02182_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02193_ ), .ZN(_02721_ ) );
OR2_X1 _10352_ ( .A1(_02347_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02722_ ) );
OAI211_X1 _10353_ ( .A(_02722_ ), .B(_02339_ ), .C1(fanout_net_23 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02723_ ) );
OR2_X1 _10354_ ( .A1(_02347_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02724_ ) );
OAI211_X1 _10355_ ( .A(_02724_ ), .B(fanout_net_28 ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02725_ ) );
NAND3_X1 _10356_ ( .A1(_02723_ ), .A2(_02725_ ), .A3(_02164_ ), .ZN(_02726_ ) );
MUX2_X1 _10357_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02727_ ) );
MUX2_X1 _10358_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02728_ ) );
MUX2_X1 _10359_ ( .A(_02727_ ), .B(_02728_ ), .S(_02141_ ), .Z(_02729_ ) );
OAI211_X1 _10360_ ( .A(_02157_ ), .B(_02726_ ), .C1(_02729_ ), .C2(_02164_ ), .ZN(_02730_ ) );
OR2_X1 _10361_ ( .A1(_02347_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02731_ ) );
OAI211_X1 _10362_ ( .A(_02731_ ), .B(fanout_net_28 ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02732_ ) );
OR2_X1 _10363_ ( .A1(_02530_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02733_ ) );
OAI211_X1 _10364_ ( .A(_02733_ ), .B(_02141_ ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02734_ ) );
NAND3_X1 _10365_ ( .A1(_02732_ ), .A2(_02734_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02735_ ) );
MUX2_X1 _10366_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02736_ ) );
MUX2_X1 _10367_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02737_ ) );
MUX2_X1 _10368_ ( .A(_02736_ ), .B(_02737_ ), .S(fanout_net_28 ), .Z(_02738_ ) );
OAI211_X1 _10369_ ( .A(fanout_net_30 ), .B(_02735_ ), .C1(_02738_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02739_ ) );
OAI211_X1 _10370_ ( .A(_02730_ ), .B(_02739_ ), .C1(_02324_ ), .C2(_02326_ ), .ZN(_02740_ ) );
NAND2_X1 _10371_ ( .A1(_02721_ ), .A2(_02740_ ), .ZN(_02741_ ) );
INV_X1 _10372_ ( .A(\ID_EX_imm [2] ), .ZN(_02742_ ) );
XNOR2_X1 _10373_ ( .A(_02741_ ), .B(_02742_ ), .ZN(_02743_ ) );
OR3_X1 _10374_ ( .A1(_02181_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02192_ ), .ZN(_02744_ ) );
OR2_X1 _10375_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02745_ ) );
OAI211_X1 _10376_ ( .A(_02745_ ), .B(_02338_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02746_ ) );
OR2_X1 _10377_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02747_ ) );
OAI211_X1 _10378_ ( .A(_02747_ ), .B(fanout_net_28 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02748_ ) );
NAND3_X1 _10379_ ( .A1(_02746_ ), .A2(_02748_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02749_ ) );
MUX2_X1 _10380_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02750_ ) );
MUX2_X1 _10381_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02751_ ) );
MUX2_X1 _10382_ ( .A(_02750_ ), .B(_02751_ ), .S(_02140_ ), .Z(_02752_ ) );
OAI211_X1 _10383_ ( .A(_02156_ ), .B(_02749_ ), .C1(_02752_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02753_ ) );
NOR2_X1 _10384_ ( .A1(_02530_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02754_ ) );
OAI21_X1 _10385_ ( .A(fanout_net_28 ), .B1(fanout_net_24 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02755_ ) );
NOR2_X1 _10386_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02756_ ) );
OAI21_X1 _10387_ ( .A(_02140_ ), .B1(_02530_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02757_ ) );
OAI221_X1 _10388_ ( .A(_02163_ ), .B1(_02754_ ), .B2(_02755_ ), .C1(_02756_ ), .C2(_02757_ ), .ZN(_02758_ ) );
MUX2_X1 _10389_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02759_ ) );
MUX2_X1 _10390_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02760_ ) );
MUX2_X1 _10391_ ( .A(_02759_ ), .B(_02760_ ), .S(fanout_net_28 ), .Z(_02761_ ) );
OAI211_X1 _10392_ ( .A(fanout_net_30 ), .B(_02758_ ), .C1(_02761_ ), .C2(_02536_ ), .ZN(_02762_ ) );
OAI211_X1 _10393_ ( .A(_02753_ ), .B(_02762_ ), .C1(_02181_ ), .C2(_02192_ ), .ZN(_02763_ ) );
NAND2_X2 _10394_ ( .A1(_02744_ ), .A2(_02763_ ), .ZN(_02764_ ) );
INV_X1 _10395_ ( .A(\ID_EX_imm [1] ), .ZN(_02765_ ) );
XNOR2_X1 _10396_ ( .A(_02764_ ), .B(_02765_ ), .ZN(_02766_ ) );
NOR2_X1 _10397_ ( .A1(_02182_ ), .A2(_02193_ ), .ZN(_02767_ ) );
NAND2_X1 _10398_ ( .A1(_02767_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_02768_ ) );
OR2_X1 _10399_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02769_ ) );
OAI211_X1 _10400_ ( .A(_02769_ ), .B(_02142_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(fanout_net_24 ), .ZN(_02770_ ) );
OR2_X1 _10401_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02771_ ) );
OAI211_X1 _10402_ ( .A(_02771_ ), .B(fanout_net_28 ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02772_ ) );
NAND3_X1 _10403_ ( .A1(_02770_ ), .A2(_02772_ ), .A3(_02164_ ), .ZN(_02773_ ) );
MUX2_X1 _10404_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02774_ ) );
MUX2_X1 _10405_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02775_ ) );
MUX2_X1 _10406_ ( .A(_02774_ ), .B(_02775_ ), .S(_02339_ ), .Z(_02776_ ) );
OAI211_X1 _10407_ ( .A(_02157_ ), .B(_02773_ ), .C1(_02776_ ), .C2(_02537_ ), .ZN(_02777_ ) );
OR2_X1 _10408_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02778_ ) );
OAI211_X1 _10409_ ( .A(_02778_ ), .B(fanout_net_28 ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02779_ ) );
OR2_X1 _10410_ ( .A1(_02133_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02780_ ) );
OAI211_X1 _10411_ ( .A(_02780_ ), .B(_02142_ ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02781_ ) );
NAND3_X1 _10412_ ( .A1(_02779_ ), .A2(_02781_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02782_ ) );
MUX2_X1 _10413_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02783_ ) );
MUX2_X1 _10414_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02784_ ) );
MUX2_X1 _10415_ ( .A(_02783_ ), .B(_02784_ ), .S(fanout_net_28 ), .Z(_02785_ ) );
OAI211_X1 _10416_ ( .A(fanout_net_30 ), .B(_02782_ ), .C1(_02785_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02786_ ) );
NAND2_X1 _10417_ ( .A1(_02777_ ), .A2(_02786_ ), .ZN(_02787_ ) );
OAI21_X1 _10418_ ( .A(_02787_ ), .B1(_02183_ ), .B2(_02194_ ), .ZN(_02788_ ) );
AND3_X1 _10419_ ( .A1(_02768_ ), .A2(\ID_EX_imm [0] ), .A3(_02788_ ), .ZN(_02789_ ) );
AND2_X1 _10420_ ( .A1(_02766_ ), .A2(_02789_ ), .ZN(_02790_ ) );
AOI21_X1 _10421_ ( .A(_02765_ ), .B1(_02744_ ), .B2(_02763_ ), .ZN(_02791_ ) );
OAI21_X1 _10422_ ( .A(_02743_ ), .B1(_02790_ ), .B2(_02791_ ), .ZN(_02792_ ) );
INV_X1 _10423_ ( .A(_02741_ ), .ZN(_02793_ ) );
OAI21_X1 _10424_ ( .A(_02792_ ), .B1(_02742_ ), .B2(_02793_ ), .ZN(_02794_ ) );
OR3_X1 _10425_ ( .A1(_02182_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02193_ ), .ZN(_02795_ ) );
OR2_X1 _10426_ ( .A1(_02347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02796_ ) );
OAI211_X1 _10427_ ( .A(_02796_ ), .B(_02339_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02797_ ) );
OR2_X1 _10428_ ( .A1(_02347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02798_ ) );
OAI211_X1 _10429_ ( .A(_02798_ ), .B(fanout_net_28 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02799_ ) );
NAND3_X1 _10430_ ( .A1(_02797_ ), .A2(_02799_ ), .A3(_02164_ ), .ZN(_02800_ ) );
MUX2_X1 _10431_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02801_ ) );
MUX2_X1 _10432_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02802_ ) );
MUX2_X1 _10433_ ( .A(_02801_ ), .B(_02802_ ), .S(_02141_ ), .Z(_02803_ ) );
OAI211_X1 _10434_ ( .A(fanout_net_30 ), .B(_02800_ ), .C1(_02803_ ), .C2(_02537_ ), .ZN(_02804_ ) );
OR2_X1 _10435_ ( .A1(_02347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02805_ ) );
OAI211_X1 _10436_ ( .A(_02805_ ), .B(_02339_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02806_ ) );
OR2_X1 _10437_ ( .A1(_02347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02807_ ) );
OAI211_X1 _10438_ ( .A(_02807_ ), .B(fanout_net_28 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02808_ ) );
NAND3_X1 _10439_ ( .A1(_02806_ ), .A2(_02808_ ), .A3(_02164_ ), .ZN(_02809_ ) );
MUX2_X1 _10440_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02810_ ) );
MUX2_X1 _10441_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02811_ ) );
MUX2_X1 _10442_ ( .A(_02810_ ), .B(_02811_ ), .S(_02141_ ), .Z(_02812_ ) );
OAI211_X1 _10443_ ( .A(_02157_ ), .B(_02809_ ), .C1(_02812_ ), .C2(_02537_ ), .ZN(_02813_ ) );
OAI211_X1 _10444_ ( .A(_02804_ ), .B(_02813_ ), .C1(_02324_ ), .C2(_02326_ ), .ZN(_02814_ ) );
NAND2_X2 _10445_ ( .A1(_02795_ ), .A2(_02814_ ), .ZN(_02815_ ) );
INV_X1 _10446_ ( .A(\ID_EX_imm [3] ), .ZN(_02816_ ) );
XNOR2_X1 _10447_ ( .A(_02815_ ), .B(_02816_ ), .ZN(_02817_ ) );
NAND2_X1 _10448_ ( .A1(_02794_ ), .A2(_02817_ ), .ZN(_02818_ ) );
INV_X1 _10449_ ( .A(_02815_ ), .ZN(_02819_ ) );
OR2_X1 _10450_ ( .A1(_02819_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02820_ ) );
NAND2_X1 _10451_ ( .A1(_02818_ ), .A2(_02820_ ), .ZN(_02821_ ) );
OR3_X1 _10452_ ( .A1(_02182_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02193_ ), .ZN(_02822_ ) );
OR2_X1 _10453_ ( .A1(_02530_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02823_ ) );
OAI211_X1 _10454_ ( .A(_02823_ ), .B(_02141_ ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02824_ ) );
OR2_X1 _10455_ ( .A1(_02530_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02825_ ) );
OAI211_X1 _10456_ ( .A(_02825_ ), .B(fanout_net_28 ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02826_ ) );
NAND3_X1 _10457_ ( .A1(_02824_ ), .A2(_02826_ ), .A3(_02536_ ), .ZN(_02827_ ) );
MUX2_X1 _10458_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02828_ ) );
MUX2_X1 _10459_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02829_ ) );
MUX2_X1 _10460_ ( .A(_02828_ ), .B(_02829_ ), .S(_02141_ ), .Z(_02830_ ) );
OAI211_X1 _10461_ ( .A(_02157_ ), .B(_02827_ ), .C1(_02830_ ), .C2(_02164_ ), .ZN(_02831_ ) );
OR2_X1 _10462_ ( .A1(_02530_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02832_ ) );
OAI211_X1 _10463_ ( .A(_02832_ ), .B(fanout_net_28 ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02833_ ) );
OR2_X1 _10464_ ( .A1(_02530_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02834_ ) );
OAI211_X1 _10465_ ( .A(_02834_ ), .B(_02141_ ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02835_ ) );
NAND3_X1 _10466_ ( .A1(_02833_ ), .A2(_02835_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02836_ ) );
MUX2_X1 _10467_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02837_ ) );
MUX2_X1 _10468_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02838_ ) );
MUX2_X1 _10469_ ( .A(_02837_ ), .B(_02838_ ), .S(fanout_net_28 ), .Z(_02839_ ) );
OAI211_X1 _10470_ ( .A(fanout_net_30 ), .B(_02836_ ), .C1(_02839_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02840_ ) );
OAI211_X1 _10471_ ( .A(_02831_ ), .B(_02840_ ), .C1(_02324_ ), .C2(_02326_ ), .ZN(_02841_ ) );
NAND2_X1 _10472_ ( .A1(_02822_ ), .A2(_02841_ ), .ZN(_02842_ ) );
INV_X1 _10473_ ( .A(\ID_EX_imm [4] ), .ZN(_02843_ ) );
XNOR2_X1 _10474_ ( .A(_02842_ ), .B(_02843_ ), .ZN(_02844_ ) );
NAND2_X1 _10475_ ( .A1(_02821_ ), .A2(_02844_ ), .ZN(_02845_ ) );
NAND2_X1 _10476_ ( .A1(_02767_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02846_ ) );
OR2_X1 _10477_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02847_ ) );
OAI211_X1 _10478_ ( .A(_02847_ ), .B(_02338_ ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02848_ ) );
OR2_X1 _10479_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02849_ ) );
OAI211_X1 _10480_ ( .A(_02849_ ), .B(fanout_net_28 ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02850_ ) );
NAND3_X1 _10481_ ( .A1(_02848_ ), .A2(_02850_ ), .A3(_02163_ ), .ZN(_02851_ ) );
MUX2_X1 _10482_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02852_ ) );
MUX2_X1 _10483_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02853_ ) );
MUX2_X1 _10484_ ( .A(_02852_ ), .B(_02853_ ), .S(_02140_ ), .Z(_02854_ ) );
OAI211_X1 _10485_ ( .A(_02156_ ), .B(_02851_ ), .C1(_02854_ ), .C2(_02536_ ), .ZN(_02855_ ) );
OR2_X1 _10486_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02856_ ) );
OAI211_X1 _10487_ ( .A(_02856_ ), .B(fanout_net_28 ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02857_ ) );
OR2_X1 _10488_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02858_ ) );
OAI211_X1 _10489_ ( .A(_02858_ ), .B(_02140_ ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02859_ ) );
NAND3_X1 _10490_ ( .A1(_02857_ ), .A2(_02859_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02860_ ) );
MUX2_X1 _10491_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02861_ ) );
MUX2_X1 _10492_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02862_ ) );
MUX2_X1 _10493_ ( .A(_02861_ ), .B(_02862_ ), .S(fanout_net_28 ), .Z(_02863_ ) );
OAI211_X1 _10494_ ( .A(fanout_net_30 ), .B(_02860_ ), .C1(_02863_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02864_ ) );
NAND2_X1 _10495_ ( .A1(_02855_ ), .A2(_02864_ ), .ZN(_02865_ ) );
OAI21_X1 _10496_ ( .A(_02865_ ), .B1(_02182_ ), .B2(_02193_ ), .ZN(_02866_ ) );
AND2_X2 _10497_ ( .A1(_02846_ ), .A2(_02866_ ), .ZN(_02867_ ) );
XNOR2_X1 _10498_ ( .A(_02867_ ), .B(\ID_EX_imm [5] ), .ZN(_02868_ ) );
NOR2_X1 _10499_ ( .A1(_02845_ ), .A2(_02868_ ), .ZN(_02869_ ) );
OR3_X1 _10500_ ( .A1(_02324_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02193_ ), .ZN(_02870_ ) );
OR2_X1 _10501_ ( .A1(_02347_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02871_ ) );
OAI211_X1 _10502_ ( .A(_02871_ ), .B(_02339_ ), .C1(fanout_net_25 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02872_ ) );
OR2_X1 _10503_ ( .A1(_02347_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02873_ ) );
OAI211_X1 _10504_ ( .A(_02873_ ), .B(fanout_net_28 ), .C1(fanout_net_25 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02874_ ) );
NAND3_X1 _10505_ ( .A1(_02872_ ), .A2(_02874_ ), .A3(_02164_ ), .ZN(_02875_ ) );
MUX2_X1 _10506_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02876_ ) );
MUX2_X1 _10507_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02877_ ) );
MUX2_X1 _10508_ ( .A(_02876_ ), .B(_02877_ ), .S(_02339_ ), .Z(_02878_ ) );
OAI211_X1 _10509_ ( .A(fanout_net_30 ), .B(_02875_ ), .C1(_02878_ ), .C2(_02537_ ), .ZN(_02879_ ) );
NOR2_X1 _10510_ ( .A1(_02531_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02880_ ) );
OAI21_X1 _10511_ ( .A(fanout_net_28 ), .B1(fanout_net_25 ), .B2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02881_ ) );
NOR2_X1 _10512_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02882_ ) );
OAI21_X1 _10513_ ( .A(_02339_ ), .B1(_02531_ ), .B2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02883_ ) );
OAI221_X1 _10514_ ( .A(_02536_ ), .B1(_02880_ ), .B2(_02881_ ), .C1(_02882_ ), .C2(_02883_ ), .ZN(_02884_ ) );
MUX2_X1 _10515_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02885_ ) );
MUX2_X1 _10516_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02886_ ) );
MUX2_X1 _10517_ ( .A(_02885_ ), .B(_02886_ ), .S(_02339_ ), .Z(_02887_ ) );
OAI211_X1 _10518_ ( .A(_02157_ ), .B(_02884_ ), .C1(_02887_ ), .C2(_02537_ ), .ZN(_02888_ ) );
OAI211_X1 _10519_ ( .A(_02879_ ), .B(_02888_ ), .C1(_02324_ ), .C2(_02326_ ), .ZN(_02889_ ) );
NAND2_X2 _10520_ ( .A1(_02870_ ), .A2(_02889_ ), .ZN(_02890_ ) );
INV_X1 _10521_ ( .A(\ID_EX_imm [6] ), .ZN(_02891_ ) );
XNOR2_X1 _10522_ ( .A(_02890_ ), .B(_02891_ ), .ZN(_02892_ ) );
INV_X1 _10523_ ( .A(_02892_ ), .ZN(_02893_ ) );
OR3_X1 _10524_ ( .A1(_02181_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02192_ ), .ZN(_02894_ ) );
OR2_X1 _10525_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02895_ ) );
OAI211_X1 _10526_ ( .A(_02895_ ), .B(_02140_ ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02896_ ) );
OR2_X1 _10527_ ( .A1(_02131_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02897_ ) );
OAI211_X1 _10528_ ( .A(_02897_ ), .B(fanout_net_28 ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02898_ ) );
NAND3_X1 _10529_ ( .A1(_02896_ ), .A2(_02898_ ), .A3(_02163_ ), .ZN(_02899_ ) );
MUX2_X1 _10530_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02900_ ) );
MUX2_X1 _10531_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02901_ ) );
MUX2_X1 _10532_ ( .A(_02900_ ), .B(_02901_ ), .S(_02140_ ), .Z(_02902_ ) );
OAI211_X1 _10533_ ( .A(_02156_ ), .B(_02899_ ), .C1(_02902_ ), .C2(_02163_ ), .ZN(_02903_ ) );
OR2_X1 _10534_ ( .A1(_02346_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02904_ ) );
OAI211_X1 _10535_ ( .A(_02904_ ), .B(fanout_net_28 ), .C1(fanout_net_25 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02905_ ) );
OR2_X1 _10536_ ( .A1(_02131_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02906_ ) );
OAI211_X1 _10537_ ( .A(_02906_ ), .B(_02140_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02907_ ) );
NAND3_X1 _10538_ ( .A1(_02905_ ), .A2(_02907_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02908_ ) );
MUX2_X1 _10539_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02909_ ) );
MUX2_X1 _10540_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02910_ ) );
MUX2_X1 _10541_ ( .A(_02909_ ), .B(_02910_ ), .S(fanout_net_28 ), .Z(_02911_ ) );
OAI211_X1 _10542_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02908_ ), .C1(_02911_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02912_ ) );
OAI211_X1 _10543_ ( .A(_02903_ ), .B(_02912_ ), .C1(_02181_ ), .C2(_02192_ ), .ZN(_02913_ ) );
NAND2_X1 _10544_ ( .A1(_02894_ ), .A2(_02913_ ), .ZN(_02914_ ) );
XNOR2_X1 _10545_ ( .A(_02914_ ), .B(\ID_EX_imm [7] ), .ZN(_02915_ ) );
NOR2_X1 _10546_ ( .A1(_02893_ ), .A2(_02915_ ), .ZN(_02916_ ) );
NAND2_X1 _10547_ ( .A1(_02869_ ), .A2(_02916_ ), .ZN(_02917_ ) );
INV_X1 _10548_ ( .A(_02890_ ), .ZN(_02918_ ) );
NOR3_X1 _10549_ ( .A1(_02915_ ), .A2(_02891_ ), .A3(_02918_ ), .ZN(_02919_ ) );
AND2_X1 _10550_ ( .A1(_02842_ ), .A2(\ID_EX_imm [4] ), .ZN(_02920_ ) );
INV_X1 _10551_ ( .A(_02920_ ), .ZN(_02921_ ) );
OR2_X1 _10552_ ( .A1(_02868_ ), .A2(_02921_ ), .ZN(_02922_ ) );
INV_X1 _10553_ ( .A(_02867_ ), .ZN(_02923_ ) );
OAI21_X1 _10554_ ( .A(_02922_ ), .B1(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_02923_ ), .ZN(_02924_ ) );
AOI221_X4 _10555_ ( .A(_02919_ ), .B1(\ID_EX_imm [7] ), .B2(_02914_ ), .C1(_02924_ ), .C2(_02916_ ), .ZN(_02925_ ) );
AOI211_X1 _10556_ ( .A(_02626_ ), .B(_02720_ ), .C1(_02917_ ), .C2(_02925_ ), .ZN(_02926_ ) );
AND2_X1 _10557_ ( .A1(_02647_ ), .A2(\ID_EX_imm [8] ), .ZN(_02927_ ) );
AND2_X1 _10558_ ( .A1(_02672_ ), .A2(_02927_ ), .ZN(_02928_ ) );
AOI21_X1 _10559_ ( .A(_02928_ ), .B1(\ID_EX_imm [9] ), .B2(_02670_ ), .ZN(_02929_ ) );
INV_X1 _10560_ ( .A(_02929_ ), .ZN(_02930_ ) );
NAND3_X1 _10561_ ( .A1(_02930_ ), .A2(_02696_ ), .A3(_02719_ ), .ZN(_02931_ ) );
AND2_X1 _10562_ ( .A1(_02718_ ), .A2(\ID_EX_imm [10] ), .ZN(_02932_ ) );
AND2_X1 _10563_ ( .A1(_02696_ ), .A2(_02932_ ), .ZN(_02933_ ) );
AOI21_X1 _10564_ ( .A(_02933_ ), .B1(\ID_EX_imm [11] ), .B2(_02694_ ), .ZN(_02934_ ) );
AND2_X1 _10565_ ( .A1(_02931_ ), .A2(_02934_ ), .ZN(_02935_ ) );
OR2_X1 _10566_ ( .A1(_02935_ ), .A2(_02626_ ), .ZN(_02936_ ) );
NAND2_X1 _10567_ ( .A1(_02553_ ), .A2(\ID_EX_imm [15] ), .ZN(_02937_ ) );
NAND3_X1 _10568_ ( .A1(_02554_ ), .A2(\ID_EX_imm [14] ), .A3(_02575_ ), .ZN(_02938_ ) );
NAND2_X1 _10569_ ( .A1(_02600_ ), .A2(\ID_EX_imm [13] ), .ZN(_02939_ ) );
NAND2_X1 _10570_ ( .A1(_02622_ ), .A2(\ID_EX_imm [12] ), .ZN(_02940_ ) );
OAI21_X1 _10571_ ( .A(_02939_ ), .B1(_02601_ ), .B2(_02940_ ), .ZN(_02941_ ) );
NAND3_X1 _10572_ ( .A1(_02941_ ), .A2(_02554_ ), .A3(_02577_ ), .ZN(_02942_ ) );
NAND4_X1 _10573_ ( .A1(_02936_ ), .A2(_02937_ ), .A3(_02938_ ), .A4(_02942_ ), .ZN(_02943_ ) );
OAI211_X1 _10574_ ( .A(_02432_ ), .B(_02528_ ), .C1(_02926_ ), .C2(_02943_ ), .ZN(_02944_ ) );
NAND3_X1 _10575_ ( .A1(_02478_ ), .A2(\ID_EX_imm [16] ), .A3(_02453_ ), .ZN(_02945_ ) );
INV_X1 _10576_ ( .A(_02476_ ), .ZN(_02946_ ) );
OAI21_X1 _10577_ ( .A(_02945_ ), .B1(_02477_ ), .B2(_02946_ ), .ZN(_02947_ ) );
AND2_X1 _10578_ ( .A1(_02947_ ), .A2(_02527_ ), .ZN(_02948_ ) );
AOI21_X1 _10579_ ( .A(_02525_ ), .B1(_02504_ ), .B2(_02523_ ), .ZN(_02949_ ) );
AND2_X1 _10580_ ( .A1(_02501_ ), .A2(\ID_EX_imm [18] ), .ZN(_02950_ ) );
AND2_X1 _10581_ ( .A1(_02526_ ), .A2(_02950_ ), .ZN(_02951_ ) );
OR3_X1 _10582_ ( .A1(_02948_ ), .A2(_02949_ ), .A3(_02951_ ), .ZN(_02952_ ) );
NAND2_X1 _10583_ ( .A1(_02952_ ), .A2(_02432_ ), .ZN(_02953_ ) );
AND2_X1 _10584_ ( .A1(_02406_ ), .A2(\ID_EX_imm [23] ), .ZN(_02954_ ) );
AND2_X1 _10585_ ( .A1(_02429_ ), .A2(\ID_EX_imm [22] ), .ZN(_02955_ ) );
AOI21_X1 _10586_ ( .A(_02954_ ), .B1(_02408_ ), .B2(_02955_ ), .ZN(_02956_ ) );
NAND2_X1 _10587_ ( .A1(_02358_ ), .A2(\ID_EX_imm [20] ), .ZN(_02957_ ) );
NOR3_X1 _10588_ ( .A1(_02957_ ), .A2(_02382_ ), .A3(_02383_ ), .ZN(_02958_ ) );
OAI211_X1 _10589_ ( .A(_02408_ ), .B(_02431_ ), .C1(_02958_ ), .C2(_02383_ ), .ZN(_02959_ ) );
AND3_X1 _10590_ ( .A1(_02953_ ), .A2(_02956_ ), .A3(_02959_ ), .ZN(_02960_ ) );
AOI211_X1 _10591_ ( .A(_02299_ ), .B(_02323_ ), .C1(_02944_ ), .C2(_02960_ ), .ZN(_02961_ ) );
INV_X1 _10592_ ( .A(_02961_ ), .ZN(_02962_ ) );
AND2_X1 _10593_ ( .A1(_02296_ ), .A2(\ID_EX_imm [24] ), .ZN(_02963_ ) );
AND2_X1 _10594_ ( .A1(_02322_ ), .A2(_02963_ ), .ZN(_02964_ ) );
AOI21_X1 _10595_ ( .A(_02964_ ), .B1(\ID_EX_imm [25] ), .B2(_02320_ ), .ZN(_02965_ ) );
AOI211_X1 _10596_ ( .A(_02250_ ), .B(_02274_ ), .C1(_02962_ ), .C2(_02965_ ), .ZN(_02966_ ) );
INV_X1 _10597_ ( .A(_02966_ ), .ZN(_02967_ ) );
AND2_X1 _10598_ ( .A1(_02271_ ), .A2(\ID_EX_imm [26] ), .ZN(_02968_ ) );
AOI21_X1 _10599_ ( .A(_02248_ ), .B1(_02249_ ), .B2(_02968_ ), .ZN(_02969_ ) );
AOI21_X1 _10600_ ( .A(_02225_ ), .B1(_02967_ ), .B2(_02969_ ), .ZN(_02970_ ) );
OR3_X1 _10601_ ( .A1(_02185_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02196_ ), .ZN(_02971_ ) );
OR2_X1 _10602_ ( .A1(_02136_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02972_ ) );
OAI211_X1 _10603_ ( .A(_02972_ ), .B(_02145_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02973_ ) );
INV_X1 _10604_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02974_ ) );
NAND2_X1 _10605_ ( .A1(_02974_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .ZN(_02975_ ) );
OAI211_X1 _10606_ ( .A(_02975_ ), .B(fanout_net_28 ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02976_ ) );
NAND3_X1 _10607_ ( .A1(_02973_ ), .A2(_02976_ ), .A3(_02167_ ), .ZN(_02977_ ) );
MUX2_X1 _10608_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02978_ ) );
MUX2_X1 _10609_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02979_ ) );
MUX2_X1 _10610_ ( .A(_02978_ ), .B(_02979_ ), .S(_02145_ ), .Z(_02980_ ) );
OAI211_X1 _10611_ ( .A(_02159_ ), .B(_02977_ ), .C1(_02980_ ), .C2(_02167_ ), .ZN(_02981_ ) );
OR2_X1 _10612_ ( .A1(_02136_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02982_ ) );
OAI211_X1 _10613_ ( .A(_02982_ ), .B(fanout_net_28 ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02983_ ) );
OR2_X1 _10614_ ( .A1(_02136_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02984_ ) );
OAI211_X1 _10615_ ( .A(_02984_ ), .B(_02145_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02985_ ) );
NAND3_X1 _10616_ ( .A1(_02983_ ), .A2(_02985_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02986_ ) );
MUX2_X1 _10617_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02987_ ) );
MUX2_X1 _10618_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02988_ ) );
MUX2_X1 _10619_ ( .A(_02987_ ), .B(_02988_ ), .S(fanout_net_28 ), .Z(_02989_ ) );
OAI211_X1 _10620_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02986_ ), .C1(_02989_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02990_ ) );
OAI211_X1 _10621_ ( .A(_02981_ ), .B(_02990_ ), .C1(_02185_ ), .C2(_02196_ ), .ZN(_02991_ ) );
NAND2_X2 _10622_ ( .A1(_02971_ ), .A2(_02991_ ), .ZN(_02992_ ) );
INV_X1 _10623_ ( .A(\ID_EX_imm [29] ), .ZN(_02993_ ) );
XNOR2_X1 _10624_ ( .A(_02992_ ), .B(_02993_ ), .ZN(_02994_ ) );
AND2_X1 _10625_ ( .A1(_02970_ ), .A2(_02994_ ), .ZN(_02995_ ) );
AOI21_X1 _10626_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02201_ ), .B2(_02223_ ), .ZN(_02996_ ) );
NAND2_X1 _10627_ ( .A1(_02994_ ), .A2(_02996_ ), .ZN(_02997_ ) );
INV_X1 _10628_ ( .A(_02992_ ), .ZN(_02998_ ) );
OAI21_X1 _10629_ ( .A(_02997_ ), .B1(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_02998_ ), .ZN(_02999_ ) );
OAI21_X1 _10630_ ( .A(_02200_ ), .B1(_02995_ ), .B2(_02999_ ), .ZN(_03000_ ) );
OR2_X1 _10631_ ( .A1(_02199_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03001_ ) );
AND2_X1 _10632_ ( .A1(_03000_ ), .A2(_03001_ ), .ZN(_03002_ ) );
NAND2_X1 _10633_ ( .A1(_02767_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_03003_ ) );
OR2_X1 _10634_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03004_ ) );
OAI211_X1 _10635_ ( .A(_03004_ ), .B(_02145_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03005_ ) );
INV_X1 _10636_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03006_ ) );
NAND2_X1 _10637_ ( .A1(_03006_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .ZN(_03007_ ) );
OAI211_X1 _10638_ ( .A(_03007_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03008_ ) );
NAND3_X1 _10639_ ( .A1(_03005_ ), .A2(_03008_ ), .A3(_02166_ ), .ZN(_03009_ ) );
MUX2_X1 _10640_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03010_ ) );
MUX2_X1 _10641_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03011_ ) );
MUX2_X1 _10642_ ( .A(_03010_ ), .B(_03011_ ), .S(_02210_ ), .Z(_03012_ ) );
OAI211_X1 _10643_ ( .A(_02159_ ), .B(_03009_ ), .C1(_03012_ ), .C2(_02167_ ), .ZN(_03013_ ) );
OR2_X1 _10644_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03014_ ) );
OAI211_X1 _10645_ ( .A(_03014_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03015_ ) );
OR2_X1 _10646_ ( .A1(_02213_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03016_ ) );
OAI211_X1 _10647_ ( .A(_03016_ ), .B(_02210_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03017_ ) );
NAND3_X1 _10648_ ( .A1(_03015_ ), .A2(_03017_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03018_ ) );
MUX2_X1 _10649_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03019_ ) );
MUX2_X1 _10650_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03020_ ) );
MUX2_X1 _10651_ ( .A(_03019_ ), .B(_03020_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03021_ ) );
OAI211_X1 _10652_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03018_ ), .C1(_03021_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03022_ ) );
NAND2_X1 _10653_ ( .A1(_03013_ ), .A2(_03022_ ), .ZN(_03023_ ) );
OAI21_X1 _10654_ ( .A(_03023_ ), .B1(_02185_ ), .B2(_02196_ ), .ZN(_03024_ ) );
AND2_X2 _10655_ ( .A1(_03003_ ), .A2(_03024_ ), .ZN(_03025_ ) );
XNOR2_X1 _10656_ ( .A(_03025_ ), .B(\ID_EX_imm [31] ), .ZN(_03026_ ) );
XNOR2_X1 _10657_ ( .A(_03002_ ), .B(_03026_ ), .ZN(_03027_ ) );
AND2_X1 _10658_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_03028_ ) );
BUF_X4 _10659_ ( .A(_03028_ ), .Z(_03029_ ) );
BUF_X4 _10660_ ( .A(_03029_ ), .Z(_03030_ ) );
NOR2_X1 _10661_ ( .A1(_03027_ ), .A2(_03030_ ), .ZN(_00097_ ) );
OR3_X1 _10662_ ( .A1(_02995_ ), .A2(_02999_ ), .A3(_02200_ ), .ZN(_03031_ ) );
INV_X1 _10663_ ( .A(_03029_ ), .ZN(_03032_ ) );
BUF_X2 _10664_ ( .A(_03032_ ), .Z(_03033_ ) );
AND3_X1 _10665_ ( .A1(_03031_ ), .A2(_03033_ ), .A3(_03000_ ), .ZN(_00098_ ) );
NOR2_X1 _10666_ ( .A1(_02926_ ), .A2(_02943_ ), .ZN(_03034_ ) );
NAND2_X1 _10667_ ( .A1(_02479_ ), .A2(_02527_ ), .ZN(_03035_ ) );
NOR2_X1 _10668_ ( .A1(_03034_ ), .A2(_03035_ ), .ZN(_03036_ ) );
OAI21_X1 _10669_ ( .A(_02360_ ), .B1(_03036_ ), .B2(_02952_ ), .ZN(_03037_ ) );
NAND2_X1 _10670_ ( .A1(_03037_ ), .A2(_02957_ ), .ZN(_03038_ ) );
XNOR2_X1 _10671_ ( .A(_03038_ ), .B(_02384_ ), .ZN(_03039_ ) );
NOR2_X1 _10672_ ( .A1(_03039_ ), .A2(_03030_ ), .ZN(_00099_ ) );
OR3_X1 _10673_ ( .A1(_03036_ ), .A2(_02360_ ), .A3(_02952_ ), .ZN(_03040_ ) );
AND3_X1 _10674_ ( .A1(_03040_ ), .A2(_03033_ ), .A3(_03037_ ), .ZN(_00100_ ) );
INV_X1 _10675_ ( .A(_02503_ ), .ZN(_03041_ ) );
OAI21_X1 _10676_ ( .A(_02479_ ), .B1(_02926_ ), .B2(_02943_ ), .ZN(_03042_ ) );
INV_X1 _10677_ ( .A(_02947_ ), .ZN(_03043_ ) );
AOI21_X1 _10678_ ( .A(_03041_ ), .B1(_03042_ ), .B2(_03043_ ), .ZN(_03044_ ) );
OR2_X1 _10679_ ( .A1(_03044_ ), .A2(_02950_ ), .ZN(_03045_ ) );
XNOR2_X1 _10680_ ( .A(_03045_ ), .B(_02526_ ), .ZN(_03046_ ) );
NOR2_X1 _10681_ ( .A1(_03046_ ), .A2(_03030_ ), .ZN(_00101_ ) );
AND3_X1 _10682_ ( .A1(_03042_ ), .A2(_03041_ ), .A3(_03043_ ), .ZN(_03047_ ) );
NOR3_X1 _10683_ ( .A1(_03047_ ), .A2(_03044_ ), .A3(_03029_ ), .ZN(_00102_ ) );
OAI21_X1 _10684_ ( .A(_02455_ ), .B1(_02926_ ), .B2(_02943_ ), .ZN(_03048_ ) );
NAND2_X1 _10685_ ( .A1(_02453_ ), .A2(\ID_EX_imm [16] ), .ZN(_03049_ ) );
NAND2_X1 _10686_ ( .A1(_03048_ ), .A2(_03049_ ), .ZN(_03050_ ) );
XNOR2_X1 _10687_ ( .A(_03050_ ), .B(_02478_ ), .ZN(_03051_ ) );
NOR2_X1 _10688_ ( .A1(_03051_ ), .A2(_03030_ ), .ZN(_00103_ ) );
XNOR2_X1 _10689_ ( .A(_03034_ ), .B(_02455_ ), .ZN(_03052_ ) );
AND2_X1 _10690_ ( .A1(_03052_ ), .A2(_03033_ ), .ZN(_00104_ ) );
AOI21_X1 _10691_ ( .A(_02720_ ), .B1(_02917_ ), .B2(_02925_ ), .ZN(_03053_ ) );
INV_X1 _10692_ ( .A(_02935_ ), .ZN(_03054_ ) );
NOR2_X1 _10693_ ( .A1(_03053_ ), .A2(_03054_ ), .ZN(_03055_ ) );
NOR3_X1 _10694_ ( .A1(_03055_ ), .A2(_02601_ ), .A3(_02625_ ), .ZN(_03056_ ) );
OAI21_X1 _10695_ ( .A(_02577_ ), .B1(_03056_ ), .B2(_02941_ ), .ZN(_03057_ ) );
NAND2_X1 _10696_ ( .A1(_02575_ ), .A2(\ID_EX_imm [14] ), .ZN(_03058_ ) );
NAND2_X1 _10697_ ( .A1(_03057_ ), .A2(_03058_ ), .ZN(_03059_ ) );
XNOR2_X1 _10698_ ( .A(_03059_ ), .B(_02554_ ), .ZN(_03060_ ) );
NOR2_X1 _10699_ ( .A1(_03060_ ), .A2(_03030_ ), .ZN(_00105_ ) );
OR3_X1 _10700_ ( .A1(_03056_ ), .A2(_02577_ ), .A3(_02941_ ), .ZN(_03061_ ) );
AND3_X1 _10701_ ( .A1(_03061_ ), .A2(_03033_ ), .A3(_03057_ ), .ZN(_00106_ ) );
OAI21_X1 _10702_ ( .A(_02624_ ), .B1(_03053_ ), .B2(_03054_ ), .ZN(_03062_ ) );
AND2_X1 _10703_ ( .A1(_03062_ ), .A2(_02940_ ), .ZN(_03063_ ) );
XNOR2_X1 _10704_ ( .A(_03063_ ), .B(_02601_ ), .ZN(_03064_ ) );
NOR2_X1 _10705_ ( .A1(_03064_ ), .A2(_03030_ ), .ZN(_00107_ ) );
XNOR2_X1 _10706_ ( .A(_03055_ ), .B(_02624_ ), .ZN(_03065_ ) );
AND2_X1 _10707_ ( .A1(_03065_ ), .A2(_03033_ ), .ZN(_00108_ ) );
OR2_X1 _10708_ ( .A1(_02970_ ), .A2(_02996_ ), .ZN(_03066_ ) );
XNOR2_X1 _10709_ ( .A(_03066_ ), .B(_02994_ ), .ZN(_03067_ ) );
NOR2_X1 _10710_ ( .A1(_03067_ ), .A2(_03030_ ), .ZN(_00109_ ) );
AND3_X1 _10711_ ( .A1(_02967_ ), .A2(_02969_ ), .A3(_02225_ ), .ZN(_03068_ ) );
NOR3_X1 _10712_ ( .A1(_03068_ ), .A2(_02970_ ), .A3(_03029_ ), .ZN(_00110_ ) );
AOI21_X1 _10713_ ( .A(_02274_ ), .B1(_02962_ ), .B2(_02965_ ), .ZN(_03069_ ) );
NOR2_X1 _10714_ ( .A1(_03069_ ), .A2(_02968_ ), .ZN(_03070_ ) );
XNOR2_X1 _10715_ ( .A(_03070_ ), .B(_02250_ ), .ZN(_03071_ ) );
NOR2_X1 _10716_ ( .A1(_03071_ ), .A2(_03030_ ), .ZN(_00111_ ) );
AND3_X1 _10717_ ( .A1(_02962_ ), .A2(_02274_ ), .A3(_02965_ ), .ZN(_03072_ ) );
NOR3_X1 _10718_ ( .A1(_03072_ ), .A2(_03069_ ), .A3(_03029_ ), .ZN(_00112_ ) );
AOI21_X1 _10719_ ( .A(_02299_ ), .B1(_02944_ ), .B2(_02960_ ), .ZN(_03073_ ) );
NOR2_X1 _10720_ ( .A1(_03073_ ), .A2(_02963_ ), .ZN(_03074_ ) );
XNOR2_X1 _10721_ ( .A(_03074_ ), .B(_02323_ ), .ZN(_03075_ ) );
NOR2_X1 _10722_ ( .A1(_03075_ ), .A2(_03030_ ), .ZN(_00113_ ) );
AND3_X1 _10723_ ( .A1(_02944_ ), .A2(_02960_ ), .A3(_02299_ ), .ZN(_03076_ ) );
NOR3_X1 _10724_ ( .A1(_03076_ ), .A2(_03073_ ), .A3(_03029_ ), .ZN(_00114_ ) );
OAI21_X1 _10725_ ( .A(_02385_ ), .B1(_03036_ ), .B2(_02952_ ), .ZN(_03077_ ) );
NOR2_X1 _10726_ ( .A1(_02958_ ), .A2(_02383_ ), .ZN(_03078_ ) );
NAND2_X1 _10727_ ( .A1(_03077_ ), .A2(_03078_ ), .ZN(_03079_ ) );
AND2_X1 _10728_ ( .A1(_03079_ ), .A2(_02431_ ), .ZN(_03080_ ) );
OR2_X1 _10729_ ( .A1(_03080_ ), .A2(_02955_ ), .ZN(_03081_ ) );
XNOR2_X1 _10730_ ( .A(_03081_ ), .B(_02408_ ), .ZN(_03082_ ) );
NOR2_X1 _10731_ ( .A1(_03082_ ), .A2(_03030_ ), .ZN(_00115_ ) );
XNOR2_X1 _10732_ ( .A(_03079_ ), .B(_02431_ ), .ZN(_03083_ ) );
NOR2_X1 _10733_ ( .A1(_03083_ ), .A2(_03029_ ), .ZN(_00116_ ) );
CLKBUF_X2 _10734_ ( .A(_02115_ ), .Z(_03084_ ) );
AND2_X1 _10735_ ( .A1(_03084_ ), .A2(\ID_EX_rd [4] ), .ZN(_00117_ ) );
AND2_X1 _10736_ ( .A1(_03084_ ), .A2(\ID_EX_rd [3] ), .ZN(_00118_ ) );
AND2_X1 _10737_ ( .A1(_03084_ ), .A2(\ID_EX_rd [2] ), .ZN(_00119_ ) );
AND2_X1 _10738_ ( .A1(_03084_ ), .A2(\ID_EX_rd [1] ), .ZN(_00120_ ) );
AND2_X1 _10739_ ( .A1(_03084_ ), .A2(\ID_EX_rd [0] ), .ZN(_00121_ ) );
INV_X2 _10740_ ( .A(_02115_ ), .ZN(_03085_ ) );
BUF_X4 _10741_ ( .A(_03085_ ), .Z(_03086_ ) );
AND2_X1 _10742_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_03087_ ) );
AND2_X1 _10743_ ( .A1(_03087_ ), .A2(\ID_EX_pc [4] ), .ZN(_03088_ ) );
AND2_X1 _10744_ ( .A1(_03088_ ), .A2(\ID_EX_pc [5] ), .ZN(_03089_ ) );
AND2_X1 _10745_ ( .A1(_03089_ ), .A2(\ID_EX_pc [6] ), .ZN(_03090_ ) );
AND2_X1 _10746_ ( .A1(_03090_ ), .A2(\ID_EX_pc [7] ), .ZN(_03091_ ) );
AND2_X1 _10747_ ( .A1(_03091_ ), .A2(\ID_EX_pc [8] ), .ZN(_03092_ ) );
AND2_X2 _10748_ ( .A1(_03092_ ), .A2(\ID_EX_pc [9] ), .ZN(_03093_ ) );
AND3_X1 _10749_ ( .A1(_03093_ ), .A2(\ID_EX_pc [11] ), .A3(\ID_EX_pc [10] ), .ZN(_03094_ ) );
AND3_X1 _10750_ ( .A1(_03094_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_03095_ ) );
AND3_X1 _10751_ ( .A1(_03095_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_03096_ ) );
AND3_X1 _10752_ ( .A1(_03096_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_03097_ ) );
AND3_X1 _10753_ ( .A1(_03097_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_03098_ ) );
AND3_X1 _10754_ ( .A1(_03098_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_03099_ ) );
AND3_X1 _10755_ ( .A1(_03099_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_03100_ ) );
AND3_X1 _10756_ ( .A1(_03100_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_03101_ ) );
AND3_X1 _10757_ ( .A1(_03101_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_03102_ ) );
NAND3_X1 _10758_ ( .A1(_03102_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_03103_ ) );
XNOR2_X1 _10759_ ( .A(_03103_ ), .B(\ID_EX_pc [30] ), .ZN(_03104_ ) );
XOR2_X1 _10760_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_03105_ ) );
AND2_X1 _10761_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_03106_ ) );
NOR2_X1 _10762_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_03107_ ) );
NOR2_X1 _10763_ ( .A1(_03106_ ), .A2(_03107_ ), .ZN(_03108_ ) );
AND2_X1 _10764_ ( .A1(_03105_ ), .A2(_03108_ ), .ZN(_03109_ ) );
XOR2_X1 _10765_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_03110_ ) );
AND2_X1 _10766_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_03111_ ) );
NOR2_X1 _10767_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_03112_ ) );
NOR2_X1 _10768_ ( .A1(_03111_ ), .A2(_03112_ ), .ZN(_03113_ ) );
AND2_X1 _10769_ ( .A1(_03110_ ), .A2(_03113_ ), .ZN(_03114_ ) );
AND2_X1 _10770_ ( .A1(_03109_ ), .A2(_03114_ ), .ZN(_03115_ ) );
XOR2_X1 _10771_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_03116_ ) );
XOR2_X1 _10772_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_03117_ ) );
AND2_X1 _10773_ ( .A1(_03116_ ), .A2(_03117_ ), .ZN(_03118_ ) );
XOR2_X1 _10774_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_03119_ ) );
AND2_X1 _10775_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_03120_ ) );
NOR2_X1 _10776_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_03121_ ) );
NOR2_X1 _10777_ ( .A1(_03120_ ), .A2(_03121_ ), .ZN(_03122_ ) );
AND2_X1 _10778_ ( .A1(_03119_ ), .A2(_03122_ ), .ZN(_03123_ ) );
AND2_X1 _10779_ ( .A1(_03118_ ), .A2(_03123_ ), .ZN(_03124_ ) );
XOR2_X1 _10780_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_03125_ ) );
XOR2_X1 _10781_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_03126_ ) );
AND2_X1 _10782_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_03127_ ) );
AND2_X1 _10783_ ( .A1(_03126_ ), .A2(_03127_ ), .ZN(_03128_ ) );
AND2_X1 _10784_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_03129_ ) );
OAI21_X1 _10785_ ( .A(_03125_ ), .B1(_03128_ ), .B2(_03129_ ), .ZN(_03130_ ) );
INV_X1 _10786_ ( .A(_03130_ ), .ZN(_03131_ ) );
AND2_X1 _10787_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_03132_ ) );
NOR2_X1 _10788_ ( .A1(_03131_ ), .A2(_03132_ ), .ZN(_03133_ ) );
NOR2_X1 _10789_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03134_ ) );
NOR2_X1 _10790_ ( .A1(_03133_ ), .A2(_03134_ ), .ZN(_03135_ ) );
AND2_X1 _10791_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03136_ ) );
NOR2_X1 _10792_ ( .A1(_03135_ ), .A2(_03136_ ), .ZN(_03137_ ) );
AND2_X1 _10793_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03138_ ) );
NOR2_X1 _10794_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03139_ ) );
NOR3_X1 _10795_ ( .A1(_03137_ ), .A2(_03138_ ), .A3(_03139_ ), .ZN(_03140_ ) );
NOR2_X1 _10796_ ( .A1(_03140_ ), .A2(_03138_ ), .ZN(_03141_ ) );
NOR2_X1 _10797_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03142_ ) );
NOR2_X1 _10798_ ( .A1(_03141_ ), .A2(_03142_ ), .ZN(_03143_ ) );
AND2_X1 _10799_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03144_ ) );
NOR2_X1 _10800_ ( .A1(_03143_ ), .A2(_03144_ ), .ZN(_03145_ ) );
AND2_X1 _10801_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03146_ ) );
NOR2_X1 _10802_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03147_ ) );
NOR3_X1 _10803_ ( .A1(_03145_ ), .A2(_03146_ ), .A3(_03147_ ), .ZN(_03148_ ) );
NOR2_X1 _10804_ ( .A1(_03148_ ), .A2(_03146_ ), .ZN(_03149_ ) );
NOR2_X1 _10805_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03150_ ) );
NOR2_X1 _10806_ ( .A1(_03149_ ), .A2(_03150_ ), .ZN(_03151_ ) );
AND2_X1 _10807_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03152_ ) );
NOR2_X1 _10808_ ( .A1(_03151_ ), .A2(_03152_ ), .ZN(_03153_ ) );
XOR2_X1 _10809_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_03154_ ) );
INV_X1 _10810_ ( .A(_03154_ ), .ZN(_03155_ ) );
XNOR2_X1 _10811_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .ZN(_03156_ ) );
NOR2_X1 _10812_ ( .A1(_03155_ ), .A2(_03156_ ), .ZN(_03157_ ) );
XOR2_X1 _10813_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_03158_ ) );
XOR2_X1 _10814_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_03159_ ) );
AND2_X1 _10815_ ( .A1(_03158_ ), .A2(_03159_ ), .ZN(_03160_ ) );
XOR2_X1 _10816_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_03161_ ) );
XOR2_X1 _10817_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_03162_ ) );
AND2_X1 _10818_ ( .A1(_03161_ ), .A2(_03162_ ), .ZN(_03163_ ) );
XOR2_X1 _10819_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_03164_ ) );
XOR2_X1 _10820_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_03165_ ) );
AND2_X1 _10821_ ( .A1(_03164_ ), .A2(_03165_ ), .ZN(_03166_ ) );
NAND4_X1 _10822_ ( .A1(_03157_ ), .A2(_03160_ ), .A3(_03163_ ), .A4(_03166_ ), .ZN(_03167_ ) );
NOR2_X1 _10823_ ( .A1(_03153_ ), .A2(_03167_ ), .ZN(_03168_ ) );
AND3_X1 _10824_ ( .A1(_03158_ ), .A2(\ID_EX_pc [14] ), .A3(\ID_EX_imm [14] ), .ZN(_03169_ ) );
AOI21_X1 _10825_ ( .A(_03169_ ), .B1(\ID_EX_pc [15] ), .B2(\ID_EX_imm [15] ), .ZN(_03170_ ) );
INV_X1 _10826_ ( .A(_03160_ ), .ZN(_03171_ ) );
NAND2_X1 _10827_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_03172_ ) );
NOR2_X1 _10828_ ( .A1(_03156_ ), .A2(_03172_ ), .ZN(_03173_ ) );
AOI21_X1 _10829_ ( .A(_03173_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_03174_ ) );
NAND3_X1 _10830_ ( .A1(_03161_ ), .A2(\ID_EX_pc [10] ), .A3(\ID_EX_imm [10] ), .ZN(_03175_ ) );
INV_X1 _10831_ ( .A(\ID_EX_pc [11] ), .ZN(_03176_ ) );
OAI21_X1 _10832_ ( .A(_03175_ ), .B1(_03176_ ), .B2(_02695_ ), .ZN(_03177_ ) );
AND2_X1 _10833_ ( .A1(\ID_EX_pc [9] ), .A2(\ID_EX_imm [9] ), .ZN(_03178_ ) );
AND2_X1 _10834_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_03179_ ) );
AOI21_X1 _10835_ ( .A(_03178_ ), .B1(_03165_ ), .B2(_03179_ ), .ZN(_03180_ ) );
INV_X1 _10836_ ( .A(_03180_ ), .ZN(_03181_ ) );
AOI21_X1 _10837_ ( .A(_03177_ ), .B1(_03163_ ), .B2(_03181_ ), .ZN(_03182_ ) );
NAND2_X1 _10838_ ( .A1(_03157_ ), .A2(_03160_ ), .ZN(_03183_ ) );
OAI221_X1 _10839_ ( .A(_03170_ ), .B1(_03171_ ), .B2(_03174_ ), .C1(_03182_ ), .C2(_03183_ ), .ZN(_03184_ ) );
OAI211_X1 _10840_ ( .A(_03115_ ), .B(_03124_ ), .C1(_03168_ ), .C2(_03184_ ), .ZN(_03185_ ) );
NAND2_X1 _10841_ ( .A1(_03105_ ), .A2(_03106_ ), .ZN(_03186_ ) );
INV_X1 _10842_ ( .A(\ID_EX_pc [23] ), .ZN(_03187_ ) );
OAI21_X1 _10843_ ( .A(_03186_ ), .B1(_03187_ ), .B2(_02407_ ), .ZN(_03188_ ) );
NAND2_X1 _10844_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_03189_ ) );
NOR3_X1 _10845_ ( .A1(_03111_ ), .A2(_03112_ ), .A3(_03189_ ), .ZN(_03190_ ) );
OR2_X1 _10846_ ( .A1(_03190_ ), .A2(_03111_ ), .ZN(_03191_ ) );
AND2_X1 _10847_ ( .A1(_03119_ ), .A2(_03120_ ), .ZN(_03192_ ) );
AOI21_X1 _10848_ ( .A(_03192_ ), .B1(\ID_EX_pc [19] ), .B2(\ID_EX_imm [19] ), .ZN(_03193_ ) );
AND2_X1 _10849_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_03194_ ) );
AND2_X1 _10850_ ( .A1(_03117_ ), .A2(_03194_ ), .ZN(_03195_ ) );
AOI21_X1 _10851_ ( .A(_03195_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_03196_ ) );
INV_X1 _10852_ ( .A(_03123_ ), .ZN(_03197_ ) );
OAI21_X1 _10853_ ( .A(_03193_ ), .B1(_03196_ ), .B2(_03197_ ), .ZN(_03198_ ) );
AOI221_X4 _10854_ ( .A(_03188_ ), .B1(_03109_ ), .B2(_03191_ ), .C1(_03198_ ), .C2(_03115_ ), .ZN(_03199_ ) );
NAND2_X1 _10855_ ( .A1(_03185_ ), .A2(_03199_ ), .ZN(_03200_ ) );
XOR2_X1 _10856_ ( .A(\ID_EX_pc [25] ), .B(\ID_EX_imm [25] ), .Z(_03201_ ) );
XOR2_X1 _10857_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_03202_ ) );
NAND3_X1 _10858_ ( .A1(_03200_ ), .A2(_03201_ ), .A3(_03202_ ), .ZN(_03203_ ) );
AND2_X1 _10859_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_03204_ ) );
AND2_X1 _10860_ ( .A1(_03201_ ), .A2(_03204_ ), .ZN(_03205_ ) );
AOI21_X1 _10861_ ( .A(_03205_ ), .B1(\ID_EX_pc [25] ), .B2(\ID_EX_imm [25] ), .ZN(_03206_ ) );
NAND2_X1 _10862_ ( .A1(_03203_ ), .A2(_03206_ ), .ZN(_03207_ ) );
XOR2_X1 _10863_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_03208_ ) );
XOR2_X1 _10864_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_03209_ ) );
NAND3_X1 _10865_ ( .A1(_03207_ ), .A2(_03208_ ), .A3(_03209_ ), .ZN(_03210_ ) );
AND3_X1 _10866_ ( .A1(_03208_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_03211_ ) );
AOI21_X1 _10867_ ( .A(_03211_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_03212_ ) );
NAND2_X1 _10868_ ( .A1(_03210_ ), .A2(_03212_ ), .ZN(_03213_ ) );
XOR2_X1 _10869_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_03214_ ) );
NAND2_X1 _10870_ ( .A1(_03213_ ), .A2(_03214_ ), .ZN(_03215_ ) );
NAND2_X1 _10871_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_03216_ ) );
INV_X1 _10872_ ( .A(\ID_EX_pc [29] ), .ZN(_03217_ ) );
AOI22_X1 _10873_ ( .A1(_03215_ ), .A2(_03216_ ), .B1(_03217_ ), .B2(_02993_ ), .ZN(_03218_ ) );
XOR2_X1 _10874_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_03219_ ) );
AND2_X1 _10875_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_03220_ ) );
OR3_X1 _10876_ ( .A1(_03218_ ), .A2(_03219_ ), .A3(_03220_ ), .ZN(_03221_ ) );
OAI21_X1 _10877_ ( .A(_03219_ ), .B1(_03218_ ), .B2(_03220_ ), .ZN(_03222_ ) );
AND2_X1 _10878_ ( .A1(_03221_ ), .A2(_03222_ ), .ZN(_03223_ ) );
NOR2_X1 _10879_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_7 ), .ZN(_03224_ ) );
AND2_X1 _10880_ ( .A1(_03224_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_03225_ ) );
INV_X1 _10881_ ( .A(_03225_ ), .ZN(_03226_ ) );
XNOR2_X1 _10882_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_03227_ ) );
NAND2_X1 _10883_ ( .A1(_02179_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_03228_ ) );
NAND4_X4 _10884_ ( .A1(_02175_ ), .A2(_02178_ ), .A3(_03227_ ), .A4(_03228_ ), .ZN(_03229_ ) );
BUF_X16 _10885_ ( .A(_03229_ ), .Z(_03230_ ) );
BUF_X16 _10886_ ( .A(_03230_ ), .Z(_03231_ ) );
XNOR2_X1 _10887_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_03232_ ) );
INV_X1 _10888_ ( .A(\ID_EX_rs2 [3] ), .ZN(_03233_ ) );
NAND2_X1 _10889_ ( .A1(_03233_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_03234_ ) );
AND3_X1 _10890_ ( .A1(_03232_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y ), .A3(_03234_ ), .ZN(_03235_ ) );
OR2_X1 _10891_ ( .A1(_03233_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_03236_ ) );
OR2_X1 _10892_ ( .A1(_02179_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_03237_ ) );
XNOR2_X1 _10893_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_03238_ ) );
NAND4_X4 _10894_ ( .A1(_03235_ ), .A2(_03236_ ), .A3(_03237_ ), .A4(_03238_ ), .ZN(_03239_ ) );
CLKBUF_X2 _10895_ ( .A(_03239_ ), .Z(_03240_ ) );
BUF_X2 _10896_ ( .A(_03240_ ), .Z(_03241_ ) );
OR3_X1 _10897_ ( .A1(_03231_ ), .A2(\EX_LS_result_reg [19] ), .A3(_03241_ ), .ZN(_03242_ ) );
INV_X1 _10898_ ( .A(fanout_net_42 ), .ZN(_03243_ ) );
BUF_X4 _10899_ ( .A(_03243_ ), .Z(_03244_ ) );
BUF_X4 _10900_ ( .A(_03244_ ), .Z(_03245_ ) );
INV_X1 _10901_ ( .A(fanout_net_31 ), .ZN(_03246_ ) );
BUF_X4 _10902_ ( .A(_03246_ ), .Z(_03247_ ) );
BUF_X4 _10903_ ( .A(_03247_ ), .Z(_03248_ ) );
BUF_X2 _10904_ ( .A(_03248_ ), .Z(_03249_ ) );
OR2_X1 _10905_ ( .A1(_03249_ ), .A2(\myreg.Reg[7][19] ), .ZN(_03250_ ) );
OAI211_X1 _10906_ ( .A(_03250_ ), .B(fanout_net_39 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[6][19] ), .ZN(_03251_ ) );
OR2_X1 _10907_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[4][19] ), .ZN(_03252_ ) );
INV_X2 _10908_ ( .A(fanout_net_39 ), .ZN(_03253_ ) );
BUF_X4 _10909_ ( .A(_03253_ ), .Z(_03254_ ) );
BUF_X4 _10910_ ( .A(_03254_ ), .Z(_03255_ ) );
BUF_X4 _10911_ ( .A(_03255_ ), .Z(_03256_ ) );
BUF_X4 _10912_ ( .A(_03247_ ), .Z(_03257_ ) );
BUF_X4 _10913_ ( .A(_03257_ ), .Z(_03258_ ) );
OAI211_X1 _10914_ ( .A(_03252_ ), .B(_03256_ ), .C1(_03258_ ), .C2(\myreg.Reg[5][19] ), .ZN(_03259_ ) );
NAND3_X1 _10915_ ( .A1(_03251_ ), .A2(fanout_net_41 ), .A3(_03259_ ), .ZN(_03260_ ) );
MUX2_X1 _10916_ ( .A(\myreg.Reg[2][19] ), .B(\myreg.Reg[3][19] ), .S(fanout_net_31 ), .Z(_03261_ ) );
MUX2_X1 _10917_ ( .A(\myreg.Reg[0][19] ), .B(\myreg.Reg[1][19] ), .S(fanout_net_31 ), .Z(_03262_ ) );
MUX2_X1 _10918_ ( .A(_03261_ ), .B(_03262_ ), .S(_03256_ ), .Z(_03263_ ) );
OAI211_X1 _10919_ ( .A(_03245_ ), .B(_03260_ ), .C1(_03263_ ), .C2(fanout_net_41 ), .ZN(_03264_ ) );
INV_X2 _10920_ ( .A(fanout_net_41 ), .ZN(_03265_ ) );
BUF_X4 _10921_ ( .A(_03265_ ), .Z(_03266_ ) );
BUF_X4 _10922_ ( .A(_03266_ ), .Z(_03267_ ) );
NOR2_X1 _10923_ ( .A1(_03258_ ), .A2(\myreg.Reg[11][19] ), .ZN(_03268_ ) );
OAI21_X1 _10924_ ( .A(fanout_net_39 ), .B1(fanout_net_31 ), .B2(\myreg.Reg[10][19] ), .ZN(_03269_ ) );
NOR2_X1 _10925_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][19] ), .ZN(_03270_ ) );
OAI21_X1 _10926_ ( .A(_03256_ ), .B1(_03258_ ), .B2(\myreg.Reg[9][19] ), .ZN(_03271_ ) );
OAI221_X1 _10927_ ( .A(_03267_ ), .B1(_03268_ ), .B2(_03269_ ), .C1(_03270_ ), .C2(_03271_ ), .ZN(_03272_ ) );
MUX2_X1 _10928_ ( .A(\myreg.Reg[12][19] ), .B(\myreg.Reg[13][19] ), .S(fanout_net_31 ), .Z(_03273_ ) );
MUX2_X1 _10929_ ( .A(\myreg.Reg[14][19] ), .B(\myreg.Reg[15][19] ), .S(fanout_net_31 ), .Z(_03274_ ) );
MUX2_X1 _10930_ ( .A(_03273_ ), .B(_03274_ ), .S(fanout_net_39 ), .Z(_03275_ ) );
OAI211_X1 _10931_ ( .A(fanout_net_42 ), .B(_03272_ ), .C1(_03275_ ), .C2(_03267_ ), .ZN(_03276_ ) );
BUF_X4 _10932_ ( .A(_03231_ ), .Z(_03277_ ) );
BUF_X4 _10933_ ( .A(_03241_ ), .Z(_03278_ ) );
OAI211_X1 _10934_ ( .A(_03264_ ), .B(_03276_ ), .C1(_03277_ ), .C2(_03278_ ), .ZN(_03279_ ) );
NAND2_X1 _10935_ ( .A1(_03242_ ), .A2(_03279_ ), .ZN(_03280_ ) );
XOR2_X1 _10936_ ( .A(_02524_ ), .B(_03280_ ), .Z(_03281_ ) );
OR2_X1 _10937_ ( .A1(_03258_ ), .A2(\myreg.Reg[11][18] ), .ZN(_03282_ ) );
OAI211_X1 _10938_ ( .A(_03282_ ), .B(fanout_net_39 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[10][18] ), .ZN(_03283_ ) );
BUF_X4 _10939_ ( .A(_03267_ ), .Z(_03284_ ) );
OR2_X1 _10940_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][18] ), .ZN(_03285_ ) );
BUF_X4 _10941_ ( .A(_03255_ ), .Z(_03286_ ) );
BUF_X4 _10942_ ( .A(_03258_ ), .Z(_03287_ ) );
OAI211_X1 _10943_ ( .A(_03285_ ), .B(_03286_ ), .C1(_03287_ ), .C2(\myreg.Reg[9][18] ), .ZN(_03288_ ) );
NAND3_X1 _10944_ ( .A1(_03283_ ), .A2(_03284_ ), .A3(_03288_ ), .ZN(_03289_ ) );
MUX2_X1 _10945_ ( .A(\myreg.Reg[14][18] ), .B(\myreg.Reg[15][18] ), .S(fanout_net_31 ), .Z(_03290_ ) );
MUX2_X1 _10946_ ( .A(\myreg.Reg[12][18] ), .B(\myreg.Reg[13][18] ), .S(fanout_net_31 ), .Z(_03291_ ) );
MUX2_X1 _10947_ ( .A(_03290_ ), .B(_03291_ ), .S(_03286_ ), .Z(_03292_ ) );
BUF_X4 _10948_ ( .A(_03267_ ), .Z(_03293_ ) );
OAI211_X1 _10949_ ( .A(fanout_net_42 ), .B(_03289_ ), .C1(_03292_ ), .C2(_03293_ ), .ZN(_03294_ ) );
MUX2_X1 _10950_ ( .A(\myreg.Reg[2][18] ), .B(\myreg.Reg[3][18] ), .S(fanout_net_31 ), .Z(_03295_ ) );
AND2_X1 _10951_ ( .A1(_03295_ ), .A2(fanout_net_39 ), .ZN(_03296_ ) );
BUF_X4 _10952_ ( .A(_03256_ ), .Z(_03297_ ) );
BUF_X4 _10953_ ( .A(_03297_ ), .Z(_03298_ ) );
MUX2_X1 _10954_ ( .A(\myreg.Reg[0][18] ), .B(\myreg.Reg[1][18] ), .S(fanout_net_31 ), .Z(_03299_ ) );
AOI211_X1 _10955_ ( .A(fanout_net_41 ), .B(_03296_ ), .C1(_03298_ ), .C2(_03299_ ), .ZN(_03300_ ) );
MUX2_X1 _10956_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_31 ), .Z(_03301_ ) );
MUX2_X1 _10957_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_31 ), .Z(_03302_ ) );
MUX2_X1 _10958_ ( .A(_03301_ ), .B(_03302_ ), .S(_03256_ ), .Z(_03303_ ) );
OAI21_X1 _10959_ ( .A(_03245_ ), .B1(_03303_ ), .B2(_03284_ ), .ZN(_03304_ ) );
BUF_X2 _10960_ ( .A(_03231_ ), .Z(_03305_ ) );
BUF_X2 _10961_ ( .A(_03241_ ), .Z(_03306_ ) );
OAI221_X1 _10962_ ( .A(_03294_ ), .B1(_03300_ ), .B2(_03304_ ), .C1(_03305_ ), .C2(_03306_ ), .ZN(_03307_ ) );
OR3_X1 _10963_ ( .A1(_03277_ ), .A2(\EX_LS_result_reg [18] ), .A3(_03278_ ), .ZN(_03308_ ) );
NAND2_X1 _10964_ ( .A1(_03307_ ), .A2(_03308_ ), .ZN(_03309_ ) );
XOR2_X1 _10965_ ( .A(_03309_ ), .B(_02500_ ), .Z(_03310_ ) );
AND2_X1 _10966_ ( .A1(_03281_ ), .A2(_03310_ ), .ZN(_03311_ ) );
OR2_X1 _10967_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[8][16] ), .ZN(_03312_ ) );
BUF_X4 _10968_ ( .A(_03258_ ), .Z(_03313_ ) );
BUF_X4 _10969_ ( .A(_03313_ ), .Z(_03314_ ) );
OAI211_X1 _10970_ ( .A(_03312_ ), .B(_03297_ ), .C1(_03314_ ), .C2(\myreg.Reg[9][16] ), .ZN(_03315_ ) );
OR2_X1 _10971_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[10][16] ), .ZN(_03316_ ) );
OAI211_X1 _10972_ ( .A(_03316_ ), .B(fanout_net_39 ), .C1(_03314_ ), .C2(\myreg.Reg[11][16] ), .ZN(_03317_ ) );
NAND3_X1 _10973_ ( .A1(_03315_ ), .A2(_03317_ ), .A3(_03284_ ), .ZN(_03318_ ) );
MUX2_X1 _10974_ ( .A(\myreg.Reg[14][16] ), .B(\myreg.Reg[15][16] ), .S(fanout_net_31 ), .Z(_03319_ ) );
MUX2_X1 _10975_ ( .A(\myreg.Reg[12][16] ), .B(\myreg.Reg[13][16] ), .S(fanout_net_31 ), .Z(_03320_ ) );
MUX2_X1 _10976_ ( .A(_03319_ ), .B(_03320_ ), .S(_03297_ ), .Z(_03321_ ) );
OAI211_X1 _10977_ ( .A(fanout_net_42 ), .B(_03318_ ), .C1(_03321_ ), .C2(_03293_ ), .ZN(_03322_ ) );
MUX2_X1 _10978_ ( .A(\myreg.Reg[2][16] ), .B(\myreg.Reg[3][16] ), .S(fanout_net_31 ), .Z(_03323_ ) );
AND2_X1 _10979_ ( .A1(_03323_ ), .A2(fanout_net_39 ), .ZN(_03324_ ) );
MUX2_X1 _10980_ ( .A(\myreg.Reg[0][16] ), .B(\myreg.Reg[1][16] ), .S(fanout_net_31 ), .Z(_03325_ ) );
AOI211_X1 _10981_ ( .A(fanout_net_41 ), .B(_03324_ ), .C1(_03298_ ), .C2(_03325_ ), .ZN(_03326_ ) );
MUX2_X1 _10982_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_31 ), .Z(_03327_ ) );
MUX2_X1 _10983_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_31 ), .Z(_03328_ ) );
MUX2_X1 _10984_ ( .A(_03327_ ), .B(_03328_ ), .S(_03286_ ), .Z(_03329_ ) );
OAI21_X1 _10985_ ( .A(_03245_ ), .B1(_03329_ ), .B2(_03284_ ), .ZN(_03330_ ) );
OAI221_X1 _10986_ ( .A(_03322_ ), .B1(_03326_ ), .B2(_03330_ ), .C1(_03305_ ), .C2(_03306_ ), .ZN(_03331_ ) );
OR3_X1 _10987_ ( .A1(_03277_ ), .A2(\EX_LS_result_reg [16] ), .A3(_03278_ ), .ZN(_03332_ ) );
NAND2_X1 _10988_ ( .A1(_03331_ ), .A2(_03332_ ), .ZN(_03333_ ) );
XOR2_X1 _10989_ ( .A(_03333_ ), .B(_02453_ ), .Z(_03334_ ) );
OR3_X1 _10990_ ( .A1(_03277_ ), .A2(\EX_LS_result_reg [17] ), .A3(_03278_ ), .ZN(_03335_ ) );
BUF_X4 _10991_ ( .A(_03245_ ), .Z(_03336_ ) );
OR2_X1 _10992_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[4][17] ), .ZN(_03337_ ) );
OAI211_X1 _10993_ ( .A(_03337_ ), .B(_03297_ ), .C1(_03287_ ), .C2(\myreg.Reg[5][17] ), .ZN(_03338_ ) );
OR2_X1 _10994_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[6][17] ), .ZN(_03339_ ) );
OAI211_X1 _10995_ ( .A(_03339_ ), .B(fanout_net_39 ), .C1(_03287_ ), .C2(\myreg.Reg[7][17] ), .ZN(_03340_ ) );
NAND3_X1 _10996_ ( .A1(_03338_ ), .A2(_03340_ ), .A3(fanout_net_41 ), .ZN(_03341_ ) );
MUX2_X1 _10997_ ( .A(\myreg.Reg[2][17] ), .B(\myreg.Reg[3][17] ), .S(fanout_net_31 ), .Z(_03342_ ) );
MUX2_X1 _10998_ ( .A(\myreg.Reg[0][17] ), .B(\myreg.Reg[1][17] ), .S(fanout_net_31 ), .Z(_03343_ ) );
MUX2_X1 _10999_ ( .A(_03342_ ), .B(_03343_ ), .S(_03297_ ), .Z(_03344_ ) );
OAI211_X1 _11000_ ( .A(_03336_ ), .B(_03341_ ), .C1(_03344_ ), .C2(fanout_net_41 ), .ZN(_03345_ ) );
NOR2_X1 _11001_ ( .A1(_03287_ ), .A2(\myreg.Reg[11][17] ), .ZN(_03346_ ) );
OAI21_X1 _11002_ ( .A(fanout_net_39 ), .B1(fanout_net_31 ), .B2(\myreg.Reg[10][17] ), .ZN(_03347_ ) );
NOR2_X1 _11003_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][17] ), .ZN(_03348_ ) );
OAI21_X1 _11004_ ( .A(_03297_ ), .B1(_03287_ ), .B2(\myreg.Reg[9][17] ), .ZN(_03349_ ) );
OAI221_X1 _11005_ ( .A(_03284_ ), .B1(_03346_ ), .B2(_03347_ ), .C1(_03348_ ), .C2(_03349_ ), .ZN(_03350_ ) );
MUX2_X1 _11006_ ( .A(\myreg.Reg[12][17] ), .B(\myreg.Reg[13][17] ), .S(fanout_net_32 ), .Z(_03351_ ) );
MUX2_X1 _11007_ ( .A(\myreg.Reg[14][17] ), .B(\myreg.Reg[15][17] ), .S(fanout_net_32 ), .Z(_03352_ ) );
MUX2_X1 _11008_ ( .A(_03351_ ), .B(_03352_ ), .S(fanout_net_39 ), .Z(_03353_ ) );
OAI211_X1 _11009_ ( .A(fanout_net_42 ), .B(_03350_ ), .C1(_03353_ ), .C2(_03293_ ), .ZN(_03354_ ) );
OAI211_X1 _11010_ ( .A(_03345_ ), .B(_03354_ ), .C1(_03305_ ), .C2(_03306_ ), .ZN(_03355_ ) );
NAND2_X1 _11011_ ( .A1(_03335_ ), .A2(_03355_ ), .ZN(_03356_ ) );
AND2_X1 _11012_ ( .A1(_03356_ ), .A2(_02476_ ), .ZN(_03357_ ) );
NOR2_X1 _11013_ ( .A1(_03356_ ), .A2(_02476_ ), .ZN(_03358_ ) );
NOR2_X1 _11014_ ( .A1(_03357_ ), .A2(_03358_ ), .ZN(_03359_ ) );
AND3_X1 _11015_ ( .A1(_03311_ ), .A2(_03334_ ), .A3(_03359_ ), .ZN(_03360_ ) );
OR3_X1 _11016_ ( .A1(_03231_ ), .A2(\EX_LS_result_reg [23] ), .A3(_03241_ ), .ZN(_03361_ ) );
OR2_X1 _11017_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][23] ), .ZN(_03362_ ) );
OAI211_X1 _11018_ ( .A(_03362_ ), .B(_03256_ ), .C1(_03313_ ), .C2(\myreg.Reg[1][23] ), .ZN(_03363_ ) );
OR2_X1 _11019_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][23] ), .ZN(_03364_ ) );
OAI211_X1 _11020_ ( .A(_03364_ ), .B(fanout_net_39 ), .C1(_03313_ ), .C2(\myreg.Reg[3][23] ), .ZN(_03365_ ) );
NAND3_X1 _11021_ ( .A1(_03363_ ), .A2(_03365_ ), .A3(_03267_ ), .ZN(_03366_ ) );
MUX2_X1 _11022_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_32 ), .Z(_03367_ ) );
MUX2_X1 _11023_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_32 ), .Z(_03368_ ) );
MUX2_X1 _11024_ ( .A(_03367_ ), .B(_03368_ ), .S(_03256_ ), .Z(_03369_ ) );
OAI211_X1 _11025_ ( .A(_03245_ ), .B(_03366_ ), .C1(_03369_ ), .C2(_03284_ ), .ZN(_03370_ ) );
OR2_X1 _11026_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[14][23] ), .ZN(_03371_ ) );
OAI211_X1 _11027_ ( .A(_03371_ ), .B(fanout_net_39 ), .C1(_03313_ ), .C2(\myreg.Reg[15][23] ), .ZN(_03372_ ) );
OR2_X1 _11028_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][23] ), .ZN(_03373_ ) );
OAI211_X1 _11029_ ( .A(_03373_ ), .B(_03256_ ), .C1(_03313_ ), .C2(\myreg.Reg[13][23] ), .ZN(_03374_ ) );
NAND3_X1 _11030_ ( .A1(_03372_ ), .A2(_03374_ ), .A3(fanout_net_41 ), .ZN(_03375_ ) );
MUX2_X1 _11031_ ( .A(\myreg.Reg[8][23] ), .B(\myreg.Reg[9][23] ), .S(fanout_net_32 ), .Z(_03376_ ) );
MUX2_X1 _11032_ ( .A(\myreg.Reg[10][23] ), .B(\myreg.Reg[11][23] ), .S(fanout_net_32 ), .Z(_03377_ ) );
MUX2_X1 _11033_ ( .A(_03376_ ), .B(_03377_ ), .S(fanout_net_39 ), .Z(_03378_ ) );
OAI211_X1 _11034_ ( .A(fanout_net_42 ), .B(_03375_ ), .C1(_03378_ ), .C2(fanout_net_41 ), .ZN(_03379_ ) );
OAI211_X1 _11035_ ( .A(_03370_ ), .B(_03379_ ), .C1(_03277_ ), .C2(_03278_ ), .ZN(_03380_ ) );
NAND2_X1 _11036_ ( .A1(_03361_ ), .A2(_03380_ ), .ZN(_03381_ ) );
XOR2_X1 _11037_ ( .A(_02406_ ), .B(_03381_ ), .Z(_03382_ ) );
OR3_X1 _11038_ ( .A1(_03277_ ), .A2(\EX_LS_result_reg [22] ), .A3(_03278_ ), .ZN(_03383_ ) );
OR2_X1 _11039_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[4][22] ), .ZN(_03384_ ) );
OAI211_X1 _11040_ ( .A(_03384_ ), .B(_03297_ ), .C1(_03287_ ), .C2(\myreg.Reg[5][22] ), .ZN(_03385_ ) );
OR2_X1 _11041_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[6][22] ), .ZN(_03386_ ) );
OAI211_X1 _11042_ ( .A(_03386_ ), .B(fanout_net_39 ), .C1(_03287_ ), .C2(\myreg.Reg[7][22] ), .ZN(_03387_ ) );
NAND3_X1 _11043_ ( .A1(_03385_ ), .A2(_03387_ ), .A3(fanout_net_41 ), .ZN(_03388_ ) );
MUX2_X1 _11044_ ( .A(\myreg.Reg[2][22] ), .B(\myreg.Reg[3][22] ), .S(fanout_net_32 ), .Z(_03389_ ) );
MUX2_X1 _11045_ ( .A(\myreg.Reg[0][22] ), .B(\myreg.Reg[1][22] ), .S(fanout_net_32 ), .Z(_03390_ ) );
MUX2_X1 _11046_ ( .A(_03389_ ), .B(_03390_ ), .S(_03286_ ), .Z(_03391_ ) );
OAI211_X1 _11047_ ( .A(_03336_ ), .B(_03388_ ), .C1(_03391_ ), .C2(fanout_net_41 ), .ZN(_03392_ ) );
NOR2_X1 _11048_ ( .A1(_03313_ ), .A2(\myreg.Reg[11][22] ), .ZN(_03393_ ) );
OAI21_X1 _11049_ ( .A(fanout_net_39 ), .B1(fanout_net_32 ), .B2(\myreg.Reg[10][22] ), .ZN(_03394_ ) );
NOR2_X1 _11050_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][22] ), .ZN(_03395_ ) );
OAI21_X1 _11051_ ( .A(_03286_ ), .B1(_03313_ ), .B2(\myreg.Reg[9][22] ), .ZN(_03396_ ) );
OAI221_X1 _11052_ ( .A(_03267_ ), .B1(_03393_ ), .B2(_03394_ ), .C1(_03395_ ), .C2(_03396_ ), .ZN(_03397_ ) );
MUX2_X1 _11053_ ( .A(\myreg.Reg[12][22] ), .B(\myreg.Reg[13][22] ), .S(fanout_net_32 ), .Z(_03398_ ) );
MUX2_X1 _11054_ ( .A(\myreg.Reg[14][22] ), .B(\myreg.Reg[15][22] ), .S(fanout_net_32 ), .Z(_03399_ ) );
MUX2_X1 _11055_ ( .A(_03398_ ), .B(_03399_ ), .S(fanout_net_39 ), .Z(_03400_ ) );
OAI211_X1 _11056_ ( .A(fanout_net_42 ), .B(_03397_ ), .C1(_03400_ ), .C2(_03293_ ), .ZN(_03401_ ) );
OAI211_X1 _11057_ ( .A(_03392_ ), .B(_03401_ ), .C1(_03305_ ), .C2(_03306_ ), .ZN(_03402_ ) );
NAND2_X1 _11058_ ( .A1(_03383_ ), .A2(_03402_ ), .ZN(_03403_ ) );
XOR2_X2 _11059_ ( .A(_03403_ ), .B(_02429_ ), .Z(_03404_ ) );
AND2_X1 _11060_ ( .A1(_03382_ ), .A2(_03404_ ), .ZN(_03405_ ) );
OR3_X1 _11061_ ( .A1(_03277_ ), .A2(\EX_LS_result_reg [20] ), .A3(_03278_ ), .ZN(_03406_ ) );
OR2_X1 _11062_ ( .A1(_03258_ ), .A2(\myreg.Reg[1][20] ), .ZN(_03407_ ) );
OAI211_X1 _11063_ ( .A(_03407_ ), .B(_03297_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[0][20] ), .ZN(_03408_ ) );
OR2_X1 _11064_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][20] ), .ZN(_03409_ ) );
OAI211_X1 _11065_ ( .A(_03409_ ), .B(fanout_net_39 ), .C1(_03287_ ), .C2(\myreg.Reg[3][20] ), .ZN(_03410_ ) );
NAND3_X1 _11066_ ( .A1(_03408_ ), .A2(_03284_ ), .A3(_03410_ ), .ZN(_03411_ ) );
MUX2_X1 _11067_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_32 ), .Z(_03412_ ) );
MUX2_X1 _11068_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_32 ), .Z(_03413_ ) );
MUX2_X1 _11069_ ( .A(_03412_ ), .B(_03413_ ), .S(_03286_ ), .Z(_03414_ ) );
OAI211_X1 _11070_ ( .A(_03336_ ), .B(_03411_ ), .C1(_03414_ ), .C2(_03293_ ), .ZN(_03415_ ) );
OR2_X1 _11071_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[14][20] ), .ZN(_03416_ ) );
OAI211_X1 _11072_ ( .A(_03416_ ), .B(fanout_net_39 ), .C1(_03287_ ), .C2(\myreg.Reg[15][20] ), .ZN(_03417_ ) );
OR2_X1 _11073_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][20] ), .ZN(_03418_ ) );
OAI211_X1 _11074_ ( .A(_03418_ ), .B(_03297_ ), .C1(_03287_ ), .C2(\myreg.Reg[13][20] ), .ZN(_03419_ ) );
NAND3_X1 _11075_ ( .A1(_03417_ ), .A2(_03419_ ), .A3(fanout_net_41 ), .ZN(_03420_ ) );
MUX2_X1 _11076_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_32 ), .Z(_03421_ ) );
MUX2_X1 _11077_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_32 ), .Z(_03422_ ) );
MUX2_X1 _11078_ ( .A(_03421_ ), .B(_03422_ ), .S(fanout_net_39 ), .Z(_03423_ ) );
OAI211_X1 _11079_ ( .A(fanout_net_42 ), .B(_03420_ ), .C1(_03423_ ), .C2(fanout_net_41 ), .ZN(_03424_ ) );
OAI211_X1 _11080_ ( .A(_03415_ ), .B(_03424_ ), .C1(_03305_ ), .C2(_03306_ ), .ZN(_03425_ ) );
NAND2_X1 _11081_ ( .A1(_03406_ ), .A2(_03425_ ), .ZN(_03426_ ) );
XOR2_X1 _11082_ ( .A(_02358_ ), .B(_03426_ ), .Z(_03427_ ) );
OR2_X1 _11083_ ( .A1(_03258_ ), .A2(\myreg.Reg[9][21] ), .ZN(_03428_ ) );
OAI211_X1 _11084_ ( .A(_03428_ ), .B(_03286_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[8][21] ), .ZN(_03429_ ) );
OR2_X1 _11085_ ( .A1(_03258_ ), .A2(\myreg.Reg[11][21] ), .ZN(_03430_ ) );
OAI211_X1 _11086_ ( .A(_03430_ ), .B(fanout_net_39 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[10][21] ), .ZN(_03431_ ) );
NAND3_X1 _11087_ ( .A1(_03429_ ), .A2(_03431_ ), .A3(_03267_ ), .ZN(_03432_ ) );
MUX2_X1 _11088_ ( .A(\myreg.Reg[14][21] ), .B(\myreg.Reg[15][21] ), .S(fanout_net_32 ), .Z(_03433_ ) );
MUX2_X1 _11089_ ( .A(\myreg.Reg[12][21] ), .B(\myreg.Reg[13][21] ), .S(fanout_net_33 ), .Z(_03434_ ) );
MUX2_X1 _11090_ ( .A(_03433_ ), .B(_03434_ ), .S(_03256_ ), .Z(_03435_ ) );
OAI211_X1 _11091_ ( .A(fanout_net_42 ), .B(_03432_ ), .C1(_03435_ ), .C2(_03284_ ), .ZN(_03436_ ) );
MUX2_X1 _11092_ ( .A(\myreg.Reg[2][21] ), .B(\myreg.Reg[3][21] ), .S(fanout_net_33 ), .Z(_03437_ ) );
AND2_X1 _11093_ ( .A1(_03437_ ), .A2(fanout_net_39 ), .ZN(_03438_ ) );
MUX2_X1 _11094_ ( .A(\myreg.Reg[0][21] ), .B(\myreg.Reg[1][21] ), .S(fanout_net_33 ), .Z(_03439_ ) );
AOI211_X1 _11095_ ( .A(fanout_net_41 ), .B(_03438_ ), .C1(_03297_ ), .C2(_03439_ ), .ZN(_03440_ ) );
MUX2_X1 _11096_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_33 ), .Z(_03441_ ) );
MUX2_X1 _11097_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_33 ), .Z(_03442_ ) );
MUX2_X1 _11098_ ( .A(_03441_ ), .B(_03442_ ), .S(_03256_ ), .Z(_03443_ ) );
OAI21_X1 _11099_ ( .A(_03245_ ), .B1(_03443_ ), .B2(_03284_ ), .ZN(_03444_ ) );
OAI221_X1 _11100_ ( .A(_03436_ ), .B1(_03440_ ), .B2(_03444_ ), .C1(_03277_ ), .C2(_03278_ ), .ZN(_03445_ ) );
OR3_X1 _11101_ ( .A1(_03277_ ), .A2(\EX_LS_result_reg [21] ), .A3(_03278_ ), .ZN(_03446_ ) );
NAND2_X1 _11102_ ( .A1(_03445_ ), .A2(_03446_ ), .ZN(_03447_ ) );
NAND2_X1 _11103_ ( .A1(_02361_ ), .A2(_02381_ ), .ZN(_03448_ ) );
AND2_X1 _11104_ ( .A1(_03447_ ), .A2(_03448_ ), .ZN(_03449_ ) );
NOR2_X1 _11105_ ( .A1(_03447_ ), .A2(_03448_ ), .ZN(_03450_ ) );
NOR2_X1 _11106_ ( .A1(_03449_ ), .A2(_03450_ ), .ZN(_03451_ ) );
AND2_X1 _11107_ ( .A1(_03427_ ), .A2(_03451_ ), .ZN(_03452_ ) );
AND2_X4 _11108_ ( .A1(_03405_ ), .A2(_03452_ ), .ZN(_03453_ ) );
AND2_X1 _11109_ ( .A1(_03360_ ), .A2(_03453_ ), .ZN(_03454_ ) );
OR3_X1 _11110_ ( .A1(_03277_ ), .A2(\EX_LS_result_reg [26] ), .A3(_03278_ ), .ZN(_03455_ ) );
NOR2_X1 _11111_ ( .A1(_03313_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03456_ ) );
OAI21_X1 _11112_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03457_ ) );
NOR2_X1 _11113_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03458_ ) );
OAI21_X1 _11114_ ( .A(_03286_ ), .B1(_03313_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03459_ ) );
OAI221_X1 _11115_ ( .A(_03267_ ), .B1(_03456_ ), .B2(_03457_ ), .C1(_03458_ ), .C2(_03459_ ), .ZN(_03460_ ) );
MUX2_X1 _11116_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03461_ ) );
MUX2_X1 _11117_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03462_ ) );
MUX2_X1 _11118_ ( .A(_03461_ ), .B(_03462_ ), .S(fanout_net_39 ), .Z(_03463_ ) );
OAI211_X1 _11119_ ( .A(fanout_net_42 ), .B(_03460_ ), .C1(_03463_ ), .C2(_03284_ ), .ZN(_03464_ ) );
OR2_X1 _11120_ ( .A1(_03258_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03465_ ) );
OAI211_X1 _11121_ ( .A(_03465_ ), .B(fanout_net_39 ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03466_ ) );
OR2_X1 _11122_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03467_ ) );
OAI211_X1 _11123_ ( .A(_03467_ ), .B(_03286_ ), .C1(_03313_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03468_ ) );
NAND3_X1 _11124_ ( .A1(_03466_ ), .A2(fanout_net_41 ), .A3(_03468_ ), .ZN(_03469_ ) );
MUX2_X1 _11125_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03470_ ) );
MUX2_X1 _11126_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03471_ ) );
MUX2_X1 _11127_ ( .A(_03470_ ), .B(_03471_ ), .S(_03286_ ), .Z(_03472_ ) );
OAI211_X1 _11128_ ( .A(_03245_ ), .B(_03469_ ), .C1(_03472_ ), .C2(fanout_net_41 ), .ZN(_03473_ ) );
NAND2_X1 _11129_ ( .A1(_03464_ ), .A2(_03473_ ), .ZN(_03474_ ) );
OAI21_X1 _11130_ ( .A(_03474_ ), .B1(_03305_ ), .B2(_03306_ ), .ZN(_03475_ ) );
AND2_X1 _11131_ ( .A1(_03455_ ), .A2(_03475_ ), .ZN(_03476_ ) );
XNOR2_X1 _11132_ ( .A(_03476_ ), .B(_02271_ ), .ZN(_03477_ ) );
NAND2_X1 _11133_ ( .A1(_02226_ ), .A2(_02246_ ), .ZN(_03478_ ) );
INV_X1 _11134_ ( .A(\EX_LS_result_reg [27] ), .ZN(_03479_ ) );
OR3_X1 _11135_ ( .A1(_03305_ ), .A2(_03479_ ), .A3(_03306_ ), .ZN(_03480_ ) );
OR2_X1 _11136_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03481_ ) );
OAI211_X1 _11137_ ( .A(_03481_ ), .B(_03298_ ), .C1(_03314_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03482_ ) );
OR2_X1 _11138_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03483_ ) );
OAI211_X1 _11139_ ( .A(_03483_ ), .B(fanout_net_39 ), .C1(_03314_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03484_ ) );
NAND3_X1 _11140_ ( .A1(_03482_ ), .A2(_03484_ ), .A3(fanout_net_41 ), .ZN(_03485_ ) );
MUX2_X1 _11141_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03486_ ) );
MUX2_X1 _11142_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03487_ ) );
MUX2_X1 _11143_ ( .A(_03486_ ), .B(_03487_ ), .S(_03298_ ), .Z(_03488_ ) );
OAI211_X1 _11144_ ( .A(_03336_ ), .B(_03485_ ), .C1(_03488_ ), .C2(fanout_net_41 ), .ZN(_03489_ ) );
NOR2_X1 _11145_ ( .A1(_03314_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03490_ ) );
OAI21_X1 _11146_ ( .A(fanout_net_39 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03491_ ) );
NOR2_X1 _11147_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03492_ ) );
OAI21_X1 _11148_ ( .A(_03298_ ), .B1(_03314_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03493_ ) );
OAI221_X1 _11149_ ( .A(_03293_ ), .B1(_03490_ ), .B2(_03491_ ), .C1(_03492_ ), .C2(_03493_ ), .ZN(_03494_ ) );
MUX2_X1 _11150_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03495_ ) );
MUX2_X1 _11151_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03496_ ) );
MUX2_X1 _11152_ ( .A(_03495_ ), .B(_03496_ ), .S(fanout_net_39 ), .Z(_03497_ ) );
OAI211_X1 _11153_ ( .A(fanout_net_42 ), .B(_03494_ ), .C1(_03497_ ), .C2(_03293_ ), .ZN(_03498_ ) );
OAI211_X1 _11154_ ( .A(_03489_ ), .B(_03498_ ), .C1(_03305_ ), .C2(_03306_ ), .ZN(_03499_ ) );
NAND3_X1 _11155_ ( .A1(_03478_ ), .A2(_03480_ ), .A3(_03499_ ), .ZN(_03500_ ) );
NAND2_X1 _11156_ ( .A1(_03480_ ), .A2(_03499_ ), .ZN(_03501_ ) );
NAND3_X1 _11157_ ( .A1(_03501_ ), .A2(_02246_ ), .A3(_02226_ ), .ZN(_03502_ ) );
AND3_X1 _11158_ ( .A1(_03477_ ), .A2(_03500_ ), .A3(_03502_ ), .ZN(_03503_ ) );
NOR2_X1 _11159_ ( .A1(_03229_ ), .A2(_03239_ ), .ZN(_03504_ ) );
NAND2_X1 _11160_ ( .A1(_03504_ ), .A2(\EX_LS_result_reg [24] ), .ZN(_03505_ ) );
OR2_X1 _11161_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03506_ ) );
BUF_X4 _11162_ ( .A(_03298_ ), .Z(_03507_ ) );
BUF_X4 _11163_ ( .A(_03314_ ), .Z(_03508_ ) );
OAI211_X1 _11164_ ( .A(_03506_ ), .B(_03507_ ), .C1(_03508_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03509_ ) );
OR2_X1 _11165_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03510_ ) );
OAI211_X1 _11166_ ( .A(_03510_ ), .B(fanout_net_39 ), .C1(_03508_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03511_ ) );
BUF_X4 _11167_ ( .A(_03293_ ), .Z(_03512_ ) );
NAND3_X1 _11168_ ( .A1(_03509_ ), .A2(_03511_ ), .A3(_03512_ ), .ZN(_03513_ ) );
MUX2_X1 _11169_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03514_ ) );
MUX2_X1 _11170_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03515_ ) );
BUF_X4 _11171_ ( .A(_03298_ ), .Z(_03516_ ) );
MUX2_X1 _11172_ ( .A(_03514_ ), .B(_03515_ ), .S(_03516_ ), .Z(_03517_ ) );
BUF_X4 _11173_ ( .A(_03293_ ), .Z(_03518_ ) );
OAI211_X1 _11174_ ( .A(fanout_net_42 ), .B(_03513_ ), .C1(_03517_ ), .C2(_03518_ ), .ZN(_03519_ ) );
OR2_X1 _11175_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03520_ ) );
OAI211_X1 _11176_ ( .A(_03520_ ), .B(_03507_ ), .C1(_03508_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03521_ ) );
OR2_X1 _11177_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03522_ ) );
OAI211_X1 _11178_ ( .A(_03522_ ), .B(fanout_net_39 ), .C1(_03508_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03523_ ) );
NAND3_X1 _11179_ ( .A1(_03521_ ), .A2(_03523_ ), .A3(_03512_ ), .ZN(_03524_ ) );
MUX2_X1 _11180_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03525_ ) );
MUX2_X1 _11181_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_03526_ ) );
MUX2_X1 _11182_ ( .A(_03525_ ), .B(_03526_ ), .S(_03516_ ), .Z(_03527_ ) );
OAI211_X1 _11183_ ( .A(_03336_ ), .B(_03524_ ), .C1(_03527_ ), .C2(_03518_ ), .ZN(_03528_ ) );
BUF_X2 _11184_ ( .A(_03305_ ), .Z(_03529_ ) );
BUF_X2 _11185_ ( .A(_03306_ ), .Z(_03530_ ) );
OAI211_X1 _11186_ ( .A(_03519_ ), .B(_03528_ ), .C1(_03529_ ), .C2(_03530_ ), .ZN(_03531_ ) );
NAND2_X1 _11187_ ( .A1(_03505_ ), .A2(_03531_ ), .ZN(_03532_ ) );
XNOR2_X1 _11188_ ( .A(_03532_ ), .B(_02296_ ), .ZN(_03533_ ) );
OR2_X1 _11189_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03534_ ) );
BUF_X4 _11190_ ( .A(_03314_ ), .Z(_03535_ ) );
OAI211_X1 _11191_ ( .A(_03534_ ), .B(_03516_ ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03536_ ) );
OR2_X1 _11192_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03537_ ) );
OAI211_X1 _11193_ ( .A(_03537_ ), .B(fanout_net_40 ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03538_ ) );
NAND3_X1 _11194_ ( .A1(_03536_ ), .A2(_03538_ ), .A3(_03293_ ), .ZN(_03539_ ) );
MUX2_X1 _11195_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03540_ ) );
MUX2_X1 _11196_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03541_ ) );
MUX2_X1 _11197_ ( .A(_03540_ ), .B(_03541_ ), .S(_03298_ ), .Z(_03542_ ) );
OAI211_X1 _11198_ ( .A(fanout_net_42 ), .B(_03539_ ), .C1(_03542_ ), .C2(_03512_ ), .ZN(_03543_ ) );
MUX2_X1 _11199_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03544_ ) );
AND2_X1 _11200_ ( .A1(_03544_ ), .A2(_03298_ ), .ZN(_03545_ ) );
MUX2_X1 _11201_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03546_ ) );
AOI211_X1 _11202_ ( .A(fanout_net_41 ), .B(_03545_ ), .C1(fanout_net_40 ), .C2(_03546_ ), .ZN(_03547_ ) );
MUX2_X1 _11203_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03548_ ) );
MUX2_X1 _11204_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03549_ ) );
MUX2_X1 _11205_ ( .A(_03548_ ), .B(_03549_ ), .S(_03298_ ), .Z(_03550_ ) );
OAI21_X1 _11206_ ( .A(_03336_ ), .B1(_03550_ ), .B2(_03512_ ), .ZN(_03551_ ) );
OAI221_X1 _11207_ ( .A(_03543_ ), .B1(_03547_ ), .B2(_03551_ ), .C1(_03529_ ), .C2(_03530_ ), .ZN(_03552_ ) );
INV_X1 _11208_ ( .A(\EX_LS_result_reg [25] ), .ZN(_03553_ ) );
OR3_X1 _11209_ ( .A1(_03305_ ), .A2(_03553_ ), .A3(_03306_ ), .ZN(_03554_ ) );
NAND2_X1 _11210_ ( .A1(_03552_ ), .A2(_03554_ ), .ZN(_03555_ ) );
XNOR2_X1 _11211_ ( .A(_03555_ ), .B(_02320_ ), .ZN(_03556_ ) );
AND2_X1 _11212_ ( .A1(_03533_ ), .A2(_03556_ ), .ZN(_03557_ ) );
AND2_X1 _11213_ ( .A1(_03503_ ), .A2(_03557_ ), .ZN(_03558_ ) );
OR3_X1 _11214_ ( .A1(_03529_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_03530_ ), .ZN(_03559_ ) );
OR2_X1 _11215_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03560_ ) );
OAI211_X1 _11216_ ( .A(_03560_ ), .B(_03507_ ), .C1(_03508_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03561_ ) );
OR2_X1 _11217_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03562_ ) );
OAI211_X1 _11218_ ( .A(_03562_ ), .B(fanout_net_40 ), .C1(_03508_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03563_ ) );
NAND3_X1 _11219_ ( .A1(_03561_ ), .A2(_03563_ ), .A3(_03518_ ), .ZN(_03564_ ) );
MUX2_X1 _11220_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03565_ ) );
MUX2_X1 _11221_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03566_ ) );
MUX2_X1 _11222_ ( .A(_03565_ ), .B(_03566_ ), .S(_03507_ ), .Z(_03567_ ) );
OAI211_X1 _11223_ ( .A(fanout_net_42 ), .B(_03564_ ), .C1(_03567_ ), .C2(_03518_ ), .ZN(_03568_ ) );
OR2_X1 _11224_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03569_ ) );
OAI211_X1 _11225_ ( .A(_03569_ ), .B(_03507_ ), .C1(_03508_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03570_ ) );
OR2_X1 _11226_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03571_ ) );
OAI211_X1 _11227_ ( .A(_03571_ ), .B(fanout_net_40 ), .C1(_03508_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03572_ ) );
NAND3_X1 _11228_ ( .A1(_03570_ ), .A2(_03572_ ), .A3(_03512_ ), .ZN(_03573_ ) );
MUX2_X1 _11229_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03574_ ) );
MUX2_X1 _11230_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03575_ ) );
MUX2_X1 _11231_ ( .A(_03574_ ), .B(_03575_ ), .S(_03507_ ), .Z(_03576_ ) );
OAI211_X1 _11232_ ( .A(_03336_ ), .B(_03573_ ), .C1(_03576_ ), .C2(_03518_ ), .ZN(_03577_ ) );
OAI211_X1 _11233_ ( .A(_03568_ ), .B(_03577_ ), .C1(_03529_ ), .C2(_03530_ ), .ZN(_03578_ ) );
NAND2_X1 _11234_ ( .A1(_03559_ ), .A2(_03578_ ), .ZN(_03579_ ) );
XNOR2_X1 _11235_ ( .A(_03579_ ), .B(_02224_ ), .ZN(_03580_ ) );
OR3_X1 _11236_ ( .A1(_03529_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03530_ ), .ZN(_03581_ ) );
OR2_X1 _11237_ ( .A1(_03314_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03582_ ) );
OAI211_X1 _11238_ ( .A(_03582_ ), .B(fanout_net_40 ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03583_ ) );
OR2_X1 _11239_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03584_ ) );
OAI211_X1 _11240_ ( .A(_03584_ ), .B(_03516_ ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03585_ ) );
NAND3_X1 _11241_ ( .A1(_03583_ ), .A2(_03512_ ), .A3(_03585_ ), .ZN(_03586_ ) );
MUX2_X1 _11242_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03587_ ) );
MUX2_X1 _11243_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03588_ ) );
MUX2_X1 _11244_ ( .A(_03587_ ), .B(_03588_ ), .S(_03516_ ), .Z(_03589_ ) );
OAI211_X1 _11245_ ( .A(fanout_net_42 ), .B(_03586_ ), .C1(_03589_ ), .C2(_03518_ ), .ZN(_03590_ ) );
OR2_X1 _11246_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03591_ ) );
OAI211_X1 _11247_ ( .A(_03591_ ), .B(_03507_ ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03592_ ) );
OR2_X1 _11248_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03593_ ) );
OAI211_X1 _11249_ ( .A(_03593_ ), .B(fanout_net_40 ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03594_ ) );
NAND3_X1 _11250_ ( .A1(_03592_ ), .A2(_03594_ ), .A3(_03512_ ), .ZN(_03595_ ) );
MUX2_X1 _11251_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03596_ ) );
MUX2_X1 _11252_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03597_ ) );
MUX2_X1 _11253_ ( .A(_03596_ ), .B(_03597_ ), .S(_03516_ ), .Z(_03598_ ) );
OAI211_X1 _11254_ ( .A(_03336_ ), .B(_03595_ ), .C1(_03598_ ), .C2(_03518_ ), .ZN(_03599_ ) );
OAI211_X1 _11255_ ( .A(_03590_ ), .B(_03599_ ), .C1(_03529_ ), .C2(_03530_ ), .ZN(_03600_ ) );
NAND2_X1 _11256_ ( .A1(_03581_ ), .A2(_03600_ ), .ZN(_03601_ ) );
XNOR2_X1 _11257_ ( .A(_02992_ ), .B(_03601_ ), .ZN(_03602_ ) );
AND2_X1 _11258_ ( .A1(_03580_ ), .A2(_03602_ ), .ZN(_03603_ ) );
OR3_X1 _11259_ ( .A1(_03529_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03530_ ), .ZN(_03604_ ) );
OR2_X1 _11260_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03605_ ) );
OAI211_X1 _11261_ ( .A(_03605_ ), .B(_03507_ ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03606_ ) );
OR2_X1 _11262_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03607_ ) );
OAI211_X1 _11263_ ( .A(_03607_ ), .B(fanout_net_40 ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03608_ ) );
NAND3_X1 _11264_ ( .A1(_03606_ ), .A2(_03608_ ), .A3(_03512_ ), .ZN(_03609_ ) );
MUX2_X1 _11265_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03610_ ) );
MUX2_X1 _11266_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03611_ ) );
MUX2_X1 _11267_ ( .A(_03610_ ), .B(_03611_ ), .S(_03516_ ), .Z(_03612_ ) );
OAI211_X1 _11268_ ( .A(fanout_net_42 ), .B(_03609_ ), .C1(_03612_ ), .C2(_03518_ ), .ZN(_03613_ ) );
OR2_X1 _11269_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03614_ ) );
OAI211_X1 _11270_ ( .A(_03614_ ), .B(_03516_ ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03615_ ) );
OR2_X1 _11271_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03616_ ) );
OAI211_X1 _11272_ ( .A(_03616_ ), .B(fanout_net_40 ), .C1(_03535_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03617_ ) );
NAND3_X1 _11273_ ( .A1(_03615_ ), .A2(_03617_ ), .A3(_03512_ ), .ZN(_03618_ ) );
MUX2_X1 _11274_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_03619_ ) );
MUX2_X1 _11275_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03620_ ) );
MUX2_X1 _11276_ ( .A(_03619_ ), .B(_03620_ ), .S(_03516_ ), .Z(_03621_ ) );
OAI211_X1 _11277_ ( .A(_03336_ ), .B(_03618_ ), .C1(_03621_ ), .C2(_03518_ ), .ZN(_03622_ ) );
OAI211_X1 _11278_ ( .A(_03613_ ), .B(_03622_ ), .C1(_03529_ ), .C2(_03530_ ), .ZN(_03623_ ) );
NAND2_X1 _11279_ ( .A1(_03604_ ), .A2(_03623_ ), .ZN(_03624_ ) );
XNOR2_X1 _11280_ ( .A(_03025_ ), .B(_03624_ ), .ZN(_03625_ ) );
OR3_X1 _11281_ ( .A1(_03529_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_03530_ ), .ZN(_03626_ ) );
OR2_X1 _11282_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03627_ ) );
OAI211_X1 _11283_ ( .A(_03627_ ), .B(_03507_ ), .C1(_03508_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03628_ ) );
OR2_X1 _11284_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03629_ ) );
OAI211_X1 _11285_ ( .A(_03629_ ), .B(fanout_net_40 ), .C1(_03508_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03630_ ) );
NAND3_X1 _11286_ ( .A1(_03628_ ), .A2(_03630_ ), .A3(_03512_ ), .ZN(_03631_ ) );
MUX2_X1 _11287_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03632_ ) );
MUX2_X1 _11288_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03633_ ) );
MUX2_X1 _11289_ ( .A(_03632_ ), .B(_03633_ ), .S(_03516_ ), .Z(_03634_ ) );
OAI211_X1 _11290_ ( .A(_03336_ ), .B(_03631_ ), .C1(_03634_ ), .C2(_03518_ ), .ZN(_03635_ ) );
OR2_X1 _11291_ ( .A1(_03314_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03636_ ) );
OAI211_X1 _11292_ ( .A(_03636_ ), .B(_03507_ ), .C1(fanout_net_35 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03637_ ) );
OR2_X1 _11293_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03638_ ) );
OAI211_X1 _11294_ ( .A(_03638_ ), .B(fanout_net_40 ), .C1(_03535_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03639_ ) );
NAND3_X1 _11295_ ( .A1(_03637_ ), .A2(fanout_net_41 ), .A3(_03639_ ), .ZN(_03640_ ) );
MUX2_X1 _11296_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03641_ ) );
MUX2_X1 _11297_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03642_ ) );
MUX2_X1 _11298_ ( .A(_03641_ ), .B(_03642_ ), .S(fanout_net_40 ), .Z(_03643_ ) );
OAI211_X1 _11299_ ( .A(fanout_net_42 ), .B(_03640_ ), .C1(_03643_ ), .C2(fanout_net_41 ), .ZN(_03644_ ) );
OAI211_X1 _11300_ ( .A(_03635_ ), .B(_03644_ ), .C1(_03529_ ), .C2(_03530_ ), .ZN(_03645_ ) );
NAND2_X1 _11301_ ( .A1(_03626_ ), .A2(_03645_ ), .ZN(_03646_ ) );
XOR2_X1 _11302_ ( .A(_02199_ ), .B(_03646_ ), .Z(_03647_ ) );
AND3_X1 _11303_ ( .A1(_03603_ ), .A2(_03625_ ), .A3(_03647_ ), .ZN(_03648_ ) );
AND2_X1 _11304_ ( .A1(_03558_ ), .A2(_03648_ ), .ZN(_03649_ ) );
NAND2_X1 _11305_ ( .A1(_03454_ ), .A2(_03649_ ), .ZN(_03650_ ) );
OR3_X1 _11306_ ( .A1(_03229_ ), .A2(\EX_LS_result_reg [7] ), .A3(_03239_ ), .ZN(_03651_ ) );
OR2_X1 _11307_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[4][7] ), .ZN(_03652_ ) );
BUF_X2 _11308_ ( .A(_03246_ ), .Z(_03653_ ) );
OAI211_X1 _11309_ ( .A(_03652_ ), .B(_03254_ ), .C1(_03653_ ), .C2(\myreg.Reg[5][7] ), .ZN(_03654_ ) );
OR2_X1 _11310_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[6][7] ), .ZN(_03655_ ) );
OAI211_X1 _11311_ ( .A(_03655_ ), .B(fanout_net_40 ), .C1(_03653_ ), .C2(\myreg.Reg[7][7] ), .ZN(_03656_ ) );
NAND3_X1 _11312_ ( .A1(_03654_ ), .A2(_03656_ ), .A3(fanout_net_41 ), .ZN(_03657_ ) );
MUX2_X1 _11313_ ( .A(\myreg.Reg[2][7] ), .B(\myreg.Reg[3][7] ), .S(fanout_net_35 ), .Z(_03658_ ) );
MUX2_X1 _11314_ ( .A(\myreg.Reg[0][7] ), .B(\myreg.Reg[1][7] ), .S(fanout_net_35 ), .Z(_03659_ ) );
MUX2_X1 _11315_ ( .A(_03658_ ), .B(_03659_ ), .S(_03253_ ), .Z(_03660_ ) );
OAI211_X1 _11316_ ( .A(_03243_ ), .B(_03657_ ), .C1(_03660_ ), .C2(fanout_net_41 ), .ZN(_03661_ ) );
NOR2_X1 _11317_ ( .A1(_03247_ ), .A2(\myreg.Reg[11][7] ), .ZN(_03662_ ) );
OAI21_X1 _11318_ ( .A(fanout_net_40 ), .B1(fanout_net_35 ), .B2(\myreg.Reg[10][7] ), .ZN(_03663_ ) );
NOR2_X1 _11319_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[8][7] ), .ZN(_03664_ ) );
OAI21_X1 _11320_ ( .A(_03253_ ), .B1(_03247_ ), .B2(\myreg.Reg[9][7] ), .ZN(_03665_ ) );
OAI221_X1 _11321_ ( .A(_03265_ ), .B1(_03662_ ), .B2(_03663_ ), .C1(_03664_ ), .C2(_03665_ ), .ZN(_03666_ ) );
MUX2_X1 _11322_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_35 ), .Z(_03667_ ) );
MUX2_X1 _11323_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_35 ), .Z(_03668_ ) );
MUX2_X1 _11324_ ( .A(_03667_ ), .B(_03668_ ), .S(fanout_net_40 ), .Z(_03669_ ) );
OAI211_X1 _11325_ ( .A(fanout_net_42 ), .B(_03666_ ), .C1(_03669_ ), .C2(_03265_ ), .ZN(_03670_ ) );
OAI211_X1 _11326_ ( .A(_03661_ ), .B(_03670_ ), .C1(_03229_ ), .C2(_03239_ ), .ZN(_03671_ ) );
NAND2_X1 _11327_ ( .A1(_03651_ ), .A2(_03671_ ), .ZN(_03672_ ) );
XOR2_X1 _11328_ ( .A(_02914_ ), .B(_03672_ ), .Z(_03673_ ) );
INV_X1 _11329_ ( .A(_03673_ ), .ZN(_03674_ ) );
OR3_X1 _11330_ ( .A1(_03230_ ), .A2(\EX_LS_result_reg [6] ), .A3(_03240_ ), .ZN(_03675_ ) );
OR2_X1 _11331_ ( .A1(_03248_ ), .A2(\myreg.Reg[3][6] ), .ZN(_03676_ ) );
OAI211_X1 _11332_ ( .A(_03676_ ), .B(fanout_net_40 ), .C1(fanout_net_35 ), .C2(\myreg.Reg[2][6] ), .ZN(_03677_ ) );
OR2_X1 _11333_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][6] ), .ZN(_03678_ ) );
BUF_X4 _11334_ ( .A(_03254_ ), .Z(_03679_ ) );
BUF_X4 _11335_ ( .A(_03248_ ), .Z(_03680_ ) );
OAI211_X1 _11336_ ( .A(_03678_ ), .B(_03679_ ), .C1(_03680_ ), .C2(\myreg.Reg[1][6] ), .ZN(_03681_ ) );
NAND3_X1 _11337_ ( .A1(_03677_ ), .A2(_03266_ ), .A3(_03681_ ), .ZN(_03682_ ) );
MUX2_X1 _11338_ ( .A(\myreg.Reg[6][6] ), .B(\myreg.Reg[7][6] ), .S(fanout_net_35 ), .Z(_03683_ ) );
MUX2_X1 _11339_ ( .A(\myreg.Reg[4][6] ), .B(\myreg.Reg[5][6] ), .S(fanout_net_35 ), .Z(_03684_ ) );
MUX2_X1 _11340_ ( .A(_03683_ ), .B(_03684_ ), .S(_03679_ ), .Z(_03685_ ) );
BUF_X4 _11341_ ( .A(_03265_ ), .Z(_03686_ ) );
BUF_X4 _11342_ ( .A(_03686_ ), .Z(_03687_ ) );
OAI211_X1 _11343_ ( .A(_03244_ ), .B(_03682_ ), .C1(_03685_ ), .C2(_03687_ ), .ZN(_03688_ ) );
OR2_X1 _11344_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[14][6] ), .ZN(_03689_ ) );
BUF_X4 _11345_ ( .A(_03248_ ), .Z(_03690_ ) );
OAI211_X1 _11346_ ( .A(_03689_ ), .B(fanout_net_40 ), .C1(_03690_ ), .C2(\myreg.Reg[15][6] ), .ZN(_03691_ ) );
OR2_X1 _11347_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[12][6] ), .ZN(_03692_ ) );
OAI211_X1 _11348_ ( .A(_03692_ ), .B(_03679_ ), .C1(_03680_ ), .C2(\myreg.Reg[13][6] ), .ZN(_03693_ ) );
NAND3_X1 _11349_ ( .A1(_03691_ ), .A2(_03693_ ), .A3(fanout_net_41 ), .ZN(_03694_ ) );
MUX2_X1 _11350_ ( .A(\myreg.Reg[8][6] ), .B(\myreg.Reg[9][6] ), .S(fanout_net_35 ), .Z(_03695_ ) );
MUX2_X1 _11351_ ( .A(\myreg.Reg[10][6] ), .B(\myreg.Reg[11][6] ), .S(fanout_net_35 ), .Z(_03696_ ) );
MUX2_X1 _11352_ ( .A(_03695_ ), .B(_03696_ ), .S(fanout_net_40 ), .Z(_03697_ ) );
OAI211_X1 _11353_ ( .A(fanout_net_42 ), .B(_03694_ ), .C1(_03697_ ), .C2(fanout_net_41 ), .ZN(_03698_ ) );
BUF_X4 _11354_ ( .A(_03229_ ), .Z(_03699_ ) );
BUF_X2 _11355_ ( .A(_03239_ ), .Z(_03700_ ) );
OAI211_X1 _11356_ ( .A(_03688_ ), .B(_03698_ ), .C1(_03699_ ), .C2(_03700_ ), .ZN(_03701_ ) );
NAND2_X1 _11357_ ( .A1(_03675_ ), .A2(_03701_ ), .ZN(_03702_ ) );
XNOR2_X2 _11358_ ( .A(_02890_ ), .B(_03702_ ), .ZN(_03703_ ) );
NOR2_X1 _11359_ ( .A1(_03674_ ), .A2(_03703_ ), .ZN(_03704_ ) );
OR3_X1 _11360_ ( .A1(_03230_ ), .A2(\EX_LS_result_reg [4] ), .A3(_03240_ ), .ZN(_03705_ ) );
OR2_X1 _11361_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][4] ), .ZN(_03706_ ) );
BUF_X4 _11362_ ( .A(_03254_ ), .Z(_03707_ ) );
OAI211_X1 _11363_ ( .A(_03706_ ), .B(_03707_ ), .C1(_03690_ ), .C2(\myreg.Reg[1][4] ), .ZN(_03708_ ) );
OR2_X1 _11364_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][4] ), .ZN(_03709_ ) );
OAI211_X1 _11365_ ( .A(_03709_ ), .B(fanout_net_40 ), .C1(_03680_ ), .C2(\myreg.Reg[3][4] ), .ZN(_03710_ ) );
NAND3_X1 _11366_ ( .A1(_03708_ ), .A2(_03710_ ), .A3(_03686_ ), .ZN(_03711_ ) );
MUX2_X1 _11367_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_35 ), .Z(_03712_ ) );
MUX2_X1 _11368_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_35 ), .Z(_03713_ ) );
MUX2_X1 _11369_ ( .A(_03712_ ), .B(_03713_ ), .S(_03679_ ), .Z(_03714_ ) );
OAI211_X1 _11370_ ( .A(_03244_ ), .B(_03711_ ), .C1(_03714_ ), .C2(_03687_ ), .ZN(_03715_ ) );
OR2_X1 _11371_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[14][4] ), .ZN(_03716_ ) );
OAI211_X1 _11372_ ( .A(_03716_ ), .B(fanout_net_40 ), .C1(_03680_ ), .C2(\myreg.Reg[15][4] ), .ZN(_03717_ ) );
OR2_X1 _11373_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[12][4] ), .ZN(_03718_ ) );
OAI211_X1 _11374_ ( .A(_03718_ ), .B(_03679_ ), .C1(_03680_ ), .C2(\myreg.Reg[13][4] ), .ZN(_03719_ ) );
NAND3_X1 _11375_ ( .A1(_03717_ ), .A2(_03719_ ), .A3(fanout_net_41 ), .ZN(_03720_ ) );
MUX2_X1 _11376_ ( .A(\myreg.Reg[8][4] ), .B(\myreg.Reg[9][4] ), .S(fanout_net_36 ), .Z(_03721_ ) );
MUX2_X1 _11377_ ( .A(\myreg.Reg[10][4] ), .B(\myreg.Reg[11][4] ), .S(fanout_net_36 ), .Z(_03722_ ) );
MUX2_X1 _11378_ ( .A(_03721_ ), .B(_03722_ ), .S(fanout_net_40 ), .Z(_03723_ ) );
OAI211_X1 _11379_ ( .A(fanout_net_42 ), .B(_03720_ ), .C1(_03723_ ), .C2(fanout_net_41 ), .ZN(_03724_ ) );
OAI211_X1 _11380_ ( .A(_03715_ ), .B(_03724_ ), .C1(_03699_ ), .C2(_03700_ ), .ZN(_03725_ ) );
NAND2_X1 _11381_ ( .A1(_03705_ ), .A2(_03725_ ), .ZN(_03726_ ) );
XOR2_X1 _11382_ ( .A(_02842_ ), .B(_03726_ ), .Z(_03727_ ) );
OR2_X1 _11383_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03728_ ) );
OAI211_X1 _11384_ ( .A(_03728_ ), .B(_03254_ ), .C1(_03653_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03729_ ) );
OR2_X1 _11385_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03730_ ) );
OAI211_X1 _11386_ ( .A(_03730_ ), .B(fanout_net_40 ), .C1(_03653_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03731_ ) );
NAND3_X1 _11387_ ( .A1(_03729_ ), .A2(_03731_ ), .A3(_03265_ ), .ZN(_03732_ ) );
MUX2_X1 _11388_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03733_ ) );
MUX2_X1 _11389_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03734_ ) );
MUX2_X1 _11390_ ( .A(_03733_ ), .B(_03734_ ), .S(_03253_ ), .Z(_03735_ ) );
OAI211_X1 _11391_ ( .A(_03243_ ), .B(_03732_ ), .C1(_03735_ ), .C2(_03265_ ), .ZN(_03736_ ) );
OR2_X1 _11392_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03737_ ) );
OAI211_X1 _11393_ ( .A(_03737_ ), .B(fanout_net_40 ), .C1(_03653_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03738_ ) );
OR2_X1 _11394_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03739_ ) );
OAI211_X1 _11395_ ( .A(_03739_ ), .B(_03253_ ), .C1(_03653_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03740_ ) );
NAND3_X1 _11396_ ( .A1(_03738_ ), .A2(_03740_ ), .A3(fanout_net_41 ), .ZN(_03741_ ) );
MUX2_X1 _11397_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03742_ ) );
MUX2_X1 _11398_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03743_ ) );
MUX2_X1 _11399_ ( .A(_03742_ ), .B(_03743_ ), .S(fanout_net_40 ), .Z(_03744_ ) );
OAI211_X1 _11400_ ( .A(fanout_net_42 ), .B(_03741_ ), .C1(_03744_ ), .C2(fanout_net_41 ), .ZN(_03745_ ) );
AOI21_X1 _11401_ ( .A(_03504_ ), .B1(_03736_ ), .B2(_03745_ ), .ZN(_03746_ ) );
AND2_X1 _11402_ ( .A1(_03504_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_03747_ ) );
NOR2_X2 _11403_ ( .A1(_03746_ ), .A2(_03747_ ), .ZN(_03748_ ) );
XNOR2_X1 _11404_ ( .A(_03748_ ), .B(_02867_ ), .ZN(_03749_ ) );
AND3_X1 _11405_ ( .A1(_03704_ ), .A2(_03727_ ), .A3(_03749_ ), .ZN(_03750_ ) );
OR3_X1 _11406_ ( .A1(_03699_ ), .A2(\EX_LS_result_reg [15] ), .A3(_03700_ ), .ZN(_03751_ ) );
OR2_X1 _11407_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[0][15] ), .ZN(_03752_ ) );
OAI211_X1 _11408_ ( .A(_03752_ ), .B(_03255_ ), .C1(_03249_ ), .C2(\myreg.Reg[1][15] ), .ZN(_03753_ ) );
OR2_X1 _11409_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[2][15] ), .ZN(_03754_ ) );
OAI211_X1 _11410_ ( .A(_03754_ ), .B(fanout_net_40 ), .C1(_03249_ ), .C2(\myreg.Reg[3][15] ), .ZN(_03755_ ) );
NAND3_X1 _11411_ ( .A1(_03753_ ), .A2(_03755_ ), .A3(_03266_ ), .ZN(_03756_ ) );
MUX2_X1 _11412_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_36 ), .Z(_03757_ ) );
MUX2_X1 _11413_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_36 ), .Z(_03758_ ) );
MUX2_X1 _11414_ ( .A(_03757_ ), .B(_03758_ ), .S(_03707_ ), .Z(_03759_ ) );
OAI211_X1 _11415_ ( .A(_03244_ ), .B(_03756_ ), .C1(_03759_ ), .C2(_03687_ ), .ZN(_03760_ ) );
OR2_X1 _11416_ ( .A1(_03248_ ), .A2(\myreg.Reg[13][15] ), .ZN(_03761_ ) );
OAI211_X1 _11417_ ( .A(_03761_ ), .B(_03255_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[12][15] ), .ZN(_03762_ ) );
OR2_X1 _11418_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][15] ), .ZN(_03763_ ) );
OAI211_X1 _11419_ ( .A(_03763_ ), .B(fanout_net_40 ), .C1(_03690_ ), .C2(\myreg.Reg[15][15] ), .ZN(_03764_ ) );
NAND3_X1 _11420_ ( .A1(_03762_ ), .A2(fanout_net_41 ), .A3(_03764_ ), .ZN(_03765_ ) );
MUX2_X1 _11421_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_36 ), .Z(_03766_ ) );
MUX2_X1 _11422_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_36 ), .Z(_03767_ ) );
MUX2_X1 _11423_ ( .A(_03766_ ), .B(_03767_ ), .S(fanout_net_40 ), .Z(_03768_ ) );
OAI211_X1 _11424_ ( .A(fanout_net_42 ), .B(_03765_ ), .C1(_03768_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03769_ ) );
OAI211_X4 _11425_ ( .A(_03760_ ), .B(_03769_ ), .C1(_03231_ ), .C2(_03241_ ), .ZN(_03770_ ) );
NAND2_X1 _11426_ ( .A1(_03751_ ), .A2(_03770_ ), .ZN(_03771_ ) );
XOR2_X1 _11427_ ( .A(_02553_ ), .B(_03771_ ), .Z(_03772_ ) );
OR3_X1 _11428_ ( .A1(_03699_ ), .A2(\EX_LS_result_reg [14] ), .A3(_03700_ ), .ZN(_03773_ ) );
OR2_X1 _11429_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[4][14] ), .ZN(_03774_ ) );
OAI211_X1 _11430_ ( .A(_03774_ ), .B(_03255_ ), .C1(_03249_ ), .C2(\myreg.Reg[5][14] ), .ZN(_03775_ ) );
OR2_X1 _11431_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[6][14] ), .ZN(_03776_ ) );
OAI211_X1 _11432_ ( .A(_03776_ ), .B(fanout_net_40 ), .C1(_03249_ ), .C2(\myreg.Reg[7][14] ), .ZN(_03777_ ) );
NAND3_X1 _11433_ ( .A1(_03775_ ), .A2(_03777_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03778_ ) );
MUX2_X1 _11434_ ( .A(\myreg.Reg[2][14] ), .B(\myreg.Reg[3][14] ), .S(fanout_net_36 ), .Z(_03779_ ) );
MUX2_X1 _11435_ ( .A(\myreg.Reg[0][14] ), .B(\myreg.Reg[1][14] ), .S(fanout_net_36 ), .Z(_03780_ ) );
MUX2_X1 _11436_ ( .A(_03779_ ), .B(_03780_ ), .S(_03707_ ), .Z(_03781_ ) );
OAI211_X1 _11437_ ( .A(_03244_ ), .B(_03778_ ), .C1(_03781_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03782_ ) );
NOR2_X1 _11438_ ( .A1(_03680_ ), .A2(\myreg.Reg[11][14] ), .ZN(_03783_ ) );
OAI21_X1 _11439_ ( .A(fanout_net_40 ), .B1(fanout_net_36 ), .B2(\myreg.Reg[10][14] ), .ZN(_03784_ ) );
NOR2_X1 _11440_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[8][14] ), .ZN(_03785_ ) );
OAI21_X1 _11441_ ( .A(_03707_ ), .B1(_03680_ ), .B2(\myreg.Reg[9][14] ), .ZN(_03786_ ) );
OAI221_X1 _11442_ ( .A(_03266_ ), .B1(_03783_ ), .B2(_03784_ ), .C1(_03785_ ), .C2(_03786_ ), .ZN(_03787_ ) );
MUX2_X1 _11443_ ( .A(\myreg.Reg[12][14] ), .B(\myreg.Reg[13][14] ), .S(fanout_net_36 ), .Z(_03788_ ) );
MUX2_X1 _11444_ ( .A(\myreg.Reg[14][14] ), .B(\myreg.Reg[15][14] ), .S(fanout_net_36 ), .Z(_03789_ ) );
MUX2_X1 _11445_ ( .A(_03788_ ), .B(_03789_ ), .S(fanout_net_40 ), .Z(_03790_ ) );
OAI211_X1 _11446_ ( .A(fanout_net_42 ), .B(_03787_ ), .C1(_03790_ ), .C2(_03687_ ), .ZN(_03791_ ) );
OAI211_X2 _11447_ ( .A(_03782_ ), .B(_03791_ ), .C1(_03231_ ), .C2(_03241_ ), .ZN(_03792_ ) );
NAND2_X1 _11448_ ( .A1(_03773_ ), .A2(_03792_ ), .ZN(_03793_ ) );
XOR2_X1 _11449_ ( .A(_03793_ ), .B(_02575_ ), .Z(_03794_ ) );
AND2_X2 _11450_ ( .A1(_03772_ ), .A2(_03794_ ), .ZN(_03795_ ) );
OR3_X1 _11451_ ( .A1(_03699_ ), .A2(\EX_LS_result_reg [12] ), .A3(_03700_ ), .ZN(_03796_ ) );
OR2_X1 _11452_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[0][12] ), .ZN(_03797_ ) );
OAI211_X1 _11453_ ( .A(_03797_ ), .B(_03255_ ), .C1(_03249_ ), .C2(\myreg.Reg[1][12] ), .ZN(_03798_ ) );
OR2_X1 _11454_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[2][12] ), .ZN(_03799_ ) );
OAI211_X1 _11455_ ( .A(_03799_ ), .B(fanout_net_40 ), .C1(_03249_ ), .C2(\myreg.Reg[3][12] ), .ZN(_03800_ ) );
NAND3_X1 _11456_ ( .A1(_03798_ ), .A2(_03800_ ), .A3(_03687_ ), .ZN(_03801_ ) );
MUX2_X1 _11457_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_36 ), .Z(_03802_ ) );
MUX2_X1 _11458_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_37 ), .Z(_03803_ ) );
MUX2_X1 _11459_ ( .A(_03802_ ), .B(_03803_ ), .S(_03255_ ), .Z(_03804_ ) );
OAI211_X1 _11460_ ( .A(_03245_ ), .B(_03801_ ), .C1(_03804_ ), .C2(_03267_ ), .ZN(_03805_ ) );
OR2_X1 _11461_ ( .A1(_03257_ ), .A2(\myreg.Reg[15][12] ), .ZN(_03806_ ) );
OAI211_X1 _11462_ ( .A(_03806_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][12] ), .ZN(_03807_ ) );
OR2_X1 _11463_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][12] ), .ZN(_03808_ ) );
OAI211_X1 _11464_ ( .A(_03808_ ), .B(_03255_ ), .C1(_03249_ ), .C2(\myreg.Reg[13][12] ), .ZN(_03809_ ) );
NAND3_X1 _11465_ ( .A1(_03807_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03809_ ), .ZN(_03810_ ) );
MUX2_X1 _11466_ ( .A(\myreg.Reg[8][12] ), .B(\myreg.Reg[9][12] ), .S(fanout_net_37 ), .Z(_03811_ ) );
MUX2_X1 _11467_ ( .A(\myreg.Reg[10][12] ), .B(\myreg.Reg[11][12] ), .S(fanout_net_37 ), .Z(_03812_ ) );
MUX2_X1 _11468_ ( .A(_03811_ ), .B(_03812_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03813_ ) );
OAI211_X1 _11469_ ( .A(fanout_net_42 ), .B(_03810_ ), .C1(_03813_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03814_ ) );
OAI211_X1 _11470_ ( .A(_03805_ ), .B(_03814_ ), .C1(_03231_ ), .C2(_03241_ ), .ZN(_03815_ ) );
NAND2_X1 _11471_ ( .A1(_03796_ ), .A2(_03815_ ), .ZN(_03816_ ) );
XOR2_X1 _11472_ ( .A(_02622_ ), .B(_03816_ ), .Z(_03817_ ) );
OR3_X1 _11473_ ( .A1(_03230_ ), .A2(\EX_LS_result_reg [13] ), .A3(_03240_ ), .ZN(_03818_ ) );
OR2_X1 _11474_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][13] ), .ZN(_03819_ ) );
OAI211_X1 _11475_ ( .A(_03819_ ), .B(_03707_ ), .C1(_03690_ ), .C2(\myreg.Reg[1][13] ), .ZN(_03820_ ) );
OR2_X1 _11476_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][13] ), .ZN(_03821_ ) );
OAI211_X1 _11477_ ( .A(_03821_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03690_ ), .C2(\myreg.Reg[3][13] ), .ZN(_03822_ ) );
NAND3_X1 _11478_ ( .A1(_03820_ ), .A2(_03822_ ), .A3(_03266_ ), .ZN(_03823_ ) );
MUX2_X1 _11479_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_37 ), .Z(_03824_ ) );
MUX2_X1 _11480_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_37 ), .Z(_03825_ ) );
MUX2_X1 _11481_ ( .A(_03824_ ), .B(_03825_ ), .S(_03679_ ), .Z(_03826_ ) );
OAI211_X1 _11482_ ( .A(_03244_ ), .B(_03823_ ), .C1(_03826_ ), .C2(_03687_ ), .ZN(_03827_ ) );
OR2_X1 _11483_ ( .A1(_03248_ ), .A2(\myreg.Reg[13][13] ), .ZN(_03828_ ) );
OAI211_X1 _11484_ ( .A(_03828_ ), .B(_03707_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[12][13] ), .ZN(_03829_ ) );
OR2_X1 _11485_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[14][13] ), .ZN(_03830_ ) );
OAI211_X1 _11486_ ( .A(_03830_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03690_ ), .C2(\myreg.Reg[15][13] ), .ZN(_03831_ ) );
NAND3_X1 _11487_ ( .A1(_03829_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03831_ ), .ZN(_03832_ ) );
MUX2_X1 _11488_ ( .A(\myreg.Reg[8][13] ), .B(\myreg.Reg[9][13] ), .S(fanout_net_37 ), .Z(_03833_ ) );
MUX2_X1 _11489_ ( .A(\myreg.Reg[10][13] ), .B(\myreg.Reg[11][13] ), .S(fanout_net_37 ), .Z(_03834_ ) );
MUX2_X1 _11490_ ( .A(_03833_ ), .B(_03834_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03835_ ) );
OAI211_X1 _11491_ ( .A(fanout_net_42 ), .B(_03832_ ), .C1(_03835_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03836_ ) );
OAI211_X1 _11492_ ( .A(_03827_ ), .B(_03836_ ), .C1(_03231_ ), .C2(_03241_ ), .ZN(_03837_ ) );
NAND2_X1 _11493_ ( .A1(_03818_ ), .A2(_03837_ ), .ZN(_03838_ ) );
AND2_X1 _11494_ ( .A1(_02600_ ), .A2(_03838_ ), .ZN(_03839_ ) );
NOR2_X1 _11495_ ( .A1(_02600_ ), .A2(_03838_ ), .ZN(_03840_ ) );
NOR2_X1 _11496_ ( .A1(_03839_ ), .A2(_03840_ ), .ZN(_03841_ ) );
AND3_X4 _11497_ ( .A1(_03795_ ), .A2(_03817_ ), .A3(_03841_ ), .ZN(_03842_ ) );
OR3_X4 _11498_ ( .A1(_03230_ ), .A2(\EX_LS_result_reg [11] ), .A3(_03240_ ), .ZN(_03843_ ) );
OR2_X1 _11499_ ( .A1(_03247_ ), .A2(\myreg.Reg[9][11] ), .ZN(_03844_ ) );
OAI211_X1 _11500_ ( .A(_03844_ ), .B(_03679_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[8][11] ), .ZN(_03845_ ) );
OR2_X1 _11501_ ( .A1(_03247_ ), .A2(\myreg.Reg[11][11] ), .ZN(_03846_ ) );
OAI211_X1 _11502_ ( .A(_03846_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[10][11] ), .ZN(_03847_ ) );
NAND3_X1 _11503_ ( .A1(_03845_ ), .A2(_03847_ ), .A3(_03686_ ), .ZN(_03848_ ) );
MUX2_X1 _11504_ ( .A(\myreg.Reg[14][11] ), .B(\myreg.Reg[15][11] ), .S(fanout_net_37 ), .Z(_03849_ ) );
MUX2_X1 _11505_ ( .A(\myreg.Reg[12][11] ), .B(\myreg.Reg[13][11] ), .S(fanout_net_37 ), .Z(_03850_ ) );
BUF_X4 _11506_ ( .A(_03253_ ), .Z(_03851_ ) );
MUX2_X1 _11507_ ( .A(_03849_ ), .B(_03850_ ), .S(_03851_ ), .Z(_03852_ ) );
OAI211_X1 _11508_ ( .A(fanout_net_42 ), .B(_03848_ ), .C1(_03852_ ), .C2(_03266_ ), .ZN(_03853_ ) );
OAI21_X1 _11509_ ( .A(_03851_ ), .B1(_03248_ ), .B2(\myreg.Reg[1][11] ), .ZN(_03854_ ) );
NOR2_X1 _11510_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][11] ), .ZN(_03855_ ) );
NOR2_X1 _11511_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][11] ), .ZN(_03856_ ) );
OAI21_X1 _11512_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(_03257_ ), .B2(\myreg.Reg[3][11] ), .ZN(_03857_ ) );
OAI221_X1 _11513_ ( .A(_03686_ ), .B1(_03854_ ), .B2(_03855_ ), .C1(_03856_ ), .C2(_03857_ ), .ZN(_03858_ ) );
MUX2_X1 _11514_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_37 ), .Z(_03859_ ) );
MUX2_X1 _11515_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_37 ), .Z(_03860_ ) );
MUX2_X1 _11516_ ( .A(_03859_ ), .B(_03860_ ), .S(_03851_ ), .Z(_03861_ ) );
OAI211_X1 _11517_ ( .A(_03244_ ), .B(_03858_ ), .C1(_03861_ ), .C2(_03266_ ), .ZN(_03862_ ) );
OAI211_X1 _11518_ ( .A(_03853_ ), .B(_03862_ ), .C1(_03699_ ), .C2(_03700_ ), .ZN(_03863_ ) );
NAND2_X1 _11519_ ( .A1(_03843_ ), .A2(_03863_ ), .ZN(_03864_ ) );
XOR2_X1 _11520_ ( .A(_02694_ ), .B(_03864_ ), .Z(_03865_ ) );
OR3_X1 _11521_ ( .A1(_03699_ ), .A2(\EX_LS_result_reg [10] ), .A3(_03700_ ), .ZN(_03866_ ) );
OR2_X1 _11522_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[4][10] ), .ZN(_03867_ ) );
OAI211_X1 _11523_ ( .A(_03867_ ), .B(_03255_ ), .C1(_03249_ ), .C2(\myreg.Reg[5][10] ), .ZN(_03868_ ) );
OR2_X1 _11524_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[6][10] ), .ZN(_03869_ ) );
OAI211_X1 _11525_ ( .A(_03869_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03249_ ), .C2(\myreg.Reg[7][10] ), .ZN(_03870_ ) );
NAND3_X1 _11526_ ( .A1(_03868_ ), .A2(_03870_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03871_ ) );
MUX2_X1 _11527_ ( .A(\myreg.Reg[2][10] ), .B(\myreg.Reg[3][10] ), .S(fanout_net_37 ), .Z(_03872_ ) );
MUX2_X1 _11528_ ( .A(\myreg.Reg[0][10] ), .B(\myreg.Reg[1][10] ), .S(fanout_net_37 ), .Z(_03873_ ) );
MUX2_X1 _11529_ ( .A(_03872_ ), .B(_03873_ ), .S(_03255_ ), .Z(_03874_ ) );
OAI211_X1 _11530_ ( .A(_03245_ ), .B(_03871_ ), .C1(_03874_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03875_ ) );
NOR2_X1 _11531_ ( .A1(_03690_ ), .A2(\myreg.Reg[11][10] ), .ZN(_03876_ ) );
OAI21_X1 _11532_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_37 ), .B2(\myreg.Reg[10][10] ), .ZN(_03877_ ) );
NOR2_X1 _11533_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][10] ), .ZN(_03878_ ) );
OAI21_X1 _11534_ ( .A(_03707_ ), .B1(_03690_ ), .B2(\myreg.Reg[9][10] ), .ZN(_03879_ ) );
OAI221_X1 _11535_ ( .A(_03266_ ), .B1(_03876_ ), .B2(_03877_ ), .C1(_03878_ ), .C2(_03879_ ), .ZN(_03880_ ) );
MUX2_X1 _11536_ ( .A(\myreg.Reg[12][10] ), .B(\myreg.Reg[13][10] ), .S(fanout_net_37 ), .Z(_03881_ ) );
MUX2_X1 _11537_ ( .A(\myreg.Reg[14][10] ), .B(\myreg.Reg[15][10] ), .S(fanout_net_37 ), .Z(_03882_ ) );
MUX2_X1 _11538_ ( .A(_03881_ ), .B(_03882_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03883_ ) );
OAI211_X1 _11539_ ( .A(fanout_net_42 ), .B(_03880_ ), .C1(_03883_ ), .C2(_03267_ ), .ZN(_03884_ ) );
OAI211_X1 _11540_ ( .A(_03875_ ), .B(_03884_ ), .C1(_03231_ ), .C2(_03241_ ), .ZN(_03885_ ) );
NAND2_X1 _11541_ ( .A1(_03866_ ), .A2(_03885_ ), .ZN(_03886_ ) );
XOR2_X1 _11542_ ( .A(_03886_ ), .B(_02717_ ), .Z(_03887_ ) );
AND2_X1 _11543_ ( .A1(_03865_ ), .A2(_03887_ ), .ZN(_03888_ ) );
OR3_X1 _11544_ ( .A1(_03229_ ), .A2(\EX_LS_result_reg [9] ), .A3(_03239_ ), .ZN(_03889_ ) );
OR2_X1 _11545_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][9] ), .ZN(_03890_ ) );
OAI211_X1 _11546_ ( .A(_03890_ ), .B(_03254_ ), .C1(_03248_ ), .C2(\myreg.Reg[9][9] ), .ZN(_03891_ ) );
OR2_X1 _11547_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[10][9] ), .ZN(_03892_ ) );
OAI211_X1 _11548_ ( .A(_03892_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03248_ ), .C2(\myreg.Reg[11][9] ), .ZN(_03893_ ) );
NAND3_X1 _11549_ ( .A1(_03891_ ), .A2(_03893_ ), .A3(_03265_ ), .ZN(_03894_ ) );
MUX2_X1 _11550_ ( .A(\myreg.Reg[14][9] ), .B(\myreg.Reg[15][9] ), .S(fanout_net_38 ), .Z(_03895_ ) );
MUX2_X1 _11551_ ( .A(\myreg.Reg[12][9] ), .B(\myreg.Reg[13][9] ), .S(fanout_net_38 ), .Z(_03896_ ) );
MUX2_X1 _11552_ ( .A(_03895_ ), .B(_03896_ ), .S(_03254_ ), .Z(_03897_ ) );
OAI211_X1 _11553_ ( .A(fanout_net_42 ), .B(_03894_ ), .C1(_03897_ ), .C2(_03686_ ), .ZN(_03898_ ) );
NOR2_X1 _11554_ ( .A1(_03247_ ), .A2(\myreg.Reg[3][9] ), .ZN(_03899_ ) );
OAI21_X1 _11555_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_38 ), .B2(\myreg.Reg[2][9] ), .ZN(_03900_ ) );
NOR2_X1 _11556_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][9] ), .ZN(_03901_ ) );
OAI21_X1 _11557_ ( .A(_03253_ ), .B1(_03653_ ), .B2(\myreg.Reg[1][9] ), .ZN(_03902_ ) );
OAI221_X1 _11558_ ( .A(_03265_ ), .B1(_03899_ ), .B2(_03900_ ), .C1(_03901_ ), .C2(_03902_ ), .ZN(_03903_ ) );
MUX2_X1 _11559_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_38 ), .Z(_03904_ ) );
MUX2_X1 _11560_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_38 ), .Z(_03905_ ) );
MUX2_X1 _11561_ ( .A(_03904_ ), .B(_03905_ ), .S(_03254_ ), .Z(_03906_ ) );
OAI211_X1 _11562_ ( .A(_03243_ ), .B(_03903_ ), .C1(_03906_ ), .C2(_03686_ ), .ZN(_03907_ ) );
OAI211_X1 _11563_ ( .A(_03898_ ), .B(_03907_ ), .C1(_03230_ ), .C2(_03240_ ), .ZN(_03908_ ) );
NAND2_X1 _11564_ ( .A1(_03889_ ), .A2(_03908_ ), .ZN(_03909_ ) );
XOR2_X1 _11565_ ( .A(_02670_ ), .B(_03909_ ), .Z(_03910_ ) );
OR3_X1 _11566_ ( .A1(_03229_ ), .A2(\EX_LS_result_reg [8] ), .A3(_03239_ ), .ZN(_03911_ ) );
OR2_X1 _11567_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][8] ), .ZN(_03912_ ) );
OAI211_X1 _11568_ ( .A(_03912_ ), .B(_03851_ ), .C1(_03257_ ), .C2(\myreg.Reg[1][8] ), .ZN(_03913_ ) );
OR2_X1 _11569_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[2][8] ), .ZN(_03914_ ) );
OAI211_X1 _11570_ ( .A(_03914_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03257_ ), .C2(\myreg.Reg[3][8] ), .ZN(_03915_ ) );
NAND3_X1 _11571_ ( .A1(_03913_ ), .A2(_03915_ ), .A3(_03265_ ), .ZN(_03916_ ) );
MUX2_X1 _11572_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_38 ), .Z(_03917_ ) );
MUX2_X1 _11573_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_38 ), .Z(_03918_ ) );
MUX2_X1 _11574_ ( .A(_03917_ ), .B(_03918_ ), .S(_03851_ ), .Z(_03919_ ) );
OAI211_X1 _11575_ ( .A(_03244_ ), .B(_03916_ ), .C1(_03919_ ), .C2(_03266_ ), .ZN(_03920_ ) );
OR2_X1 _11576_ ( .A1(_03247_ ), .A2(\myreg.Reg[15][8] ), .ZN(_03921_ ) );
OAI211_X1 _11577_ ( .A(_03921_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myreg.Reg[14][8] ), .ZN(_03922_ ) );
OR2_X1 _11578_ ( .A1(_03247_ ), .A2(\myreg.Reg[13][8] ), .ZN(_03923_ ) );
OAI211_X1 _11579_ ( .A(_03923_ ), .B(_03851_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[12][8] ), .ZN(_03924_ ) );
NAND3_X1 _11580_ ( .A1(_03922_ ), .A2(_03924_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03925_ ) );
MUX2_X1 _11581_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_38 ), .Z(_03926_ ) );
MUX2_X1 _11582_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_38 ), .Z(_03927_ ) );
MUX2_X1 _11583_ ( .A(_03926_ ), .B(_03927_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03928_ ) );
OAI211_X1 _11584_ ( .A(fanout_net_42 ), .B(_03925_ ), .C1(_03928_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03929_ ) );
OAI211_X1 _11585_ ( .A(_03920_ ), .B(_03929_ ), .C1(_03230_ ), .C2(_03240_ ), .ZN(_03930_ ) );
NAND2_X1 _11586_ ( .A1(_03911_ ), .A2(_03930_ ), .ZN(_03931_ ) );
XOR2_X1 _11587_ ( .A(_02647_ ), .B(_03931_ ), .Z(_03932_ ) );
AND3_X1 _11588_ ( .A1(_03888_ ), .A2(_03910_ ), .A3(_03932_ ), .ZN(_03933_ ) );
NAND3_X1 _11589_ ( .A1(_03750_ ), .A2(_03842_ ), .A3(_03933_ ), .ZN(_03934_ ) );
NOR2_X1 _11590_ ( .A1(_03650_ ), .A2(_03934_ ), .ZN(_03935_ ) );
OR3_X1 _11591_ ( .A1(_03699_ ), .A2(\EX_LS_result_reg [2] ), .A3(_03700_ ), .ZN(_03936_ ) );
OR2_X1 _11592_ ( .A1(_03248_ ), .A2(\myreg.Reg[7][2] ), .ZN(_03937_ ) );
OAI211_X1 _11593_ ( .A(_03937_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myreg.Reg[6][2] ), .ZN(_03938_ ) );
OR2_X1 _11594_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[4][2] ), .ZN(_03939_ ) );
OAI211_X1 _11595_ ( .A(_03939_ ), .B(_03707_ ), .C1(_03690_ ), .C2(\myreg.Reg[5][2] ), .ZN(_03940_ ) );
NAND3_X1 _11596_ ( .A1(_03938_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03940_ ), .ZN(_03941_ ) );
MUX2_X1 _11597_ ( .A(\myreg.Reg[2][2] ), .B(\myreg.Reg[3][2] ), .S(fanout_net_38 ), .Z(_03942_ ) );
MUX2_X1 _11598_ ( .A(\myreg.Reg[0][2] ), .B(\myreg.Reg[1][2] ), .S(fanout_net_38 ), .Z(_03943_ ) );
MUX2_X1 _11599_ ( .A(_03942_ ), .B(_03943_ ), .S(_03707_ ), .Z(_03944_ ) );
OAI211_X1 _11600_ ( .A(_03245_ ), .B(_03941_ ), .C1(_03944_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03945_ ) );
NOR2_X1 _11601_ ( .A1(_03680_ ), .A2(\myreg.Reg[11][2] ), .ZN(_03946_ ) );
OAI21_X1 _11602_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_38 ), .B2(\myreg.Reg[10][2] ), .ZN(_03947_ ) );
NOR2_X1 _11603_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[8][2] ), .ZN(_03948_ ) );
OAI21_X1 _11604_ ( .A(_03707_ ), .B1(_03690_ ), .B2(\myreg.Reg[9][2] ), .ZN(_03949_ ) );
OAI221_X1 _11605_ ( .A(_03266_ ), .B1(_03946_ ), .B2(_03947_ ), .C1(_03948_ ), .C2(_03949_ ), .ZN(_03950_ ) );
MUX2_X1 _11606_ ( .A(\myreg.Reg[12][2] ), .B(\myreg.Reg[13][2] ), .S(fanout_net_38 ), .Z(_03951_ ) );
MUX2_X1 _11607_ ( .A(\myreg.Reg[14][2] ), .B(\myreg.Reg[15][2] ), .S(fanout_net_38 ), .Z(_03952_ ) );
MUX2_X1 _11608_ ( .A(_03951_ ), .B(_03952_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03953_ ) );
OAI211_X1 _11609_ ( .A(fanout_net_42 ), .B(_03950_ ), .C1(_03953_ ), .C2(_03687_ ), .ZN(_03954_ ) );
OAI211_X1 _11610_ ( .A(_03945_ ), .B(_03954_ ), .C1(_03231_ ), .C2(_03241_ ), .ZN(_03955_ ) );
NAND2_X1 _11611_ ( .A1(_03936_ ), .A2(_03955_ ), .ZN(_03956_ ) );
XOR2_X2 _11612_ ( .A(_03956_ ), .B(_02741_ ), .Z(_03957_ ) );
OR3_X1 _11613_ ( .A1(_03230_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03240_ ), .ZN(_03958_ ) );
OR2_X1 _11614_ ( .A1(fanout_net_38 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03959_ ) );
OAI211_X1 _11615_ ( .A(_03959_ ), .B(_03679_ ), .C1(_03680_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03960_ ) );
OR2_X1 _11616_ ( .A1(fanout_net_38 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03961_ ) );
OAI211_X1 _11617_ ( .A(_03961_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03257_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03962_ ) );
NAND3_X1 _11618_ ( .A1(_03960_ ), .A2(_03962_ ), .A3(_03686_ ), .ZN(_03963_ ) );
MUX2_X1 _11619_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_38 ), .Z(_03964_ ) );
MUX2_X1 _11620_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_38 ), .Z(_03965_ ) );
MUX2_X1 _11621_ ( .A(_03964_ ), .B(_03965_ ), .S(_03851_ ), .Z(_03966_ ) );
OAI211_X1 _11622_ ( .A(_03244_ ), .B(_03963_ ), .C1(_03966_ ), .C2(_03687_ ), .ZN(_03967_ ) );
OR2_X1 _11623_ ( .A1(fanout_net_38 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03968_ ) );
OAI211_X1 _11624_ ( .A(_03968_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03680_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03969_ ) );
OR2_X1 _11625_ ( .A1(fanout_net_38 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03970_ ) );
OAI211_X1 _11626_ ( .A(_03970_ ), .B(_03679_ ), .C1(_03257_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03971_ ) );
NAND3_X1 _11627_ ( .A1(_03969_ ), .A2(_03971_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03972_ ) );
MUX2_X1 _11628_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_38 ), .Z(_03973_ ) );
MUX2_X1 _11629_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03974_ ) );
MUX2_X1 _11630_ ( .A(_03973_ ), .B(_03974_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03975_ ) );
OAI211_X1 _11631_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03972_ ), .C1(_03975_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03976_ ) );
OAI211_X1 _11632_ ( .A(_03967_ ), .B(_03976_ ), .C1(_03699_ ), .C2(_03700_ ), .ZN(_03977_ ) );
NAND2_X1 _11633_ ( .A1(_03958_ ), .A2(_03977_ ), .ZN(_03978_ ) );
XNOR2_X1 _11634_ ( .A(_02815_ ), .B(_03978_ ), .ZN(_03979_ ) );
AND2_X1 _11635_ ( .A1(_03957_ ), .A2(_03979_ ), .ZN(_03980_ ) );
OR3_X1 _11636_ ( .A1(_03229_ ), .A2(\EX_LS_result_reg [1] ), .A3(_03239_ ), .ZN(_03981_ ) );
OR2_X1 _11637_ ( .A1(_03247_ ), .A2(\myreg.Reg[3][1] ), .ZN(_03982_ ) );
OAI211_X1 _11638_ ( .A(_03982_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[2][1] ), .ZN(_03983_ ) );
OR2_X1 _11639_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[0][1] ), .ZN(_03984_ ) );
OAI211_X1 _11640_ ( .A(_03984_ ), .B(_03254_ ), .C1(_03653_ ), .C2(\myreg.Reg[1][1] ), .ZN(_03985_ ) );
NAND3_X1 _11641_ ( .A1(_03983_ ), .A2(_03265_ ), .A3(_03985_ ), .ZN(_03986_ ) );
MUX2_X1 _11642_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03987_ ) );
MUX2_X1 _11643_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03988_ ) );
MUX2_X1 _11644_ ( .A(_03987_ ), .B(_03988_ ), .S(_03253_ ), .Z(_03989_ ) );
OAI211_X1 _11645_ ( .A(_03243_ ), .B(_03986_ ), .C1(_03989_ ), .C2(_03686_ ), .ZN(_03990_ ) );
OR2_X1 _11646_ ( .A1(_03246_ ), .A2(\myreg.Reg[13][1] ), .ZN(_03991_ ) );
OAI211_X1 _11647_ ( .A(_03991_ ), .B(_03254_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[12][1] ), .ZN(_03992_ ) );
OR2_X1 _11648_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[14][1] ), .ZN(_03993_ ) );
OAI211_X1 _11649_ ( .A(_03993_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03653_ ), .C2(\myreg.Reg[15][1] ), .ZN(_03994_ ) );
NAND3_X1 _11650_ ( .A1(_03992_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03994_ ), .ZN(_03995_ ) );
MUX2_X1 _11651_ ( .A(\myreg.Reg[8][1] ), .B(\myreg.Reg[9][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03996_ ) );
MUX2_X1 _11652_ ( .A(\myreg.Reg[10][1] ), .B(\myreg.Reg[11][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03997_ ) );
MUX2_X1 _11653_ ( .A(_03996_ ), .B(_03997_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03998_ ) );
OAI211_X1 _11654_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03995_ ), .C1(_03998_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03999_ ) );
OAI211_X1 _11655_ ( .A(_03990_ ), .B(_03999_ ), .C1(_03230_ ), .C2(_03240_ ), .ZN(_04000_ ) );
NAND2_X2 _11656_ ( .A1(_03981_ ), .A2(_04000_ ), .ZN(_04001_ ) );
XOR2_X1 _11657_ ( .A(_02764_ ), .B(_04001_ ), .Z(_04002_ ) );
INV_X1 _11658_ ( .A(_04002_ ), .ZN(_04003_ ) );
AND2_X2 _11659_ ( .A1(_02768_ ), .A2(_02788_ ), .ZN(_04004_ ) );
OR3_X1 _11660_ ( .A1(_03230_ ), .A2(\EX_LS_result_reg [0] ), .A3(_03240_ ), .ZN(_04005_ ) );
OR2_X1 _11661_ ( .A1(_03653_ ), .A2(\myreg.Reg[9][0] ), .ZN(_04006_ ) );
OAI211_X1 _11662_ ( .A(_04006_ ), .B(_03679_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[8][0] ), .ZN(_04007_ ) );
OR2_X1 _11663_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[10][0] ), .ZN(_04008_ ) );
OAI211_X1 _11664_ ( .A(_04008_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03257_ ), .C2(\myreg.Reg[11][0] ), .ZN(_04009_ ) );
NAND3_X1 _11665_ ( .A1(_04007_ ), .A2(_03686_ ), .A3(_04009_ ), .ZN(_04010_ ) );
MUX2_X1 _11666_ ( .A(\myreg.Reg[14][0] ), .B(\myreg.Reg[15][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04011_ ) );
MUX2_X1 _11667_ ( .A(\myreg.Reg[12][0] ), .B(\myreg.Reg[13][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04012_ ) );
MUX2_X1 _11668_ ( .A(_04011_ ), .B(_04012_ ), .S(_03851_ ), .Z(_04013_ ) );
OAI211_X1 _11669_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04010_ ), .C1(_04013_ ), .C2(_03687_ ), .ZN(_04014_ ) );
OAI21_X1 _11670_ ( .A(_03851_ ), .B1(_03257_ ), .B2(\myreg.Reg[1][0] ), .ZN(_04015_ ) );
NOR2_X1 _11671_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[0][0] ), .ZN(_04016_ ) );
NOR2_X1 _11672_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[2][0] ), .ZN(_04017_ ) );
OAI21_X1 _11673_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(_03257_ ), .B2(\myreg.Reg[3][0] ), .ZN(_04018_ ) );
OAI221_X1 _11674_ ( .A(_03686_ ), .B1(_04015_ ), .B2(_04016_ ), .C1(_04017_ ), .C2(_04018_ ), .ZN(_04019_ ) );
MUX2_X1 _11675_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04020_ ) );
MUX2_X1 _11676_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04021_ ) );
MUX2_X1 _11677_ ( .A(_04020_ ), .B(_04021_ ), .S(_03851_ ), .Z(_04022_ ) );
OAI211_X1 _11678_ ( .A(_03244_ ), .B(_04019_ ), .C1(_04022_ ), .C2(_03687_ ), .ZN(_04023_ ) );
OAI211_X1 _11679_ ( .A(_04014_ ), .B(_04023_ ), .C1(_03699_ ), .C2(_03700_ ), .ZN(_04024_ ) );
NAND2_X1 _11680_ ( .A1(_04005_ ), .A2(_04024_ ), .ZN(_04025_ ) );
XNOR2_X1 _11681_ ( .A(_04004_ ), .B(_04025_ ), .ZN(_04026_ ) );
NOR2_X1 _11682_ ( .A1(_04003_ ), .A2(_04026_ ), .ZN(_04027_ ) );
AND3_X1 _11683_ ( .A1(_03935_ ), .A2(_03980_ ), .A3(_04027_ ), .ZN(_04028_ ) );
INV_X1 _11684_ ( .A(fanout_net_7 ), .ZN(_04029_ ) );
NOR2_X1 _11685_ ( .A1(_04029_ ), .A2(\ID_EX_typ [1] ), .ZN(_04030_ ) );
AND2_X1 _11686_ ( .A1(_04030_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04031_ ) );
INV_X1 _11687_ ( .A(_04031_ ), .ZN(_04032_ ) );
OR2_X1 _11688_ ( .A1(_03476_ ), .A2(fanout_net_8 ), .ZN(_04033_ ) );
NAND2_X1 _11689_ ( .A1(_02272_ ), .A2(fanout_net_8 ), .ZN(_04034_ ) );
NAND2_X1 _11690_ ( .A1(_04033_ ), .A2(_04034_ ), .ZN(_04035_ ) );
INV_X1 _11691_ ( .A(_02271_ ), .ZN(_04036_ ) );
NOR2_X1 _11692_ ( .A1(_04035_ ), .A2(_04036_ ), .ZN(_04037_ ) );
AOI21_X1 _11693_ ( .A(_02271_ ), .B1(_04033_ ), .B2(_04034_ ), .ZN(_04038_ ) );
NOR2_X1 _11694_ ( .A1(_04037_ ), .A2(_04038_ ), .ZN(_04039_ ) );
INV_X2 _11695_ ( .A(fanout_net_8 ), .ZN(_04040_ ) );
BUF_X4 _11696_ ( .A(_04040_ ), .Z(_04041_ ) );
BUF_X4 _11697_ ( .A(_04041_ ), .Z(_04042_ ) );
NAND3_X1 _11698_ ( .A1(_03480_ ), .A2(_04042_ ), .A3(_03499_ ), .ZN(_04043_ ) );
NAND2_X1 _11699_ ( .A1(_02227_ ), .A2(fanout_net_8 ), .ZN(_04044_ ) );
NAND2_X1 _11700_ ( .A1(_04043_ ), .A2(_04044_ ), .ZN(_04045_ ) );
XNOR2_X1 _11701_ ( .A(_04045_ ), .B(_03478_ ), .ZN(_04046_ ) );
NOR2_X1 _11702_ ( .A1(_04039_ ), .A2(_04046_ ), .ZN(_04047_ ) );
INV_X1 _11703_ ( .A(_04047_ ), .ZN(_04048_ ) );
BUF_X2 _11704_ ( .A(_04042_ ), .Z(_04049_ ) );
NAND3_X1 _11705_ ( .A1(_03505_ ), .A2(_04049_ ), .A3(_03531_ ), .ZN(_04050_ ) );
NAND2_X1 _11706_ ( .A1(_02297_ ), .A2(fanout_net_8 ), .ZN(_04051_ ) );
NAND2_X1 _11707_ ( .A1(_04050_ ), .A2(_04051_ ), .ZN(_04052_ ) );
NAND3_X1 _11708_ ( .A1(_03552_ ), .A2(_03554_ ), .A3(_04049_ ), .ZN(_04053_ ) );
NAND2_X1 _11709_ ( .A1(_02321_ ), .A2(fanout_net_8 ), .ZN(_04054_ ) );
NAND2_X1 _11710_ ( .A1(_04053_ ), .A2(_04054_ ), .ZN(_04055_ ) );
INV_X1 _11711_ ( .A(_02320_ ), .ZN(_04056_ ) );
AND2_X1 _11712_ ( .A1(_04055_ ), .A2(_04056_ ), .ZN(_04057_ ) );
NOR2_X1 _11713_ ( .A1(_04055_ ), .A2(_04056_ ), .ZN(_04058_ ) );
OAI211_X1 _11714_ ( .A(_04052_ ), .B(_02296_ ), .C1(_04057_ ), .C2(_04058_ ), .ZN(_04059_ ) );
NAND2_X1 _11715_ ( .A1(_04055_ ), .A2(_02320_ ), .ZN(_04060_ ) );
AOI21_X1 _11716_ ( .A(_04048_ ), .B1(_04059_ ), .B2(_04060_ ), .ZN(_04061_ ) );
INV_X1 _11717_ ( .A(_04046_ ), .ZN(_04062_ ) );
AND3_X1 _11718_ ( .A1(_04062_ ), .A2(_02271_ ), .A3(_04035_ ), .ZN(_04063_ ) );
INV_X1 _11719_ ( .A(_03478_ ), .ZN(_04064_ ) );
AOI21_X1 _11720_ ( .A(_04064_ ), .B1(_04043_ ), .B2(_04044_ ), .ZN(_04065_ ) );
NOR3_X1 _11721_ ( .A1(_04061_ ), .A2(_04063_ ), .A3(_04065_ ), .ZN(_04066_ ) );
NAND3_X1 _11722_ ( .A1(_03773_ ), .A2(_03792_ ), .A3(_04040_ ), .ZN(_04067_ ) );
NAND2_X1 _11723_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [14] ), .ZN(_04068_ ) );
AND2_X1 _11724_ ( .A1(_04067_ ), .A2(_04068_ ), .ZN(_04069_ ) );
XNOR2_X1 _11725_ ( .A(_04069_ ), .B(_02575_ ), .ZN(_04070_ ) );
NAND3_X1 _11726_ ( .A1(_03751_ ), .A2(_04040_ ), .A3(_03770_ ), .ZN(_04071_ ) );
NAND2_X1 _11727_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [15] ), .ZN(_04072_ ) );
AND2_X2 _11728_ ( .A1(_04071_ ), .A2(_04072_ ), .ZN(_04073_ ) );
XNOR2_X2 _11729_ ( .A(_04073_ ), .B(_02553_ ), .ZN(_04074_ ) );
NOR2_X2 _11730_ ( .A1(_04070_ ), .A2(_04074_ ), .ZN(_04075_ ) );
NAND3_X1 _11731_ ( .A1(_03866_ ), .A2(_03885_ ), .A3(_04041_ ), .ZN(_04076_ ) );
NAND2_X1 _11732_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [10] ), .ZN(_04077_ ) );
AND2_X4 _11733_ ( .A1(_04076_ ), .A2(_04077_ ), .ZN(_04078_ ) );
XNOR2_X1 _11734_ ( .A(_04078_ ), .B(_02718_ ), .ZN(_04079_ ) );
NAND3_X1 _11735_ ( .A1(_03843_ ), .A2(_04040_ ), .A3(_03863_ ), .ZN(_04080_ ) );
NAND2_X1 _11736_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [11] ), .ZN(_04081_ ) );
AND2_X1 _11737_ ( .A1(_04080_ ), .A2(_04081_ ), .ZN(_04082_ ) );
INV_X4 _11738_ ( .A(_02694_ ), .ZN(_04083_ ) );
NOR2_X1 _11739_ ( .A1(_04082_ ), .A2(_04083_ ), .ZN(_04084_ ) );
AND3_X1 _11740_ ( .A1(_04083_ ), .A2(_04081_ ), .A3(_04080_ ), .ZN(_04085_ ) );
NOR2_X2 _11741_ ( .A1(_04084_ ), .A2(_04085_ ), .ZN(_04086_ ) );
NOR2_X1 _11742_ ( .A1(_04079_ ), .A2(_04086_ ), .ZN(_04087_ ) );
NAND3_X1 _11743_ ( .A1(_03796_ ), .A2(_03815_ ), .A3(_04041_ ), .ZN(_04088_ ) );
NAND2_X1 _11744_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [12] ), .ZN(_04089_ ) );
AND2_X2 _11745_ ( .A1(_04088_ ), .A2(_04089_ ), .ZN(_04090_ ) );
XNOR2_X1 _11746_ ( .A(_04090_ ), .B(_02622_ ), .ZN(_04091_ ) );
INV_X1 _11747_ ( .A(_04091_ ), .ZN(_04092_ ) );
NAND3_X1 _11748_ ( .A1(_03818_ ), .A2(_04040_ ), .A3(_03837_ ), .ZN(_04093_ ) );
NAND2_X1 _11749_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [13] ), .ZN(_04094_ ) );
AND2_X4 _11750_ ( .A1(_04093_ ), .A2(_04094_ ), .ZN(_04095_ ) );
XNOR2_X1 _11751_ ( .A(_04095_ ), .B(_02599_ ), .ZN(_04096_ ) );
INV_X1 _11752_ ( .A(_04096_ ), .ZN(_04097_ ) );
AND4_X2 _11753_ ( .A1(_04075_ ), .A2(_04087_ ), .A3(_04092_ ), .A4(_04097_ ), .ZN(_04098_ ) );
NAND3_X1 _11754_ ( .A1(_03911_ ), .A2(_03930_ ), .A3(_04042_ ), .ZN(_04099_ ) );
NAND2_X1 _11755_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [8] ), .ZN(_04100_ ) );
AND2_X2 _11756_ ( .A1(_04099_ ), .A2(_04100_ ), .ZN(_04101_ ) );
XNOR2_X1 _11757_ ( .A(_04101_ ), .B(_02647_ ), .ZN(_04102_ ) );
INV_X1 _11758_ ( .A(_04102_ ), .ZN(_04103_ ) );
NAND3_X1 _11759_ ( .A1(_03889_ ), .A2(_04041_ ), .A3(_03908_ ), .ZN(_04104_ ) );
NAND2_X1 _11760_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [9] ), .ZN(_04105_ ) );
AND2_X1 _11761_ ( .A1(_04104_ ), .A2(_04105_ ), .ZN(_04106_ ) );
INV_X1 _11762_ ( .A(_02670_ ), .ZN(_04107_ ) );
NOR2_X1 _11763_ ( .A1(_04106_ ), .A2(_04107_ ), .ZN(_04108_ ) );
AND2_X1 _11764_ ( .A1(_04106_ ), .A2(_04107_ ), .ZN(_04109_ ) );
OAI211_X1 _11765_ ( .A(_04098_ ), .B(_04103_ ), .C1(_04108_ ), .C2(_04109_ ), .ZN(_04110_ ) );
NAND3_X1 _11766_ ( .A1(_03651_ ), .A2(_04040_ ), .A3(_03671_ ), .ZN(_04111_ ) );
NAND2_X1 _11767_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [7] ), .ZN(_04112_ ) );
AND2_X1 _11768_ ( .A1(_04111_ ), .A2(_04112_ ), .ZN(_04113_ ) );
INV_X1 _11769_ ( .A(_02914_ ), .ZN(_04114_ ) );
NOR2_X1 _11770_ ( .A1(_04113_ ), .A2(_04114_ ), .ZN(_04115_ ) );
AND3_X1 _11771_ ( .A1(_04114_ ), .A2(_04112_ ), .A3(_04111_ ), .ZN(_04116_ ) );
NOR2_X2 _11772_ ( .A1(_04115_ ), .A2(_04116_ ), .ZN(_04117_ ) );
INV_X1 _11773_ ( .A(_04117_ ), .ZN(_04118_ ) );
NAND3_X1 _11774_ ( .A1(_03675_ ), .A2(_03701_ ), .A3(_04041_ ), .ZN(_04119_ ) );
NAND2_X1 _11775_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [6] ), .ZN(_04120_ ) );
AND2_X2 _11776_ ( .A1(_04119_ ), .A2(_04120_ ), .ZN(_04121_ ) );
AND3_X1 _11777_ ( .A1(_04118_ ), .A2(_02890_ ), .A3(_04121_ ), .ZN(_04122_ ) );
NAND2_X1 _11778_ ( .A1(_03748_ ), .A2(_04040_ ), .ZN(_04123_ ) );
OR2_X1 _11779_ ( .A1(_04040_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04124_ ) );
NAND2_X2 _11780_ ( .A1(_04123_ ), .A2(_04124_ ), .ZN(_04125_ ) );
XNOR2_X2 _11781_ ( .A(_04125_ ), .B(_02923_ ), .ZN(_04126_ ) );
INV_X1 _11782_ ( .A(_04126_ ), .ZN(_04127_ ) );
NAND2_X1 _11783_ ( .A1(_03726_ ), .A2(_04042_ ), .ZN(_04128_ ) );
NAND2_X1 _11784_ ( .A1(_02843_ ), .A2(fanout_net_8 ), .ZN(_04129_ ) );
NAND2_X1 _11785_ ( .A1(_04128_ ), .A2(_04129_ ), .ZN(_04130_ ) );
NAND3_X1 _11786_ ( .A1(_04127_ ), .A2(_02842_ ), .A3(_04130_ ), .ZN(_04131_ ) );
OAI21_X1 _11787_ ( .A(_04131_ ), .B1(_02923_ ), .B2(_04125_ ), .ZN(_04132_ ) );
XNOR2_X1 _11788_ ( .A(_04121_ ), .B(_02890_ ), .ZN(_04133_ ) );
NOR2_X1 _11789_ ( .A1(_04133_ ), .A2(_04117_ ), .ZN(_04134_ ) );
AOI221_X1 _11790_ ( .A(_04122_ ), .B1(_02914_ ), .B2(_04113_ ), .C1(_04132_ ), .C2(_04134_ ), .ZN(_04135_ ) );
NAND3_X1 _11791_ ( .A1(_03958_ ), .A2(_04040_ ), .A3(_03977_ ), .ZN(_04136_ ) );
NAND2_X1 _11792_ ( .A1(fanout_net_8 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_04137_ ) );
AND2_X4 _11793_ ( .A1(_04136_ ), .A2(_04137_ ), .ZN(_04138_ ) );
XNOR2_X1 _11794_ ( .A(_04138_ ), .B(_02819_ ), .ZN(_04139_ ) );
NAND3_X1 _11795_ ( .A1(_03936_ ), .A2(_03955_ ), .A3(_04040_ ), .ZN(_04140_ ) );
NAND2_X1 _11796_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [2] ), .ZN(_04141_ ) );
AND2_X2 _11797_ ( .A1(_04140_ ), .A2(_04141_ ), .ZN(_04142_ ) );
XNOR2_X1 _11798_ ( .A(_04142_ ), .B(_02741_ ), .ZN(_04143_ ) );
NAND2_X1 _11799_ ( .A1(_04001_ ), .A2(_04041_ ), .ZN(_04144_ ) );
NAND2_X1 _11800_ ( .A1(_02765_ ), .A2(fanout_net_8 ), .ZN(_04145_ ) );
NAND2_X1 _11801_ ( .A1(_04144_ ), .A2(_04145_ ), .ZN(_04146_ ) );
NAND2_X1 _11802_ ( .A1(_04146_ ), .A2(_02764_ ), .ZN(_04147_ ) );
AND3_X1 _11803_ ( .A1(_04144_ ), .A2(_02764_ ), .A3(_04145_ ), .ZN(_04148_ ) );
AOI21_X1 _11804_ ( .A(_02764_ ), .B1(_04144_ ), .B2(_04145_ ), .ZN(_04149_ ) );
NAND2_X1 _11805_ ( .A1(_04025_ ), .A2(_04041_ ), .ZN(_04150_ ) );
OR2_X2 _11806_ ( .A1(_04041_ ), .A2(\ID_EX_imm [0] ), .ZN(_04151_ ) );
NAND2_X1 _11807_ ( .A1(_04150_ ), .A2(_04151_ ), .ZN(_04152_ ) );
OAI22_X1 _11808_ ( .A1(_04148_ ), .A2(_04149_ ), .B1(_04004_ ), .B2(_04152_ ), .ZN(_04153_ ) );
AOI211_X1 _11809_ ( .A(_04139_ ), .B(_04143_ ), .C1(_04147_ ), .C2(_04153_ ), .ZN(_04154_ ) );
AOI21_X1 _11810_ ( .A(_02819_ ), .B1(_04137_ ), .B2(_04136_ ), .ZN(_04155_ ) );
INV_X2 _11811_ ( .A(_04142_ ), .ZN(_04156_ ) );
NOR3_X1 _11812_ ( .A1(_04139_ ), .A2(_02793_ ), .A3(_04156_ ), .ZN(_04157_ ) );
OR3_X2 _11813_ ( .A1(_04154_ ), .A2(_04155_ ), .A3(_04157_ ), .ZN(_04158_ ) );
INV_X1 _11814_ ( .A(_02842_ ), .ZN(_04159_ ) );
NOR2_X1 _11815_ ( .A1(_04130_ ), .A2(_04159_ ), .ZN(_04160_ ) );
AOI21_X1 _11816_ ( .A(_02842_ ), .B1(_04128_ ), .B2(_04129_ ), .ZN(_04161_ ) );
NOR2_X1 _11817_ ( .A1(_04160_ ), .A2(_04161_ ), .ZN(_04162_ ) );
INV_X1 _11818_ ( .A(_04162_ ), .ZN(_04163_ ) );
NAND4_X1 _11819_ ( .A1(_04158_ ), .A2(_04134_ ), .A3(_04127_ ), .A4(_04163_ ), .ZN(_04164_ ) );
AOI21_X1 _11820_ ( .A(_04110_ ), .B1(_04135_ ), .B2(_04164_ ), .ZN(_04165_ ) );
INV_X1 _11821_ ( .A(_02575_ ), .ZN(_04166_ ) );
INV_X1 _11822_ ( .A(_04069_ ), .ZN(_04167_ ) );
NOR3_X1 _11823_ ( .A1(_04074_ ), .A2(_04166_ ), .A3(_04167_ ), .ZN(_04168_ ) );
AND3_X1 _11824_ ( .A1(_04075_ ), .A2(_04092_ ), .A3(_04097_ ), .ZN(_04169_ ) );
INV_X1 _11825_ ( .A(_04087_ ), .ZN(_04170_ ) );
NAND3_X1 _11826_ ( .A1(_04104_ ), .A2(_02670_ ), .A3(_04105_ ), .ZN(_04171_ ) );
OAI211_X1 _11827_ ( .A(_02647_ ), .B(_04101_ ), .C1(_04109_ ), .C2(_04108_ ), .ZN(_04172_ ) );
AOI21_X1 _11828_ ( .A(_04170_ ), .B1(_04171_ ), .B2(_04172_ ), .ZN(_04173_ ) );
INV_X1 _11829_ ( .A(_04086_ ), .ZN(_04174_ ) );
NAND3_X1 _11830_ ( .A1(_04174_ ), .A2(_02718_ ), .A3(_04078_ ), .ZN(_04175_ ) );
INV_X1 _11831_ ( .A(_04082_ ), .ZN(_04176_ ) );
OAI21_X1 _11832_ ( .A(_04175_ ), .B1(_04083_ ), .B2(_04176_ ), .ZN(_04177_ ) );
OAI21_X1 _11833_ ( .A(_04169_ ), .B1(_04173_ ), .B2(_04177_ ), .ZN(_04178_ ) );
INV_X1 _11834_ ( .A(_02622_ ), .ZN(_04179_ ) );
INV_X1 _11835_ ( .A(_04090_ ), .ZN(_04180_ ) );
NOR3_X1 _11836_ ( .A1(_04096_ ), .A2(_04179_ ), .A3(_04180_ ), .ZN(_04181_ ) );
AND3_X1 _11837_ ( .A1(_04093_ ), .A2(_02600_ ), .A3(_04094_ ), .ZN(_04182_ ) );
OAI21_X1 _11838_ ( .A(_04075_ ), .B1(_04181_ ), .B2(_04182_ ), .ZN(_04183_ ) );
INV_X1 _11839_ ( .A(_02553_ ), .ZN(_04184_ ) );
INV_X1 _11840_ ( .A(_04073_ ), .ZN(_04185_ ) );
OAI211_X1 _11841_ ( .A(_04178_ ), .B(_04183_ ), .C1(_04184_ ), .C2(_04185_ ), .ZN(_04186_ ) );
OR3_X2 _11842_ ( .A1(_04165_ ), .A2(_04168_ ), .A3(_04186_ ), .ZN(_04187_ ) );
NAND3_X1 _11843_ ( .A1(_03383_ ), .A2(_03402_ ), .A3(_04042_ ), .ZN(_04188_ ) );
NAND2_X1 _11844_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [22] ), .ZN(_04189_ ) );
AND2_X1 _11845_ ( .A1(_04188_ ), .A2(_04189_ ), .ZN(_04190_ ) );
XNOR2_X1 _11846_ ( .A(_04190_ ), .B(_02429_ ), .ZN(_04191_ ) );
NAND3_X1 _11847_ ( .A1(_03361_ ), .A2(_04041_ ), .A3(_03380_ ), .ZN(_04192_ ) );
NAND2_X1 _11848_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [23] ), .ZN(_04193_ ) );
AND2_X1 _11849_ ( .A1(_04192_ ), .A2(_04193_ ), .ZN(_04194_ ) );
INV_X1 _11850_ ( .A(_02406_ ), .ZN(_04195_ ) );
NOR2_X1 _11851_ ( .A1(_04194_ ), .A2(_04195_ ), .ZN(_04196_ ) );
AND3_X1 _11852_ ( .A1(_04195_ ), .A2(_04193_ ), .A3(_04192_ ), .ZN(_04197_ ) );
NOR2_X1 _11853_ ( .A1(_04196_ ), .A2(_04197_ ), .ZN(_04198_ ) );
NOR2_X1 _11854_ ( .A1(_04191_ ), .A2(_04198_ ), .ZN(_04199_ ) );
NAND3_X1 _11855_ ( .A1(_03406_ ), .A2(_03425_ ), .A3(_04042_ ), .ZN(_04200_ ) );
NAND2_X1 _11856_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [20] ), .ZN(_04201_ ) );
AND2_X2 _11857_ ( .A1(_04200_ ), .A2(_04201_ ), .ZN(_04202_ ) );
XNOR2_X1 _11858_ ( .A(_04202_ ), .B(_02358_ ), .ZN(_04203_ ) );
INV_X1 _11859_ ( .A(_04203_ ), .ZN(_04204_ ) );
AOI21_X1 _11860_ ( .A(fanout_net_8 ), .B1(_03445_ ), .B2(_03446_ ), .ZN(_04205_ ) );
NOR2_X1 _11861_ ( .A1(_04042_ ), .A2(\ID_EX_imm [21] ), .ZN(_04206_ ) );
NOR2_X2 _11862_ ( .A1(_04205_ ), .A2(_04206_ ), .ZN(_04207_ ) );
INV_X1 _11863_ ( .A(_03448_ ), .ZN(_04208_ ) );
XNOR2_X1 _11864_ ( .A(_04207_ ), .B(_04208_ ), .ZN(_04209_ ) );
INV_X1 _11865_ ( .A(_04209_ ), .ZN(_04210_ ) );
AND3_X1 _11866_ ( .A1(_04199_ ), .A2(_04204_ ), .A3(_04210_ ), .ZN(_04211_ ) );
NAND3_X1 _11867_ ( .A1(_03307_ ), .A2(_03308_ ), .A3(_04042_ ), .ZN(_04212_ ) );
NAND2_X1 _11868_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [18] ), .ZN(_04213_ ) );
AND2_X2 _11869_ ( .A1(_04212_ ), .A2(_04213_ ), .ZN(_04214_ ) );
XNOR2_X1 _11870_ ( .A(_04214_ ), .B(_02501_ ), .ZN(_04215_ ) );
NAND3_X1 _11871_ ( .A1(_03331_ ), .A2(_03332_ ), .A3(_04042_ ), .ZN(_04216_ ) );
NAND2_X1 _11872_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [16] ), .ZN(_04217_ ) );
AND2_X1 _11873_ ( .A1(_04216_ ), .A2(_04217_ ), .ZN(_04218_ ) );
INV_X1 _11874_ ( .A(_02453_ ), .ZN(_04219_ ) );
NOR2_X1 _11875_ ( .A1(_04218_ ), .A2(_04219_ ), .ZN(_04220_ ) );
AND3_X1 _11876_ ( .A1(_04219_ ), .A2(_04217_ ), .A3(_04216_ ), .ZN(_04221_ ) );
NOR2_X1 _11877_ ( .A1(_04220_ ), .A2(_04221_ ), .ZN(_04222_ ) );
NAND3_X1 _11878_ ( .A1(_03335_ ), .A2(_04042_ ), .A3(_03355_ ), .ZN(_04223_ ) );
NAND2_X1 _11879_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [17] ), .ZN(_04224_ ) );
AND2_X4 _11880_ ( .A1(_04223_ ), .A2(_04224_ ), .ZN(_04225_ ) );
XNOR2_X1 _11881_ ( .A(_04225_ ), .B(_02476_ ), .ZN(_04226_ ) );
NAND3_X1 _11882_ ( .A1(_03242_ ), .A2(_04041_ ), .A3(_03279_ ), .ZN(_04227_ ) );
NAND2_X1 _11883_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [19] ), .ZN(_04228_ ) );
AND2_X1 _11884_ ( .A1(_04227_ ), .A2(_04228_ ), .ZN(_04229_ ) );
INV_X1 _11885_ ( .A(_02524_ ), .ZN(_04230_ ) );
NOR2_X1 _11886_ ( .A1(_04229_ ), .A2(_04230_ ), .ZN(_04231_ ) );
AND3_X1 _11887_ ( .A1(_04230_ ), .A2(_04228_ ), .A3(_04227_ ), .ZN(_04232_ ) );
NOR2_X4 _11888_ ( .A1(_04231_ ), .A2(_04232_ ), .ZN(_04233_ ) );
NOR4_X1 _11889_ ( .A1(_04215_ ), .A2(_04222_ ), .A3(_04226_ ), .A4(_04233_ ), .ZN(_04234_ ) );
AND2_X1 _11890_ ( .A1(_04211_ ), .A2(_04234_ ), .ZN(_04235_ ) );
AND2_X2 _11891_ ( .A1(_04187_ ), .A2(_04235_ ), .ZN(_04236_ ) );
NAND3_X1 _11892_ ( .A1(_04199_ ), .A2(_04204_ ), .A3(_04210_ ), .ZN(_04237_ ) );
OR2_X1 _11893_ ( .A1(_04215_ ), .A2(_04233_ ), .ZN(_04238_ ) );
NAND3_X1 _11894_ ( .A1(_04223_ ), .A2(_02476_ ), .A3(_04224_ ), .ZN(_04239_ ) );
AND2_X1 _11895_ ( .A1(_04225_ ), .A2(_02946_ ), .ZN(_04240_ ) );
NOR2_X1 _11896_ ( .A1(_04225_ ), .A2(_02946_ ), .ZN(_04241_ ) );
OAI211_X1 _11897_ ( .A(_02453_ ), .B(_04218_ ), .C1(_04240_ ), .C2(_04241_ ), .ZN(_04242_ ) );
AOI21_X1 _11898_ ( .A(_04238_ ), .B1(_04239_ ), .B2(_04242_ ), .ZN(_04243_ ) );
AOI21_X1 _11899_ ( .A(_04243_ ), .B1(_02524_ ), .B2(_04229_ ), .ZN(_04244_ ) );
INV_X1 _11900_ ( .A(_04233_ ), .ZN(_04245_ ) );
NAND3_X1 _11901_ ( .A1(_04245_ ), .A2(_02501_ ), .A3(_04214_ ), .ZN(_04246_ ) );
AOI21_X1 _11902_ ( .A(_04237_ ), .B1(_04244_ ), .B2(_04246_ ), .ZN(_04247_ ) );
INV_X1 _11903_ ( .A(_02429_ ), .ZN(_04248_ ) );
INV_X1 _11904_ ( .A(_04190_ ), .ZN(_04249_ ) );
NOR3_X1 _11905_ ( .A1(_04198_ ), .A2(_04248_ ), .A3(_04249_ ), .ZN(_04250_ ) );
INV_X1 _11906_ ( .A(_02358_ ), .ZN(_04251_ ) );
INV_X1 _11907_ ( .A(_04202_ ), .ZN(_04252_ ) );
NOR3_X1 _11908_ ( .A1(_04209_ ), .A2(_04251_ ), .A3(_04252_ ), .ZN(_04253_ ) );
NOR2_X1 _11909_ ( .A1(_04207_ ), .A2(_04208_ ), .ZN(_04254_ ) );
OAI21_X1 _11910_ ( .A(_04199_ ), .B1(_04253_ ), .B2(_04254_ ), .ZN(_04255_ ) );
INV_X1 _11911_ ( .A(_04194_ ), .ZN(_04256_ ) );
OAI21_X1 _11912_ ( .A(_04255_ ), .B1(_04195_ ), .B2(_04256_ ), .ZN(_04257_ ) );
NOR4_X2 _11913_ ( .A1(_04236_ ), .A2(_04247_ ), .A3(_04250_ ), .A4(_04257_ ), .ZN(_04258_ ) );
XNOR2_X1 _11914_ ( .A(_04055_ ), .B(_02320_ ), .ZN(_04259_ ) );
INV_X1 _11915_ ( .A(_04259_ ), .ZN(_04260_ ) );
INV_X1 _11916_ ( .A(_02296_ ), .ZN(_04261_ ) );
NOR2_X1 _11917_ ( .A1(_04052_ ), .A2(_04261_ ), .ZN(_04262_ ) );
AOI21_X1 _11918_ ( .A(_02296_ ), .B1(_04050_ ), .B2(_04051_ ), .ZN(_04263_ ) );
NOR2_X1 _11919_ ( .A1(_04262_ ), .A2(_04263_ ), .ZN(_04264_ ) );
INV_X1 _11920_ ( .A(_04264_ ), .ZN(_04265_ ) );
NAND3_X1 _11921_ ( .A1(_04047_ ), .A2(_04260_ ), .A3(_04265_ ), .ZN(_04266_ ) );
OAI21_X2 _11922_ ( .A(_04066_ ), .B1(_04258_ ), .B2(_04266_ ), .ZN(_04267_ ) );
NAND3_X1 _11923_ ( .A1(_03626_ ), .A2(_04049_ ), .A3(_03645_ ), .ZN(_04268_ ) );
NAND2_X1 _11924_ ( .A1(fanout_net_8 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04269_ ) );
AND2_X1 _11925_ ( .A1(_04268_ ), .A2(_04269_ ), .ZN(_04270_ ) );
XNOR2_X1 _11926_ ( .A(_04270_ ), .B(_02199_ ), .ZN(_04271_ ) );
INV_X1 _11927_ ( .A(_03025_ ), .ZN(_04272_ ) );
NAND3_X1 _11928_ ( .A1(_03604_ ), .A2(_04049_ ), .A3(_03623_ ), .ZN(_04273_ ) );
INV_X1 _11929_ ( .A(\ID_EX_imm [31] ), .ZN(_04274_ ) );
NAND2_X1 _11930_ ( .A1(_04274_ ), .A2(fanout_net_8 ), .ZN(_04275_ ) );
NAND2_X1 _11931_ ( .A1(_04273_ ), .A2(_04275_ ), .ZN(_04276_ ) );
NAND2_X1 _11932_ ( .A1(_04272_ ), .A2(_04276_ ), .ZN(_04277_ ) );
NAND3_X1 _11933_ ( .A1(_03025_ ), .A2(_04273_ ), .A3(_04275_ ), .ZN(_04278_ ) );
NAND2_X1 _11934_ ( .A1(_04277_ ), .A2(_04278_ ), .ZN(_04279_ ) );
INV_X1 _11935_ ( .A(_04279_ ), .ZN(_04280_ ) );
NOR2_X1 _11936_ ( .A1(_04271_ ), .A2(_04280_ ), .ZN(_04281_ ) );
NAND3_X1 _11937_ ( .A1(_03581_ ), .A2(_04049_ ), .A3(_03600_ ), .ZN(_04282_ ) );
NAND2_X1 _11938_ ( .A1(\ID_EX_typ [4] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04283_ ) );
AND2_X2 _11939_ ( .A1(_04282_ ), .A2(_04283_ ), .ZN(_04284_ ) );
XNOR2_X1 _11940_ ( .A(_04284_ ), .B(_02998_ ), .ZN(_04285_ ) );
INV_X1 _11941_ ( .A(_04285_ ), .ZN(_04286_ ) );
NAND3_X1 _11942_ ( .A1(_03559_ ), .A2(_04049_ ), .A3(_03578_ ), .ZN(_04287_ ) );
NAND2_X1 _11943_ ( .A1(\ID_EX_typ [4] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04288_ ) );
AND2_X1 _11944_ ( .A1(_04287_ ), .A2(_04288_ ), .ZN(_04289_ ) );
INV_X1 _11945_ ( .A(_02224_ ), .ZN(_04290_ ) );
XNOR2_X1 _11946_ ( .A(_04289_ ), .B(_04290_ ), .ZN(_04291_ ) );
INV_X1 _11947_ ( .A(_04291_ ), .ZN(_04292_ ) );
AND3_X1 _11948_ ( .A1(_04281_ ), .A2(_04286_ ), .A3(_04292_ ), .ZN(_04293_ ) );
AND2_X2 _11949_ ( .A1(_04267_ ), .A2(_04293_ ), .ZN(_04294_ ) );
INV_X1 _11950_ ( .A(_04289_ ), .ZN(_04295_ ) );
AND2_X1 _11951_ ( .A1(_04284_ ), .A2(_02992_ ), .ZN(_04296_ ) );
NOR2_X1 _11952_ ( .A1(_04284_ ), .A2(_02992_ ), .ZN(_04297_ ) );
OAI211_X1 _11953_ ( .A(_04295_ ), .B(_02224_ ), .C1(_04296_ ), .C2(_04297_ ), .ZN(_04298_ ) );
OAI21_X1 _11954_ ( .A(_04298_ ), .B1(_02998_ ), .B2(_04284_ ), .ZN(_04299_ ) );
AND2_X1 _11955_ ( .A1(_04299_ ), .A2(_04281_ ), .ZN(_04300_ ) );
AOI21_X1 _11956_ ( .A(_02199_ ), .B1(_04268_ ), .B2(_04269_ ), .ZN(_04301_ ) );
AOI21_X1 _11957_ ( .A(_04300_ ), .B1(_04279_ ), .B2(_04301_ ), .ZN(_04302_ ) );
OAI21_X1 _11958_ ( .A(_04302_ ), .B1(_03025_ ), .B2(_04276_ ), .ZN(_04303_ ) );
INV_X1 _11959_ ( .A(\ID_EX_typ [1] ), .ZN(_04304_ ) );
NAND3_X1 _11960_ ( .A1(_04304_ ), .A2(_04029_ ), .A3(\ID_EX_typ [2] ), .ZN(_04305_ ) );
NOR3_X4 _11961_ ( .A1(_04294_ ), .A2(_04303_ ), .A3(_04305_ ), .ZN(_04306_ ) );
AND2_X1 _11962_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_7 ), .ZN(_04307_ ) );
AND2_X1 _11963_ ( .A1(_04307_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04308_ ) );
INV_X1 _11964_ ( .A(_04308_ ), .ZN(_04309_ ) );
AND2_X1 _11965_ ( .A1(_02647_ ), .A2(_03931_ ), .ZN(_04310_ ) );
AND2_X1 _11966_ ( .A1(_03910_ ), .A2(_04310_ ), .ZN(_04311_ ) );
AOI21_X1 _11967_ ( .A(_04311_ ), .B1(_02670_ ), .B2(_03909_ ), .ZN(_04312_ ) );
INV_X1 _11968_ ( .A(_04312_ ), .ZN(_04313_ ) );
AND2_X1 _11969_ ( .A1(_04313_ ), .A2(_03888_ ), .ZN(_04314_ ) );
AND2_X1 _11970_ ( .A1(_03864_ ), .A2(_02694_ ), .ZN(_04315_ ) );
AND2_X1 _11971_ ( .A1(_03886_ ), .A2(_02718_ ), .ZN(_04316_ ) );
AND2_X1 _11972_ ( .A1(_03865_ ), .A2(_04316_ ), .ZN(_04317_ ) );
NOR3_X1 _11973_ ( .A1(_04314_ ), .A2(_04315_ ), .A3(_04317_ ), .ZN(_04318_ ) );
INV_X1 _11974_ ( .A(_04318_ ), .ZN(_04319_ ) );
NAND2_X1 _11975_ ( .A1(_04319_ ), .A2(_03842_ ), .ZN(_04320_ ) );
AND3_X1 _11976_ ( .A1(_03841_ ), .A2(_02622_ ), .A3(_03816_ ), .ZN(_04321_ ) );
OAI21_X1 _11977_ ( .A(_03795_ ), .B1(_04321_ ), .B2(_03839_ ), .ZN(_04322_ ) );
AND2_X1 _11978_ ( .A1(_03793_ ), .A2(_02575_ ), .ZN(_04323_ ) );
AND2_X1 _11979_ ( .A1(_03772_ ), .A2(_04323_ ), .ZN(_04324_ ) );
AOI21_X1 _11980_ ( .A(_04324_ ), .B1(_02553_ ), .B2(_03771_ ), .ZN(_04325_ ) );
AND3_X1 _11981_ ( .A1(_04320_ ), .A2(_04322_ ), .A3(_04325_ ), .ZN(_04326_ ) );
NAND2_X1 _11982_ ( .A1(_02764_ ), .A2(_04001_ ), .ZN(_04327_ ) );
AOI21_X1 _11983_ ( .A(_04025_ ), .B1(_02788_ ), .B2(_02768_ ), .ZN(_04328_ ) );
OAI21_X2 _11984_ ( .A(_04327_ ), .B1(_04003_ ), .B2(_04328_ ), .ZN(_04329_ ) );
NAND2_X1 _11985_ ( .A1(_04329_ ), .A2(_03957_ ), .ZN(_04330_ ) );
AND2_X1 _11986_ ( .A1(_03956_ ), .A2(_02741_ ), .ZN(_04331_ ) );
INV_X1 _11987_ ( .A(_04331_ ), .ZN(_04332_ ) );
OAI211_X2 _11988_ ( .A(_04330_ ), .B(_04332_ ), .C1(_02819_ ), .C2(_03978_ ), .ZN(_04333_ ) );
NAND3_X1 _11989_ ( .A1(_03978_ ), .A2(_02795_ ), .A3(_02814_ ), .ZN(_04334_ ) );
NAND3_X1 _11990_ ( .A1(_04333_ ), .A2(_04334_ ), .A3(_03750_ ), .ZN(_04335_ ) );
AND3_X1 _11991_ ( .A1(_03673_ ), .A2(_02890_ ), .A3(_03702_ ), .ZN(_04336_ ) );
AND2_X1 _11992_ ( .A1(_02842_ ), .A2(_03726_ ), .ZN(_04337_ ) );
NAND2_X1 _11993_ ( .A1(_03749_ ), .A2(_04337_ ), .ZN(_04338_ ) );
OAI21_X1 _11994_ ( .A(_04338_ ), .B1(_02923_ ), .B2(_03748_ ), .ZN(_04339_ ) );
AOI221_X4 _11995_ ( .A(_04336_ ), .B1(_02914_ ), .B2(_03672_ ), .C1(_04339_ ), .C2(_03704_ ), .ZN(_04340_ ) );
AND2_X4 _11996_ ( .A1(_04335_ ), .A2(_04340_ ), .ZN(_04341_ ) );
INV_X4 _11997_ ( .A(_04341_ ), .ZN(_04342_ ) );
AND2_X4 _11998_ ( .A1(_03842_ ), .A2(_03933_ ), .ZN(_04343_ ) );
NAND2_X4 _11999_ ( .A1(_04342_ ), .A2(_04343_ ), .ZN(_04344_ ) );
AND2_X4 _12000_ ( .A1(_04326_ ), .A2(_04344_ ), .ZN(_04345_ ) );
INV_X2 _12001_ ( .A(_04345_ ), .ZN(_04346_ ) );
AND3_X4 _12002_ ( .A1(_04346_ ), .A2(_03453_ ), .A3(_03360_ ), .ZN(_04347_ ) );
INV_X1 _12003_ ( .A(_03357_ ), .ZN(_04348_ ) );
NAND2_X1 _12004_ ( .A1(_03333_ ), .A2(_02453_ ), .ZN(_04349_ ) );
AOI21_X1 _12005_ ( .A(_03358_ ), .B1(_04348_ ), .B2(_04349_ ), .ZN(_04350_ ) );
AND3_X1 _12006_ ( .A1(_04350_ ), .A2(_03281_ ), .A3(_03310_ ), .ZN(_04351_ ) );
AND2_X1 _12007_ ( .A1(_03280_ ), .A2(_02524_ ), .ZN(_04352_ ) );
AND3_X1 _12008_ ( .A1(_03281_ ), .A2(_02501_ ), .A3(_03309_ ), .ZN(_04353_ ) );
NOR3_X1 _12009_ ( .A1(_04351_ ), .A2(_04352_ ), .A3(_04353_ ), .ZN(_04354_ ) );
INV_X1 _12010_ ( .A(_03453_ ), .ZN(_04355_ ) );
NOR2_X1 _12011_ ( .A1(_04354_ ), .A2(_04355_ ), .ZN(_04356_ ) );
INV_X1 _12012_ ( .A(_04356_ ), .ZN(_04357_ ) );
INV_X1 _12013_ ( .A(_03405_ ), .ZN(_04358_ ) );
AOI21_X1 _12014_ ( .A(_03449_ ), .B1(_02358_ ), .B2(_03426_ ), .ZN(_04359_ ) );
NOR3_X1 _12015_ ( .A1(_04358_ ), .A2(_03450_ ), .A3(_04359_ ), .ZN(_04360_ ) );
INV_X1 _12016_ ( .A(_04360_ ), .ZN(_04361_ ) );
AND2_X1 _12017_ ( .A1(_03403_ ), .A2(_02429_ ), .ZN(_04362_ ) );
AND2_X1 _12018_ ( .A1(_03382_ ), .A2(_04362_ ), .ZN(_04363_ ) );
AOI21_X1 _12019_ ( .A(_04363_ ), .B1(_02406_ ), .B2(_03381_ ), .ZN(_04364_ ) );
AND3_X1 _12020_ ( .A1(_04357_ ), .A2(_04361_ ), .A3(_04364_ ), .ZN(_04365_ ) );
INV_X1 _12021_ ( .A(_04365_ ), .ZN(_04366_ ) );
OAI21_X1 _12022_ ( .A(_03649_ ), .B1(_04347_ ), .B2(_04366_ ), .ZN(_04367_ ) );
AND3_X1 _12023_ ( .A1(_02320_ ), .A2(_03554_ ), .A3(_03552_ ), .ZN(_04368_ ) );
NOR2_X1 _12024_ ( .A1(_04261_ ), .A2(_03532_ ), .ZN(_04369_ ) );
AND2_X1 _12025_ ( .A1(_03556_ ), .A2(_04369_ ), .ZN(_04370_ ) );
OAI21_X1 _12026_ ( .A(_03503_ ), .B1(_04368_ ), .B2(_04370_ ), .ZN(_04371_ ) );
INV_X1 _12027_ ( .A(_03476_ ), .ZN(_04372_ ) );
NAND4_X1 _12028_ ( .A1(_03500_ ), .A2(_04372_ ), .A3(_03502_ ), .A4(_02271_ ), .ZN(_04373_ ) );
AND3_X1 _12029_ ( .A1(_04371_ ), .A2(_03500_ ), .A3(_04373_ ), .ZN(_04374_ ) );
INV_X1 _12030_ ( .A(_03648_ ), .ZN(_04375_ ) );
NOR2_X1 _12031_ ( .A1(_04374_ ), .A2(_04375_ ), .ZN(_04376_ ) );
NOR2_X1 _12032_ ( .A1(_02199_ ), .A2(_03646_ ), .ZN(_04377_ ) );
NAND2_X1 _12033_ ( .A1(_03625_ ), .A2(_04377_ ), .ZN(_04378_ ) );
OAI21_X1 _12034_ ( .A(_04378_ ), .B1(_04272_ ), .B2(_03624_ ), .ZN(_04379_ ) );
NOR2_X1 _12035_ ( .A1(_04290_ ), .A2(_03579_ ), .ZN(_04380_ ) );
AOI21_X1 _12036_ ( .A(_03601_ ), .B1(_02971_ ), .B2(_02991_ ), .ZN(_04381_ ) );
NOR2_X1 _12037_ ( .A1(_04380_ ), .A2(_04381_ ), .ZN(_04382_ ) );
AOI21_X1 _12038_ ( .A(_02992_ ), .B1(_03581_ ), .B2(_03600_ ), .ZN(_04383_ ) );
NOR2_X1 _12039_ ( .A1(_04382_ ), .A2(_04383_ ), .ZN(_04384_ ) );
AND3_X1 _12040_ ( .A1(_04384_ ), .A2(_03625_ ), .A3(_03647_ ), .ZN(_04385_ ) );
NOR3_X1 _12041_ ( .A1(_04376_ ), .A2(_04379_ ), .A3(_04385_ ), .ZN(_04386_ ) );
AOI21_X1 _12042_ ( .A(_04309_ ), .B1(_04367_ ), .B2(_04386_ ), .ZN(_04387_ ) );
AND2_X1 _12043_ ( .A1(_04030_ ), .A2(\ID_EX_typ [2] ), .ZN(_04388_ ) );
AND3_X2 _12044_ ( .A1(_04367_ ), .A2(_04386_ ), .A3(_04388_ ), .ZN(_04389_ ) );
OR4_X4 _12045_ ( .A1(_04306_ ), .A2(_04387_ ), .A3(_04031_ ), .A4(_04389_ ), .ZN(_04390_ ) );
AOI21_X1 _12046_ ( .A(_04303_ ), .B1(_04267_ ), .B2(_04293_ ), .ZN(_04391_ ) );
NOR2_X1 _12047_ ( .A1(_04304_ ), .A2(fanout_net_7 ), .ZN(_04392_ ) );
INV_X1 _12048_ ( .A(\ID_EX_typ [2] ), .ZN(_04393_ ) );
AND2_X2 _12049_ ( .A1(_04392_ ), .A2(_04393_ ), .ZN(_04394_ ) );
INV_X1 _12050_ ( .A(_04394_ ), .ZN(_04395_ ) );
NOR2_X1 _12051_ ( .A1(_04391_ ), .A2(_04395_ ), .ZN(_04396_ ) );
OAI221_X2 _12052_ ( .A(_03226_ ), .B1(_04028_ ), .B2(_04032_ ), .C1(_04390_ ), .C2(_04396_ ), .ZN(_04397_ ) );
NAND4_X1 _12053_ ( .A1(_04343_ ), .A2(_03980_ ), .A3(_04027_ ), .A4(_03750_ ), .ZN(_04398_ ) );
OAI21_X1 _12054_ ( .A(_03225_ ), .B1(_04398_ ), .B2(_03650_ ), .ZN(_04399_ ) );
AND2_X4 _12055_ ( .A1(_04397_ ), .A2(_04399_ ), .ZN(_04400_ ) );
BUF_X8 _12056_ ( .A(_04400_ ), .Z(_04401_ ) );
MUX2_X1 _12057_ ( .A(_03104_ ), .B(_03223_ ), .S(_04401_ ), .Z(_04402_ ) );
OR2_X1 _12058_ ( .A1(_04402_ ), .A2(\ID_EX_typ [3] ), .ZN(_04403_ ) );
INV_X1 _12059_ ( .A(_02127_ ), .ZN(_04404_ ) );
BUF_X4 _12060_ ( .A(_04404_ ), .Z(_04405_ ) );
BUF_X4 _12061_ ( .A(_04405_ ), .Z(_04406_ ) );
INV_X1 _12062_ ( .A(\ID_EX_typ [3] ), .ZN(_04407_ ) );
BUF_X4 _12063_ ( .A(_04407_ ), .Z(_04408_ ) );
BUF_X4 _12064_ ( .A(_04408_ ), .Z(_04409_ ) );
XNOR2_X1 _12065_ ( .A(\EX_LS_dest_csreg_mem [8] ), .B(\ID_EX_csr [8] ), .ZN(_04410_ ) );
XNOR2_X1 _12066_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_04411_ ) );
INV_X1 _12067_ ( .A(\ID_EX_csr [6] ), .ZN(_04412_ ) );
NAND2_X1 _12068_ ( .A1(_04412_ ), .A2(\EX_LS_dest_csreg_mem [6] ), .ZN(_04413_ ) );
INV_X1 _12069_ ( .A(\ID_EX_csr [3] ), .ZN(_04414_ ) );
NAND2_X1 _12070_ ( .A1(_04414_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .ZN(_04415_ ) );
AND3_X1 _12071_ ( .A1(_04411_ ), .A2(_04413_ ), .A3(_04415_ ), .ZN(_04416_ ) );
INV_X1 _12072_ ( .A(\ID_EX_csr [1] ), .ZN(_04417_ ) );
INV_X1 _12073_ ( .A(\ID_EX_csr [5] ), .ZN(_04418_ ) );
AOI22_X1 _12074_ ( .A1(fanout_net_6 ), .A2(_04417_ ), .B1(_04418_ ), .B2(\EX_LS_dest_csreg_mem [5] ), .ZN(_04419_ ) );
INV_X1 _12075_ ( .A(fanout_net_6 ), .ZN(_04420_ ) );
INV_X1 _12076_ ( .A(\EX_LS_dest_csreg_mem [5] ), .ZN(_04421_ ) );
AOI22_X1 _12077_ ( .A1(_04420_ ), .A2(\ID_EX_csr [1] ), .B1(_04421_ ), .B2(\ID_EX_csr [5] ), .ZN(_04422_ ) );
AND3_X1 _12078_ ( .A1(_04416_ ), .A2(_04419_ ), .A3(_04422_ ), .ZN(_04423_ ) );
INV_X1 _12079_ ( .A(\EX_LS_dest_csreg_mem [6] ), .ZN(_04424_ ) );
NAND2_X1 _12080_ ( .A1(_04424_ ), .A2(\ID_EX_csr [6] ), .ZN(_04425_ ) );
INV_X1 _12081_ ( .A(\EX_LS_dest_csreg_mem [3] ), .ZN(_04426_ ) );
NAND2_X1 _12082_ ( .A1(_04426_ ), .A2(\ID_EX_csr [3] ), .ZN(_04427_ ) );
AND4_X2 _12083_ ( .A1(_04410_ ), .A2(_04423_ ), .A3(_04425_ ), .A4(_04427_ ), .ZN(_04428_ ) );
BUF_X2 _12084_ ( .A(_04428_ ), .Z(_04429_ ) );
INV_X1 _12085_ ( .A(\EX_LS_result_csreg_mem [30] ), .ZN(_04430_ ) );
XNOR2_X1 _12086_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .ZN(_04431_ ) );
XNOR2_X1 _12087_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_04432_ ) );
XNOR2_X1 _12088_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_04433_ ) );
XNOR2_X1 _12089_ ( .A(fanout_net_5 ), .B(\ID_EX_csr [0] ), .ZN(_04434_ ) );
AND4_X1 _12090_ ( .A1(_04431_ ), .A2(_04432_ ), .A3(_04433_ ), .A4(_04434_ ), .ZN(_04435_ ) );
XNOR2_X1 _12091_ ( .A(\EX_LS_dest_csreg_mem [9] ), .B(\ID_EX_csr [9] ), .ZN(_04436_ ) );
XNOR2_X1 _12092_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_04437_ ) );
AND4_X2 _12093_ ( .A1(_02173_ ), .A2(_04435_ ), .A3(_04436_ ), .A4(_04437_ ), .ZN(_04438_ ) );
BUF_X2 _12094_ ( .A(_04438_ ), .Z(_04439_ ) );
AND3_X1 _12095_ ( .A1(_04429_ ), .A2(_04430_ ), .A3(_04439_ ), .ZN(_04440_ ) );
AND2_X2 _12096_ ( .A1(_04428_ ), .A2(_04438_ ), .ZN(_04441_ ) );
AND4_X1 _12097_ ( .A1(\ID_EX_csr [10] ), .A2(_04418_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_04442_ ) );
AND2_X1 _12098_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_04443_ ) );
NOR2_X2 _12099_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_04444_ ) );
AND3_X1 _12100_ ( .A1(_04442_ ), .A2(_04443_ ), .A3(_04444_ ), .ZN(_04445_ ) );
INV_X1 _12101_ ( .A(\ID_EX_csr [2] ), .ZN(_04446_ ) );
NAND2_X1 _12102_ ( .A1(_04414_ ), .A2(_04446_ ), .ZN(_04447_ ) );
NAND2_X1 _12103_ ( .A1(_04417_ ), .A2(\ID_EX_csr [0] ), .ZN(_04448_ ) );
NOR2_X1 _12104_ ( .A1(_04447_ ), .A2(_04448_ ), .ZN(_04449_ ) );
AND2_X1 _12105_ ( .A1(_04445_ ), .A2(_04449_ ), .ZN(_04450_ ) );
NOR2_X1 _12106_ ( .A1(_04441_ ), .A2(_04450_ ), .ZN(_04451_ ) );
NOR4_X1 _12107_ ( .A1(\ID_EX_csr [10] ), .A2(\ID_EX_csr [5] ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_04452_ ) );
AND2_X2 _12108_ ( .A1(_04452_ ), .A2(_04443_ ), .ZN(_04453_ ) );
NOR3_X1 _12109_ ( .A1(_04447_ ), .A2(\ID_EX_csr [1] ), .A3(\ID_EX_csr [0] ), .ZN(_04454_ ) );
BUF_X2 _12110_ ( .A(_04454_ ), .Z(_04455_ ) );
BUF_X2 _12111_ ( .A(_04455_ ), .Z(_04456_ ) );
NAND4_X1 _12112_ ( .A1(_04453_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_04444_ ), .A4(_04456_ ), .ZN(_04457_ ) );
INV_X1 _12113_ ( .A(\ID_EX_csr [7] ), .ZN(_04458_ ) );
AND3_X1 _12114_ ( .A1(_04453_ ), .A2(_04458_ ), .A3(\ID_EX_csr [6] ), .ZN(_04459_ ) );
BUF_X4 _12115_ ( .A(_04459_ ), .Z(_04460_ ) );
BUF_X4 _12116_ ( .A(_04460_ ), .Z(_04461_ ) );
BUF_X4 _12117_ ( .A(_04461_ ), .Z(_04462_ ) );
BUF_X4 _12118_ ( .A(_04449_ ), .Z(_04463_ ) );
BUF_X4 _12119_ ( .A(_04463_ ), .Z(_04464_ ) );
NAND3_X1 _12120_ ( .A1(_04462_ ), .A2(\mepc [30] ), .A3(_04464_ ), .ZN(_04465_ ) );
NAND3_X1 _12121_ ( .A1(_04414_ ), .A2(_04446_ ), .A3(\ID_EX_csr [1] ), .ZN(_04466_ ) );
NOR2_X1 _12122_ ( .A1(_04466_ ), .A2(\ID_EX_csr [0] ), .ZN(_04467_ ) );
BUF_X4 _12123_ ( .A(_04467_ ), .Z(_04468_ ) );
BUF_X4 _12124_ ( .A(_04468_ ), .Z(_04469_ ) );
NAND3_X1 _12125_ ( .A1(_04462_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_04469_ ), .ZN(_04470_ ) );
AND3_X1 _12126_ ( .A1(_04452_ ), .A2(_04443_ ), .A3(_04444_ ), .ZN(_04471_ ) );
BUF_X4 _12127_ ( .A(_04471_ ), .Z(_04472_ ) );
BUF_X2 _12128_ ( .A(_04472_ ), .Z(_04473_ ) );
NOR3_X1 _12129_ ( .A1(_04448_ ), .A2(\ID_EX_csr [3] ), .A3(_04446_ ), .ZN(_04474_ ) );
BUF_X2 _12130_ ( .A(_04474_ ), .Z(_04475_ ) );
BUF_X4 _12131_ ( .A(_04475_ ), .Z(_04476_ ) );
NAND3_X1 _12132_ ( .A1(_04473_ ), .A2(\mtvec [30] ), .A3(_04476_ ), .ZN(_04477_ ) );
AND4_X1 _12133_ ( .A1(_04457_ ), .A2(_04465_ ), .A3(_04470_ ), .A4(_04477_ ), .ZN(_04478_ ) );
AOI21_X1 _12134_ ( .A(_04440_ ), .B1(_04451_ ), .B2(_04478_ ), .ZN(_04479_ ) );
OAI211_X1 _12135_ ( .A(_04403_ ), .B(_04406_ ), .C1(_04409_ ), .C2(_04479_ ), .ZN(_04480_ ) );
AND3_X1 _12136_ ( .A1(_03031_ ), .A2(_02128_ ), .A3(_03000_ ), .ZN(_04481_ ) );
BUF_X4 _12137_ ( .A(_04029_ ), .Z(_04482_ ) );
AND2_X1 _12138_ ( .A1(_02127_ ), .A2(_04482_ ), .ZN(_04483_ ) );
BUF_X4 _12139_ ( .A(_04483_ ), .Z(_04484_ ) );
BUF_X4 _12140_ ( .A(_04484_ ), .Z(_04485_ ) );
AOI21_X1 _12141_ ( .A(_04481_ ), .B1(_03223_ ), .B2(_04485_ ), .ZN(_04486_ ) );
AOI21_X1 _12142_ ( .A(_03086_ ), .B1(_04480_ ), .B2(_04486_ ), .ZN(_00122_ ) );
BUF_X4 _12143_ ( .A(_02127_ ), .Z(_04487_ ) );
BUF_X2 _12144_ ( .A(_04460_ ), .Z(_04488_ ) );
BUF_X4 _12145_ ( .A(_04449_ ), .Z(_04489_ ) );
NAND3_X1 _12146_ ( .A1(_04488_ ), .A2(\mepc [29] ), .A3(_04489_ ), .ZN(_04490_ ) );
BUF_X2 _12147_ ( .A(_04454_ ), .Z(_04491_ ) );
NAND4_X1 _12148_ ( .A1(_04453_ ), .A2(_04491_ ), .A3(\mycsreg.CSReg[0][29] ), .A4(_04444_ ), .ZN(_04492_ ) );
AND2_X1 _12149_ ( .A1(_04490_ ), .A2(_04492_ ), .ZN(_04493_ ) );
BUF_X2 _12150_ ( .A(_04467_ ), .Z(_04494_ ) );
NAND3_X1 _12151_ ( .A1(_04488_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_04494_ ), .ZN(_04495_ ) );
INV_X1 _12152_ ( .A(_04450_ ), .ZN(_04496_ ) );
BUF_X2 _12153_ ( .A(_04496_ ), .Z(_04497_ ) );
AND2_X1 _12154_ ( .A1(_04495_ ), .A2(_04497_ ), .ZN(_04498_ ) );
AND3_X1 _12155_ ( .A1(_04472_ ), .A2(\mtvec [29] ), .A3(_04475_ ), .ZN(_04499_ ) );
AND4_X1 _12156_ ( .A1(_04425_ ), .A2(_04437_ ), .A3(_04433_ ), .A4(_04413_ ), .ZN(_04500_ ) );
AND4_X2 _12157_ ( .A1(_04427_ ), .A2(_04500_ ), .A3(_04415_ ), .A4(_04432_ ), .ZN(_04501_ ) );
BUF_X2 _12158_ ( .A(_04501_ ), .Z(_04502_ ) );
AND4_X1 _12159_ ( .A1(_02173_ ), .A2(_04410_ ), .A3(_04436_ ), .A4(_04431_ ), .ZN(_04503_ ) );
XNOR2_X1 _12160_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_04504_ ) );
XNOR2_X1 _12161_ ( .A(fanout_net_6 ), .B(\ID_EX_csr [1] ), .ZN(_04505_ ) );
AND4_X1 _12162_ ( .A1(_04411_ ), .A2(_04434_ ), .A3(_04504_ ), .A4(_04505_ ), .ZN(_04506_ ) );
AND2_X2 _12163_ ( .A1(_04503_ ), .A2(_04506_ ), .ZN(_04507_ ) );
BUF_X2 _12164_ ( .A(_04507_ ), .Z(_04508_ ) );
AOI21_X1 _12165_ ( .A(_04499_ ), .B1(_04502_ ), .B2(_04508_ ), .ZN(_04509_ ) );
NAND3_X1 _12166_ ( .A1(_04493_ ), .A2(_04498_ ), .A3(_04509_ ), .ZN(_04510_ ) );
BUF_X2 _12167_ ( .A(_04507_ ), .Z(_04511_ ) );
INV_X1 _12168_ ( .A(\EX_LS_result_csreg_mem [29] ), .ZN(_04512_ ) );
BUF_X2 _12169_ ( .A(_04501_ ), .Z(_04513_ ) );
NAND3_X1 _12170_ ( .A1(_04511_ ), .A2(_04512_ ), .A3(_04513_ ), .ZN(_04514_ ) );
NAND2_X1 _12171_ ( .A1(_04510_ ), .A2(_04514_ ), .ZN(_04515_ ) );
AOI21_X1 _12172_ ( .A(_04487_ ), .B1(_04515_ ), .B2(\ID_EX_typ [3] ), .ZN(_04516_ ) );
AND4_X1 _12173_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_04517_ ) );
AND2_X1 _12174_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_04518_ ) );
AND4_X1 _12175_ ( .A1(\ID_EX_pc [13] ), .A2(_04517_ ), .A3(\ID_EX_pc [12] ), .A4(_04518_ ), .ZN(_04519_ ) );
AND2_X1 _12176_ ( .A1(_03093_ ), .A2(_04519_ ), .ZN(_04520_ ) );
AND4_X1 _12177_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_04521_ ) );
AND2_X1 _12178_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_04522_ ) );
AND4_X1 _12179_ ( .A1(\ID_EX_pc [21] ), .A2(_04521_ ), .A3(\ID_EX_pc [20] ), .A4(_04522_ ), .ZN(_04523_ ) );
AND2_X1 _12180_ ( .A1(_04520_ ), .A2(_04523_ ), .ZN(_04524_ ) );
NAND3_X1 _12181_ ( .A1(_04524_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_04525_ ) );
INV_X1 _12182_ ( .A(\ID_EX_pc [28] ), .ZN(_04526_ ) );
NOR2_X1 _12183_ ( .A1(_04525_ ), .A2(_04526_ ), .ZN(_04527_ ) );
XNOR2_X1 _12184_ ( .A(_04527_ ), .B(_03217_ ), .ZN(_04528_ ) );
NAND2_X1 _12185_ ( .A1(_03215_ ), .A2(_03216_ ), .ZN(_04529_ ) );
XNOR2_X1 _12186_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .ZN(_04530_ ) );
XOR2_X1 _12187_ ( .A(_04529_ ), .B(_04530_ ), .Z(_04531_ ) );
INV_X1 _12188_ ( .A(_04531_ ), .ZN(_04532_ ) );
MUX2_X1 _12189_ ( .A(_04528_ ), .B(_04532_ ), .S(_04401_ ), .Z(_04533_ ) );
OAI21_X1 _12190_ ( .A(_04516_ ), .B1(_04533_ ), .B2(\ID_EX_typ [3] ), .ZN(_04534_ ) );
OR2_X1 _12191_ ( .A1(_03067_ ), .A2(_02129_ ), .ZN(_04535_ ) );
AND2_X1 _12192_ ( .A1(_04534_ ), .A2(_04535_ ), .ZN(_04536_ ) );
INV_X1 _12193_ ( .A(_04484_ ), .ZN(_04537_ ) );
OR2_X1 _12194_ ( .A1(_04531_ ), .A2(_04537_ ), .ZN(_04538_ ) );
AOI21_X1 _12195_ ( .A(_03086_ ), .B1(_04536_ ), .B2(_04538_ ), .ZN(_00123_ ) );
NAND3_X1 _12196_ ( .A1(_03093_ ), .A2(_04519_ ), .A3(_04522_ ), .ZN(_04539_ ) );
XNOR2_X1 _12197_ ( .A(_04539_ ), .B(\ID_EX_pc [20] ), .ZN(_04540_ ) );
NOR2_X1 _12198_ ( .A1(_03168_ ), .A2(_03184_ ), .ZN(_04541_ ) );
INV_X1 _12199_ ( .A(_04541_ ), .ZN(_04542_ ) );
AND2_X1 _12200_ ( .A1(_04542_ ), .A2(_03124_ ), .ZN(_04543_ ) );
NOR2_X1 _12201_ ( .A1(_04543_ ), .A2(_03198_ ), .ZN(_04544_ ) );
XNOR2_X1 _12202_ ( .A(_04544_ ), .B(_03110_ ), .ZN(_04545_ ) );
MUX2_X1 _12203_ ( .A(_04540_ ), .B(_04545_ ), .S(_04401_ ), .Z(_04546_ ) );
OR2_X1 _12204_ ( .A1(_04546_ ), .A2(\ID_EX_typ [3] ), .ZN(_04547_ ) );
AND2_X2 _12205_ ( .A1(_04445_ ), .A2(_04467_ ), .ZN(_04548_ ) );
NOR2_X1 _12206_ ( .A1(_04450_ ), .A2(_04548_ ), .ZN(_04549_ ) );
NAND3_X1 _12207_ ( .A1(_04461_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_04468_ ), .ZN(_04550_ ) );
AND2_X1 _12208_ ( .A1(_04549_ ), .A2(_04550_ ), .ZN(_04551_ ) );
BUF_X4 _12209_ ( .A(_04460_ ), .Z(_04552_ ) );
NAND3_X1 _12210_ ( .A1(_04552_ ), .A2(\mepc [20] ), .A3(_04463_ ), .ZN(_04553_ ) );
BUF_X2 _12211_ ( .A(_04471_ ), .Z(_04554_ ) );
NAND3_X1 _12212_ ( .A1(_04554_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_04455_ ), .ZN(_04555_ ) );
AND2_X1 _12213_ ( .A1(_04553_ ), .A2(_04555_ ), .ZN(_04556_ ) );
CLKBUF_X2 _12214_ ( .A(_04471_ ), .Z(_04557_ ) );
AND3_X1 _12215_ ( .A1(_04557_ ), .A2(\mtvec [20] ), .A3(_04475_ ), .ZN(_04558_ ) );
AOI21_X1 _12216_ ( .A(_04558_ ), .B1(_04502_ ), .B2(_04507_ ), .ZN(_04559_ ) );
NAND3_X1 _12217_ ( .A1(_04551_ ), .A2(_04556_ ), .A3(_04559_ ), .ZN(_04560_ ) );
INV_X1 _12218_ ( .A(\EX_LS_result_csreg_mem [20] ), .ZN(_04561_ ) );
NAND3_X1 _12219_ ( .A1(_04511_ ), .A2(_04561_ ), .A3(_04513_ ), .ZN(_04562_ ) );
AND2_X1 _12220_ ( .A1(_04560_ ), .A2(_04562_ ), .ZN(_04563_ ) );
OAI211_X1 _12221_ ( .A(_04547_ ), .B(_04406_ ), .C1(_04409_ ), .C2(_04563_ ), .ZN(_04564_ ) );
AND3_X1 _12222_ ( .A1(_03040_ ), .A2(_02128_ ), .A3(_03037_ ), .ZN(_04565_ ) );
BUF_X4 _12223_ ( .A(_04484_ ), .Z(_04566_ ) );
AOI21_X1 _12224_ ( .A(_04565_ ), .B1(_04566_ ), .B2(_04545_ ), .ZN(_04567_ ) );
AOI21_X1 _12225_ ( .A(_03086_ ), .B1(_04564_ ), .B2(_04567_ ), .ZN(_00124_ ) );
BUF_X4 _12226_ ( .A(_04401_ ), .Z(_04568_ ) );
OAI21_X1 _12227_ ( .A(_03118_ ), .B1(_03168_ ), .B2(_03184_ ), .ZN(_04569_ ) );
AND2_X1 _12228_ ( .A1(_04569_ ), .A2(_03196_ ), .ZN(_04570_ ) );
NOR3_X1 _12229_ ( .A1(_04570_ ), .A2(_03120_ ), .A3(_03121_ ), .ZN(_04571_ ) );
NOR2_X1 _12230_ ( .A1(_04571_ ), .A2(_03120_ ), .ZN(_04572_ ) );
XNOR2_X1 _12231_ ( .A(_04572_ ), .B(_03119_ ), .ZN(_04573_ ) );
AOI21_X1 _12232_ ( .A(\ID_EX_typ [3] ), .B1(_04568_ ), .B2(_04573_ ), .ZN(_04574_ ) );
NAND3_X1 _12233_ ( .A1(_03093_ ), .A2(\ID_EX_pc [18] ), .A3(_04519_ ), .ZN(_04575_ ) );
INV_X1 _12234_ ( .A(\ID_EX_pc [19] ), .ZN(_04576_ ) );
XNOR2_X1 _12235_ ( .A(_04575_ ), .B(_04576_ ), .ZN(_04577_ ) );
OAI21_X1 _12236_ ( .A(_04574_ ), .B1(_04568_ ), .B2(_04577_ ), .ZN(_04578_ ) );
INV_X2 _12237_ ( .A(_04441_ ), .ZN(_04579_ ) );
BUF_X4 _12238_ ( .A(_04552_ ), .Z(_04580_ ) );
NAND3_X1 _12239_ ( .A1(_04580_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_04469_ ), .ZN(_04581_ ) );
BUF_X4 _12240_ ( .A(_04472_ ), .Z(_04582_ ) );
NAND3_X1 _12241_ ( .A1(_04582_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_04491_ ), .ZN(_04583_ ) );
NAND3_X1 _12242_ ( .A1(_04582_ ), .A2(\mtvec [19] ), .A3(_04476_ ), .ZN(_04584_ ) );
NAND3_X1 _12243_ ( .A1(_04581_ ), .A2(_04583_ ), .A3(_04584_ ), .ZN(_04585_ ) );
NAND3_X1 _12244_ ( .A1(_04580_ ), .A2(\mepc [19] ), .A3(_04489_ ), .ZN(_04586_ ) );
INV_X1 _12245_ ( .A(_04548_ ), .ZN(_04587_ ) );
BUF_X4 _12246_ ( .A(_04587_ ), .Z(_04588_ ) );
NAND2_X1 _12247_ ( .A1(_04586_ ), .A2(_04588_ ), .ZN(_04589_ ) );
OAI21_X1 _12248_ ( .A(_04579_ ), .B1(_04585_ ), .B2(_04589_ ), .ZN(_04590_ ) );
BUF_X2 _12249_ ( .A(_04428_ ), .Z(_04591_ ) );
BUF_X2 _12250_ ( .A(_04438_ ), .Z(_04592_ ) );
NAND3_X1 _12251_ ( .A1(_04591_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_04592_ ), .ZN(_04593_ ) );
AND2_X1 _12252_ ( .A1(_04590_ ), .A2(_04593_ ), .ZN(_04594_ ) );
INV_X1 _12253_ ( .A(_04594_ ), .ZN(_04595_ ) );
OAI211_X1 _12254_ ( .A(_04578_ ), .B(_04406_ ), .C1(_04409_ ), .C2(_04595_ ), .ZN(_04596_ ) );
NOR2_X1 _12255_ ( .A1(_03046_ ), .A2(_02130_ ), .ZN(_04597_ ) );
AOI21_X1 _12256_ ( .A(_04597_ ), .B1(_04566_ ), .B2(_04573_ ), .ZN(_04598_ ) );
AOI21_X1 _12257_ ( .A(_03086_ ), .B1(_04596_ ), .B2(_04598_ ), .ZN(_00125_ ) );
BUF_X4 _12258_ ( .A(_04407_ ), .Z(_04599_ ) );
BUF_X4 _12259_ ( .A(_04397_ ), .Z(_04600_ ) );
BUF_X4 _12260_ ( .A(_04399_ ), .Z(_04601_ ) );
XNOR2_X1 _12261_ ( .A(_04570_ ), .B(_03122_ ), .ZN(_04602_ ) );
NAND3_X1 _12262_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_04602_ ), .ZN(_04603_ ) );
XNOR2_X1 _12263_ ( .A(_04520_ ), .B(\ID_EX_pc [18] ), .ZN(_04604_ ) );
OAI211_X1 _12264_ ( .A(_04599_ ), .B(_04603_ ), .C1(_04568_ ), .C2(_04604_ ), .ZN(_04605_ ) );
BUF_X4 _12265_ ( .A(_04405_ ), .Z(_04606_ ) );
NAND3_X1 _12266_ ( .A1(_04580_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_04469_ ), .ZN(_04607_ ) );
NAND3_X1 _12267_ ( .A1(_04582_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_04491_ ), .ZN(_04608_ ) );
NAND3_X1 _12268_ ( .A1(_04582_ ), .A2(\mtvec [18] ), .A3(_04476_ ), .ZN(_04609_ ) );
NAND3_X1 _12269_ ( .A1(_04607_ ), .A2(_04608_ ), .A3(_04609_ ), .ZN(_04610_ ) );
BUF_X4 _12270_ ( .A(_04552_ ), .Z(_04611_ ) );
NAND3_X1 _12271_ ( .A1(_04611_ ), .A2(\mepc [18] ), .A3(_04489_ ), .ZN(_04612_ ) );
NAND2_X1 _12272_ ( .A1(_04612_ ), .A2(_04588_ ), .ZN(_04613_ ) );
OAI21_X1 _12273_ ( .A(_04579_ ), .B1(_04610_ ), .B2(_04613_ ), .ZN(_04614_ ) );
NAND3_X1 _12274_ ( .A1(_04591_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_04592_ ), .ZN(_04615_ ) );
AND2_X1 _12275_ ( .A1(_04614_ ), .A2(_04615_ ), .ZN(_04616_ ) );
INV_X1 _12276_ ( .A(_04616_ ), .ZN(_04617_ ) );
OAI211_X1 _12277_ ( .A(_04605_ ), .B(_04606_ ), .C1(_04409_ ), .C2(_04617_ ), .ZN(_04618_ ) );
NOR3_X1 _12278_ ( .A1(_03047_ ), .A2(_03044_ ), .A3(_02129_ ), .ZN(_04619_ ) );
AOI21_X1 _12279_ ( .A(_04619_ ), .B1(_04566_ ), .B2(_04602_ ), .ZN(_04620_ ) );
AOI21_X1 _12280_ ( .A(_03086_ ), .B1(_04618_ ), .B2(_04620_ ), .ZN(_00126_ ) );
AND3_X1 _12281_ ( .A1(_04518_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_04621_ ) );
NAND2_X1 _12282_ ( .A1(_03093_ ), .A2(_04621_ ), .ZN(_04622_ ) );
INV_X1 _12283_ ( .A(\ID_EX_pc [15] ), .ZN(_04623_ ) );
INV_X1 _12284_ ( .A(\ID_EX_pc [14] ), .ZN(_04624_ ) );
NOR3_X1 _12285_ ( .A1(_04622_ ), .A2(_04623_ ), .A3(_04624_ ), .ZN(_04625_ ) );
NAND2_X1 _12286_ ( .A1(_04625_ ), .A2(\ID_EX_pc [16] ), .ZN(_04626_ ) );
INV_X1 _12287_ ( .A(\ID_EX_pc [17] ), .ZN(_04627_ ) );
XNOR2_X1 _12288_ ( .A(_04626_ ), .B(_04627_ ), .ZN(_04628_ ) );
AND2_X1 _12289_ ( .A1(_04542_ ), .A2(_03116_ ), .ZN(_04629_ ) );
NOR2_X1 _12290_ ( .A1(_04629_ ), .A2(_03194_ ), .ZN(_04630_ ) );
XOR2_X1 _12291_ ( .A(_04630_ ), .B(_03117_ ), .Z(_04631_ ) );
MUX2_X1 _12292_ ( .A(_04628_ ), .B(_04631_ ), .S(_04401_ ), .Z(_04632_ ) );
NAND2_X1 _12293_ ( .A1(_04632_ ), .A2(_04599_ ), .ZN(_04633_ ) );
NAND3_X1 _12294_ ( .A1(_04488_ ), .A2(\mepc [17] ), .A3(_04463_ ), .ZN(_04634_ ) );
NAND3_X1 _12295_ ( .A1(_04461_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_04494_ ), .ZN(_04635_ ) );
BUF_X2 _12296_ ( .A(_04474_ ), .Z(_04636_ ) );
NAND3_X1 _12297_ ( .A1(_04554_ ), .A2(\mtvec [17] ), .A3(_04636_ ), .ZN(_04637_ ) );
NAND4_X1 _12298_ ( .A1(_04549_ ), .A2(_04634_ ), .A3(_04635_ ), .A4(_04637_ ), .ZN(_04638_ ) );
AND2_X1 _12299_ ( .A1(_04501_ ), .A2(_04507_ ), .ZN(_04639_ ) );
BUF_X2 _12300_ ( .A(_04557_ ), .Z(_04640_ ) );
AND3_X1 _12301_ ( .A1(_04640_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_04455_ ), .ZN(_04641_ ) );
NOR3_X1 _12302_ ( .A1(_04638_ ), .A2(_04639_ ), .A3(_04641_ ), .ZN(_04642_ ) );
INV_X1 _12303_ ( .A(\EX_LS_result_csreg_mem [17] ), .ZN(_04643_ ) );
AND3_X1 _12304_ ( .A1(_04508_ ), .A2(_04643_ ), .A3(_04502_ ), .ZN(_04644_ ) );
NOR2_X1 _12305_ ( .A1(_04642_ ), .A2(_04644_ ), .ZN(_04645_ ) );
OAI211_X1 _12306_ ( .A(_04633_ ), .B(_04606_ ), .C1(_04409_ ), .C2(_04645_ ), .ZN(_04646_ ) );
NOR2_X1 _12307_ ( .A1(_03051_ ), .A2(_02130_ ), .ZN(_04647_ ) );
NOR2_X1 _12308_ ( .A1(_04631_ ), .A2(_04537_ ), .ZN(_04648_ ) );
NOR2_X1 _12309_ ( .A1(_04647_ ), .A2(_04648_ ), .ZN(_04649_ ) );
AOI21_X1 _12310_ ( .A(_03086_ ), .B1(_04646_ ), .B2(_04649_ ), .ZN(_00127_ ) );
INV_X1 _12311_ ( .A(\ID_EX_pc [16] ), .ZN(_04650_ ) );
XNOR2_X1 _12312_ ( .A(_04625_ ), .B(_04650_ ), .ZN(_04651_ ) );
XNOR2_X1 _12313_ ( .A(_04541_ ), .B(_03116_ ), .ZN(_04652_ ) );
MUX2_X1 _12314_ ( .A(_04651_ ), .B(_04652_ ), .S(_04401_ ), .Z(_04653_ ) );
OR2_X1 _12315_ ( .A1(_04653_ ), .A2(\ID_EX_typ [3] ), .ZN(_04654_ ) );
NAND3_X1 _12316_ ( .A1(_04472_ ), .A2(\mtvec [16] ), .A3(_04475_ ), .ZN(_04655_ ) );
NAND3_X1 _12317_ ( .A1(_04552_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_04468_ ), .ZN(_04656_ ) );
AND3_X1 _12318_ ( .A1(_04549_ ), .A2(_04655_ ), .A3(_04656_ ), .ZN(_04657_ ) );
INV_X1 _12319_ ( .A(_04639_ ), .ZN(_04658_ ) );
NAND3_X1 _12320_ ( .A1(_04552_ ), .A2(\mepc [16] ), .A3(_04463_ ), .ZN(_04659_ ) );
AND3_X1 _12321_ ( .A1(_04557_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_04454_ ), .ZN(_04660_ ) );
INV_X1 _12322_ ( .A(_04660_ ), .ZN(_04661_ ) );
AND2_X1 _12323_ ( .A1(_04659_ ), .A2(_04661_ ), .ZN(_04662_ ) );
NAND3_X1 _12324_ ( .A1(_04657_ ), .A2(_04658_ ), .A3(_04662_ ), .ZN(_04663_ ) );
INV_X1 _12325_ ( .A(\EX_LS_result_csreg_mem [16] ), .ZN(_04664_ ) );
NAND3_X1 _12326_ ( .A1(_04511_ ), .A2(_04664_ ), .A3(_04513_ ), .ZN(_04665_ ) );
AND2_X1 _12327_ ( .A1(_04663_ ), .A2(_04665_ ), .ZN(_04666_ ) );
OAI211_X1 _12328_ ( .A(_04654_ ), .B(_04606_ ), .C1(_04409_ ), .C2(_04666_ ), .ZN(_04667_ ) );
BUF_X4 _12329_ ( .A(_02128_ ), .Z(_04668_ ) );
AOI22_X1 _12330_ ( .A1(_03052_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04652_ ), .ZN(_04669_ ) );
AOI21_X1 _12331_ ( .A(_03086_ ), .B1(_04667_ ), .B2(_04669_ ), .ZN(_00128_ ) );
NAND3_X1 _12332_ ( .A1(_04591_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_04592_ ), .ZN(_04670_ ) );
NAND3_X1 _12333_ ( .A1(_04611_ ), .A2(\mepc [15] ), .A3(_04489_ ), .ZN(_04671_ ) );
NAND4_X1 _12334_ ( .A1(_04453_ ), .A2(_04491_ ), .A3(\mycsreg.CSReg[0][15] ), .A4(_04444_ ), .ZN(_04672_ ) );
NAND3_X1 _12335_ ( .A1(_04640_ ), .A2(\mtvec [15] ), .A3(_04636_ ), .ZN(_04673_ ) );
NAND3_X1 _12336_ ( .A1(_04671_ ), .A2(_04672_ ), .A3(_04673_ ), .ZN(_04674_ ) );
NAND3_X1 _12337_ ( .A1(_04611_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_04494_ ), .ZN(_04675_ ) );
NAND2_X1 _12338_ ( .A1(_04675_ ), .A2(_04587_ ), .ZN(_04676_ ) );
NOR2_X1 _12339_ ( .A1(_04674_ ), .A2(_04676_ ), .ZN(_04677_ ) );
OAI21_X1 _12340_ ( .A(_04670_ ), .B1(_04677_ ), .B2(_04441_ ), .ZN(_04678_ ) );
NAND3_X1 _12341_ ( .A1(_03093_ ), .A2(\ID_EX_pc [14] ), .A3(_04621_ ), .ZN(_04679_ ) );
XNOR2_X1 _12342_ ( .A(_04679_ ), .B(\ID_EX_pc [15] ), .ZN(_04680_ ) );
OAI211_X1 _12343_ ( .A(_03163_ ), .B(_03166_ ), .C1(_03151_ ), .C2(_03152_ ), .ZN(_04681_ ) );
NAND2_X1 _12344_ ( .A1(_04681_ ), .A2(_03182_ ), .ZN(_04682_ ) );
NAND2_X1 _12345_ ( .A1(_04682_ ), .A2(_03157_ ), .ZN(_04683_ ) );
NAND2_X1 _12346_ ( .A1(_04683_ ), .A2(_03174_ ), .ZN(_04684_ ) );
NAND2_X1 _12347_ ( .A1(_04684_ ), .A2(_03159_ ), .ZN(_04685_ ) );
NAND2_X1 _12348_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04686_ ) );
AND2_X1 _12349_ ( .A1(_04685_ ), .A2(_04686_ ), .ZN(_04687_ ) );
XNOR2_X1 _12350_ ( .A(_04687_ ), .B(_03158_ ), .ZN(_04688_ ) );
BUF_X8 _12351_ ( .A(_04400_ ), .Z(_04689_ ) );
MUX2_X1 _12352_ ( .A(_04680_ ), .B(_04688_ ), .S(_04689_ ), .Z(_04690_ ) );
MUX2_X1 _12353_ ( .A(_04678_ ), .B(_04690_ ), .S(_04408_ ), .Z(_04691_ ) );
NAND2_X1 _12354_ ( .A1(_04691_ ), .A2(_04406_ ), .ZN(_04692_ ) );
NOR2_X1 _12355_ ( .A1(_03060_ ), .A2(_02130_ ), .ZN(_04693_ ) );
AOI21_X1 _12356_ ( .A(_04693_ ), .B1(_04566_ ), .B2(_04688_ ), .ZN(_04694_ ) );
AOI21_X1 _12357_ ( .A(_03086_ ), .B1(_04692_ ), .B2(_04694_ ), .ZN(_00129_ ) );
BUF_X4 _12358_ ( .A(_03085_ ), .Z(_04695_ ) );
XOR2_X1 _12359_ ( .A(_04684_ ), .B(_03159_ ), .Z(_04696_ ) );
NAND3_X1 _12360_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_04696_ ), .ZN(_04697_ ) );
XNOR2_X1 _12361_ ( .A(_04622_ ), .B(_04624_ ), .ZN(_04698_ ) );
OAI211_X1 _12362_ ( .A(_04599_ ), .B(_04697_ ), .C1(_04568_ ), .C2(_04698_ ), .ZN(_04699_ ) );
NAND3_X1 _12363_ ( .A1(_04472_ ), .A2(\mtvec [14] ), .A3(_04475_ ), .ZN(_04700_ ) );
NAND3_X1 _12364_ ( .A1(_04552_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_04468_ ), .ZN(_04701_ ) );
AND3_X1 _12365_ ( .A1(_04549_ ), .A2(_04700_ ), .A3(_04701_ ), .ZN(_04702_ ) );
NAND3_X1 _12366_ ( .A1(_04552_ ), .A2(\mepc [14] ), .A3(_04463_ ), .ZN(_04703_ ) );
AND3_X1 _12367_ ( .A1(_04557_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_04454_ ), .ZN(_04704_ ) );
INV_X1 _12368_ ( .A(_04704_ ), .ZN(_04705_ ) );
AND2_X1 _12369_ ( .A1(_04703_ ), .A2(_04705_ ), .ZN(_04706_ ) );
NAND3_X1 _12370_ ( .A1(_04702_ ), .A2(_04658_ ), .A3(_04706_ ), .ZN(_04707_ ) );
INV_X1 _12371_ ( .A(\EX_LS_result_csreg_mem [14] ), .ZN(_04708_ ) );
NAND3_X1 _12372_ ( .A1(_04508_ ), .A2(_04708_ ), .A3(_04513_ ), .ZN(_04709_ ) );
AND2_X1 _12373_ ( .A1(_04707_ ), .A2(_04709_ ), .ZN(_04710_ ) );
OAI211_X1 _12374_ ( .A(_04699_ ), .B(_04606_ ), .C1(_04409_ ), .C2(_04710_ ), .ZN(_04711_ ) );
AND3_X1 _12375_ ( .A1(_03061_ ), .A2(_02128_ ), .A3(_03057_ ), .ZN(_04712_ ) );
AOI21_X1 _12376_ ( .A(_04712_ ), .B1(_04566_ ), .B2(_04696_ ), .ZN(_04713_ ) );
AOI21_X1 _12377_ ( .A(_04695_ ), .B1(_04711_ ), .B2(_04713_ ), .ZN(_00130_ ) );
NAND3_X1 _12378_ ( .A1(_03092_ ), .A2(\ID_EX_pc [9] ), .A3(_04518_ ), .ZN(_04714_ ) );
INV_X1 _12379_ ( .A(\ID_EX_pc [12] ), .ZN(_04715_ ) );
NOR2_X1 _12380_ ( .A1(_04714_ ), .A2(_04715_ ), .ZN(_04716_ ) );
INV_X1 _12381_ ( .A(\ID_EX_pc [13] ), .ZN(_04717_ ) );
XNOR2_X1 _12382_ ( .A(_04716_ ), .B(_04717_ ), .ZN(_04718_ ) );
NAND2_X1 _12383_ ( .A1(_04682_ ), .A2(_03154_ ), .ZN(_04719_ ) );
NAND2_X1 _12384_ ( .A1(_04719_ ), .A2(_03172_ ), .ZN(_04720_ ) );
XNOR2_X1 _12385_ ( .A(_04720_ ), .B(_03156_ ), .ZN(_04721_ ) );
MUX2_X1 _12386_ ( .A(_04718_ ), .B(_04721_ ), .S(_04689_ ), .Z(_04722_ ) );
OR2_X1 _12387_ ( .A1(_04722_ ), .A2(\ID_EX_typ [3] ), .ZN(_04723_ ) );
BUF_X4 _12388_ ( .A(_04579_ ), .Z(_04724_ ) );
BUF_X2 _12389_ ( .A(_04497_ ), .Z(_04725_ ) );
AND3_X1 _12390_ ( .A1(_04473_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_04456_ ), .ZN(_04726_ ) );
AND3_X1 _12391_ ( .A1(_04557_ ), .A2(\mtvec [13] ), .A3(_04475_ ), .ZN(_04727_ ) );
NOR2_X1 _12392_ ( .A1(_04726_ ), .A2(_04727_ ), .ZN(_04728_ ) );
NAND3_X1 _12393_ ( .A1(_04461_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_04468_ ), .ZN(_04729_ ) );
NAND3_X1 _12394_ ( .A1(_04461_ ), .A2(\mepc [13] ), .A3(_04463_ ), .ZN(_04730_ ) );
AND2_X1 _12395_ ( .A1(_04729_ ), .A2(_04730_ ), .ZN(_04731_ ) );
NAND4_X1 _12396_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04728_ ), .A4(_04731_ ), .ZN(_04732_ ) );
INV_X1 _12397_ ( .A(\EX_LS_result_csreg_mem [13] ), .ZN(_04733_ ) );
NAND3_X1 _12398_ ( .A1(_04429_ ), .A2(_04733_ ), .A3(_04439_ ), .ZN(_04734_ ) );
AND2_X1 _12399_ ( .A1(_04732_ ), .A2(_04734_ ), .ZN(_04735_ ) );
OAI211_X1 _12400_ ( .A(_04723_ ), .B(_04606_ ), .C1(_04409_ ), .C2(_04735_ ), .ZN(_04736_ ) );
NOR2_X1 _12401_ ( .A1(_03064_ ), .A2(_02129_ ), .ZN(_04737_ ) );
AOI21_X1 _12402_ ( .A(_04737_ ), .B1(_04566_ ), .B2(_04721_ ), .ZN(_04738_ ) );
AOI21_X1 _12403_ ( .A(_04695_ ), .B1(_04736_ ), .B2(_04738_ ), .ZN(_00131_ ) );
XNOR2_X1 _12404_ ( .A(_04714_ ), .B(\ID_EX_pc [12] ), .ZN(_04739_ ) );
XNOR2_X1 _12405_ ( .A(_04682_ ), .B(_03155_ ), .ZN(_04740_ ) );
MUX2_X1 _12406_ ( .A(_04739_ ), .B(_04740_ ), .S(_04401_ ), .Z(_04741_ ) );
AND2_X1 _12407_ ( .A1(_04741_ ), .A2(_04408_ ), .ZN(_04742_ ) );
NAND4_X1 _12408_ ( .A1(_04453_ ), .A2(_04455_ ), .A3(\mycsreg.CSReg[0][12] ), .A4(_04444_ ), .ZN(_04743_ ) );
NAND3_X1 _12409_ ( .A1(_04460_ ), .A2(\mepc [12] ), .A3(_04449_ ), .ZN(_04744_ ) );
NAND3_X1 _12410_ ( .A1(_04460_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_04467_ ), .ZN(_04745_ ) );
NAND3_X1 _12411_ ( .A1(_04557_ ), .A2(\mtvec [12] ), .A3(_04474_ ), .ZN(_04746_ ) );
AND4_X1 _12412_ ( .A1(_04743_ ), .A2(_04744_ ), .A3(_04745_ ), .A4(_04746_ ), .ZN(_04747_ ) );
NAND4_X1 _12413_ ( .A1(_04579_ ), .A2(_04497_ ), .A3(_04587_ ), .A4(_04747_ ), .ZN(_04748_ ) );
INV_X1 _12414_ ( .A(\EX_LS_result_csreg_mem [12] ), .ZN(_04749_ ) );
NAND3_X1 _12415_ ( .A1(_04428_ ), .A2(_04749_ ), .A3(_04438_ ), .ZN(_04750_ ) );
AND3_X1 _12416_ ( .A1(_04748_ ), .A2(\ID_EX_typ [3] ), .A3(_04750_ ), .ZN(_04751_ ) );
OAI21_X1 _12417_ ( .A(_04406_ ), .B1(_04742_ ), .B2(_04751_ ), .ZN(_04752_ ) );
AOI22_X1 _12418_ ( .A1(_03065_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04740_ ), .ZN(_04753_ ) );
AOI21_X1 _12419_ ( .A(_04695_ ), .B1(_04752_ ), .B2(_04753_ ), .ZN(_00132_ ) );
AND2_X1 _12420_ ( .A1(_03093_ ), .A2(\ID_EX_pc [10] ), .ZN(_04754_ ) );
XNOR2_X1 _12421_ ( .A(_04754_ ), .B(_03176_ ), .ZN(_04755_ ) );
OAI21_X1 _12422_ ( .A(_03166_ ), .B1(_03151_ ), .B2(_03152_ ), .ZN(_04756_ ) );
NAND2_X1 _12423_ ( .A1(_04756_ ), .A2(_03180_ ), .ZN(_04757_ ) );
NAND2_X1 _12424_ ( .A1(_04757_ ), .A2(_03162_ ), .ZN(_04758_ ) );
NAND2_X1 _12425_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_04759_ ) );
AND2_X1 _12426_ ( .A1(_04758_ ), .A2(_04759_ ), .ZN(_04760_ ) );
XNOR2_X1 _12427_ ( .A(_04760_ ), .B(_03161_ ), .ZN(_04761_ ) );
MUX2_X1 _12428_ ( .A(_04755_ ), .B(_04761_ ), .S(_04689_ ), .Z(_04762_ ) );
OR2_X1 _12429_ ( .A1(_04762_ ), .A2(\ID_EX_typ [3] ), .ZN(_04763_ ) );
NAND3_X1 _12430_ ( .A1(_04611_ ), .A2(\mepc [11] ), .A3(_04489_ ), .ZN(_04764_ ) );
NAND4_X1 _12431_ ( .A1(_04453_ ), .A2(_04491_ ), .A3(\mycsreg.CSReg[0][11] ), .A4(_04444_ ), .ZN(_04765_ ) );
NAND2_X1 _12432_ ( .A1(_04764_ ), .A2(_04765_ ), .ZN(_04766_ ) );
AND3_X1 _12433_ ( .A1(_04488_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_04494_ ), .ZN(_04767_ ) );
AND3_X1 _12434_ ( .A1(_04640_ ), .A2(\mtvec [11] ), .A3(_04636_ ), .ZN(_04768_ ) );
NOR3_X1 _12435_ ( .A1(_04766_ ), .A2(_04767_ ), .A3(_04768_ ), .ZN(_04769_ ) );
NAND4_X1 _12436_ ( .A1(_04579_ ), .A2(_04497_ ), .A3(_04588_ ), .A4(_04769_ ), .ZN(_04770_ ) );
INV_X1 _12437_ ( .A(\EX_LS_result_csreg_mem [11] ), .ZN(_04771_ ) );
NAND3_X1 _12438_ ( .A1(_04429_ ), .A2(_04771_ ), .A3(_04439_ ), .ZN(_04772_ ) );
AND2_X1 _12439_ ( .A1(_04770_ ), .A2(_04772_ ), .ZN(_04773_ ) );
OAI211_X1 _12440_ ( .A(_04763_ ), .B(_04606_ ), .C1(_04409_ ), .C2(_04773_ ), .ZN(_04774_ ) );
NAND2_X1 _12441_ ( .A1(_02917_ ), .A2(_02925_ ), .ZN(_04775_ ) );
AOI21_X1 _12442_ ( .A(_02930_ ), .B1(_04775_ ), .B2(_02673_ ), .ZN(_04776_ ) );
NOR2_X1 _12443_ ( .A1(_02718_ ), .A2(\ID_EX_imm [10] ), .ZN(_04777_ ) );
NOR3_X1 _12444_ ( .A1(_04776_ ), .A2(_02932_ ), .A3(_04777_ ), .ZN(_04778_ ) );
NOR2_X1 _12445_ ( .A1(_04778_ ), .A2(_02932_ ), .ZN(_04779_ ) );
XNOR2_X1 _12446_ ( .A(_04779_ ), .B(_02696_ ), .ZN(_04780_ ) );
AOI22_X1 _12447_ ( .A1(_04780_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04761_ ), .ZN(_04781_ ) );
AOI21_X1 _12448_ ( .A(_04695_ ), .B1(_04774_ ), .B2(_04781_ ), .ZN(_00133_ ) );
XNOR2_X1 _12449_ ( .A(_04525_ ), .B(\ID_EX_pc [28] ), .ZN(_04782_ ) );
XOR2_X1 _12450_ ( .A(_03213_ ), .B(_03214_ ), .Z(_04783_ ) );
MUX2_X1 _12451_ ( .A(_04782_ ), .B(_04783_ ), .S(_04689_ ), .Z(_04784_ ) );
OR2_X1 _12452_ ( .A1(_04784_ ), .A2(\ID_EX_typ [3] ), .ZN(_04785_ ) );
BUF_X4 _12453_ ( .A(_04408_ ), .Z(_04786_ ) );
NAND3_X1 _12454_ ( .A1(_04461_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_04468_ ), .ZN(_04787_ ) );
NAND3_X1 _12455_ ( .A1(_04554_ ), .A2(\mtvec [28] ), .A3(_04636_ ), .ZN(_04788_ ) );
AND3_X1 _12456_ ( .A1(_04787_ ), .A2(_04496_ ), .A3(_04788_ ), .ZN(_04789_ ) );
NAND3_X1 _12457_ ( .A1(_04580_ ), .A2(\mepc [28] ), .A3(_04464_ ), .ZN(_04790_ ) );
NAND3_X1 _12458_ ( .A1(_04473_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_04456_ ), .ZN(_04791_ ) );
NAND4_X1 _12459_ ( .A1(_04658_ ), .A2(_04789_ ), .A3(_04790_ ), .A4(_04791_ ), .ZN(_04792_ ) );
INV_X1 _12460_ ( .A(\EX_LS_result_csreg_mem [28] ), .ZN(_04793_ ) );
NAND3_X1 _12461_ ( .A1(_04511_ ), .A2(_04793_ ), .A3(_04513_ ), .ZN(_04794_ ) );
AND2_X1 _12462_ ( .A1(_04792_ ), .A2(_04794_ ), .ZN(_04795_ ) );
OAI211_X1 _12463_ ( .A(_04785_ ), .B(_04606_ ), .C1(_04786_ ), .C2(_04795_ ), .ZN(_04796_ ) );
NOR3_X1 _12464_ ( .A1(_03068_ ), .A2(_02970_ ), .A3(_02129_ ), .ZN(_04797_ ) );
AOI21_X1 _12465_ ( .A(_04797_ ), .B1(_04566_ ), .B2(_04783_ ), .ZN(_04798_ ) );
AOI21_X1 _12466_ ( .A(_04695_ ), .B1(_04796_ ), .B2(_04798_ ), .ZN(_00134_ ) );
XOR2_X1 _12467_ ( .A(_04757_ ), .B(_03162_ ), .Z(_04799_ ) );
NAND3_X1 _12468_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_04799_ ), .ZN(_04800_ ) );
XNOR2_X1 _12469_ ( .A(_03093_ ), .B(\ID_EX_pc [10] ), .ZN(_04801_ ) );
OAI211_X1 _12470_ ( .A(_04599_ ), .B(_04800_ ), .C1(_04568_ ), .C2(_04801_ ), .ZN(_04802_ ) );
NAND3_X1 _12471_ ( .A1(_04580_ ), .A2(\mepc [10] ), .A3(_04464_ ), .ZN(_04803_ ) );
NAND4_X1 _12472_ ( .A1(_04453_ ), .A2(_04491_ ), .A3(\mycsreg.CSReg[0][10] ), .A4(_04444_ ), .ZN(_04804_ ) );
NAND3_X1 _12473_ ( .A1(_04640_ ), .A2(\mtvec [10] ), .A3(_04476_ ), .ZN(_04805_ ) );
NAND3_X1 _12474_ ( .A1(_04803_ ), .A2(_04804_ ), .A3(_04805_ ), .ZN(_04806_ ) );
NAND3_X1 _12475_ ( .A1(_04611_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_04469_ ), .ZN(_04807_ ) );
NAND2_X1 _12476_ ( .A1(_04807_ ), .A2(_04588_ ), .ZN(_04808_ ) );
OAI21_X1 _12477_ ( .A(_04579_ ), .B1(_04806_ ), .B2(_04808_ ), .ZN(_04809_ ) );
NAND3_X1 _12478_ ( .A1(_04591_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_04592_ ), .ZN(_04810_ ) );
AND2_X1 _12479_ ( .A1(_04809_ ), .A2(_04810_ ), .ZN(_04811_ ) );
INV_X1 _12480_ ( .A(_04811_ ), .ZN(_04812_ ) );
OAI211_X1 _12481_ ( .A(_04802_ ), .B(_04606_ ), .C1(_04786_ ), .C2(_04812_ ), .ZN(_04813_ ) );
XNOR2_X1 _12482_ ( .A(_04776_ ), .B(_02719_ ), .ZN(_04814_ ) );
AOI22_X1 _12483_ ( .A1(_04814_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04799_ ), .ZN(_04815_ ) );
AOI21_X1 _12484_ ( .A(_04695_ ), .B1(_04813_ ), .B2(_04815_ ), .ZN(_00135_ ) );
OAI21_X1 _12485_ ( .A(_03164_ ), .B1(_03151_ ), .B2(_03152_ ), .ZN(_04816_ ) );
INV_X1 _12486_ ( .A(_03179_ ), .ZN(_04817_ ) );
AND2_X1 _12487_ ( .A1(_04816_ ), .A2(_04817_ ), .ZN(_04818_ ) );
XNOR2_X1 _12488_ ( .A(_04818_ ), .B(_03165_ ), .ZN(_04819_ ) );
NAND3_X1 _12489_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_04819_ ), .ZN(_04820_ ) );
XNOR2_X1 _12490_ ( .A(_03092_ ), .B(\ID_EX_pc [9] ), .ZN(_04821_ ) );
OAI211_X1 _12491_ ( .A(_04599_ ), .B(_04820_ ), .C1(_04568_ ), .C2(_04821_ ), .ZN(_04822_ ) );
AND3_X1 _12492_ ( .A1(_04554_ ), .A2(\mtvec [9] ), .A3(_04636_ ), .ZN(_04823_ ) );
NOR2_X1 _12493_ ( .A1(_04823_ ), .A2(_04548_ ), .ZN(_04824_ ) );
NAND3_X1 _12494_ ( .A1(_04580_ ), .A2(\mepc [9] ), .A3(_04464_ ), .ZN(_04825_ ) );
NAND3_X1 _12495_ ( .A1(_04580_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_04469_ ), .ZN(_04826_ ) );
NAND3_X1 _12496_ ( .A1(_04473_ ), .A2(\mycsreg.CSReg[0][9] ), .A3(_04456_ ), .ZN(_04827_ ) );
NAND4_X1 _12497_ ( .A1(_04824_ ), .A2(_04825_ ), .A3(_04826_ ), .A4(_04827_ ), .ZN(_04828_ ) );
NAND2_X1 _12498_ ( .A1(_04579_ ), .A2(_04828_ ), .ZN(_04829_ ) );
AND3_X1 _12499_ ( .A1(_04428_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_04438_ ), .ZN(_04830_ ) );
INV_X1 _12500_ ( .A(_04830_ ), .ZN(_04831_ ) );
AND2_X1 _12501_ ( .A1(_04829_ ), .A2(_04831_ ), .ZN(_04832_ ) );
INV_X1 _12502_ ( .A(_04832_ ), .ZN(_04833_ ) );
OAI211_X1 _12503_ ( .A(_04822_ ), .B(_04606_ ), .C1(_04786_ ), .C2(_04833_ ), .ZN(_04834_ ) );
INV_X1 _12504_ ( .A(_02649_ ), .ZN(_04835_ ) );
AOI21_X1 _12505_ ( .A(_04835_ ), .B1(_02917_ ), .B2(_02925_ ), .ZN(_04836_ ) );
OR2_X1 _12506_ ( .A1(_04836_ ), .A2(_02927_ ), .ZN(_04837_ ) );
XNOR2_X1 _12507_ ( .A(_04837_ ), .B(_02672_ ), .ZN(_04838_ ) );
NOR2_X1 _12508_ ( .A1(_04838_ ), .A2(_02129_ ), .ZN(_04839_ ) );
AOI21_X1 _12509_ ( .A(_04839_ ), .B1(_04566_ ), .B2(_04819_ ), .ZN(_04840_ ) );
AOI21_X1 _12510_ ( .A(_04695_ ), .B1(_04834_ ), .B2(_04840_ ), .ZN(_00136_ ) );
INV_X1 _12511_ ( .A(\ID_EX_pc [8] ), .ZN(_04841_ ) );
XNOR2_X1 _12512_ ( .A(_03091_ ), .B(_04841_ ), .ZN(_04842_ ) );
XNOR2_X1 _12513_ ( .A(_03153_ ), .B(_03164_ ), .ZN(_04843_ ) );
MUX2_X1 _12514_ ( .A(_04842_ ), .B(_04843_ ), .S(_04689_ ), .Z(_04844_ ) );
OR2_X1 _12515_ ( .A1(_04844_ ), .A2(\ID_EX_typ [3] ), .ZN(_04845_ ) );
NAND3_X1 _12516_ ( .A1(_04472_ ), .A2(\mtvec [8] ), .A3(_04475_ ), .ZN(_04846_ ) );
NAND3_X1 _12517_ ( .A1(_04460_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_04468_ ), .ZN(_04847_ ) );
AND3_X1 _12518_ ( .A1(_04549_ ), .A2(_04846_ ), .A3(_04847_ ), .ZN(_04848_ ) );
NAND3_X1 _12519_ ( .A1(_04552_ ), .A2(\mepc [8] ), .A3(_04463_ ), .ZN(_04849_ ) );
AND3_X1 _12520_ ( .A1(_04557_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_04454_ ), .ZN(_04850_ ) );
INV_X1 _12521_ ( .A(_04850_ ), .ZN(_04851_ ) );
AND2_X1 _12522_ ( .A1(_04849_ ), .A2(_04851_ ), .ZN(_04852_ ) );
NAND3_X1 _12523_ ( .A1(_04848_ ), .A2(_04658_ ), .A3(_04852_ ), .ZN(_04853_ ) );
INV_X1 _12524_ ( .A(\EX_LS_result_csreg_mem [8] ), .ZN(_04854_ ) );
NAND3_X1 _12525_ ( .A1(_04508_ ), .A2(_04854_ ), .A3(_04502_ ), .ZN(_04855_ ) );
AND2_X1 _12526_ ( .A1(_04853_ ), .A2(_04855_ ), .ZN(_04856_ ) );
OAI211_X1 _12527_ ( .A(_04845_ ), .B(_04606_ ), .C1(_04786_ ), .C2(_04856_ ), .ZN(_04857_ ) );
XNOR2_X1 _12528_ ( .A(_04775_ ), .B(_04835_ ), .ZN(_04858_ ) );
AOI22_X1 _12529_ ( .A1(_04858_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04843_ ), .ZN(_04859_ ) );
AOI21_X1 _12530_ ( .A(_04695_ ), .B1(_04857_ ), .B2(_04859_ ), .ZN(_00137_ ) );
NOR2_X1 _12531_ ( .A1(_03152_ ), .A2(_03150_ ), .ZN(_04860_ ) );
XNOR2_X1 _12532_ ( .A(_03149_ ), .B(_04860_ ), .ZN(_04861_ ) );
NAND3_X1 _12533_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_04861_ ), .ZN(_04862_ ) );
XNOR2_X1 _12534_ ( .A(_03090_ ), .B(\ID_EX_pc [7] ), .ZN(_04863_ ) );
OAI211_X1 _12535_ ( .A(_04408_ ), .B(_04862_ ), .C1(_04568_ ), .C2(_04863_ ), .ZN(_04864_ ) );
BUF_X4 _12536_ ( .A(_04405_ ), .Z(_04865_ ) );
NAND3_X1 _12537_ ( .A1(_04611_ ), .A2(\mepc [7] ), .A3(_04489_ ), .ZN(_04866_ ) );
NAND3_X1 _12538_ ( .A1(_04640_ ), .A2(\mtvec [7] ), .A3(_04636_ ), .ZN(_04867_ ) );
AND2_X1 _12539_ ( .A1(_04866_ ), .A2(_04867_ ), .ZN(_04868_ ) );
NAND3_X1 _12540_ ( .A1(_04488_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_04494_ ), .ZN(_04869_ ) );
NAND3_X1 _12541_ ( .A1(_04640_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_04491_ ), .ZN(_04870_ ) );
AND2_X1 _12542_ ( .A1(_04869_ ), .A2(_04870_ ), .ZN(_04871_ ) );
AOI22_X1 _12543_ ( .A1(_04868_ ), .A2(_04871_ ), .B1(_04591_ ), .B2(_04592_ ), .ZN(_04872_ ) );
AND3_X1 _12544_ ( .A1(_04591_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_04592_ ), .ZN(_04873_ ) );
NOR2_X1 _12545_ ( .A1(_04872_ ), .A2(_04873_ ), .ZN(_04874_ ) );
INV_X1 _12546_ ( .A(_04874_ ), .ZN(_04875_ ) );
OAI211_X1 _12547_ ( .A(_04864_ ), .B(_04865_ ), .C1(_04786_ ), .C2(_04875_ ), .ZN(_04876_ ) );
NOR2_X1 _12548_ ( .A1(_02869_ ), .A2(_02924_ ), .ZN(_04877_ ) );
NOR2_X1 _12549_ ( .A1(_04877_ ), .A2(_02893_ ), .ZN(_04878_ ) );
AND2_X1 _12550_ ( .A1(_02890_ ), .A2(\ID_EX_imm [6] ), .ZN(_04879_ ) );
OR2_X1 _12551_ ( .A1(_04878_ ), .A2(_04879_ ), .ZN(_04880_ ) );
XNOR2_X1 _12552_ ( .A(_04880_ ), .B(_02915_ ), .ZN(_04881_ ) );
AOI22_X1 _12553_ ( .A1(_04881_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04861_ ), .ZN(_04882_ ) );
AOI21_X1 _12554_ ( .A(_04695_ ), .B1(_04876_ ), .B2(_04882_ ), .ZN(_00138_ ) );
INV_X1 _12555_ ( .A(\ID_EX_pc [6] ), .ZN(_04883_ ) );
XNOR2_X1 _12556_ ( .A(_03089_ ), .B(_04883_ ), .ZN(_04884_ ) );
XOR2_X1 _12557_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_04885_ ) );
XNOR2_X1 _12558_ ( .A(_03145_ ), .B(_04885_ ), .ZN(_04886_ ) );
MUX2_X1 _12559_ ( .A(_04884_ ), .B(_04886_ ), .S(_04689_ ), .Z(_04887_ ) );
OR2_X1 _12560_ ( .A1(_04887_ ), .A2(\ID_EX_typ [3] ), .ZN(_04888_ ) );
NAND3_X1 _12561_ ( .A1(_04552_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_04468_ ), .ZN(_04889_ ) );
AND2_X1 _12562_ ( .A1(_04889_ ), .A2(_04496_ ), .ZN(_04890_ ) );
NAND3_X1 _12563_ ( .A1(_04640_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_04491_ ), .ZN(_04891_ ) );
NAND3_X1 _12564_ ( .A1(_04488_ ), .A2(\mepc [6] ), .A3(_04489_ ), .ZN(_04892_ ) );
AND3_X1 _12565_ ( .A1(_04557_ ), .A2(\mtvec [6] ), .A3(_04474_ ), .ZN(_04893_ ) );
AOI21_X1 _12566_ ( .A(_04893_ ), .B1(_04501_ ), .B2(_04507_ ), .ZN(_04894_ ) );
NAND4_X1 _12567_ ( .A1(_04890_ ), .A2(_04891_ ), .A3(_04892_ ), .A4(_04894_ ), .ZN(_04895_ ) );
INV_X1 _12568_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_04896_ ) );
NAND3_X1 _12569_ ( .A1(_04508_ ), .A2(_04896_ ), .A3(_04502_ ), .ZN(_04897_ ) );
AND2_X1 _12570_ ( .A1(_04895_ ), .A2(_04897_ ), .ZN(_04898_ ) );
OAI211_X1 _12571_ ( .A(_04888_ ), .B(_04865_ ), .C1(_04786_ ), .C2(_04898_ ), .ZN(_04899_ ) );
XNOR2_X1 _12572_ ( .A(_04877_ ), .B(_02892_ ), .ZN(_04900_ ) );
AOI22_X1 _12573_ ( .A1(_04900_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04886_ ), .ZN(_04901_ ) );
AOI21_X1 _12574_ ( .A(_04695_ ), .B1(_04899_ ), .B2(_04901_ ), .ZN(_00139_ ) );
BUF_X4 _12575_ ( .A(_03085_ ), .Z(_04902_ ) );
NOR2_X1 _12576_ ( .A1(_03144_ ), .A2(_03142_ ), .ZN(_04903_ ) );
XNOR2_X1 _12577_ ( .A(_03141_ ), .B(_04903_ ), .ZN(_04904_ ) );
NAND3_X1 _12578_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_04904_ ), .ZN(_04905_ ) );
XNOR2_X1 _12579_ ( .A(_03088_ ), .B(\ID_EX_pc [5] ), .ZN(_04906_ ) );
OAI211_X1 _12580_ ( .A(_04408_ ), .B(_04905_ ), .C1(_04568_ ), .C2(_04906_ ), .ZN(_04907_ ) );
NAND3_X1 _12581_ ( .A1(_04488_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_04494_ ), .ZN(_04908_ ) );
NAND3_X1 _12582_ ( .A1(_04488_ ), .A2(\mepc [5] ), .A3(_04489_ ), .ZN(_04909_ ) );
AND3_X1 _12583_ ( .A1(_04640_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_04491_ ), .ZN(_04910_ ) );
INV_X1 _12584_ ( .A(_04910_ ), .ZN(_04911_ ) );
NAND3_X1 _12585_ ( .A1(_04640_ ), .A2(\mtvec [5] ), .A3(_04636_ ), .ZN(_04912_ ) );
NAND4_X1 _12586_ ( .A1(_04908_ ), .A2(_04909_ ), .A3(_04911_ ), .A4(_04912_ ), .ZN(_04913_ ) );
NOR3_X1 _12587_ ( .A1(_04441_ ), .A2(_04450_ ), .A3(_04913_ ), .ZN(_04914_ ) );
INV_X1 _12588_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_04915_ ) );
AND3_X1 _12589_ ( .A1(_04429_ ), .A2(_04915_ ), .A3(_04439_ ), .ZN(_04916_ ) );
NOR2_X1 _12590_ ( .A1(_04914_ ), .A2(_04916_ ), .ZN(_04917_ ) );
OAI211_X1 _12591_ ( .A(_04907_ ), .B(_04865_ ), .C1(_04786_ ), .C2(_04917_ ), .ZN(_04918_ ) );
NAND2_X1 _12592_ ( .A1(_02845_ ), .A2(_02921_ ), .ZN(_04919_ ) );
XNOR2_X1 _12593_ ( .A(_04919_ ), .B(_02868_ ), .ZN(_04920_ ) );
AOI22_X1 _12594_ ( .A1(_04920_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04904_ ), .ZN(_04921_ ) );
AOI21_X1 _12595_ ( .A(_04902_ ), .B1(_04918_ ), .B2(_04921_ ), .ZN(_00140_ ) );
INV_X1 _12596_ ( .A(\ID_EX_pc [4] ), .ZN(_04922_ ) );
XNOR2_X1 _12597_ ( .A(_03087_ ), .B(_04922_ ), .ZN(_04923_ ) );
XOR2_X1 _12598_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_04924_ ) );
XNOR2_X1 _12599_ ( .A(_03137_ ), .B(_04924_ ), .ZN(_04925_ ) );
MUX2_X1 _12600_ ( .A(_04923_ ), .B(_04925_ ), .S(_04689_ ), .Z(_04926_ ) );
OR2_X1 _12601_ ( .A1(_04926_ ), .A2(\ID_EX_typ [3] ), .ZN(_04927_ ) );
NAND3_X1 _12602_ ( .A1(_04488_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_04494_ ), .ZN(_04928_ ) );
NAND3_X1 _12603_ ( .A1(_04488_ ), .A2(\mepc [4] ), .A3(_04463_ ), .ZN(_04929_ ) );
NAND3_X1 _12604_ ( .A1(_04640_ ), .A2(\mtvec [4] ), .A3(_04636_ ), .ZN(_04930_ ) );
NAND4_X1 _12605_ ( .A1(_04928_ ), .A2(_04929_ ), .A3(_04930_ ), .A4(_04497_ ), .ZN(_04931_ ) );
AND3_X1 _12606_ ( .A1(_04554_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_04455_ ), .ZN(_04932_ ) );
NOR3_X1 _12607_ ( .A1(_04931_ ), .A2(_04639_ ), .A3(_04932_ ), .ZN(_04933_ ) );
INV_X1 _12608_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_04934_ ) );
AND3_X1 _12609_ ( .A1(_04508_ ), .A2(_04934_ ), .A3(_04502_ ), .ZN(_04935_ ) );
NOR2_X1 _12610_ ( .A1(_04933_ ), .A2(_04935_ ), .ZN(_04936_ ) );
OAI211_X1 _12611_ ( .A(_04927_ ), .B(_04865_ ), .C1(_04786_ ), .C2(_04936_ ), .ZN(_04937_ ) );
XOR2_X1 _12612_ ( .A(_02821_ ), .B(_02844_ ), .Z(_04938_ ) );
AOI22_X1 _12613_ ( .A1(_04938_ ), .A2(_04668_ ), .B1(_04485_ ), .B2(_04925_ ), .ZN(_04939_ ) );
AOI21_X1 _12614_ ( .A(_04902_ ), .B1(_04937_ ), .B2(_04939_ ), .ZN(_00141_ ) );
XOR2_X1 _12615_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .Z(_04940_ ) );
NOR2_X1 _12616_ ( .A1(_03136_ ), .A2(_03134_ ), .ZN(_04941_ ) );
XNOR2_X1 _12617_ ( .A(_03133_ ), .B(_04941_ ), .ZN(_04942_ ) );
MUX2_X1 _12618_ ( .A(_04940_ ), .B(_04942_ ), .S(_04689_ ), .Z(_04943_ ) );
OR2_X1 _12619_ ( .A1(_04943_ ), .A2(\ID_EX_typ [3] ), .ZN(_04944_ ) );
INV_X1 _12620_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_04945_ ) );
AND3_X1 _12621_ ( .A1(_04591_ ), .A2(_04945_ ), .A3(_04592_ ), .ZN(_04946_ ) );
NAND3_X1 _12622_ ( .A1(_04582_ ), .A2(\mtvec [3] ), .A3(_04476_ ), .ZN(_04947_ ) );
NAND3_X1 _12623_ ( .A1(_04473_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_04456_ ), .ZN(_04948_ ) );
AND2_X1 _12624_ ( .A1(_04947_ ), .A2(_04948_ ), .ZN(_04949_ ) );
NAND3_X1 _12625_ ( .A1(_04580_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_04469_ ), .ZN(_04950_ ) );
NAND3_X1 _12626_ ( .A1(_04580_ ), .A2(\mepc [3] ), .A3(_04464_ ), .ZN(_04951_ ) );
AND3_X1 _12627_ ( .A1(_04949_ ), .A2(_04950_ ), .A3(_04951_ ), .ZN(_04952_ ) );
AOI21_X1 _12628_ ( .A(_04946_ ), .B1(_04451_ ), .B2(_04952_ ), .ZN(_04953_ ) );
OAI211_X1 _12629_ ( .A(_04944_ ), .B(_04865_ ), .C1(_04786_ ), .C2(_04953_ ), .ZN(_04954_ ) );
XOR2_X1 _12630_ ( .A(_02794_ ), .B(_02817_ ), .Z(_04955_ ) );
AOI22_X1 _12631_ ( .A1(_04955_ ), .A2(_04668_ ), .B1(_04484_ ), .B2(_04942_ ), .ZN(_04956_ ) );
AOI21_X1 _12632_ ( .A(_04902_ ), .B1(_04954_ ), .B2(_04956_ ), .ZN(_00142_ ) );
AOI211_X1 _12633_ ( .A(_03129_ ), .B(_03125_ ), .C1(_03127_ ), .C2(_03126_ ), .ZN(_04957_ ) );
NOR2_X1 _12634_ ( .A1(_03131_ ), .A2(_04957_ ), .ZN(_04958_ ) );
MUX2_X1 _12635_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B(_04958_ ), .S(_04689_ ), .Z(_04959_ ) );
OR2_X1 _12636_ ( .A1(_04959_ ), .A2(\ID_EX_typ [3] ), .ZN(_04960_ ) );
AND3_X1 _12637_ ( .A1(_04471_ ), .A2(\mtvec [2] ), .A3(_04474_ ), .ZN(_04961_ ) );
NOR2_X1 _12638_ ( .A1(_04961_ ), .A2(_04548_ ), .ZN(_04962_ ) );
NAND3_X1 _12639_ ( .A1(_04460_ ), .A2(\mepc [2] ), .A3(_04449_ ), .ZN(_04963_ ) );
NAND3_X1 _12640_ ( .A1(_04460_ ), .A2(\mycsreg.CSReg[3][2] ), .A3(_04467_ ), .ZN(_04964_ ) );
NAND3_X1 _12641_ ( .A1(_04557_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_04454_ ), .ZN(_04965_ ) );
NAND4_X1 _12642_ ( .A1(_04962_ ), .A2(_04963_ ), .A3(_04964_ ), .A4(_04965_ ), .ZN(_04966_ ) );
NAND2_X1 _12643_ ( .A1(_04579_ ), .A2(_04966_ ), .ZN(_04967_ ) );
NAND3_X1 _12644_ ( .A1(_04428_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_04438_ ), .ZN(_04968_ ) );
AND2_X1 _12645_ ( .A1(_04967_ ), .A2(_04968_ ), .ZN(_04969_ ) );
INV_X1 _12646_ ( .A(_04969_ ), .ZN(_04970_ ) );
OAI211_X1 _12647_ ( .A(_04960_ ), .B(_04865_ ), .C1(_04786_ ), .C2(_04970_ ), .ZN(_04971_ ) );
OR3_X1 _12648_ ( .A1(_02790_ ), .A2(_02791_ ), .A3(_02743_ ), .ZN(_04972_ ) );
AND2_X1 _12649_ ( .A1(_04972_ ), .A2(_02792_ ), .ZN(_04973_ ) );
AOI22_X1 _12650_ ( .A1(_04973_ ), .A2(_02128_ ), .B1(_04484_ ), .B2(_04958_ ), .ZN(_04974_ ) );
AOI21_X1 _12651_ ( .A(_04902_ ), .B1(_04971_ ), .B2(_04974_ ), .ZN(_00143_ ) );
XOR2_X1 _12652_ ( .A(_03126_ ), .B(_03127_ ), .Z(_04975_ ) );
AOI21_X1 _12653_ ( .A(\ID_EX_typ [3] ), .B1(_04401_ ), .B2(_04975_ ), .ZN(_04976_ ) );
INV_X1 _12654_ ( .A(\ID_EX_pc [1] ), .ZN(_04977_ ) );
OAI21_X1 _12655_ ( .A(_04976_ ), .B1(_04977_ ), .B2(_04568_ ), .ZN(_04978_ ) );
AND3_X1 _12656_ ( .A1(_04591_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_04592_ ), .ZN(_04979_ ) );
INV_X1 _12657_ ( .A(_04979_ ), .ZN(_04980_ ) );
NAND3_X1 _12658_ ( .A1(_04462_ ), .A2(\mepc [1] ), .A3(_04464_ ), .ZN(_04981_ ) );
NAND3_X1 _12659_ ( .A1(_04462_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_04469_ ), .ZN(_04982_ ) );
NAND3_X1 _12660_ ( .A1(_04473_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_04456_ ), .ZN(_04983_ ) );
NAND3_X1 _12661_ ( .A1(_04582_ ), .A2(\mtvec [1] ), .A3(_04476_ ), .ZN(_04984_ ) );
AND4_X1 _12662_ ( .A1(_04981_ ), .A2(_04982_ ), .A3(_04983_ ), .A4(_04984_ ), .ZN(_04985_ ) );
OAI21_X1 _12663_ ( .A(_04980_ ), .B1(_04441_ ), .B2(_04985_ ), .ZN(_04986_ ) );
OAI211_X1 _12664_ ( .A(_04978_ ), .B(_04865_ ), .C1(_04599_ ), .C2(_04986_ ), .ZN(_04987_ ) );
XOR2_X1 _12665_ ( .A(_02766_ ), .B(_02789_ ), .Z(_04988_ ) );
AOI22_X1 _12666_ ( .A1(_04988_ ), .A2(_02128_ ), .B1(_04484_ ), .B2(_04975_ ), .ZN(_04989_ ) );
AOI21_X1 _12667_ ( .A(_04902_ ), .B1(_04987_ ), .B2(_04989_ ), .ZN(_00144_ ) );
INV_X4 _12668_ ( .A(_04400_ ), .ZN(_04990_ ) );
NAND3_X1 _12669_ ( .A1(_04520_ ), .A2(\ID_EX_pc [26] ), .A3(_04523_ ), .ZN(_04991_ ) );
XNOR2_X1 _12670_ ( .A(_04991_ ), .B(\ID_EX_pc [27] ), .ZN(_04992_ ) );
NAND2_X1 _12671_ ( .A1(_04990_ ), .A2(_04992_ ), .ZN(_04993_ ) );
NAND2_X1 _12672_ ( .A1(_03207_ ), .A2(_03209_ ), .ZN(_04994_ ) );
NAND2_X1 _12673_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_04995_ ) );
NAND2_X1 _12674_ ( .A1(_04994_ ), .A2(_04995_ ), .ZN(_04996_ ) );
XNOR2_X1 _12675_ ( .A(_04996_ ), .B(_03208_ ), .ZN(_04997_ ) );
OAI211_X1 _12676_ ( .A(_04993_ ), .B(_04408_ ), .C1(_04990_ ), .C2(_04997_ ), .ZN(_04998_ ) );
NAND3_X1 _12677_ ( .A1(_04461_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_04468_ ), .ZN(_04999_ ) );
AND2_X1 _12678_ ( .A1(_04999_ ), .A2(_04496_ ), .ZN(_05000_ ) );
NAND3_X1 _12679_ ( .A1(_04611_ ), .A2(\mepc [27] ), .A3(_04489_ ), .ZN(_05001_ ) );
NAND4_X1 _12680_ ( .A1(_04453_ ), .A2(_04491_ ), .A3(\mycsreg.CSReg[0][27] ), .A4(_04444_ ), .ZN(_05002_ ) );
AND3_X1 _12681_ ( .A1(_04557_ ), .A2(\mtvec [27] ), .A3(_04474_ ), .ZN(_05003_ ) );
AOI21_X1 _12682_ ( .A(_05003_ ), .B1(_04501_ ), .B2(_04507_ ), .ZN(_05004_ ) );
NAND4_X1 _12683_ ( .A1(_05000_ ), .A2(_05001_ ), .A3(_05002_ ), .A4(_05004_ ), .ZN(_05005_ ) );
INV_X1 _12684_ ( .A(\EX_LS_result_csreg_mem [27] ), .ZN(_05006_ ) );
NAND3_X1 _12685_ ( .A1(_04511_ ), .A2(_05006_ ), .A3(_04513_ ), .ZN(_05007_ ) );
AND2_X1 _12686_ ( .A1(_05005_ ), .A2(_05007_ ), .ZN(_05008_ ) );
OAI211_X1 _12687_ ( .A(_04998_ ), .B(_04865_ ), .C1(_04599_ ), .C2(_05008_ ), .ZN(_05009_ ) );
NOR2_X1 _12688_ ( .A1(_03071_ ), .A2(_02130_ ), .ZN(_05010_ ) );
NOR2_X1 _12689_ ( .A1(_04997_ ), .A2(_04537_ ), .ZN(_05011_ ) );
NOR2_X1 _12690_ ( .A1(_05010_ ), .A2(_05011_ ), .ZN(_05012_ ) );
AOI21_X1 _12691_ ( .A(_04902_ ), .B1(_05009_ ), .B2(_05012_ ), .ZN(_00145_ ) );
XOR2_X1 _12692_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05013_ ) );
OAI21_X1 _12693_ ( .A(_04407_ ), .B1(_04990_ ), .B2(_05013_ ), .ZN(_05014_ ) );
INV_X1 _12694_ ( .A(\ID_EX_pc [0] ), .ZN(_05015_ ) );
AOI21_X1 _12695_ ( .A(_05014_ ), .B1(_05015_ ), .B2(_04990_ ), .ZN(_05016_ ) );
AND3_X1 _12696_ ( .A1(_04554_ ), .A2(\mtvec [0] ), .A3(_04636_ ), .ZN(_05017_ ) );
NOR2_X1 _12697_ ( .A1(_05017_ ), .A2(_04548_ ), .ZN(_05018_ ) );
NAND3_X1 _12698_ ( .A1(_04462_ ), .A2(\mepc [0] ), .A3(_04464_ ), .ZN(_05019_ ) );
NAND3_X1 _12699_ ( .A1(_04462_ ), .A2(\mycsreg.CSReg[3][0] ), .A3(_04469_ ), .ZN(_05020_ ) );
NAND3_X1 _12700_ ( .A1(_04473_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_04456_ ), .ZN(_05021_ ) );
NAND4_X1 _12701_ ( .A1(_05018_ ), .A2(_05019_ ), .A3(_05020_ ), .A4(_05021_ ), .ZN(_05022_ ) );
NAND2_X1 _12702_ ( .A1(_04579_ ), .A2(_05022_ ), .ZN(_05023_ ) );
NAND3_X1 _12703_ ( .A1(_04591_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_04592_ ), .ZN(_05024_ ) );
AOI21_X1 _12704_ ( .A(_04408_ ), .B1(_05023_ ), .B2(_05024_ ), .ZN(_05025_ ) );
OAI21_X1 _12705_ ( .A(_04406_ ), .B1(_05016_ ), .B2(_05025_ ), .ZN(_05026_ ) );
BUF_X4 _12706_ ( .A(_04482_ ), .Z(_05027_ ) );
BUF_X4 _12707_ ( .A(_05027_ ), .Z(_05028_ ) );
BUF_X4 _12708_ ( .A(_04487_ ), .Z(_05029_ ) );
NAND3_X1 _12709_ ( .A1(_05013_ ), .A2(_05028_ ), .A3(_05029_ ), .ZN(_05030_ ) );
AOI21_X1 _12710_ ( .A(_04902_ ), .B1(_05026_ ), .B2(_05030_ ), .ZN(_00146_ ) );
INV_X1 _12711_ ( .A(\ID_EX_pc [26] ), .ZN(_05031_ ) );
XNOR2_X1 _12712_ ( .A(_04524_ ), .B(_05031_ ), .ZN(_05032_ ) );
XOR2_X1 _12713_ ( .A(_03207_ ), .B(_03209_ ), .Z(_05033_ ) );
MUX2_X1 _12714_ ( .A(_05032_ ), .B(_05033_ ), .S(_04689_ ), .Z(_05034_ ) );
OR2_X1 _12715_ ( .A1(_05034_ ), .A2(\ID_EX_typ [3] ), .ZN(_05035_ ) );
NAND3_X1 _12716_ ( .A1(_04429_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_04439_ ), .ZN(_05036_ ) );
NAND3_X1 _12717_ ( .A1(_04462_ ), .A2(\mepc [26] ), .A3(_04464_ ), .ZN(_05037_ ) );
NAND3_X1 _12718_ ( .A1(_04462_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_04469_ ), .ZN(_05038_ ) );
NAND3_X1 _12719_ ( .A1(_04473_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_04456_ ), .ZN(_05039_ ) );
NAND3_X1 _12720_ ( .A1(_04582_ ), .A2(\mtvec [26] ), .A3(_04476_ ), .ZN(_05040_ ) );
AND4_X1 _12721_ ( .A1(_05037_ ), .A2(_05038_ ), .A3(_05039_ ), .A4(_05040_ ), .ZN(_05041_ ) );
OAI21_X1 _12722_ ( .A(_05036_ ), .B1(_04441_ ), .B2(_05041_ ), .ZN(_05042_ ) );
OAI211_X1 _12723_ ( .A(_05035_ ), .B(_04865_ ), .C1(_04599_ ), .C2(_05042_ ), .ZN(_05043_ ) );
NOR3_X1 _12724_ ( .A1(_03072_ ), .A2(_03069_ ), .A3(_02129_ ), .ZN(_05044_ ) );
AOI21_X1 _12725_ ( .A(_05044_ ), .B1(_04566_ ), .B2(_05033_ ), .ZN(_05045_ ) );
AOI21_X1 _12726_ ( .A(_04902_ ), .B1(_05043_ ), .B2(_05045_ ), .ZN(_00147_ ) );
AND3_X1 _12727_ ( .A1(_04522_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05046_ ) );
AND2_X1 _12728_ ( .A1(_04520_ ), .A2(_05046_ ), .ZN(_05047_ ) );
NAND3_X1 _12729_ ( .A1(_05047_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05048_ ) );
INV_X1 _12730_ ( .A(\ID_EX_pc [24] ), .ZN(_05049_ ) );
NOR2_X1 _12731_ ( .A1(_05048_ ), .A2(_05049_ ), .ZN(_05050_ ) );
INV_X1 _12732_ ( .A(\ID_EX_pc [25] ), .ZN(_05051_ ) );
XNOR2_X1 _12733_ ( .A(_05050_ ), .B(_05051_ ), .ZN(_05052_ ) );
AOI21_X1 _12734_ ( .A(_05052_ ), .B1(_04600_ ), .B2(_04601_ ), .ZN(_05053_ ) );
AND2_X1 _12735_ ( .A1(_03200_ ), .A2(_03202_ ), .ZN(_05054_ ) );
OR2_X1 _12736_ ( .A1(_05054_ ), .A2(_03204_ ), .ZN(_05055_ ) );
XNOR2_X1 _12737_ ( .A(_05055_ ), .B(_03201_ ), .ZN(_05056_ ) );
AOI21_X1 _12738_ ( .A(_05053_ ), .B1(_04401_ ), .B2(_05056_ ), .ZN(_05057_ ) );
OR2_X1 _12739_ ( .A1(_05057_ ), .A2(\ID_EX_typ [3] ), .ZN(_05058_ ) );
NAND3_X1 _12740_ ( .A1(_04429_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_04439_ ), .ZN(_05059_ ) );
NAND3_X1 _12741_ ( .A1(_04580_ ), .A2(\mepc [25] ), .A3(_04464_ ), .ZN(_05060_ ) );
NAND3_X1 _12742_ ( .A1(_04611_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_04494_ ), .ZN(_05061_ ) );
NAND3_X1 _12743_ ( .A1(_04582_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_04456_ ), .ZN(_05062_ ) );
NAND3_X1 _12744_ ( .A1(_04582_ ), .A2(\mtvec [25] ), .A3(_04476_ ), .ZN(_05063_ ) );
AND4_X1 _12745_ ( .A1(_05060_ ), .A2(_05061_ ), .A3(_05062_ ), .A4(_05063_ ), .ZN(_05064_ ) );
OAI21_X1 _12746_ ( .A(_05059_ ), .B1(_04441_ ), .B2(_05064_ ), .ZN(_05065_ ) );
OAI211_X1 _12747_ ( .A(_05058_ ), .B(_04865_ ), .C1(_04599_ ), .C2(_05065_ ), .ZN(_05066_ ) );
NOR2_X1 _12748_ ( .A1(_03075_ ), .A2(_02130_ ), .ZN(_05067_ ) );
NOR2_X1 _12749_ ( .A1(_05056_ ), .A2(_04537_ ), .ZN(_05068_ ) );
NOR2_X1 _12750_ ( .A1(_05067_ ), .A2(_05068_ ), .ZN(_05069_ ) );
AOI21_X1 _12751_ ( .A(_04902_ ), .B1(_05066_ ), .B2(_05069_ ), .ZN(_00148_ ) );
NOR3_X1 _12752_ ( .A1(_03076_ ), .A2(_03073_ ), .A3(_02129_ ), .ZN(_05070_ ) );
XOR2_X1 _12753_ ( .A(_03200_ ), .B(_03202_ ), .Z(_05071_ ) );
NAND3_X1 _12754_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_05071_ ), .ZN(_05072_ ) );
XNOR2_X1 _12755_ ( .A(_05048_ ), .B(_05049_ ), .ZN(_05073_ ) );
OAI211_X1 _12756_ ( .A(_04407_ ), .B(_05072_ ), .C1(_04401_ ), .C2(_05073_ ), .ZN(_05074_ ) );
NAND3_X1 _12757_ ( .A1(_04460_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_04467_ ), .ZN(_05075_ ) );
NAND3_X1 _12758_ ( .A1(_04460_ ), .A2(\mepc [24] ), .A3(_04449_ ), .ZN(_05076_ ) );
NAND3_X1 _12759_ ( .A1(_04472_ ), .A2(\mtvec [24] ), .A3(_04475_ ), .ZN(_05077_ ) );
NAND4_X1 _12760_ ( .A1(_04549_ ), .A2(_05075_ ), .A3(_05076_ ), .A4(_05077_ ), .ZN(_05078_ ) );
AND3_X1 _12761_ ( .A1(_04472_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_04455_ ), .ZN(_05079_ ) );
NOR3_X1 _12762_ ( .A1(_05078_ ), .A2(_04639_ ), .A3(_05079_ ), .ZN(_05080_ ) );
INV_X1 _12763_ ( .A(\EX_LS_result_csreg_mem [24] ), .ZN(_05081_ ) );
AND3_X1 _12764_ ( .A1(_04507_ ), .A2(_05081_ ), .A3(_04501_ ), .ZN(_05082_ ) );
NOR2_X1 _12765_ ( .A1(_05080_ ), .A2(_05082_ ), .ZN(_05083_ ) );
INV_X1 _12766_ ( .A(_05083_ ), .ZN(_05084_ ) );
AOI21_X1 _12767_ ( .A(_04487_ ), .B1(_05084_ ), .B2(\ID_EX_typ [3] ), .ZN(_05085_ ) );
AOI221_X1 _12768_ ( .A(_05070_ ), .B1(_04484_ ), .B2(_05071_ ), .C1(_05074_ ), .C2(_05085_ ), .ZN(_05086_ ) );
NOR2_X1 _12769_ ( .A1(_05086_ ), .A2(_03086_ ), .ZN(_00149_ ) );
NAND3_X1 _12770_ ( .A1(_04520_ ), .A2(\ID_EX_pc [22] ), .A3(_05046_ ), .ZN(_05087_ ) );
XNOR2_X1 _12771_ ( .A(_05087_ ), .B(\ID_EX_pc [23] ), .ZN(_05088_ ) );
NAND2_X1 _12772_ ( .A1(_04990_ ), .A2(_05088_ ), .ZN(_05089_ ) );
INV_X1 _12773_ ( .A(_03114_ ), .ZN(_05090_ ) );
NOR2_X1 _12774_ ( .A1(_04544_ ), .A2(_05090_ ), .ZN(_05091_ ) );
NOR2_X1 _12775_ ( .A1(_05091_ ), .A2(_03191_ ), .ZN(_05092_ ) );
NOR3_X1 _12776_ ( .A1(_05092_ ), .A2(_03106_ ), .A3(_03107_ ), .ZN(_05093_ ) );
OR2_X1 _12777_ ( .A1(_05093_ ), .A2(_03106_ ), .ZN(_05094_ ) );
XNOR2_X1 _12778_ ( .A(_05094_ ), .B(_03105_ ), .ZN(_05095_ ) );
OAI211_X1 _12779_ ( .A(_05089_ ), .B(_04408_ ), .C1(_04990_ ), .C2(_05095_ ), .ZN(_05096_ ) );
BUF_X4 _12780_ ( .A(_04405_ ), .Z(_05097_ ) );
NAND3_X1 _12781_ ( .A1(_04429_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_04439_ ), .ZN(_05098_ ) );
NAND3_X1 _12782_ ( .A1(_04462_ ), .A2(\mepc [23] ), .A3(_04464_ ), .ZN(_05099_ ) );
NAND3_X1 _12783_ ( .A1(_04462_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_04469_ ), .ZN(_05100_ ) );
NAND3_X1 _12784_ ( .A1(_04473_ ), .A2(\mtvec [23] ), .A3(_04476_ ), .ZN(_05101_ ) );
NAND3_X1 _12785_ ( .A1(_04582_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_04456_ ), .ZN(_05102_ ) );
AND4_X1 _12786_ ( .A1(_05099_ ), .A2(_05100_ ), .A3(_05101_ ), .A4(_05102_ ), .ZN(_05103_ ) );
OAI21_X1 _12787_ ( .A(_05098_ ), .B1(_04441_ ), .B2(_05103_ ), .ZN(_05104_ ) );
OAI211_X1 _12788_ ( .A(_05096_ ), .B(_05097_ ), .C1(_04599_ ), .C2(_05104_ ), .ZN(_05105_ ) );
NOR2_X1 _12789_ ( .A1(_03082_ ), .A2(_02130_ ), .ZN(_05106_ ) );
NOR2_X1 _12790_ ( .A1(_05095_ ), .A2(_04537_ ), .ZN(_05107_ ) );
NOR2_X1 _12791_ ( .A1(_05106_ ), .A2(_05107_ ), .ZN(_05108_ ) );
AOI21_X1 _12792_ ( .A(_04902_ ), .B1(_05105_ ), .B2(_05108_ ), .ZN(_00150_ ) );
XNOR2_X1 _12793_ ( .A(_05092_ ), .B(_03108_ ), .ZN(_05109_ ) );
NAND2_X1 _12794_ ( .A1(_05109_ ), .A2(_04484_ ), .ZN(_05110_ ) );
INV_X1 _12795_ ( .A(\ID_EX_pc [22] ), .ZN(_05111_ ) );
XNOR2_X1 _12796_ ( .A(_05047_ ), .B(_05111_ ), .ZN(_05112_ ) );
AND2_X4 _12797_ ( .A1(_04990_ ), .A2(_05112_ ), .ZN(_05113_ ) );
AOI211_X2 _12798_ ( .A(\ID_EX_typ [3] ), .B(_05113_ ), .C1(_04568_ ), .C2(_05109_ ), .ZN(_05114_ ) );
NAND3_X1 _12799_ ( .A1(_04461_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_04494_ ), .ZN(_05115_ ) );
AND2_X1 _12800_ ( .A1(_04549_ ), .A2(_05115_ ), .ZN(_05116_ ) );
NAND3_X1 _12801_ ( .A1(_04461_ ), .A2(\mepc [22] ), .A3(_04463_ ), .ZN(_05117_ ) );
NAND3_X1 _12802_ ( .A1(_04554_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_04455_ ), .ZN(_05118_ ) );
AND2_X1 _12803_ ( .A1(_05117_ ), .A2(_05118_ ), .ZN(_05119_ ) );
AND3_X1 _12804_ ( .A1(_04472_ ), .A2(\mtvec [22] ), .A3(_04475_ ), .ZN(_05120_ ) );
AOI21_X1 _12805_ ( .A(_05120_ ), .B1(_04502_ ), .B2(_04508_ ), .ZN(_05121_ ) );
NAND3_X1 _12806_ ( .A1(_05116_ ), .A2(_05119_ ), .A3(_05121_ ), .ZN(_05122_ ) );
INV_X1 _12807_ ( .A(\EX_LS_result_csreg_mem [22] ), .ZN(_05123_ ) );
NAND3_X1 _12808_ ( .A1(_04511_ ), .A2(_05123_ ), .A3(_04513_ ), .ZN(_05124_ ) );
AND2_X1 _12809_ ( .A1(_05122_ ), .A2(_05124_ ), .ZN(_05125_ ) );
OAI21_X1 _12810_ ( .A(_04405_ ), .B1(_05125_ ), .B2(_04408_ ), .ZN(_05126_ ) );
OAI221_X1 _12811_ ( .A(_05110_ ), .B1(_02130_ ), .B2(_03083_ ), .C1(_05114_ ), .C2(_05126_ ), .ZN(_05127_ ) );
AND2_X1 _12812_ ( .A1(_05127_ ), .A2(_02115_ ), .ZN(_00151_ ) );
OAI21_X1 _12813_ ( .A(_03110_ ), .B1(_04543_ ), .B2(_03198_ ), .ZN(_05128_ ) );
NAND2_X1 _12814_ ( .A1(_05128_ ), .A2(_03189_ ), .ZN(_05129_ ) );
XNOR2_X1 _12815_ ( .A(_05129_ ), .B(_03113_ ), .ZN(_05130_ ) );
NAND3_X1 _12816_ ( .A1(_04461_ ), .A2(\mepc [21] ), .A3(_04463_ ), .ZN(_05131_ ) );
NAND4_X1 _12817_ ( .A1(_04453_ ), .A2(_04455_ ), .A3(\mycsreg.CSReg[0][21] ), .A4(_04444_ ), .ZN(_05132_ ) );
AND2_X1 _12818_ ( .A1(_05131_ ), .A2(_05132_ ), .ZN(_05133_ ) );
NAND3_X1 _12819_ ( .A1(_04552_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_04468_ ), .ZN(_05134_ ) );
NAND3_X1 _12820_ ( .A1(_04472_ ), .A2(\mtvec [21] ), .A3(_04475_ ), .ZN(_05135_ ) );
AND3_X1 _12821_ ( .A1(_05134_ ), .A2(_04496_ ), .A3(_05135_ ), .ZN(_05136_ ) );
NAND3_X1 _12822_ ( .A1(_04658_ ), .A2(_05133_ ), .A3(_05136_ ), .ZN(_05137_ ) );
INV_X1 _12823_ ( .A(\EX_LS_result_csreg_mem [21] ), .ZN(_05138_ ) );
NAND3_X1 _12824_ ( .A1(_04511_ ), .A2(_05138_ ), .A3(_04513_ ), .ZN(_05139_ ) );
NAND2_X1 _12825_ ( .A1(_05137_ ), .A2(_05139_ ), .ZN(_05140_ ) );
AOI21_X1 _12826_ ( .A(_04487_ ), .B1(_05140_ ), .B2(\ID_EX_typ [3] ), .ZN(_05141_ ) );
NAND3_X1 _12827_ ( .A1(_04600_ ), .A2(_04601_ ), .A3(_05141_ ), .ZN(_05142_ ) );
AOI21_X1 _12828_ ( .A(_05130_ ), .B1(_05142_ ), .B2(_04537_ ), .ZN(_05143_ ) );
NOR2_X1 _12829_ ( .A1(_03039_ ), .A2(_02130_ ), .ZN(_05144_ ) );
NOR2_X1 _12830_ ( .A1(_05143_ ), .A2(_05144_ ), .ZN(_05145_ ) );
INV_X1 _12831_ ( .A(\ID_EX_pc [20] ), .ZN(_05146_ ) );
NOR2_X1 _12832_ ( .A1(_04539_ ), .A2(_05146_ ), .ZN(_05147_ ) );
XNOR2_X1 _12833_ ( .A(_05147_ ), .B(\ID_EX_pc [21] ), .ZN(_05148_ ) );
AOI21_X1 _12834_ ( .A(_05148_ ), .B1(_04600_ ), .B2(_04601_ ), .ZN(_05149_ ) );
OAI21_X1 _12835_ ( .A(_05141_ ), .B1(_05149_ ), .B2(\ID_EX_typ [3] ), .ZN(_05150_ ) );
AOI21_X1 _12836_ ( .A(_03085_ ), .B1(_05145_ ), .B2(_05150_ ), .ZN(_00152_ ) );
BUF_X2 _12837_ ( .A(_04658_ ), .Z(_05151_ ) );
NOR2_X1 _12838_ ( .A1(_05151_ ), .A2(\EX_LS_result_csreg_mem [31] ), .ZN(_05152_ ) );
NAND3_X1 _12839_ ( .A1(_04554_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04455_ ), .ZN(_05153_ ) );
NAND3_X1 _12840_ ( .A1(_04554_ ), .A2(\mtvec [31] ), .A3(_04636_ ), .ZN(_05154_ ) );
AND2_X1 _12841_ ( .A1(_05153_ ), .A2(_05154_ ), .ZN(_05155_ ) );
NAND3_X1 _12842_ ( .A1(_04611_ ), .A2(\mepc [31] ), .A3(_04489_ ), .ZN(_05156_ ) );
NAND3_X1 _12843_ ( .A1(_04611_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_04494_ ), .ZN(_05157_ ) );
NAND3_X1 _12844_ ( .A1(_05155_ ), .A2(_05156_ ), .A3(_05157_ ), .ZN(_05158_ ) );
BUF_X2 _12845_ ( .A(_04639_ ), .Z(_05159_ ) );
NOR2_X1 _12846_ ( .A1(_05158_ ), .A2(_05159_ ), .ZN(_05160_ ) );
NOR2_X1 _12847_ ( .A1(_05152_ ), .A2(_05160_ ), .ZN(_05161_ ) );
INV_X1 _12848_ ( .A(\ID_EX_pc [30] ), .ZN(_05162_ ) );
NOR2_X1 _12849_ ( .A1(_03103_ ), .A2(_05162_ ), .ZN(_05163_ ) );
INV_X1 _12850_ ( .A(\ID_EX_pc [31] ), .ZN(_05164_ ) );
XNOR2_X1 _12851_ ( .A(_05163_ ), .B(_05164_ ), .ZN(_05165_ ) );
NAND2_X1 _12852_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_05166_ ) );
NAND2_X1 _12853_ ( .A1(_03222_ ), .A2(_05166_ ), .ZN(_05167_ ) );
XNOR2_X1 _12854_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_05168_ ) );
XNOR2_X1 _12855_ ( .A(_05167_ ), .B(_05168_ ), .ZN(_05169_ ) );
MUX2_X1 _12856_ ( .A(_05165_ ), .B(_05169_ ), .S(_04400_ ), .Z(_05170_ ) );
MUX2_X1 _12857_ ( .A(_05161_ ), .B(_05170_ ), .S(_04407_ ), .Z(_05171_ ) );
NAND2_X1 _12858_ ( .A1(_05171_ ), .A2(_04406_ ), .ZN(_05172_ ) );
OR2_X1 _12859_ ( .A1(_03027_ ), .A2(_02130_ ), .ZN(_05173_ ) );
NAND2_X1 _12860_ ( .A1(_05169_ ), .A2(_04566_ ), .ZN(_05174_ ) );
NAND4_X1 _12861_ ( .A1(_05172_ ), .A2(_03084_ ), .A3(_05173_ ), .A4(_05174_ ), .ZN(_00153_ ) );
NOR3_X1 _12862_ ( .A1(_05164_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00154_ ) );
NOR3_X1 _12863_ ( .A1(_05162_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00155_ ) );
AND2_X1 _12864_ ( .A1(_03084_ ), .A2(\ID_EX_pc [21] ), .ZN(_00156_ ) );
NOR3_X1 _12865_ ( .A1(_05146_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00157_ ) );
NOR3_X1 _12866_ ( .A1(_04576_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00158_ ) );
INV_X1 _12867_ ( .A(\ID_EX_pc [18] ), .ZN(_05175_ ) );
NOR3_X1 _12868_ ( .A1(_05175_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00159_ ) );
NOR3_X1 _12869_ ( .A1(_04627_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00160_ ) );
NOR3_X1 _12870_ ( .A1(_04650_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00161_ ) );
NOR3_X1 _12871_ ( .A1(_04623_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00162_ ) );
NOR3_X1 _12872_ ( .A1(_04624_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00163_ ) );
NOR3_X1 _12873_ ( .A1(_04717_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00164_ ) );
NOR3_X1 _12874_ ( .A1(_04715_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00165_ ) );
NOR3_X1 _12875_ ( .A1(_03217_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00166_ ) );
NOR3_X1 _12876_ ( .A1(_03176_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00167_ ) );
INV_X1 _12877_ ( .A(\ID_EX_pc [10] ), .ZN(_05176_ ) );
NOR3_X1 _12878_ ( .A1(_05176_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00168_ ) );
INV_X1 _12879_ ( .A(\ID_EX_pc [9] ), .ZN(_05177_ ) );
NOR3_X1 _12880_ ( .A1(_05177_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00169_ ) );
NOR3_X1 _12881_ ( .A1(_04841_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00170_ ) );
INV_X1 _12882_ ( .A(\ID_EX_pc [7] ), .ZN(_05178_ ) );
NOR3_X1 _12883_ ( .A1(_05178_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00171_ ) );
NOR3_X1 _12884_ ( .A1(_04883_ ), .A2(fanout_net_2 ), .A3(fanout_net_17 ), .ZN(_00172_ ) );
AND2_X1 _12885_ ( .A1(_03084_ ), .A2(\ID_EX_pc [5] ), .ZN(_00173_ ) );
NOR3_X1 _12886_ ( .A1(_04922_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00174_ ) );
AND2_X1 _12887_ ( .A1(_03084_ ), .A2(\ID_EX_pc [3] ), .ZN(_00175_ ) );
AND2_X1 _12888_ ( .A1(_03084_ ), .A2(\ID_EX_pc [2] ), .ZN(_00176_ ) );
NOR3_X1 _12889_ ( .A1(_04526_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00177_ ) );
NOR3_X1 _12890_ ( .A1(_04977_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00178_ ) );
NOR3_X1 _12891_ ( .A1(_05015_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00179_ ) );
AND2_X1 _12892_ ( .A1(_02115_ ), .A2(\ID_EX_pc [27] ), .ZN(_00180_ ) );
NOR3_X1 _12893_ ( .A1(_05031_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00181_ ) );
NOR3_X1 _12894_ ( .A1(_05051_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00182_ ) );
NOR3_X1 _12895_ ( .A1(_05049_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00183_ ) );
NOR3_X1 _12896_ ( .A1(_03187_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00184_ ) );
NOR3_X1 _12897_ ( .A1(_05111_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00185_ ) );
INV_X1 _12898_ ( .A(\ID_EX_typ [7] ), .ZN(_05179_ ) );
NOR3_X1 _12899_ ( .A1(_05179_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00186_ ) );
INV_X1 _12900_ ( .A(_02091_ ), .ZN(_05180_ ) );
AND2_X4 _12901_ ( .A1(_02014_ ), .A2(_02084_ ), .ZN(_05181_ ) );
OAI21_X1 _12902_ ( .A(_05180_ ), .B1(_05181_ ), .B2(io_master_arready ), .ZN(_05182_ ) );
INV_X1 _12903_ ( .A(_02000_ ), .ZN(_05183_ ) );
BUF_X4 _12904_ ( .A(_05183_ ), .Z(_05184_ ) );
BUF_X4 _12905_ ( .A(_05184_ ), .Z(_05185_ ) );
NOR2_X1 _12906_ ( .A1(_05182_ ), .A2(_05185_ ), .ZN(_05186_ ) );
BUF_X2 _12907_ ( .A(_02005_ ), .Z(_05187_ ) );
INV_X1 _12908_ ( .A(_02021_ ), .ZN(_05188_ ) );
OR3_X1 _12909_ ( .A1(_05186_ ), .A2(_05187_ ), .A3(_05188_ ), .ZN(_05189_ ) );
OR2_X1 _12910_ ( .A1(\mylsu.state [4] ), .A2(\mylsu.state [0] ), .ZN(_05190_ ) );
INV_X1 _12911_ ( .A(_02040_ ), .ZN(_05191_ ) );
OAI21_X1 _12912_ ( .A(_05190_ ), .B1(_05191_ ), .B2(io_master_awready ), .ZN(_05192_ ) );
AOI21_X1 _12913_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .B1(_05192_ ), .B2(EXU_valid_LSU ), .ZN(_05193_ ) );
AOI21_X1 _12914_ ( .A(_03085_ ), .B1(_05189_ ), .B2(_05193_ ), .ZN(_00187_ ) );
NOR3_X1 _12915_ ( .A1(_02121_ ), .A2(fanout_net_3 ), .A3(fanout_net_17 ), .ZN(_00188_ ) );
NOR3_X1 _12916_ ( .A1(_02126_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00189_ ) );
NOR3_X1 _12917_ ( .A1(_04049_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00190_ ) );
NOR3_X1 _12918_ ( .A1(_04409_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00191_ ) );
BUF_X2 _12919_ ( .A(_04393_ ), .Z(_05194_ ) );
BUF_X2 _12920_ ( .A(_05194_ ), .Z(_05195_ ) );
NOR3_X1 _12921_ ( .A1(_05195_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00192_ ) );
NOR3_X1 _12922_ ( .A1(_04304_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00193_ ) );
NOR3_X1 _12923_ ( .A1(_05028_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00194_ ) );
INV_X1 _12924_ ( .A(\IF_ID_inst [6] ), .ZN(_05196_ ) );
NOR2_X1 _12925_ ( .A1(_05196_ ), .A2(\IF_ID_inst [12] ), .ZN(_05197_ ) );
AND2_X1 _12926_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05198_ ) );
AND3_X1 _12927_ ( .A1(_05197_ ), .A2(\IF_ID_inst [13] ), .A3(_05198_ ), .ZN(_05199_ ) );
AND2_X1 _12928_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_05200_ ) );
NOR2_X1 _12929_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_05201_ ) );
AND2_X2 _12930_ ( .A1(_05200_ ), .A2(_05201_ ), .ZN(_05202_ ) );
BUF_X2 _12931_ ( .A(_05202_ ), .Z(_05203_ ) );
AND2_X2 _12932_ ( .A1(_05199_ ), .A2(_05203_ ), .ZN(_05204_ ) );
AND4_X1 _12933_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_05205_ ) );
AND2_X2 _12934_ ( .A1(_05203_ ), .A2(_05205_ ), .ZN(_05206_ ) );
NOR2_X1 _12935_ ( .A1(_05204_ ), .A2(_05206_ ), .ZN(_05207_ ) );
BUF_X4 _12936_ ( .A(_05207_ ), .Z(_05208_ ) );
INV_X1 _12937_ ( .A(\IF_ID_inst [31] ), .ZN(_05209_ ) );
AND2_X1 _12938_ ( .A1(_02106_ ), .A2(_02115_ ), .ZN(_05210_ ) );
INV_X1 _12939_ ( .A(_05210_ ), .ZN(_05211_ ) );
BUF_X4 _12940_ ( .A(_05211_ ), .Z(_05212_ ) );
NOR3_X1 _12941_ ( .A1(_05208_ ), .A2(_05209_ ), .A3(_05212_ ), .ZN(_00195_ ) );
INV_X1 _12942_ ( .A(\IF_ID_inst [30] ), .ZN(_05213_ ) );
NOR3_X1 _12943_ ( .A1(_05208_ ), .A2(_05213_ ), .A3(_05212_ ), .ZN(_00196_ ) );
INV_X1 _12944_ ( .A(\IF_ID_inst [21] ), .ZN(_05214_ ) );
NOR3_X1 _12945_ ( .A1(_05208_ ), .A2(_05214_ ), .A3(_05212_ ), .ZN(_00197_ ) );
BUF_X4 _12946_ ( .A(_05211_ ), .Z(_05215_ ) );
INV_X1 _12947_ ( .A(_05207_ ), .ZN(_05216_ ) );
INV_X1 _12948_ ( .A(\IF_ID_inst [20] ), .ZN(_05217_ ) );
AOI21_X1 _12949_ ( .A(_05215_ ), .B1(_05216_ ), .B2(_05217_ ), .ZN(_00198_ ) );
INV_X1 _12950_ ( .A(\IF_ID_inst [29] ), .ZN(_05218_ ) );
AOI21_X1 _12951_ ( .A(_05215_ ), .B1(_05216_ ), .B2(_05218_ ), .ZN(_00199_ ) );
INV_X1 _12952_ ( .A(\IF_ID_inst [28] ), .ZN(_05219_ ) );
AOI21_X1 _12953_ ( .A(_05215_ ), .B1(_05216_ ), .B2(_05219_ ), .ZN(_00200_ ) );
INV_X1 _12954_ ( .A(\IF_ID_inst [27] ), .ZN(_05220_ ) );
BUF_X4 _12955_ ( .A(_05211_ ), .Z(_05221_ ) );
NOR3_X1 _12956_ ( .A1(_05208_ ), .A2(_05220_ ), .A3(_05221_ ), .ZN(_00201_ ) );
INV_X1 _12957_ ( .A(\IF_ID_inst [26] ), .ZN(_05222_ ) );
AOI21_X1 _12958_ ( .A(_05215_ ), .B1(_05216_ ), .B2(_05222_ ), .ZN(_00202_ ) );
INV_X1 _12959_ ( .A(\IF_ID_inst [25] ), .ZN(_05223_ ) );
NOR3_X1 _12960_ ( .A1(_05208_ ), .A2(_05223_ ), .A3(_05221_ ), .ZN(_00203_ ) );
INV_X1 _12961_ ( .A(\IF_ID_inst [24] ), .ZN(_05224_ ) );
NOR3_X1 _12962_ ( .A1(_05208_ ), .A2(_05224_ ), .A3(_05221_ ), .ZN(_00204_ ) );
INV_X1 _12963_ ( .A(\IF_ID_inst [23] ), .ZN(_05225_ ) );
NOR3_X1 _12964_ ( .A1(_05208_ ), .A2(_05225_ ), .A3(_05221_ ), .ZN(_00205_ ) );
INV_X1 _12965_ ( .A(\IF_ID_inst [22] ), .ZN(_05226_ ) );
NOR3_X1 _12966_ ( .A1(_05208_ ), .A2(_05226_ ), .A3(_05221_ ), .ZN(_00206_ ) );
AND3_X1 _12967_ ( .A1(_02106_ ), .A2(_02115_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00207_ ) );
AND3_X1 _12968_ ( .A1(_02106_ ), .A2(_02115_ ), .A3(\myidu.state [2] ), .ZN(_00208_ ) );
NOR2_X1 _12969_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_05227_ ) );
NOR2_X1 _12970_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05228_ ) );
AND4_X1 _12971_ ( .A1(\IF_ID_inst [12] ), .A2(_05227_ ), .A3(_05228_ ), .A4(_05196_ ), .ZN(_05229_ ) );
AND3_X1 _12972_ ( .A1(_05200_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_05230_ ) );
CLKBUF_X2 _12973_ ( .A(_05230_ ), .Z(_05231_ ) );
AND2_X1 _12974_ ( .A1(_05229_ ), .A2(_05231_ ), .ZN(_05232_ ) );
BUF_X2 _12975_ ( .A(_05227_ ), .Z(_05233_ ) );
INV_X1 _12976_ ( .A(\IF_ID_inst [5] ), .ZN(_05234_ ) );
NOR2_X1 _12977_ ( .A1(_05234_ ), .A2(\IF_ID_inst [4] ), .ZN(_05235_ ) );
AND2_X1 _12978_ ( .A1(_05197_ ), .A2(_05235_ ), .ZN(_05236_ ) );
CLKBUF_X2 _12979_ ( .A(_05203_ ), .Z(_05237_ ) );
AND2_X1 _12980_ ( .A1(_05236_ ), .A2(_05237_ ), .ZN(_05238_ ) );
INV_X1 _12981_ ( .A(\IF_ID_inst [12] ), .ZN(_05239_ ) );
INV_X1 _12982_ ( .A(\IF_ID_inst [7] ), .ZN(_05240_ ) );
INV_X1 _12983_ ( .A(\IF_ID_inst [15] ), .ZN(_05241_ ) );
AND4_X1 _12984_ ( .A1(_05239_ ), .A2(_05240_ ), .A3(_05241_ ), .A4(\IF_ID_inst [6] ), .ZN(_05242_ ) );
BUF_X2 _12985_ ( .A(_05198_ ), .Z(_05243_ ) );
AND3_X1 _12986_ ( .A1(_05242_ ), .A2(_05243_ ), .A3(_05233_ ), .ZN(_05244_ ) );
INV_X1 _12987_ ( .A(\IF_ID_inst [11] ), .ZN(_05245_ ) );
INV_X1 _12988_ ( .A(\IF_ID_inst [10] ), .ZN(_05246_ ) );
INV_X1 _12989_ ( .A(\IF_ID_inst [9] ), .ZN(_05247_ ) );
NAND3_X1 _12990_ ( .A1(_05245_ ), .A2(_05246_ ), .A3(_05247_ ), .ZN(_05248_ ) );
NOR2_X1 _12991_ ( .A1(_05248_ ), .A2(\IF_ID_inst [8] ), .ZN(_05249_ ) );
AND3_X1 _12992_ ( .A1(_05244_ ), .A2(_05237_ ), .A3(_05249_ ), .ZN(_05250_ ) );
NOR2_X1 _12993_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [18] ), .ZN(_05251_ ) );
NOR2_X1 _12994_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_05252_ ) );
AND2_X1 _12995_ ( .A1(_05251_ ), .A2(_05252_ ), .ZN(_05253_ ) );
NAND2_X1 _12996_ ( .A1(_05213_ ), .A2(\IF_ID_inst [29] ), .ZN(_05254_ ) );
NOR3_X1 _12997_ ( .A1(_05254_ ), .A2(_05219_ ), .A3(\IF_ID_inst [31] ), .ZN(_05255_ ) );
NOR2_X1 _12998_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_05256_ ) );
AND3_X1 _12999_ ( .A1(_05256_ ), .A2(\IF_ID_inst [21] ), .A3(_05217_ ), .ZN(_05257_ ) );
NOR2_X1 _13000_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_05258_ ) );
NOR2_X1 _13001_ ( .A1(\IF_ID_inst [27] ), .A2(\IF_ID_inst [24] ), .ZN(_05259_ ) );
AND2_X1 _13002_ ( .A1(_05258_ ), .A2(_05259_ ), .ZN(_05260_ ) );
AND4_X1 _13003_ ( .A1(_05253_ ), .A2(_05255_ ), .A3(_05257_ ), .A4(_05260_ ), .ZN(_05261_ ) );
AOI221_X4 _13004_ ( .A(_05232_ ), .B1(_05233_ ), .B2(_05238_ ), .C1(_05250_ ), .C2(_05261_ ), .ZN(_05262_ ) );
NOR2_X1 _13005_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_05263_ ) );
AND3_X1 _13006_ ( .A1(_05203_ ), .A2(_05235_ ), .A3(_05263_ ), .ZN(_05264_ ) );
INV_X1 _13007_ ( .A(\IF_ID_inst [13] ), .ZN(_05265_ ) );
NOR2_X1 _13008_ ( .A1(_05265_ ), .A2(\IF_ID_inst [14] ), .ZN(_05266_ ) );
AND2_X1 _13009_ ( .A1(_05264_ ), .A2(_05266_ ), .ZN(_05267_ ) );
INV_X1 _13010_ ( .A(_05267_ ), .ZN(_05268_ ) );
NOR2_X1 _13011_ ( .A1(_05239_ ), .A2(\IF_ID_inst [6] ), .ZN(_05269_ ) );
AND3_X1 _13012_ ( .A1(_05203_ ), .A2(_05235_ ), .A3(_05269_ ), .ZN(_05270_ ) );
OAI21_X1 _13013_ ( .A(_05227_ ), .B1(_05264_ ), .B2(_05270_ ), .ZN(_05271_ ) );
AND2_X1 _13014_ ( .A1(_05268_ ), .A2(_05271_ ), .ZN(_05272_ ) );
AND3_X1 _13015_ ( .A1(_05251_ ), .A2(_05252_ ), .A3(_05256_ ), .ZN(_05273_ ) );
AND3_X1 _13016_ ( .A1(_05273_ ), .A2(_05214_ ), .A3(\IF_ID_inst [20] ), .ZN(_05274_ ) );
INV_X1 _13017_ ( .A(_05274_ ), .ZN(_05275_ ) );
NOR4_X1 _13018_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .A4(\IF_ID_inst [31] ), .ZN(_05276_ ) );
AND2_X1 _13019_ ( .A1(_05276_ ), .A2(_05260_ ), .ZN(_05277_ ) );
NAND2_X1 _13020_ ( .A1(_05250_ ), .A2(_05277_ ), .ZN(_05278_ ) );
OAI211_X1 _13021_ ( .A(_05262_ ), .B(_05272_ ), .C1(_05275_ ), .C2(_05278_ ), .ZN(_05279_ ) );
INV_X1 _13022_ ( .A(_05203_ ), .ZN(_05280_ ) );
INV_X1 _13023_ ( .A(\IF_ID_inst [4] ), .ZN(_05281_ ) );
NAND4_X1 _13024_ ( .A1(_05281_ ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_05282_ ) );
NOR2_X1 _13025_ ( .A1(_05280_ ), .A2(_05282_ ), .ZN(_05283_ ) );
AND2_X1 _13026_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_05284_ ) );
AND2_X1 _13027_ ( .A1(_05283_ ), .A2(_05284_ ), .ZN(_05285_ ) );
INV_X1 _13028_ ( .A(_05285_ ), .ZN(_05286_ ) );
NAND2_X1 _13029_ ( .A1(_05238_ ), .A2(\IF_ID_inst [14] ), .ZN(_05287_ ) );
AND3_X1 _13030_ ( .A1(_05200_ ), .A2(\IF_ID_inst [12] ), .A3(_05201_ ), .ZN(_05288_ ) );
NAND4_X1 _13031_ ( .A1(_05288_ ), .A2(_05265_ ), .A3(\IF_ID_inst [6] ), .A4(_05235_ ), .ZN(_05289_ ) );
NAND3_X1 _13032_ ( .A1(_05286_ ), .A2(_05287_ ), .A3(_05289_ ), .ZN(_05290_ ) );
NOR4_X1 _13033_ ( .A1(_05279_ ), .A2(_05245_ ), .A3(_05221_ ), .A4(_05290_ ), .ZN(_00209_ ) );
NOR4_X1 _13034_ ( .A1(_05279_ ), .A2(_05246_ ), .A3(_05221_ ), .A4(_05290_ ), .ZN(_00210_ ) );
NOR4_X1 _13035_ ( .A1(_05279_ ), .A2(_05247_ ), .A3(_05221_ ), .A4(_05290_ ), .ZN(_00211_ ) );
INV_X1 _13036_ ( .A(\IF_ID_inst [8] ), .ZN(_05291_ ) );
NOR4_X1 _13037_ ( .A1(_05279_ ), .A2(_05291_ ), .A3(_05221_ ), .A4(_05290_ ), .ZN(_00212_ ) );
NOR4_X1 _13038_ ( .A1(_05279_ ), .A2(_05240_ ), .A3(_05221_ ), .A4(_05290_ ), .ZN(_00213_ ) );
AND4_X1 _13039_ ( .A1(\IF_ID_inst [6] ), .A2(_05203_ ), .A3(_05240_ ), .A4(_05243_ ), .ZN(_05292_ ) );
NOR4_X1 _13040_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_05293_ ) );
AND3_X1 _13041_ ( .A1(_05292_ ), .A2(_05249_ ), .A3(_05293_ ), .ZN(_05294_ ) );
AND2_X1 _13042_ ( .A1(_05274_ ), .A2(_05277_ ), .ZN(_05295_ ) );
NAND2_X1 _13043_ ( .A1(_05294_ ), .A2(_05295_ ), .ZN(_05296_ ) );
INV_X1 _13044_ ( .A(_05233_ ), .ZN(_05297_ ) );
AND3_X1 _13045_ ( .A1(_05228_ ), .A2(\IF_ID_inst [12] ), .A3(_05196_ ), .ZN(_05298_ ) );
NAND2_X1 _13046_ ( .A1(_05231_ ), .A2(_05298_ ), .ZN(_05299_ ) );
OAI21_X1 _13047_ ( .A(_05296_ ), .B1(_05297_ ), .B2(_05299_ ), .ZN(_05300_ ) );
INV_X1 _13048_ ( .A(\IF_ID_inst [19] ), .ZN(_05301_ ) );
INV_X1 _13049_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_05302_ ) );
AND2_X1 _13050_ ( .A1(_05235_ ), .A2(_05302_ ), .ZN(_05303_ ) );
AND2_X1 _13051_ ( .A1(_05303_ ), .A2(_05230_ ), .ZN(_05304_ ) );
BUF_X2 _13052_ ( .A(_05304_ ), .Z(_05305_ ) );
NAND3_X1 _13053_ ( .A1(\IF_ID_inst [2] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [1] ), .ZN(_05306_ ) );
NOR2_X1 _13054_ ( .A1(_05306_ ), .A2(\IF_ID_inst [3] ), .ZN(_05307_ ) );
NOR2_X1 _13055_ ( .A1(_05281_ ), .A2(\IF_ID_inst [6] ), .ZN(_05308_ ) );
AND2_X1 _13056_ ( .A1(_05307_ ), .A2(_05308_ ), .ZN(_05309_ ) );
NOR2_X1 _13057_ ( .A1(_05305_ ), .A2(_05309_ ), .ZN(_05310_ ) );
NAND4_X1 _13058_ ( .A1(_05203_ ), .A2(_05242_ ), .A3(_05243_ ), .A4(_05227_ ), .ZN(_05311_ ) );
NOR3_X1 _13059_ ( .A1(_05311_ ), .A2(\IF_ID_inst [8] ), .A3(_05248_ ), .ZN(_05312_ ) );
INV_X1 _13060_ ( .A(_05312_ ), .ZN(_05313_ ) );
AND4_X1 _13061_ ( .A1(_05253_ ), .A2(_05255_ ), .A3(_05257_ ), .A4(_05260_ ), .ZN(_05314_ ) );
INV_X1 _13062_ ( .A(_05314_ ), .ZN(_05315_ ) );
OAI21_X1 _13063_ ( .A(_05310_ ), .B1(_05313_ ), .B2(_05315_ ), .ZN(_05316_ ) );
BUF_X4 _13064_ ( .A(_05211_ ), .Z(_05317_ ) );
NOR4_X1 _13065_ ( .A1(_05300_ ), .A2(_05301_ ), .A3(_05316_ ), .A4(_05317_ ), .ZN(_00214_ ) );
INV_X1 _13066_ ( .A(\IF_ID_inst [18] ), .ZN(_05318_ ) );
NOR4_X1 _13067_ ( .A1(_05300_ ), .A2(_05318_ ), .A3(_05316_ ), .A4(_05317_ ), .ZN(_00215_ ) );
INV_X1 _13068_ ( .A(\IF_ID_inst [17] ), .ZN(_05319_ ) );
NOR4_X1 _13069_ ( .A1(_05300_ ), .A2(_05319_ ), .A3(_05316_ ), .A4(_05317_ ), .ZN(_00216_ ) );
AND2_X2 _13070_ ( .A1(_05203_ ), .A2(_05263_ ), .ZN(_05320_ ) );
NOR2_X1 _13071_ ( .A1(_05281_ ), .A2(\IF_ID_inst [5] ), .ZN(_05321_ ) );
AND2_X2 _13072_ ( .A1(_05320_ ), .A2(_05321_ ), .ZN(_05322_ ) );
INV_X1 _13073_ ( .A(_05322_ ), .ZN(_05323_ ) );
OAI211_X1 _13074_ ( .A(_05236_ ), .B(_05233_ ), .C1(_05307_ ), .C2(_05237_ ), .ZN(_05324_ ) );
AND4_X1 _13075_ ( .A1(\IF_ID_inst [4] ), .A2(_05234_ ), .A3(_05196_ ), .A4(\IF_ID_inst [12] ), .ZN(_05325_ ) );
AND2_X2 _13076_ ( .A1(_05203_ ), .A2(_05325_ ), .ZN(_05326_ ) );
NAND2_X1 _13077_ ( .A1(_05326_ ), .A2(\IF_ID_inst [13] ), .ZN(_05327_ ) );
AND3_X1 _13078_ ( .A1(_05323_ ), .A2(_05324_ ), .A3(_05327_ ), .ZN(_05328_ ) );
INV_X1 _13079_ ( .A(\IF_ID_inst [14] ), .ZN(_05329_ ) );
NOR2_X1 _13080_ ( .A1(_05329_ ), .A2(\IF_ID_inst [13] ), .ZN(_05330_ ) );
AND2_X1 _13081_ ( .A1(_05330_ ), .A2(_05258_ ), .ZN(_05331_ ) );
NOR3_X1 _13082_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_05332_ ) );
AND3_X1 _13083_ ( .A1(_05332_ ), .A2(_05220_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05333_ ) );
NAND3_X1 _13084_ ( .A1(_05219_ ), .A2(_05220_ ), .A3(\IF_ID_inst [30] ), .ZN(_05334_ ) );
INV_X1 _13085_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05335_ ) );
NOR3_X1 _13086_ ( .A1(_05334_ ), .A2(\IF_ID_inst [29] ), .A3(_05335_ ), .ZN(_05336_ ) );
OAI21_X1 _13087_ ( .A(_05331_ ), .B1(_05333_ ), .B2(_05336_ ), .ZN(_05337_ ) );
INV_X1 _13088_ ( .A(_05326_ ), .ZN(_05338_ ) );
NOR2_X1 _13089_ ( .A1(_05337_ ), .A2(_05338_ ), .ZN(_05339_ ) );
INV_X1 _13090_ ( .A(_05339_ ), .ZN(_05340_ ) );
AND2_X1 _13091_ ( .A1(_05320_ ), .A2(_05228_ ), .ZN(_05341_ ) );
AND2_X1 _13092_ ( .A1(_05341_ ), .A2(_05266_ ), .ZN(_05342_ ) );
INV_X1 _13093_ ( .A(_05342_ ), .ZN(_05343_ ) );
AND4_X1 _13094_ ( .A1(_05272_ ), .A2(_05328_ ), .A3(_05340_ ), .A4(_05343_ ), .ZN(_05344_ ) );
AND3_X1 _13095_ ( .A1(_05286_ ), .A2(_05287_ ), .A3(_05289_ ), .ZN(_05345_ ) );
NOR2_X1 _13096_ ( .A1(_05300_ ), .A2(_05316_ ), .ZN(_05346_ ) );
NAND2_X1 _13097_ ( .A1(_05341_ ), .A2(_05265_ ), .ZN(_05347_ ) );
AND2_X2 _13098_ ( .A1(_05320_ ), .A2(_05243_ ), .ZN(_05348_ ) );
AND2_X1 _13099_ ( .A1(_05332_ ), .A2(_05220_ ), .ZN(_05349_ ) );
AND4_X1 _13100_ ( .A1(_05329_ ), .A2(_05258_ ), .A3(\IF_ID_inst [13] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05350_ ) );
AND2_X1 _13101_ ( .A1(_05349_ ), .A2(_05350_ ), .ZN(_05351_ ) );
NAND2_X1 _13102_ ( .A1(_05348_ ), .A2(_05351_ ), .ZN(_05352_ ) );
AND3_X1 _13103_ ( .A1(_05298_ ), .A2(_05237_ ), .A3(_05265_ ), .ZN(_05353_ ) );
INV_X1 _13104_ ( .A(_05353_ ), .ZN(_05354_ ) );
AND2_X1 _13105_ ( .A1(_05227_ ), .A2(_05258_ ), .ZN(_05355_ ) );
NAND4_X1 _13106_ ( .A1(_05320_ ), .A2(_05243_ ), .A3(_05336_ ), .A4(_05355_ ), .ZN(_05356_ ) );
NAND4_X1 _13107_ ( .A1(_05347_ ), .A2(_05352_ ), .A3(_05354_ ), .A4(_05356_ ), .ZN(_05357_ ) );
AND3_X1 _13108_ ( .A1(_05326_ ), .A2(_05333_ ), .A3(_05355_ ), .ZN(_05358_ ) );
NOR3_X1 _13109_ ( .A1(_05357_ ), .A2(_05216_ ), .A3(_05358_ ), .ZN(_05359_ ) );
NAND4_X1 _13110_ ( .A1(_05344_ ), .A2(_05345_ ), .A3(_05346_ ), .A4(_05359_ ), .ZN(_05360_ ) );
AND2_X1 _13111_ ( .A1(_05333_ ), .A2(_05331_ ), .ZN(_05361_ ) );
AND2_X1 _13112_ ( .A1(_05348_ ), .A2(_05361_ ), .ZN(_05362_ ) );
INV_X1 _13113_ ( .A(_05362_ ), .ZN(_05363_ ) );
AND2_X2 _13114_ ( .A1(_05333_ ), .A2(_05355_ ), .ZN(_05364_ ) );
NAND3_X1 _13115_ ( .A1(_05364_ ), .A2(_05243_ ), .A3(_05320_ ), .ZN(_05365_ ) );
AND3_X1 _13116_ ( .A1(_05349_ ), .A2(_05284_ ), .A3(_05258_ ), .ZN(_05366_ ) );
AND3_X1 _13117_ ( .A1(_05196_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_05367_ ) );
AND2_X1 _13118_ ( .A1(_05288_ ), .A2(_05367_ ), .ZN(_05368_ ) );
OAI211_X1 _13119_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B(_05366_ ), .C1(_05348_ ), .C2(_05368_ ), .ZN(_05369_ ) );
AND3_X1 _13120_ ( .A1(_05363_ ), .A2(_05365_ ), .A3(_05369_ ), .ZN(_05370_ ) );
AND3_X1 _13121_ ( .A1(_05368_ ), .A2(_05331_ ), .A3(_05336_ ), .ZN(_05371_ ) );
INV_X1 _13122_ ( .A(_05371_ ), .ZN(_05372_ ) );
NOR3_X1 _13123_ ( .A1(_05361_ ), .A2(_05364_ ), .A3(_05351_ ), .ZN(_05373_ ) );
INV_X1 _13124_ ( .A(_05368_ ), .ZN(_05374_ ) );
NOR2_X1 _13125_ ( .A1(_05373_ ), .A2(_05374_ ), .ZN(_05375_ ) );
INV_X1 _13126_ ( .A(_05375_ ), .ZN(_05376_ ) );
NAND3_X1 _13127_ ( .A1(_05370_ ), .A2(_05372_ ), .A3(_05376_ ), .ZN(_05377_ ) );
NOR2_X1 _13128_ ( .A1(_05360_ ), .A2(_05377_ ), .ZN(_05378_ ) );
XNOR2_X1 _13129_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_05379_ ) );
XNOR2_X1 _13130_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_05380_ ) );
XNOR2_X1 _13131_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_05381_ ) );
XNOR2_X1 _13132_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_05382_ ) );
AND4_X1 _13133_ ( .A1(_05379_ ), .A2(_05380_ ), .A3(_05381_ ), .A4(_05382_ ), .ZN(_05383_ ) );
XNOR2_X1 _13134_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_05384_ ) );
XNOR2_X1 _13135_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_05385_ ) );
XNOR2_X1 _13136_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_05386_ ) );
XNOR2_X1 _13137_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_05387_ ) );
AND4_X1 _13138_ ( .A1(_05384_ ), .A2(_05385_ ), .A3(_05386_ ), .A4(_05387_ ), .ZN(_05388_ ) );
XNOR2_X1 _13139_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_05389_ ) );
XNOR2_X1 _13140_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_05390_ ) );
XNOR2_X1 _13141_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_05391_ ) );
XNOR2_X1 _13142_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_05392_ ) );
AND4_X1 _13143_ ( .A1(_05389_ ), .A2(_05390_ ), .A3(_05391_ ), .A4(_05392_ ), .ZN(_05393_ ) );
XNOR2_X1 _13144_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_05394_ ) );
XNOR2_X1 _13145_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_05395_ ) );
XNOR2_X1 _13146_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_05396_ ) );
XNOR2_X1 _13147_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_05397_ ) );
AND4_X1 _13148_ ( .A1(_05394_ ), .A2(_05395_ ), .A3(_05396_ ), .A4(_05397_ ), .ZN(_05398_ ) );
AND4_X1 _13149_ ( .A1(_05383_ ), .A2(_05388_ ), .A3(_05393_ ), .A4(_05398_ ), .ZN(_05399_ ) );
XNOR2_X1 _13150_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_05400_ ) );
XNOR2_X1 _13151_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_05401_ ) );
XNOR2_X1 _13152_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_05402_ ) );
XNOR2_X1 _13153_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_05403_ ) );
AND4_X1 _13154_ ( .A1(_05400_ ), .A2(_05401_ ), .A3(_05402_ ), .A4(_05403_ ), .ZN(_05404_ ) );
XNOR2_X1 _13155_ ( .A(fanout_net_9 ), .B(\myexu.pc_jump [3] ), .ZN(_05405_ ) );
XNOR2_X1 _13156_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_05406_ ) );
XNOR2_X1 _13157_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_05407_ ) );
INV_X1 _13158_ ( .A(\IF_ID_pc [2] ), .ZN(_05408_ ) );
AOI22_X1 _13159_ ( .A1(_01829_ ), .A2(\myexu.pc_jump [25] ), .B1(_05408_ ), .B2(\myexu.pc_jump [2] ), .ZN(_05409_ ) );
AND4_X1 _13160_ ( .A1(_05405_ ), .A2(_05406_ ), .A3(_05407_ ), .A4(_05409_ ), .ZN(_05410_ ) );
INV_X1 _13161_ ( .A(\myexu.pc_jump [1] ), .ZN(_05411_ ) );
NOR2_X1 _13162_ ( .A1(_05411_ ), .A2(\IF_ID_pc [1] ), .ZN(_05412_ ) );
INV_X1 _13163_ ( .A(fanout_net_13 ), .ZN(_05413_ ) );
AOI21_X1 _13164_ ( .A(_05412_ ), .B1(_05413_ ), .B2(\myexu.pc_jump [4] ), .ZN(_05414_ ) );
XNOR2_X1 _13165_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_05415_ ) );
XNOR2_X1 _13166_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_05416_ ) );
INV_X1 _13167_ ( .A(\myexu.pc_jump [2] ), .ZN(_05417_ ) );
AOI22_X1 _13168_ ( .A1(_05411_ ), .A2(\IF_ID_pc [1] ), .B1(_05417_ ), .B2(\IF_ID_pc [2] ), .ZN(_05418_ ) );
NAND4_X1 _13169_ ( .A1(_05414_ ), .A2(_05415_ ), .A3(_05416_ ), .A4(_05418_ ), .ZN(_05419_ ) );
XNOR2_X1 _13170_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_05420_ ) );
INV_X1 _13171_ ( .A(\myexu.pc_jump [21] ), .ZN(_05421_ ) );
OAI221_X1 _13172_ ( .A(_05420_ ), .B1(\IF_ID_pc [21] ), .B2(_05421_ ), .C1(_01829_ ), .C2(\myexu.pc_jump [25] ), .ZN(_05422_ ) );
AOI22_X1 _13173_ ( .A1(_02074_ ), .A2(\myexu.pc_jump [29] ), .B1(_05421_ ), .B2(\IF_ID_pc [21] ), .ZN(_05423_ ) );
OAI221_X1 _13174_ ( .A(_05423_ ), .B1(_05413_ ), .B2(\myexu.pc_jump [4] ), .C1(_02074_ ), .C2(\myexu.pc_jump [29] ), .ZN(_05424_ ) );
NOR3_X1 _13175_ ( .A1(_05419_ ), .A2(_05422_ ), .A3(_05424_ ), .ZN(_05425_ ) );
AND4_X2 _13176_ ( .A1(_05399_ ), .A2(_05404_ ), .A3(_05410_ ), .A4(_05425_ ), .ZN(_05426_ ) );
NOR2_X2 _13177_ ( .A1(_05426_ ), .A2(_02117_ ), .ZN(_05427_ ) );
INV_X1 _13178_ ( .A(\myifu.state [1] ), .ZN(_05428_ ) );
NOR2_X1 _13179_ ( .A1(_05428_ ), .A2(fanout_net_44 ), .ZN(_05429_ ) );
INV_X1 _13180_ ( .A(_05429_ ), .ZN(_05430_ ) );
NOR2_X1 _13181_ ( .A1(_05427_ ), .A2(_05430_ ), .ZN(_05431_ ) );
AND2_X2 _13182_ ( .A1(_05431_ ), .A2(IDU_ready_IFU ), .ZN(_05432_ ) );
INV_X1 _13183_ ( .A(_05432_ ), .ZN(_05433_ ) );
BUF_X4 _13184_ ( .A(_05433_ ), .Z(_05434_ ) );
AOI211_X1 _13185_ ( .A(_05378_ ), .B(_05434_ ), .C1(\IF_ID_inst [18] ), .C2(_05346_ ), .ZN(_05435_ ) );
NOR2_X1 _13186_ ( .A1(_05433_ ), .A2(_05378_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _13187_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_05436_ ) );
AOI211_X1 _13188_ ( .A(_05317_ ), .B(_05435_ ), .C1(_02187_ ), .C2(_05436_ ), .ZN(_00217_ ) );
INV_X1 _13189_ ( .A(\IF_ID_inst [16] ), .ZN(_05437_ ) );
NOR4_X1 _13190_ ( .A1(_05300_ ), .A2(_05437_ ), .A3(_05316_ ), .A4(_05317_ ), .ZN(_00218_ ) );
BUF_X4 _13191_ ( .A(_05378_ ), .Z(_05438_ ) );
INV_X1 _13192_ ( .A(_05438_ ), .ZN(_05439_ ) );
NAND4_X1 _13193_ ( .A1(_05439_ ), .A2(\IF_ID_inst [17] ), .A3(_05346_ ), .A4(_05432_ ), .ZN(_05440_ ) );
OAI21_X1 _13194_ ( .A(\ID_EX_rs1 [2] ), .B1(_05434_ ), .B2(_05438_ ), .ZN(_05441_ ) );
AOI21_X1 _13195_ ( .A(_05215_ ), .B1(_05440_ ), .B2(_05441_ ), .ZN(_00219_ ) );
NOR4_X1 _13196_ ( .A1(_05300_ ), .A2(_05241_ ), .A3(_05316_ ), .A4(_05317_ ), .ZN(_00220_ ) );
OAI21_X1 _13197_ ( .A(_05210_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [1] ), .ZN(_05442_ ) );
OR3_X1 _13198_ ( .A1(_05300_ ), .A2(_05437_ ), .A3(_05316_ ), .ZN(_05443_ ) );
AOI21_X1 _13199_ ( .A(_05442_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(_05443_ ), .ZN(_00221_ ) );
AND2_X1 _13200_ ( .A1(_05322_ ), .A2(_05266_ ), .ZN(_05444_ ) );
NOR2_X1 _13201_ ( .A1(_05444_ ), .A2(_05309_ ), .ZN(_05445_ ) );
NOR2_X1 _13202_ ( .A1(_05339_ ), .A2(_05358_ ), .ZN(_05446_ ) );
AND2_X1 _13203_ ( .A1(_05445_ ), .A2(_05446_ ), .ZN(_05447_ ) );
AND3_X1 _13204_ ( .A1(_05321_ ), .A2(_05200_ ), .A3(_05201_ ), .ZN(_05448_ ) );
AND2_X2 _13205_ ( .A1(_05448_ ), .A2(_05269_ ), .ZN(_05449_ ) );
AOI22_X1 _13206_ ( .A1(_05322_ ), .A2(\IF_ID_inst [14] ), .B1(\IF_ID_inst [13] ), .B2(_05449_ ), .ZN(_05450_ ) );
AND3_X1 _13207_ ( .A1(_05450_ ), .A2(_05347_ ), .A3(_05354_ ), .ZN(_05451_ ) );
AND3_X1 _13208_ ( .A1(_05197_ ), .A2(_05235_ ), .A3(_05227_ ), .ZN(_05452_ ) );
AND2_X1 _13209_ ( .A1(_05452_ ), .A2(_05307_ ), .ZN(_05453_ ) );
NOR2_X1 _13210_ ( .A1(_05453_ ), .A2(_05305_ ), .ZN(_05454_ ) );
INV_X1 _13211_ ( .A(_05454_ ), .ZN(_05455_ ) );
NOR2_X1 _13212_ ( .A1(_05342_ ), .A2(_05455_ ), .ZN(_05456_ ) );
AOI21_X1 _13213_ ( .A(_05232_ ), .B1(_05312_ ), .B2(_05314_ ), .ZN(_05457_ ) );
AND4_X1 _13214_ ( .A1(_05447_ ), .A2(_05451_ ), .A3(_05456_ ), .A4(_05457_ ), .ZN(_05458_ ) );
BUF_X2 _13215_ ( .A(_05210_ ), .Z(_05459_ ) );
NAND3_X1 _13216_ ( .A1(_05312_ ), .A2(_05274_ ), .A3(_05277_ ), .ZN(_05460_ ) );
OAI211_X1 _13217_ ( .A(_05460_ ), .B(_05207_ ), .C1(_05297_ ), .C2(_05323_ ), .ZN(_05461_ ) );
INV_X1 _13218_ ( .A(_05461_ ), .ZN(_05462_ ) );
AND4_X1 _13219_ ( .A1(\IF_ID_inst [24] ), .A2(_05458_ ), .A3(_05459_ ), .A4(_05462_ ), .ZN(_00222_ ) );
AOI211_X1 _13220_ ( .A(_05434_ ), .B(_05438_ ), .C1(\IF_ID_inst [15] ), .C2(_05346_ ), .ZN(_05463_ ) );
AOI21_X1 _13221_ ( .A(\ID_EX_rs1 [0] ), .B1(_05439_ ), .B2(_05432_ ), .ZN(_05464_ ) );
NOR3_X1 _13222_ ( .A1(_05463_ ), .A2(_05215_ ), .A3(_05464_ ), .ZN(_00223_ ) );
AND4_X1 _13223_ ( .A1(\IF_ID_inst [23] ), .A2(_05458_ ), .A3(_05459_ ), .A4(_05462_ ), .ZN(_00224_ ) );
AND4_X1 _13224_ ( .A1(\IF_ID_inst [22] ), .A2(_05458_ ), .A3(_05459_ ), .A4(_05462_ ), .ZN(_00225_ ) );
AND2_X1 _13225_ ( .A1(_05458_ ), .A2(_05462_ ), .ZN(_05465_ ) );
AOI211_X1 _13226_ ( .A(_05378_ ), .B(_05434_ ), .C1(_05465_ ), .C2(\IF_ID_inst [23] ), .ZN(_05466_ ) );
AOI211_X1 _13227_ ( .A(_05317_ ), .B(_05466_ ), .C1(_03233_ ), .C2(_05436_ ), .ZN(_00226_ ) );
AND4_X1 _13228_ ( .A1(\IF_ID_inst [21] ), .A2(_05458_ ), .A3(_05459_ ), .A4(_05462_ ), .ZN(_00227_ ) );
AOI211_X1 _13229_ ( .A(_05438_ ), .B(_05434_ ), .C1(\IF_ID_inst [22] ), .C2(_05465_ ), .ZN(_05467_ ) );
AOI21_X1 _13230_ ( .A(\ID_EX_rs2 [2] ), .B1(_05439_ ), .B2(_05432_ ), .ZN(_05468_ ) );
NOR3_X1 _13231_ ( .A1(_05467_ ), .A2(_05215_ ), .A3(_05468_ ), .ZN(_00228_ ) );
AND4_X1 _13232_ ( .A1(\IF_ID_inst [20] ), .A2(_05458_ ), .A3(_05459_ ), .A4(_05462_ ), .ZN(_00229_ ) );
AOI211_X1 _13233_ ( .A(_05438_ ), .B(_05434_ ), .C1(\IF_ID_inst [21] ), .C2(_05465_ ), .ZN(_05469_ ) );
AOI21_X1 _13234_ ( .A(\ID_EX_rs2 [1] ), .B1(_05439_ ), .B2(_05432_ ), .ZN(_05470_ ) );
NOR3_X1 _13235_ ( .A1(_05469_ ), .A2(_05215_ ), .A3(_05470_ ), .ZN(_00230_ ) );
AND4_X1 _13236_ ( .A1(_02116_ ), .A2(_05229_ ), .A3(_05210_ ), .A4(_05231_ ), .ZN(_00231_ ) );
AOI211_X1 _13237_ ( .A(_05438_ ), .B(_05434_ ), .C1(\IF_ID_inst [20] ), .C2(_05465_ ), .ZN(_05471_ ) );
AOI21_X1 _13238_ ( .A(\ID_EX_rs2 [0] ), .B1(_05439_ ), .B2(_05432_ ), .ZN(_05472_ ) );
NOR3_X1 _13239_ ( .A1(_05471_ ), .A2(_05215_ ), .A3(_05472_ ), .ZN(_00232_ ) );
XNOR2_X1 _13240_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_05473_ ) );
XNOR2_X1 _13241_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_05474_ ) );
XNOR2_X1 _13242_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_05475_ ) );
XNOR2_X1 _13243_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_05476_ ) );
NAND4_X1 _13244_ ( .A1(_05473_ ), .A2(_05474_ ), .A3(_05475_ ), .A4(_05476_ ), .ZN(_05477_ ) );
XOR2_X1 _13245_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .Z(_05478_ ) );
NOR2_X1 _13246_ ( .A1(_05477_ ), .A2(_05478_ ), .ZN(_05479_ ) );
AND2_X1 _13247_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_05480_ ) );
AND2_X1 _13248_ ( .A1(_05480_ ), .A2(_05179_ ), .ZN(_05481_ ) );
AND2_X1 _13249_ ( .A1(_05479_ ), .A2(_05481_ ), .ZN(_05482_ ) );
XNOR2_X1 _13250_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_05483_ ) );
XNOR2_X1 _13251_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_05484_ ) );
XNOR2_X1 _13252_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_05485_ ) );
AND4_X1 _13253_ ( .A1(_05481_ ), .A2(_05483_ ), .A3(_05484_ ), .A4(_05485_ ), .ZN(_05486_ ) );
XNOR2_X1 _13254_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_05487_ ) );
XNOR2_X1 _13255_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_05488_ ) );
AND3_X1 _13256_ ( .A1(_05486_ ), .A2(_05487_ ), .A3(_05488_ ), .ZN(_05489_ ) );
OR2_X1 _13257_ ( .A1(_05482_ ), .A2(_05489_ ), .ZN(_05490_ ) );
AND2_X1 _13258_ ( .A1(_05346_ ), .A2(_05490_ ), .ZN(_05491_ ) );
INV_X1 _13259_ ( .A(_05444_ ), .ZN(_05492_ ) );
NAND2_X1 _13260_ ( .A1(_05326_ ), .A2(_05266_ ), .ZN(_05493_ ) );
NAND2_X1 _13261_ ( .A1(_05326_ ), .A2(_05284_ ), .ZN(_05494_ ) );
INV_X1 _13262_ ( .A(_05284_ ), .ZN(_05495_ ) );
NAND2_X1 _13263_ ( .A1(_05341_ ), .A2(_05495_ ), .ZN(_05496_ ) );
NAND4_X1 _13264_ ( .A1(_05492_ ), .A2(_05493_ ), .A3(_05494_ ), .A4(_05496_ ), .ZN(_05497_ ) );
INV_X1 _13265_ ( .A(_05266_ ), .ZN(_05498_ ) );
NAND2_X1 _13266_ ( .A1(_05322_ ), .A2(_05498_ ), .ZN(_05499_ ) );
INV_X1 _13267_ ( .A(_05453_ ), .ZN(_05500_ ) );
NAND3_X1 _13268_ ( .A1(_05499_ ), .A2(_05500_ ), .A3(_05354_ ), .ZN(_05501_ ) );
NOR2_X1 _13269_ ( .A1(_05497_ ), .A2(_05501_ ), .ZN(_05502_ ) );
INV_X1 _13270_ ( .A(_05502_ ), .ZN(_05503_ ) );
NOR3_X1 _13271_ ( .A1(_05491_ ), .A2(_05503_ ), .A3(_05216_ ), .ZN(_05504_ ) );
BUF_X2 _13272_ ( .A(_05502_ ), .Z(_05505_ ) );
AOI21_X1 _13273_ ( .A(_05482_ ), .B1(_05505_ ), .B2(_05208_ ), .ZN(_05506_ ) );
INV_X1 _13274_ ( .A(IDU_ready_IFU ), .ZN(_05507_ ) );
NOR4_X1 _13275_ ( .A1(_05504_ ), .A2(_05506_ ), .A3(_05507_ ), .A4(_05317_ ), .ZN(_00233_ ) );
AND2_X1 _13276_ ( .A1(_05250_ ), .A2(_05261_ ), .ZN(_05508_ ) );
AND3_X1 _13277_ ( .A1(_05236_ ), .A2(_05237_ ), .A3(_05233_ ), .ZN(_05509_ ) );
AOI21_X1 _13278_ ( .A(_05509_ ), .B1(_05233_ ), .B2(_05283_ ), .ZN(_05510_ ) );
OAI21_X1 _13279_ ( .A(\IF_ID_inst [14] ), .B1(_05283_ ), .B2(_05238_ ), .ZN(_05511_ ) );
NAND2_X1 _13280_ ( .A1(_05510_ ), .A2(_05511_ ), .ZN(_05512_ ) );
NOR4_X1 _13281_ ( .A1(_05508_ ), .A2(_05512_ ), .A3(_05232_ ), .A4(_05455_ ), .ZN(_05513_ ) );
NAND4_X1 _13282_ ( .A1(_05244_ ), .A2(_05217_ ), .A3(_05237_ ), .A4(_05249_ ), .ZN(_05514_ ) );
NAND4_X1 _13283_ ( .A1(_05273_ ), .A2(_05260_ ), .A3(_05276_ ), .A4(_05214_ ), .ZN(_05515_ ) );
NOR2_X1 _13284_ ( .A1(_05514_ ), .A2(_05515_ ), .ZN(_05516_ ) );
NOR2_X1 _13285_ ( .A1(_05516_ ), .A2(_05216_ ), .ZN(_05517_ ) );
AOI21_X1 _13286_ ( .A(_05215_ ), .B1(_05513_ ), .B2(_05517_ ), .ZN(_00234_ ) );
AND2_X1 _13287_ ( .A1(_05298_ ), .A2(_05237_ ), .ZN(_05518_ ) );
NAND2_X1 _13288_ ( .A1(_05518_ ), .A2(_05233_ ), .ZN(_05519_ ) );
AND3_X1 _13289_ ( .A1(_05518_ ), .A2(\IF_ID_inst [14] ), .A3(_05265_ ), .ZN(_05520_ ) );
INV_X1 _13290_ ( .A(_05520_ ), .ZN(_05521_ ) );
AND4_X1 _13291_ ( .A1(_05272_ ), .A2(_05519_ ), .A3(_05496_ ), .A4(_05521_ ), .ZN(_05522_ ) );
AOI21_X1 _13292_ ( .A(_05212_ ), .B1(_05522_ ), .B2(_05517_ ), .ZN(_00235_ ) );
OAI211_X1 _13293_ ( .A(_05243_ ), .B(_05320_ ), .C1(_05361_ ), .C2(_05364_ ), .ZN(_05523_ ) );
AND3_X1 _13294_ ( .A1(_05243_ ), .A2(_05200_ ), .A3(_05201_ ), .ZN(_05524_ ) );
AND2_X1 _13295_ ( .A1(_05524_ ), .A2(_05269_ ), .ZN(_05525_ ) );
INV_X1 _13296_ ( .A(_05525_ ), .ZN(_05526_ ) );
OAI21_X1 _13297_ ( .A(_05523_ ), .B1(_05373_ ), .B2(_05526_ ), .ZN(_05527_ ) );
OAI211_X1 _13298_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B(_05366_ ), .C1(_05348_ ), .C2(_05525_ ), .ZN(_05528_ ) );
INV_X1 _13299_ ( .A(_05528_ ), .ZN(_05529_ ) );
OR2_X1 _13300_ ( .A1(_05527_ ), .A2(_05529_ ), .ZN(_05530_ ) );
NAND4_X1 _13301_ ( .A1(_05320_ ), .A2(_05243_ ), .A3(_05336_ ), .A4(_05355_ ), .ZN(_05531_ ) );
AND2_X1 _13302_ ( .A1(_05352_ ), .A2(_05531_ ), .ZN(_05532_ ) );
NAND4_X1 _13303_ ( .A1(_05456_ ), .A2(_05532_ ), .A3(_05347_ ), .A4(_05354_ ), .ZN(_05533_ ) );
AND3_X1 _13304_ ( .A1(_05525_ ), .A2(_05331_ ), .A3(_05336_ ), .ZN(_05534_ ) );
INV_X1 _13305_ ( .A(_05534_ ), .ZN(_05535_ ) );
AND4_X1 _13306_ ( .A1(_05214_ ), .A2(_05273_ ), .A3(_05260_ ), .A4(_05276_ ), .ZN(_05536_ ) );
NAND3_X1 _13307_ ( .A1(_05312_ ), .A2(_05217_ ), .A3(_05536_ ), .ZN(_05537_ ) );
NAND2_X1 _13308_ ( .A1(_05535_ ), .A2(_05537_ ), .ZN(_05538_ ) );
INV_X1 _13309_ ( .A(_05449_ ), .ZN(_05539_ ) );
OAI21_X1 _13310_ ( .A(_05499_ ), .B1(_05265_ ), .B2(_05539_ ), .ZN(_05540_ ) );
NOR4_X1 _13311_ ( .A1(_05530_ ), .A2(_05533_ ), .A3(_05538_ ), .A4(_05540_ ), .ZN(_05541_ ) );
AOI21_X1 _13312_ ( .A(_05212_ ), .B1(_05541_ ), .B2(_05447_ ), .ZN(_00236_ ) );
AOI221_X4 _13313_ ( .A(_05232_ ), .B1(\IF_ID_inst [13] ), .B2(_05326_ ), .C1(_05322_ ), .C2(_05498_ ), .ZN(_05542_ ) );
AOI21_X1 _13314_ ( .A(_05212_ ), .B1(_05447_ ), .B2(_05542_ ), .ZN(_00237_ ) );
AND2_X1 _13315_ ( .A1(_05348_ ), .A2(_05351_ ), .ZN(_05543_ ) );
AND4_X1 _13316_ ( .A1(_05243_ ), .A2(_05320_ ), .A3(_05336_ ), .A4(_05355_ ), .ZN(_05544_ ) );
NOR4_X1 _13317_ ( .A1(_05508_ ), .A2(_05543_ ), .A3(_05267_ ), .A4(_05544_ ), .ZN(_05545_ ) );
AOI21_X1 _13318_ ( .A(_05212_ ), .B1(_05545_ ), .B2(_05445_ ), .ZN(_00238_ ) );
NAND2_X1 _13319_ ( .A1(_05364_ ), .A2(_05449_ ), .ZN(_05546_ ) );
AND2_X1 _13320_ ( .A1(_05336_ ), .A2(_05331_ ), .ZN(_05547_ ) );
NAND2_X1 _13321_ ( .A1(_05547_ ), .A2(_05449_ ), .ZN(_05548_ ) );
NAND4_X1 _13322_ ( .A1(_05333_ ), .A2(_05448_ ), .A3(_05269_ ), .A4(_05331_ ), .ZN(_05549_ ) );
NAND3_X1 _13323_ ( .A1(_05546_ ), .A2(_05548_ ), .A3(_05549_ ), .ZN(_05550_ ) );
AND2_X1 _13324_ ( .A1(_05283_ ), .A2(\IF_ID_inst [14] ), .ZN(_05551_ ) );
AND3_X1 _13325_ ( .A1(_05237_ ), .A2(\IF_ID_inst [13] ), .A3(_05205_ ), .ZN(_05552_ ) );
NOR3_X1 _13326_ ( .A1(_05550_ ), .A2(_05551_ ), .A3(_05552_ ), .ZN(_05553_ ) );
INV_X1 _13327_ ( .A(_05309_ ), .ZN(_05554_ ) );
OAI21_X1 _13328_ ( .A(_05266_ ), .B1(_05341_ ), .B2(_05449_ ), .ZN(_05555_ ) );
AND4_X1 _13329_ ( .A1(_05268_ ), .A2(_05553_ ), .A3(_05554_ ), .A4(_05555_ ), .ZN(_05556_ ) );
NOR2_X1 _13330_ ( .A1(_05373_ ), .A2(_05526_ ), .ZN(_05557_ ) );
NOR2_X1 _13331_ ( .A1(_05557_ ), .A2(_05534_ ), .ZN(_05558_ ) );
AOI21_X1 _13332_ ( .A(_05212_ ), .B1(_05556_ ), .B2(_05558_ ), .ZN(_00239_ ) );
AOI21_X1 _13333_ ( .A(_05337_ ), .B1(_05374_ ), .B2(_05338_ ), .ZN(_05559_ ) );
AND2_X1 _13334_ ( .A1(_05366_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05560_ ) );
AND2_X1 _13335_ ( .A1(_05560_ ), .A2(_05348_ ), .ZN(_05561_ ) );
OR2_X1 _13336_ ( .A1(_05561_ ), .A2(_05520_ ), .ZN(_05562_ ) );
AOI211_X1 _13337_ ( .A(_05559_ ), .B(_05562_ ), .C1(\IF_ID_inst [14] ), .C2(_05322_ ), .ZN(_05563_ ) );
AND2_X1 _13338_ ( .A1(_05270_ ), .A2(_05233_ ), .ZN(_05564_ ) );
INV_X1 _13339_ ( .A(_05564_ ), .ZN(_05565_ ) );
AOI221_X4 _13340_ ( .A(_05204_ ), .B1(_05264_ ), .B2(_05266_ ), .C1(\IF_ID_inst [14] ), .C2(_05238_ ), .ZN(_05566_ ) );
AOI22_X1 _13341_ ( .A1(_05518_ ), .A2(_05233_ ), .B1(_05307_ ), .B2(_05367_ ), .ZN(_05567_ ) );
AND4_X1 _13342_ ( .A1(_05565_ ), .A2(_05363_ ), .A3(_05566_ ), .A4(_05567_ ), .ZN(_05568_ ) );
AOI21_X1 _13343_ ( .A(_05212_ ), .B1(_05563_ ), .B2(_05568_ ), .ZN(_00240_ ) );
AOI21_X1 _13344_ ( .A(_05204_ ), .B1(_05341_ ), .B2(_05265_ ), .ZN(_05569_ ) );
NAND3_X1 _13345_ ( .A1(_05237_ ), .A2(_05265_ ), .A3(_05205_ ), .ZN(_05570_ ) );
AOI21_X1 _13346_ ( .A(_05329_ ), .B1(_05569_ ), .B2(_05570_ ), .ZN(_05571_ ) );
OAI21_X1 _13347_ ( .A(_05271_ ), .B1(_05278_ ), .B2(_05275_ ), .ZN(_05572_ ) );
NAND3_X1 _13348_ ( .A1(_05366_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_05368_ ), .ZN(_05573_ ) );
NAND4_X1 _13349_ ( .A1(_05268_ ), .A2(_05352_ ), .A3(_05573_ ), .A4(_05500_ ), .ZN(_05574_ ) );
AOI22_X1 _13350_ ( .A1(_05348_ ), .A2(_05361_ ), .B1(_05364_ ), .B2(_05326_ ), .ZN(_05575_ ) );
NAND2_X1 _13351_ ( .A1(_05283_ ), .A2(_05233_ ), .ZN(_05576_ ) );
NAND2_X1 _13352_ ( .A1(_05575_ ), .A2(_05576_ ), .ZN(_05577_ ) );
NOR4_X1 _13353_ ( .A1(_05571_ ), .A2(_05572_ ), .A3(_05574_ ), .A4(_05577_ ), .ZN(_05578_ ) );
OAI21_X1 _13354_ ( .A(_05368_ ), .B1(_05364_ ), .B2(_05547_ ), .ZN(_05579_ ) );
OAI21_X1 _13355_ ( .A(_05284_ ), .B1(_05238_ ), .B2(_05206_ ), .ZN(_05580_ ) );
AND2_X1 _13356_ ( .A1(_05579_ ), .A2(_05580_ ), .ZN(_05581_ ) );
AOI22_X1 _13357_ ( .A1(_05353_ ), .A2(\IF_ID_inst [14] ), .B1(_05326_ ), .B2(_05284_ ), .ZN(_05582_ ) );
AND4_X1 _13358_ ( .A1(_05237_ ), .A2(_05336_ ), .A3(_05331_ ), .A4(_05325_ ), .ZN(_05583_ ) );
AOI21_X1 _13359_ ( .A(_05583_ ), .B1(_05322_ ), .B2(_05330_ ), .ZN(_05584_ ) );
AND4_X1 _13360_ ( .A1(_05286_ ), .A2(_05581_ ), .A3(_05582_ ), .A4(_05584_ ), .ZN(_05585_ ) );
AOI21_X1 _13361_ ( .A(_05212_ ), .B1(_05578_ ), .B2(_05585_ ), .ZN(_00241_ ) );
INV_X1 _13362_ ( .A(_05426_ ), .ZN(_05586_ ) );
INV_X1 _13363_ ( .A(fanout_net_44 ), .ZN(_05587_ ) );
BUF_X4 _13364_ ( .A(_05587_ ), .Z(_05588_ ) );
NAND4_X1 _13365_ ( .A1(_05586_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_05588_ ), .ZN(_05589_ ) );
NAND2_X1 _13366_ ( .A1(\mtvec [0] ), .A2(fanout_net_44 ), .ZN(_05590_ ) );
AOI21_X1 _13367_ ( .A(fanout_net_3 ), .B1(_05589_ ), .B2(_05590_ ), .ZN(_00245_ ) );
AND4_X2 _13368_ ( .A1(\IF_ID_inst [31] ), .A2(_05281_ ), .A3(_05302_ ), .A4(\IF_ID_inst [5] ), .ZN(_05591_ ) );
AND2_X1 _13369_ ( .A1(_05202_ ), .A2(_05591_ ), .ZN(_05592_ ) );
AND2_X1 _13370_ ( .A1(_05592_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05593_ ) );
CLKBUF_X2 _13371_ ( .A(_05303_ ), .Z(_05594_ ) );
OAI211_X1 _13372_ ( .A(_05594_ ), .B(\IF_ID_inst [31] ), .C1(_05231_ ), .C2(_05202_ ), .ZN(_05595_ ) );
NOR2_X1 _13373_ ( .A1(_05593_ ), .A2(_05595_ ), .ZN(_05596_ ) );
BUF_X4 _13374_ ( .A(_05596_ ), .Z(_05597_ ) );
BUF_X4 _13375_ ( .A(_05597_ ), .Z(_05598_ ) );
XNOR2_X1 _13376_ ( .A(_05598_ ), .B(\IF_ID_pc [29] ), .ZN(_05599_ ) );
XNOR2_X1 _13377_ ( .A(_05597_ ), .B(_01829_ ), .ZN(_05600_ ) );
AND3_X1 _13378_ ( .A1(_05594_ ), .A2(_05231_ ), .A3(\IF_ID_inst [18] ), .ZN(_05601_ ) );
BUF_X4 _13379_ ( .A(_05592_ ), .Z(_05602_ ) );
MUX2_X1 _13380_ ( .A(_05601_ ), .B(_05335_ ), .S(_05602_ ), .Z(_05603_ ) );
XNOR2_X1 _13381_ ( .A(_05603_ ), .B(_02067_ ), .ZN(_05604_ ) );
AND3_X1 _13382_ ( .A1(_05594_ ), .A2(_05231_ ), .A3(\IF_ID_inst [17] ), .ZN(_05605_ ) );
MUX2_X1 _13383_ ( .A(_05605_ ), .B(_05335_ ), .S(_05602_ ), .Z(_05606_ ) );
XNOR2_X1 _13384_ ( .A(_05606_ ), .B(_02011_ ), .ZN(_05607_ ) );
AND2_X1 _13385_ ( .A1(_05604_ ), .A2(_05607_ ), .ZN(_05608_ ) );
INV_X1 _13386_ ( .A(_05608_ ), .ZN(_05609_ ) );
AND3_X1 _13387_ ( .A1(_05594_ ), .A2(_05231_ ), .A3(\IF_ID_inst [19] ), .ZN(_05610_ ) );
MUX2_X1 _13388_ ( .A(_05610_ ), .B(_05335_ ), .S(_05602_ ), .Z(_05611_ ) );
XNOR2_X1 _13389_ ( .A(_05611_ ), .B(_02061_ ), .ZN(_05612_ ) );
XNOR2_X1 _13390_ ( .A(_05596_ ), .B(_02064_ ), .ZN(_05613_ ) );
AND2_X1 _13391_ ( .A1(_05612_ ), .A2(_05613_ ), .ZN(_05614_ ) );
INV_X1 _13392_ ( .A(_05614_ ), .ZN(_05615_ ) );
AND3_X1 _13393_ ( .A1(_05594_ ), .A2(_05230_ ), .A3(\IF_ID_inst [15] ), .ZN(_05616_ ) );
MUX2_X1 _13394_ ( .A(_05616_ ), .B(_05335_ ), .S(_05602_ ), .Z(_05617_ ) );
XOR2_X1 _13395_ ( .A(_05617_ ), .B(\IF_ID_pc [15] ), .Z(_05618_ ) );
INV_X1 _13396_ ( .A(_05602_ ), .ZN(_05619_ ) );
INV_X1 _13397_ ( .A(_05304_ ), .ZN(_05620_ ) );
OAI21_X1 _13398_ ( .A(_05619_ ), .B1(_05620_ ), .B2(_05437_ ), .ZN(_05621_ ) );
INV_X1 _13399_ ( .A(_05593_ ), .ZN(_05622_ ) );
AND3_X1 _13400_ ( .A1(_05621_ ), .A2(\IF_ID_pc [16] ), .A3(_05622_ ), .ZN(_05623_ ) );
AOI21_X1 _13401_ ( .A(\IF_ID_pc [16] ), .B1(_05621_ ), .B2(_05622_ ), .ZN(_05624_ ) );
NOR2_X1 _13402_ ( .A1(_05623_ ), .A2(_05624_ ), .ZN(_05625_ ) );
AND2_X1 _13403_ ( .A1(_05618_ ), .A2(_05625_ ), .ZN(_05626_ ) );
AND3_X1 _13404_ ( .A1(_05594_ ), .A2(_05231_ ), .A3(\IF_ID_inst [13] ), .ZN(_05627_ ) );
MUX2_X1 _13405_ ( .A(_05627_ ), .B(_05335_ ), .S(_05602_ ), .Z(_05628_ ) );
XOR2_X1 _13406_ ( .A(_05628_ ), .B(\IF_ID_pc [13] ), .Z(_05629_ ) );
OAI21_X1 _13407_ ( .A(_05619_ ), .B1(_05620_ ), .B2(_05329_ ), .ZN(_05630_ ) );
AND3_X1 _13408_ ( .A1(_05630_ ), .A2(\IF_ID_pc [14] ), .A3(_05622_ ), .ZN(_05631_ ) );
AOI21_X1 _13409_ ( .A(\IF_ID_pc [14] ), .B1(_05630_ ), .B2(_05622_ ), .ZN(_05632_ ) );
NOR2_X1 _13410_ ( .A1(_05631_ ), .A2(_05632_ ), .ZN(_05633_ ) );
AND2_X1 _13411_ ( .A1(_05629_ ), .A2(_05633_ ), .ZN(_05634_ ) );
AND2_X1 _13412_ ( .A1(_05626_ ), .A2(_05634_ ), .ZN(_05635_ ) );
INV_X1 _13413_ ( .A(_05635_ ), .ZN(_05636_ ) );
OAI21_X1 _13414_ ( .A(_05619_ ), .B1(_05620_ ), .B2(_05239_ ), .ZN(_05637_ ) );
NAND2_X1 _13415_ ( .A1(_05637_ ), .A2(_05622_ ), .ZN(_05638_ ) );
XNOR2_X1 _13416_ ( .A(_05638_ ), .B(\IF_ID_pc [12] ), .ZN(_05639_ ) );
INV_X1 _13417_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05640_ ) );
AND3_X1 _13418_ ( .A1(_05202_ ), .A2(_05591_ ), .A3(_05640_ ), .ZN(_05641_ ) );
AOI21_X1 _13419_ ( .A(_05641_ ), .B1(\IF_ID_inst [20] ), .B2(_05305_ ), .ZN(_05642_ ) );
XNOR2_X1 _13420_ ( .A(_05642_ ), .B(\IF_ID_pc [11] ), .ZN(_05643_ ) );
AND2_X1 _13421_ ( .A1(_05639_ ), .A2(_05643_ ), .ZN(_05644_ ) );
AND2_X1 _13422_ ( .A1(_05305_ ), .A2(\IF_ID_inst [29] ), .ZN(_05645_ ) );
INV_X1 _13423_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05646_ ) );
AOI21_X1 _13424_ ( .A(_05645_ ), .B1(_05646_ ), .B2(_05602_ ), .ZN(_05647_ ) );
XNOR2_X1 _13425_ ( .A(_05647_ ), .B(\IF_ID_pc [9] ), .ZN(_05648_ ) );
AND2_X1 _13426_ ( .A1(_05305_ ), .A2(\IF_ID_inst [30] ), .ZN(_05649_ ) );
INV_X1 _13427_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05650_ ) );
AOI21_X1 _13428_ ( .A(_05649_ ), .B1(_05650_ ), .B2(_05602_ ), .ZN(_05651_ ) );
XNOR2_X1 _13429_ ( .A(_05651_ ), .B(\IF_ID_pc [10] ), .ZN(_05652_ ) );
NAND3_X1 _13430_ ( .A1(_05644_ ), .A2(_05648_ ), .A3(_05652_ ), .ZN(_05653_ ) );
AND2_X1 _13431_ ( .A1(_05305_ ), .A2(\IF_ID_inst [26] ), .ZN(_05654_ ) );
INV_X1 _13432_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05655_ ) );
AOI21_X1 _13433_ ( .A(_05654_ ), .B1(_05655_ ), .B2(_05602_ ), .ZN(_05656_ ) );
OR2_X1 _13434_ ( .A1(_05656_ ), .A2(_01955_ ), .ZN(_05657_ ) );
AND2_X1 _13435_ ( .A1(_05305_ ), .A2(\IF_ID_inst [25] ), .ZN(_05658_ ) );
INV_X1 _13436_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_05659_ ) );
AND3_X1 _13437_ ( .A1(_05202_ ), .A2(_05591_ ), .A3(_05659_ ), .ZN(_05660_ ) );
NOR2_X1 _13438_ ( .A1(_05658_ ), .A2(_05660_ ), .ZN(_05661_ ) );
NAND3_X1 _13439_ ( .A1(_05594_ ), .A2(_05231_ ), .A3(\IF_ID_inst [24] ), .ZN(_05662_ ) );
INV_X1 _13440_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05663_ ) );
NAND3_X1 _13441_ ( .A1(_05202_ ), .A2(_05591_ ), .A3(_05663_ ), .ZN(_05664_ ) );
NAND2_X1 _13442_ ( .A1(_05662_ ), .A2(_05664_ ), .ZN(_05665_ ) );
NAND2_X1 _13443_ ( .A1(_05665_ ), .A2(fanout_net_13 ), .ZN(_05666_ ) );
NAND3_X1 _13444_ ( .A1(_05594_ ), .A2(_05230_ ), .A3(\IF_ID_inst [23] ), .ZN(_05667_ ) );
INV_X1 _13445_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_05668_ ) );
NAND3_X1 _13446_ ( .A1(_05202_ ), .A2(_05591_ ), .A3(_05668_ ), .ZN(_05669_ ) );
NAND2_X1 _13447_ ( .A1(_05667_ ), .A2(_05669_ ), .ZN(_05670_ ) );
INV_X1 _13448_ ( .A(_05670_ ), .ZN(_05671_ ) );
OR2_X1 _13449_ ( .A1(_05671_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05672_ ) );
NAND3_X1 _13450_ ( .A1(_05303_ ), .A2(_05230_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_05673_ ) );
NAND3_X1 _13451_ ( .A1(_05202_ ), .A2(_05591_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_05674_ ) );
AND3_X1 _13452_ ( .A1(_05673_ ), .A2(\IF_ID_pc [2] ), .A3(_05674_ ), .ZN(_05675_ ) );
AOI21_X1 _13453_ ( .A(\IF_ID_pc [2] ), .B1(_05673_ ), .B2(_05674_ ), .ZN(_05676_ ) );
NOR2_X1 _13454_ ( .A1(_05675_ ), .A2(_05676_ ), .ZN(_05677_ ) );
NAND3_X1 _13455_ ( .A1(_05594_ ), .A2(_05230_ ), .A3(\IF_ID_inst [21] ), .ZN(_05678_ ) );
INV_X1 _13456_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_05679_ ) );
NAND3_X1 _13457_ ( .A1(_05202_ ), .A2(_05591_ ), .A3(_05679_ ), .ZN(_05680_ ) );
NAND2_X1 _13458_ ( .A1(_05678_ ), .A2(_05680_ ), .ZN(_05681_ ) );
AND2_X1 _13459_ ( .A1(_05681_ ), .A2(\IF_ID_pc [1] ), .ZN(_05682_ ) );
AND2_X1 _13460_ ( .A1(_05677_ ), .A2(_05682_ ), .ZN(_05683_ ) );
NOR2_X1 _13461_ ( .A1(_05683_ ), .A2(_05675_ ), .ZN(_05684_ ) );
XNOR2_X1 _13462_ ( .A(_05670_ ), .B(fanout_net_9 ), .ZN(_05685_ ) );
OAI211_X1 _13463_ ( .A(_05666_ ), .B(_05672_ ), .C1(_05684_ ), .C2(_05685_ ), .ZN(_05686_ ) );
NAND3_X1 _13464_ ( .A1(_05662_ ), .A2(_05413_ ), .A3(_05664_ ), .ZN(_05687_ ) );
NAND2_X1 _13465_ ( .A1(_05686_ ), .A2(_05687_ ), .ZN(_05688_ ) );
INV_X1 _13466_ ( .A(\IF_ID_pc [5] ), .ZN(_05689_ ) );
XNOR2_X1 _13467_ ( .A(_05661_ ), .B(_05689_ ), .ZN(_05690_ ) );
OAI221_X1 _13468_ ( .A(_05657_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_05661_ ), .C1(_05688_ ), .C2(_05690_ ), .ZN(_05691_ ) );
INV_X1 _13469_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05692_ ) );
AND3_X1 _13470_ ( .A1(_05202_ ), .A2(_05591_ ), .A3(_05692_ ), .ZN(_05693_ ) );
AOI21_X1 _13471_ ( .A(_05693_ ), .B1(\IF_ID_inst [27] ), .B2(_05305_ ), .ZN(_05694_ ) );
XNOR2_X1 _13472_ ( .A(_05694_ ), .B(\IF_ID_pc [7] ), .ZN(_05695_ ) );
NAND2_X1 _13473_ ( .A1(_05656_ ), .A2(_01955_ ), .ZN(_05696_ ) );
AND3_X1 _13474_ ( .A1(_05691_ ), .A2(_05695_ ), .A3(_05696_ ), .ZN(_05697_ ) );
INV_X1 _13475_ ( .A(_05694_ ), .ZN(_05698_ ) );
AND2_X1 _13476_ ( .A1(_05698_ ), .A2(\IF_ID_pc [7] ), .ZN(_05699_ ) );
AND2_X1 _13477_ ( .A1(_05305_ ), .A2(\IF_ID_inst [28] ), .ZN(_05700_ ) );
INV_X1 _13478_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05701_ ) );
AOI21_X1 _13479_ ( .A(_05700_ ), .B1(_05701_ ), .B2(_05602_ ), .ZN(_05702_ ) );
INV_X1 _13480_ ( .A(_05702_ ), .ZN(_05703_ ) );
OAI22_X1 _13481_ ( .A1(_05697_ ), .A2(_05699_ ), .B1(\IF_ID_pc [8] ), .B2(_05703_ ), .ZN(_05704_ ) );
INV_X1 _13482_ ( .A(\IF_ID_pc [8] ), .ZN(_05705_ ) );
OR2_X1 _13483_ ( .A1(_05702_ ), .A2(_05705_ ), .ZN(_05706_ ) );
AOI211_X1 _13484_ ( .A(_05636_ ), .B(_05653_ ), .C1(_05704_ ), .C2(_05706_ ), .ZN(_05707_ ) );
INV_X1 _13485_ ( .A(_05707_ ), .ZN(_05708_ ) );
INV_X1 _13486_ ( .A(_05623_ ), .ZN(_05709_ ) );
AND2_X1 _13487_ ( .A1(_05617_ ), .A2(\IF_ID_pc [15] ), .ZN(_05710_ ) );
INV_X1 _13488_ ( .A(_05710_ ), .ZN(_05711_ ) );
OAI21_X1 _13489_ ( .A(_05709_ ), .B1(_05711_ ), .B2(_05624_ ), .ZN(_05712_ ) );
AND2_X1 _13490_ ( .A1(_05628_ ), .A2(\IF_ID_pc [13] ), .ZN(_05713_ ) );
INV_X1 _13491_ ( .A(_05713_ ), .ZN(_05714_ ) );
INV_X1 _13492_ ( .A(_05631_ ), .ZN(_05715_ ) );
AOI21_X1 _13493_ ( .A(_05632_ ), .B1(_05714_ ), .B2(_05715_ ), .ZN(_05716_ ) );
INV_X1 _13494_ ( .A(\IF_ID_pc [10] ), .ZN(_05717_ ) );
AND2_X1 _13495_ ( .A1(_05651_ ), .A2(_05717_ ), .ZN(_05718_ ) );
NOR2_X1 _13496_ ( .A1(_05651_ ), .A2(_05717_ ), .ZN(_05719_ ) );
INV_X1 _13497_ ( .A(\IF_ID_pc [9] ), .ZN(_05720_ ) );
NOR4_X1 _13498_ ( .A1(_05718_ ), .A2(_05719_ ), .A3(_05720_ ), .A4(_05647_ ), .ZN(_05721_ ) );
OAI21_X1 _13499_ ( .A(_05644_ ), .B1(_05721_ ), .B2(_05719_ ), .ZN(_05722_ ) );
AND3_X1 _13500_ ( .A1(_05637_ ), .A2(\IF_ID_pc [12] ), .A3(_05622_ ), .ZN(_05723_ ) );
INV_X1 _13501_ ( .A(\IF_ID_pc [11] ), .ZN(_05724_ ) );
NOR2_X1 _13502_ ( .A1(_05642_ ), .A2(_05724_ ), .ZN(_05725_ ) );
AOI21_X1 _13503_ ( .A(_05723_ ), .B1(_05639_ ), .B2(_05725_ ), .ZN(_05726_ ) );
AND2_X1 _13504_ ( .A1(_05722_ ), .A2(_05726_ ), .ZN(_05727_ ) );
INV_X1 _13505_ ( .A(_05727_ ), .ZN(_05728_ ) );
AOI221_X4 _13506_ ( .A(_05712_ ), .B1(_05626_ ), .B2(_05716_ ), .C1(_05728_ ), .C2(_05635_ ), .ZN(_05729_ ) );
AOI211_X1 _13507_ ( .A(_05609_ ), .B(_05615_ ), .C1(_05708_ ), .C2(_05729_ ), .ZN(_05730_ ) );
AND2_X1 _13508_ ( .A1(_05611_ ), .A2(\IF_ID_pc [19] ), .ZN(_05731_ ) );
AND2_X1 _13509_ ( .A1(_05613_ ), .A2(_05731_ ), .ZN(_05732_ ) );
AOI21_X1 _13510_ ( .A(_05732_ ), .B1(\IF_ID_pc [20] ), .B2(_05596_ ), .ZN(_05733_ ) );
AND2_X1 _13511_ ( .A1(_05603_ ), .A2(\IF_ID_pc [18] ), .ZN(_05734_ ) );
AND2_X1 _13512_ ( .A1(_05606_ ), .A2(\IF_ID_pc [17] ), .ZN(_05735_ ) );
AOI21_X1 _13513_ ( .A(_05734_ ), .B1(_05604_ ), .B2(_05735_ ), .ZN(_05736_ ) );
OAI21_X1 _13514_ ( .A(_05733_ ), .B1(_05736_ ), .B2(_05615_ ), .ZN(_05737_ ) );
OR2_X1 _13515_ ( .A1(_05730_ ), .A2(_05737_ ), .ZN(_05738_ ) );
XNOR2_X1 _13516_ ( .A(_05596_ ), .B(_01997_ ), .ZN(_05739_ ) );
XNOR2_X1 _13517_ ( .A(_05596_ ), .B(_01831_ ), .ZN(_05740_ ) );
AND2_X1 _13518_ ( .A1(_05739_ ), .A2(_05740_ ), .ZN(_05741_ ) );
XNOR2_X1 _13519_ ( .A(_05596_ ), .B(_02070_ ), .ZN(_05742_ ) );
INV_X1 _13520_ ( .A(_05742_ ), .ZN(_05743_ ) );
XNOR2_X1 _13521_ ( .A(_05597_ ), .B(\IF_ID_pc [22] ), .ZN(_05744_ ) );
NOR2_X1 _13522_ ( .A1(_05743_ ), .A2(_05744_ ), .ZN(_05745_ ) );
AND3_X1 _13523_ ( .A1(_05738_ ), .A2(_05741_ ), .A3(_05745_ ), .ZN(_05746_ ) );
AND2_X1 _13524_ ( .A1(_05597_ ), .A2(\IF_ID_pc [22] ), .ZN(_05747_ ) );
AND2_X1 _13525_ ( .A1(_05597_ ), .A2(\IF_ID_pc [21] ), .ZN(_05748_ ) );
OAI21_X1 _13526_ ( .A(_05741_ ), .B1(_05747_ ), .B2(_05748_ ), .ZN(_05749_ ) );
NAND2_X1 _13527_ ( .A1(_05597_ ), .A2(\IF_ID_pc [24] ), .ZN(_05750_ ) );
NAND2_X1 _13528_ ( .A1(_05597_ ), .A2(\IF_ID_pc [23] ), .ZN(_05751_ ) );
NAND3_X1 _13529_ ( .A1(_05749_ ), .A2(_05750_ ), .A3(_05751_ ), .ZN(_05752_ ) );
OAI21_X1 _13530_ ( .A(_05600_ ), .B1(_05746_ ), .B2(_05752_ ), .ZN(_05753_ ) );
INV_X1 _13531_ ( .A(_05753_ ), .ZN(_05754_ ) );
XNOR2_X1 _13532_ ( .A(_05597_ ), .B(_01993_ ), .ZN(_05755_ ) );
XNOR2_X1 _13533_ ( .A(_05597_ ), .B(_01900_ ), .ZN(_05756_ ) );
XOR2_X1 _13534_ ( .A(_05598_ ), .B(\IF_ID_pc [26] ), .Z(_05757_ ) );
NAND4_X1 _13535_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(_05756_ ), .A4(_05757_ ), .ZN(_05758_ ) );
OAI21_X1 _13536_ ( .A(_05597_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_05759_ ) );
INV_X1 _13537_ ( .A(_05759_ ), .ZN(_05760_ ) );
NAND3_X1 _13538_ ( .A1(_05755_ ), .A2(_05756_ ), .A3(_05760_ ), .ZN(_05761_ ) );
NAND2_X1 _13539_ ( .A1(_05598_ ), .A2(\IF_ID_pc [28] ), .ZN(_05762_ ) );
NAND2_X1 _13540_ ( .A1(_05598_ ), .A2(\IF_ID_pc [27] ), .ZN(_05763_ ) );
AND3_X1 _13541_ ( .A1(_05761_ ), .A2(_05762_ ), .A3(_05763_ ), .ZN(_05764_ ) );
AOI21_X1 _13542_ ( .A(_05599_ ), .B1(_05758_ ), .B2(_05764_ ), .ZN(_05765_ ) );
NOR3_X1 _13543_ ( .A1(_05593_ ), .A2(_02074_ ), .A3(_05595_ ), .ZN(_05766_ ) );
NOR2_X1 _13544_ ( .A1(_05765_ ), .A2(_05766_ ), .ZN(_05767_ ) );
XNOR2_X1 _13545_ ( .A(_05598_ ), .B(\IF_ID_pc [30] ), .ZN(_05768_ ) );
OR2_X1 _13546_ ( .A1(_05767_ ), .A2(_05768_ ), .ZN(_05769_ ) );
AOI21_X1 _13547_ ( .A(_05427_ ), .B1(_05767_ ), .B2(_05768_ ), .ZN(_05770_ ) );
AOI221_X4 _13548_ ( .A(fanout_net_44 ), .B1(\myexu.pc_jump [30] ), .B2(_05427_ ), .C1(_05769_ ), .C2(_05770_ ), .ZN(_05771_ ) );
BUF_X4 _13549_ ( .A(_05588_ ), .Z(_05772_ ) );
NOR2_X1 _13550_ ( .A1(_05772_ ), .A2(\mtvec [30] ), .ZN(_05773_ ) );
NOR3_X1 _13551_ ( .A1(_05771_ ), .A2(fanout_net_3 ), .A3(_05773_ ), .ZN(_00246_ ) );
INV_X1 _13552_ ( .A(_05427_ ), .ZN(_05774_ ) );
BUF_X4 _13553_ ( .A(_05774_ ), .Z(_05775_ ) );
BUF_X4 _13554_ ( .A(_05775_ ), .Z(_05776_ ) );
AND2_X1 _13555_ ( .A1(_05738_ ), .A2(_05742_ ), .ZN(_05777_ ) );
NOR3_X1 _13556_ ( .A1(_05730_ ), .A2(_05742_ ), .A3(_05737_ ), .ZN(_05778_ ) );
OAI21_X1 _13557_ ( .A(_05776_ ), .B1(_05777_ ), .B2(_05778_ ), .ZN(_05779_ ) );
BUF_X4 _13558_ ( .A(_05587_ ), .Z(_05780_ ) );
BUF_X4 _13559_ ( .A(_05775_ ), .Z(_05781_ ) );
OAI211_X1 _13560_ ( .A(_05779_ ), .B(_05780_ ), .C1(\myexu.pc_jump [21] ), .C2(_05781_ ), .ZN(_05782_ ) );
NAND2_X1 _13561_ ( .A1(\mtvec [21] ), .A2(fanout_net_44 ), .ZN(_05783_ ) );
AOI21_X1 _13562_ ( .A(fanout_net_3 ), .B1(_05782_ ), .B2(_05783_ ), .ZN(_00247_ ) );
AOI21_X1 _13563_ ( .A(_05609_ ), .B1(_05708_ ), .B2(_05729_ ), .ZN(_05784_ ) );
INV_X1 _13564_ ( .A(_05736_ ), .ZN(_05785_ ) );
NOR2_X1 _13565_ ( .A1(_05784_ ), .A2(_05785_ ), .ZN(_05786_ ) );
INV_X1 _13566_ ( .A(_05786_ ), .ZN(_05787_ ) );
AND2_X1 _13567_ ( .A1(_05787_ ), .A2(_05612_ ), .ZN(_05788_ ) );
OR3_X1 _13568_ ( .A1(_05788_ ), .A2(_05731_ ), .A3(_05613_ ), .ZN(_05789_ ) );
OAI21_X1 _13569_ ( .A(_05613_ ), .B1(_05788_ ), .B2(_05731_ ), .ZN(_05790_ ) );
AND3_X1 _13570_ ( .A1(_05789_ ), .A2(_05774_ ), .A3(_05790_ ), .ZN(_05791_ ) );
BUF_X4 _13571_ ( .A(_05427_ ), .Z(_05792_ ) );
BUF_X4 _13572_ ( .A(_05792_ ), .Z(_05793_ ) );
AOI211_X1 _13573_ ( .A(fanout_net_44 ), .B(_05791_ ), .C1(\myexu.pc_jump [20] ), .C2(_05793_ ), .ZN(_05794_ ) );
NOR2_X1 _13574_ ( .A1(_05772_ ), .A2(\mtvec [20] ), .ZN(_05795_ ) );
NOR3_X1 _13575_ ( .A1(_05794_ ), .A2(fanout_net_3 ), .A3(_05795_ ), .ZN(_00248_ ) );
NOR3_X1 _13576_ ( .A1(_05784_ ), .A2(_05785_ ), .A3(_05612_ ), .ZN(_05796_ ) );
OAI21_X1 _13577_ ( .A(_05775_ ), .B1(_05788_ ), .B2(_05796_ ), .ZN(_05797_ ) );
OAI211_X1 _13578_ ( .A(_05797_ ), .B(_05780_ ), .C1(\myexu.pc_jump [19] ), .C2(_05781_ ), .ZN(_05798_ ) );
NAND2_X1 _13579_ ( .A1(\mtvec [19] ), .A2(fanout_net_44 ), .ZN(_05799_ ) );
AOI21_X1 _13580_ ( .A(fanout_net_3 ), .B1(_05798_ ), .B2(_05799_ ), .ZN(_00249_ ) );
INV_X1 _13581_ ( .A(_05607_ ), .ZN(_05800_ ) );
AOI21_X1 _13582_ ( .A(_05800_ ), .B1(_05708_ ), .B2(_05729_ ), .ZN(_05801_ ) );
OR3_X1 _13583_ ( .A1(_05801_ ), .A2(_05604_ ), .A3(_05735_ ), .ZN(_05802_ ) );
OAI21_X1 _13584_ ( .A(_05604_ ), .B1(_05801_ ), .B2(_05735_ ), .ZN(_05803_ ) );
AND3_X1 _13585_ ( .A1(_05802_ ), .A2(_05774_ ), .A3(_05803_ ), .ZN(_05804_ ) );
AOI211_X1 _13586_ ( .A(fanout_net_44 ), .B(_05804_ ), .C1(\myexu.pc_jump [18] ), .C2(_05793_ ), .ZN(_05805_ ) );
NOR2_X1 _13587_ ( .A1(_05772_ ), .A2(\mtvec [18] ), .ZN(_05806_ ) );
NOR3_X1 _13588_ ( .A1(_05805_ ), .A2(fanout_net_3 ), .A3(_05806_ ), .ZN(_00250_ ) );
AND3_X1 _13589_ ( .A1(_05708_ ), .A2(_05729_ ), .A3(_05800_ ), .ZN(_05807_ ) );
OAI21_X1 _13590_ ( .A(_05775_ ), .B1(_05807_ ), .B2(_05801_ ), .ZN(_05808_ ) );
OAI211_X1 _13591_ ( .A(_05808_ ), .B(_05780_ ), .C1(\myexu.pc_jump [17] ), .C2(_05781_ ), .ZN(_05809_ ) );
NAND2_X1 _13592_ ( .A1(\mtvec [17] ), .A2(fanout_net_44 ), .ZN(_05810_ ) );
AOI21_X1 _13593_ ( .A(fanout_net_3 ), .B1(_05809_ ), .B2(_05810_ ), .ZN(_00251_ ) );
AOI21_X1 _13594_ ( .A(_05653_ ), .B1(_05704_ ), .B2(_05706_ ), .ZN(_05811_ ) );
OR2_X1 _13595_ ( .A1(_05811_ ), .A2(_05728_ ), .ZN(_05812_ ) );
AND2_X1 _13596_ ( .A1(_05812_ ), .A2(_05634_ ), .ZN(_05813_ ) );
OR2_X1 _13597_ ( .A1(_05813_ ), .A2(_05716_ ), .ZN(_05814_ ) );
AOI211_X1 _13598_ ( .A(_05625_ ), .B(_05710_ ), .C1(_05814_ ), .C2(_05618_ ), .ZN(_05815_ ) );
OAI21_X1 _13599_ ( .A(_05618_ ), .B1(_05813_ ), .B2(_05716_ ), .ZN(_05816_ ) );
AOI211_X1 _13600_ ( .A(_05623_ ), .B(_05624_ ), .C1(_05816_ ), .C2(_05711_ ), .ZN(_05817_ ) );
NOR3_X1 _13601_ ( .A1(_05815_ ), .A2(_05817_ ), .A3(_05792_ ), .ZN(_05818_ ) );
AOI211_X1 _13602_ ( .A(fanout_net_44 ), .B(_05818_ ), .C1(\myexu.pc_jump [16] ), .C2(_05793_ ), .ZN(_05819_ ) );
NOR2_X1 _13603_ ( .A1(_05772_ ), .A2(\mtvec [16] ), .ZN(_05820_ ) );
NOR3_X1 _13604_ ( .A1(_05819_ ), .A2(fanout_net_3 ), .A3(_05820_ ), .ZN(_00252_ ) );
XNOR2_X1 _13605_ ( .A(_05814_ ), .B(_05618_ ), .ZN(_05821_ ) );
NOR2_X1 _13606_ ( .A1(_05821_ ), .A2(_05792_ ), .ZN(_05822_ ) );
AOI211_X1 _13607_ ( .A(fanout_net_44 ), .B(_05822_ ), .C1(\myexu.pc_jump [15] ), .C2(_05793_ ), .ZN(_05823_ ) );
NOR2_X1 _13608_ ( .A1(_05772_ ), .A2(\mtvec [15] ), .ZN(_05824_ ) );
NOR3_X1 _13609_ ( .A1(_05823_ ), .A2(fanout_net_3 ), .A3(_05824_ ), .ZN(_00253_ ) );
OAI21_X1 _13610_ ( .A(_05629_ ), .B1(_05811_ ), .B2(_05728_ ), .ZN(_05825_ ) );
AND2_X1 _13611_ ( .A1(_05825_ ), .A2(_05714_ ), .ZN(_05826_ ) );
XNOR2_X1 _13612_ ( .A(_05826_ ), .B(_05633_ ), .ZN(_05827_ ) );
MUX2_X1 _13613_ ( .A(\myexu.pc_jump [14] ), .B(_05827_ ), .S(_05774_ ), .Z(_05828_ ) );
MUX2_X1 _13614_ ( .A(\mtvec [14] ), .B(_05828_ ), .S(_05587_ ), .Z(_05829_ ) );
AND2_X1 _13615_ ( .A1(_05829_ ), .A2(_01585_ ), .ZN(_00254_ ) );
XNOR2_X1 _13616_ ( .A(_05812_ ), .B(_05629_ ), .ZN(_05830_ ) );
NAND2_X1 _13617_ ( .A1(_05830_ ), .A2(_05776_ ), .ZN(_05831_ ) );
OAI211_X1 _13618_ ( .A(_05831_ ), .B(_05780_ ), .C1(\myexu.pc_jump [13] ), .C2(_05781_ ), .ZN(_05832_ ) );
NAND2_X1 _13619_ ( .A1(\mtvec [13] ), .A2(fanout_net_44 ), .ZN(_05833_ ) );
AOI21_X1 _13620_ ( .A(fanout_net_3 ), .B1(_05832_ ), .B2(_05833_ ), .ZN(_00255_ ) );
NAND2_X1 _13621_ ( .A1(_05704_ ), .A2(_05706_ ), .ZN(_05834_ ) );
NAND3_X1 _13622_ ( .A1(_05834_ ), .A2(_05648_ ), .A3(_05652_ ), .ZN(_05835_ ) );
INV_X1 _13623_ ( .A(_05718_ ), .ZN(_05836_ ) );
NOR2_X1 _13624_ ( .A1(_05647_ ), .A2(_05720_ ), .ZN(_05837_ ) );
AOI21_X1 _13625_ ( .A(_05719_ ), .B1(_05836_ ), .B2(_05837_ ), .ZN(_05838_ ) );
AND2_X1 _13626_ ( .A1(_05835_ ), .A2(_05838_ ), .ZN(_05839_ ) );
INV_X1 _13627_ ( .A(_05643_ ), .ZN(_05840_ ) );
NOR2_X1 _13628_ ( .A1(_05839_ ), .A2(_05840_ ), .ZN(_05841_ ) );
OR3_X1 _13629_ ( .A1(_05841_ ), .A2(_05725_ ), .A3(_05639_ ), .ZN(_05842_ ) );
OAI21_X1 _13630_ ( .A(_05639_ ), .B1(_05841_ ), .B2(_05725_ ), .ZN(_05843_ ) );
AND3_X1 _13631_ ( .A1(_05842_ ), .A2(_05774_ ), .A3(_05843_ ), .ZN(_05844_ ) );
AOI211_X1 _13632_ ( .A(fanout_net_44 ), .B(_05844_ ), .C1(\myexu.pc_jump [12] ), .C2(_05793_ ), .ZN(_05845_ ) );
NOR2_X1 _13633_ ( .A1(_05772_ ), .A2(\mtvec [12] ), .ZN(_05846_ ) );
NOR3_X1 _13634_ ( .A1(_05845_ ), .A2(fanout_net_3 ), .A3(_05846_ ), .ZN(_00256_ ) );
AND3_X1 _13635_ ( .A1(_05758_ ), .A2(_05764_ ), .A3(_05599_ ), .ZN(_05847_ ) );
OAI21_X1 _13636_ ( .A(_05775_ ), .B1(_05847_ ), .B2(_05765_ ), .ZN(_05848_ ) );
OAI211_X1 _13637_ ( .A(_05848_ ), .B(_05780_ ), .C1(\myexu.pc_jump [29] ), .C2(_05781_ ), .ZN(_05849_ ) );
NAND2_X1 _13638_ ( .A1(\mtvec [29] ), .A2(fanout_net_44 ), .ZN(_05850_ ) );
AOI21_X1 _13639_ ( .A(fanout_net_3 ), .B1(_05849_ ), .B2(_05850_ ), .ZN(_00257_ ) );
AND3_X1 _13640_ ( .A1(_05835_ ), .A2(_05840_ ), .A3(_05838_ ), .ZN(_05851_ ) );
OAI21_X1 _13641_ ( .A(_05775_ ), .B1(_05841_ ), .B2(_05851_ ), .ZN(_05852_ ) );
OAI211_X1 _13642_ ( .A(_05852_ ), .B(_05780_ ), .C1(\myexu.pc_jump [11] ), .C2(_05781_ ), .ZN(_05853_ ) );
NAND2_X1 _13643_ ( .A1(\mtvec [11] ), .A2(fanout_net_44 ), .ZN(_05854_ ) );
AOI21_X1 _13644_ ( .A(fanout_net_3 ), .B1(_05853_ ), .B2(_05854_ ), .ZN(_00258_ ) );
INV_X1 _13645_ ( .A(_05648_ ), .ZN(_05855_ ) );
AOI21_X1 _13646_ ( .A(_05855_ ), .B1(_05704_ ), .B2(_05706_ ), .ZN(_05856_ ) );
NOR2_X1 _13647_ ( .A1(_05856_ ), .A2(_05837_ ), .ZN(_05857_ ) );
INV_X1 _13648_ ( .A(_05857_ ), .ZN(_05858_ ) );
OAI21_X1 _13649_ ( .A(_05774_ ), .B1(_05858_ ), .B2(_05652_ ), .ZN(_05859_ ) );
AOI21_X1 _13650_ ( .A(_05859_ ), .B1(_05858_ ), .B2(_05652_ ), .ZN(_05860_ ) );
AOI211_X1 _13651_ ( .A(fanout_net_44 ), .B(_05860_ ), .C1(\myexu.pc_jump [10] ), .C2(_05793_ ), .ZN(_05861_ ) );
NOR2_X1 _13652_ ( .A1(_05772_ ), .A2(\mtvec [10] ), .ZN(_05862_ ) );
NOR3_X1 _13653_ ( .A1(_05861_ ), .A2(fanout_net_4 ), .A3(_05862_ ), .ZN(_00259_ ) );
OR3_X1 _13654_ ( .A1(_05426_ ), .A2(_02117_ ), .A3(\myexu.pc_jump [9] ), .ZN(_05863_ ) );
XNOR2_X1 _13655_ ( .A(_05834_ ), .B(_05855_ ), .ZN(_05864_ ) );
OAI211_X1 _13656_ ( .A(_05780_ ), .B(_05863_ ), .C1(_05864_ ), .C2(_05793_ ), .ZN(_05865_ ) );
NAND2_X1 _13657_ ( .A1(\mtvec [9] ), .A2(fanout_net_44 ), .ZN(_05866_ ) );
AOI21_X1 _13658_ ( .A(fanout_net_4 ), .B1(_05865_ ), .B2(_05866_ ), .ZN(_00260_ ) );
NOR2_X1 _13659_ ( .A1(_05697_ ), .A2(_05699_ ), .ZN(_05867_ ) );
XNOR2_X1 _13660_ ( .A(_05702_ ), .B(_05705_ ), .ZN(_05868_ ) );
OR2_X1 _13661_ ( .A1(_05867_ ), .A2(_05868_ ), .ZN(_05869_ ) );
AOI21_X1 _13662_ ( .A(_05427_ ), .B1(_05867_ ), .B2(_05868_ ), .ZN(_05870_ ) );
AOI221_X4 _13663_ ( .A(fanout_net_44 ), .B1(\myexu.pc_jump [8] ), .B2(_05427_ ), .C1(_05869_ ), .C2(_05870_ ), .ZN(_05871_ ) );
NOR2_X1 _13664_ ( .A1(_05772_ ), .A2(\mtvec [8] ), .ZN(_05872_ ) );
NOR3_X1 _13665_ ( .A1(_05871_ ), .A2(fanout_net_4 ), .A3(_05872_ ), .ZN(_00261_ ) );
AOI21_X1 _13666_ ( .A(_05695_ ), .B1(_05691_ ), .B2(_05696_ ), .ZN(_05873_ ) );
OAI21_X1 _13667_ ( .A(_05775_ ), .B1(_05697_ ), .B2(_05873_ ), .ZN(_05874_ ) );
OAI211_X1 _13668_ ( .A(_05874_ ), .B(_05588_ ), .C1(\myexu.pc_jump [7] ), .C2(_05781_ ), .ZN(_05875_ ) );
NAND2_X1 _13669_ ( .A1(\mtvec [7] ), .A2(fanout_net_44 ), .ZN(_05876_ ) );
AOI21_X1 _13670_ ( .A(fanout_net_4 ), .B1(_05875_ ), .B2(_05876_ ), .ZN(_00262_ ) );
NOR2_X1 _13671_ ( .A1(_05688_ ), .A2(_05690_ ), .ZN(_05877_ ) );
NOR2_X1 _13672_ ( .A1(_05661_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05878_ ) );
XNOR2_X1 _13673_ ( .A(_05656_ ), .B(_01955_ ), .ZN(_05879_ ) );
OR3_X1 _13674_ ( .A1(_05877_ ), .A2(_05878_ ), .A3(_05879_ ), .ZN(_05880_ ) );
OAI21_X1 _13675_ ( .A(_05879_ ), .B1(_05877_ ), .B2(_05878_ ), .ZN(_05881_ ) );
NAND3_X1 _13676_ ( .A1(_05880_ ), .A2(_05776_ ), .A3(_05881_ ), .ZN(_05882_ ) );
OAI211_X1 _13677_ ( .A(_05882_ ), .B(_05588_ ), .C1(\myexu.pc_jump [6] ), .C2(_05781_ ), .ZN(_05883_ ) );
NAND2_X1 _13678_ ( .A1(\mtvec [6] ), .A2(fanout_net_44 ), .ZN(_05884_ ) );
AOI21_X1 _13679_ ( .A(fanout_net_4 ), .B1(_05883_ ), .B2(_05884_ ), .ZN(_00263_ ) );
AND2_X1 _13680_ ( .A1(_05688_ ), .A2(_05690_ ), .ZN(_05885_ ) );
NOR3_X1 _13681_ ( .A1(_05885_ ), .A2(_05877_ ), .A3(_05792_ ), .ZN(_05886_ ) );
AOI211_X1 _13682_ ( .A(fanout_net_44 ), .B(_05886_ ), .C1(\myexu.pc_jump [5] ), .C2(_05792_ ), .ZN(_05887_ ) );
NOR2_X1 _13683_ ( .A1(_05772_ ), .A2(\mtvec [5] ), .ZN(_05888_ ) );
NOR3_X1 _13684_ ( .A1(_05887_ ), .A2(fanout_net_4 ), .A3(_05888_ ), .ZN(_00264_ ) );
OR2_X1 _13685_ ( .A1(_05684_ ), .A2(_05685_ ), .ZN(_05889_ ) );
AND2_X1 _13686_ ( .A1(_05666_ ), .A2(_05687_ ), .ZN(_05890_ ) );
AND3_X1 _13687_ ( .A1(_05889_ ), .A2(_05672_ ), .A3(_05890_ ), .ZN(_05891_ ) );
AOI21_X1 _13688_ ( .A(_05890_ ), .B1(_05889_ ), .B2(_05672_ ), .ZN(_05892_ ) );
OR3_X1 _13689_ ( .A1(_05891_ ), .A2(_05892_ ), .A3(_05427_ ), .ZN(_05893_ ) );
OAI211_X1 _13690_ ( .A(_05893_ ), .B(_05587_ ), .C1(\myexu.pc_jump [4] ), .C2(_05774_ ), .ZN(_05894_ ) );
NAND2_X1 _13691_ ( .A1(\mtvec [4] ), .A2(fanout_net_44 ), .ZN(_05895_ ) );
AOI21_X1 _13692_ ( .A(fanout_net_4 ), .B1(_05894_ ), .B2(_05895_ ), .ZN(_00265_ ) );
AND2_X1 _13693_ ( .A1(_05889_ ), .A2(_05774_ ), .ZN(_05896_ ) );
NAND2_X1 _13694_ ( .A1(_05684_ ), .A2(_05685_ ), .ZN(_05897_ ) );
AOI22_X1 _13695_ ( .A1(_05896_ ), .A2(_05897_ ), .B1(\myexu.pc_jump [3] ), .B2(_05427_ ), .ZN(_05898_ ) );
NOR2_X1 _13696_ ( .A1(_05898_ ), .A2(fanout_net_44 ), .ZN(_05899_ ) );
AOI21_X1 _13697_ ( .A(_05899_ ), .B1(\mtvec [3] ), .B2(fanout_net_44 ), .ZN(_05900_ ) );
NOR2_X1 _13698_ ( .A1(_05900_ ), .A2(fanout_net_4 ), .ZN(_00266_ ) );
AND2_X1 _13699_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
AND3_X1 _13700_ ( .A1(_05894_ ), .A2(_05895_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_05901_ ) );
BUF_X4 _13701_ ( .A(_05413_ ), .Z(_05902_ ) );
BUF_X4 _13702_ ( .A(_05902_ ), .Z(_05903_ ) );
BUF_X4 _13703_ ( .A(_05903_ ), .Z(_05904_ ) );
BUF_X2 _13704_ ( .A(_05904_ ), .Z(_05905_ ) );
INV_X1 _13705_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_05906_ ) );
AOI211_X1 _13706_ ( .A(fanout_net_4 ), .B(_05901_ ), .C1(_05905_ ), .C2(_05906_ ), .ZN(_00267_ ) );
NAND3_X1 _13707_ ( .A1(_05425_ ), .A2(_05404_ ), .A3(_05410_ ), .ZN(_05907_ ) );
INV_X1 _13708_ ( .A(_05399_ ), .ZN(_05908_ ) );
OAI211_X1 _13709_ ( .A(check_quest ), .B(_05417_ ), .C1(_05907_ ), .C2(_05908_ ), .ZN(_05909_ ) );
XOR2_X1 _13710_ ( .A(_05677_ ), .B(_05682_ ), .Z(_05910_ ) );
OAI211_X1 _13711_ ( .A(_05780_ ), .B(_05909_ ), .C1(_05910_ ), .C2(_05793_ ), .ZN(_05911_ ) );
NAND2_X1 _13712_ ( .A1(\mtvec [2] ), .A2(fanout_net_44 ), .ZN(_05912_ ) );
AOI21_X1 _13713_ ( .A(fanout_net_4 ), .B1(_05911_ ), .B2(_05912_ ), .ZN(_00268_ ) );
AOI211_X1 _13714_ ( .A(_05906_ ), .B(_05899_ ), .C1(\mtvec [3] ), .C2(fanout_net_44 ), .ZN(_05913_ ) );
INV_X2 _13715_ ( .A(fanout_net_9 ), .ZN(_05914_ ) );
BUF_X4 _13716_ ( .A(_05914_ ), .Z(_05915_ ) );
BUF_X2 _13717_ ( .A(_05915_ ), .Z(_05916_ ) );
AOI211_X1 _13718_ ( .A(fanout_net_4 ), .B(_05913_ ), .C1(_05916_ ), .C2(_05906_ ), .ZN(_00269_ ) );
AND2_X1 _13719_ ( .A1(_05754_ ), .A2(_05757_ ), .ZN(_05917_ ) );
OAI21_X1 _13720_ ( .A(_05756_ ), .B1(_05917_ ), .B2(_05760_ ), .ZN(_05918_ ) );
NAND2_X1 _13721_ ( .A1(_05918_ ), .A2(_05763_ ), .ZN(_05919_ ) );
XNOR2_X1 _13722_ ( .A(_05919_ ), .B(_05755_ ), .ZN(_05920_ ) );
NOR2_X1 _13723_ ( .A1(_05920_ ), .A2(_05792_ ), .ZN(_05921_ ) );
AOI211_X1 _13724_ ( .A(fanout_net_44 ), .B(_05921_ ), .C1(\myexu.pc_jump [28] ), .C2(_05792_ ), .ZN(_05922_ ) );
NOR2_X1 _13725_ ( .A1(_05780_ ), .A2(\mtvec [28] ), .ZN(_05923_ ) );
NOR3_X1 _13726_ ( .A1(_05922_ ), .A2(fanout_net_4 ), .A3(_05923_ ), .ZN(_00270_ ) );
NOR2_X1 _13727_ ( .A1(_05588_ ), .A2(\mtvec [1] ), .ZN(_05924_ ) );
XNOR2_X1 _13728_ ( .A(_05681_ ), .B(\IF_ID_pc [1] ), .ZN(_05925_ ) );
MUX2_X1 _13729_ ( .A(_05925_ ), .B(_05411_ ), .S(_05792_ ), .Z(_05926_ ) );
AOI211_X1 _13730_ ( .A(fanout_net_4 ), .B(_05924_ ), .C1(_05926_ ), .C2(_05772_ ), .ZN(_00271_ ) );
NOR2_X1 _13731_ ( .A1(_05917_ ), .A2(_05760_ ), .ZN(_05927_ ) );
XOR2_X1 _13732_ ( .A(_05927_ ), .B(_05756_ ), .Z(_05928_ ) );
NAND2_X1 _13733_ ( .A1(_05928_ ), .A2(_05776_ ), .ZN(_05929_ ) );
OAI211_X1 _13734_ ( .A(_05929_ ), .B(_05588_ ), .C1(\myexu.pc_jump [27] ), .C2(_05781_ ), .ZN(_05930_ ) );
NAND2_X1 _13735_ ( .A1(\mtvec [27] ), .A2(fanout_net_44 ), .ZN(_05931_ ) );
AOI21_X1 _13736_ ( .A(fanout_net_4 ), .B1(_05930_ ), .B2(_05931_ ), .ZN(_00272_ ) );
NAND2_X1 _13737_ ( .A1(_05598_ ), .A2(\IF_ID_pc [25] ), .ZN(_05932_ ) );
AND2_X1 _13738_ ( .A1(_05753_ ), .A2(_05932_ ), .ZN(_05933_ ) );
XNOR2_X1 _13739_ ( .A(_05933_ ), .B(_05757_ ), .ZN(_05934_ ) );
AND2_X1 _13740_ ( .A1(_05934_ ), .A2(_05775_ ), .ZN(_05935_ ) );
AOI211_X1 _13741_ ( .A(fanout_net_44 ), .B(_05935_ ), .C1(\myexu.pc_jump [26] ), .C2(_05792_ ), .ZN(_05936_ ) );
NOR2_X1 _13742_ ( .A1(_05780_ ), .A2(\mtvec [26] ), .ZN(_05937_ ) );
NOR3_X1 _13743_ ( .A1(_05936_ ), .A2(fanout_net_4 ), .A3(_05937_ ), .ZN(_00273_ ) );
NOR3_X1 _13744_ ( .A1(_05746_ ), .A2(_05752_ ), .A3(_05600_ ), .ZN(_05938_ ) );
OAI21_X1 _13745_ ( .A(_05775_ ), .B1(_05754_ ), .B2(_05938_ ), .ZN(_05939_ ) );
OAI211_X1 _13746_ ( .A(_05939_ ), .B(_05588_ ), .C1(\myexu.pc_jump [25] ), .C2(_05776_ ), .ZN(_05940_ ) );
NAND2_X1 _13747_ ( .A1(\mtvec [25] ), .A2(fanout_net_44 ), .ZN(_05941_ ) );
AOI21_X1 _13748_ ( .A(fanout_net_4 ), .B1(_05940_ ), .B2(_05941_ ), .ZN(_00274_ ) );
OAI21_X1 _13749_ ( .A(_05745_ ), .B1(_05730_ ), .B2(_05737_ ), .ZN(_05942_ ) );
OAI21_X1 _13750_ ( .A(_05598_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_05943_ ) );
NAND2_X1 _13751_ ( .A1(_05942_ ), .A2(_05943_ ), .ZN(_05944_ ) );
NAND2_X1 _13752_ ( .A1(_05944_ ), .A2(_05740_ ), .ZN(_05945_ ) );
AND3_X1 _13753_ ( .A1(_05945_ ), .A2(_05739_ ), .A3(_05751_ ), .ZN(_05946_ ) );
AOI21_X1 _13754_ ( .A(_05739_ ), .B1(_05945_ ), .B2(_05751_ ), .ZN(_05947_ ) );
OR3_X1 _13755_ ( .A1(_05946_ ), .A2(_05947_ ), .A3(_05427_ ), .ZN(_05948_ ) );
OAI211_X1 _13756_ ( .A(_05948_ ), .B(_05588_ ), .C1(\myexu.pc_jump [24] ), .C2(_05776_ ), .ZN(_05949_ ) );
NAND2_X1 _13757_ ( .A1(\mtvec [24] ), .A2(\myifu.to_reset ), .ZN(_05950_ ) );
AOI21_X1 _13758_ ( .A(fanout_net_4 ), .B1(_05949_ ), .B2(_05950_ ), .ZN(_00275_ ) );
XNOR2_X1 _13759_ ( .A(_05944_ ), .B(_05740_ ), .ZN(_05951_ ) );
NAND2_X1 _13760_ ( .A1(_05951_ ), .A2(_05776_ ), .ZN(_05952_ ) );
OAI211_X1 _13761_ ( .A(_05952_ ), .B(_05588_ ), .C1(\myexu.pc_jump [23] ), .C2(_05776_ ), .ZN(_05953_ ) );
NAND2_X1 _13762_ ( .A1(\mtvec [23] ), .A2(\myifu.to_reset ), .ZN(_05954_ ) );
AOI21_X1 _13763_ ( .A(fanout_net_4 ), .B1(_05953_ ), .B2(_05954_ ), .ZN(_00276_ ) );
OR3_X1 _13764_ ( .A1(_05777_ ), .A2(_05748_ ), .A3(_05744_ ), .ZN(_05955_ ) );
OAI21_X1 _13765_ ( .A(_05744_ ), .B1(_05777_ ), .B2(_05748_ ), .ZN(_05956_ ) );
NAND3_X1 _13766_ ( .A1(_05955_ ), .A2(_05776_ ), .A3(_05956_ ), .ZN(_05957_ ) );
OAI211_X1 _13767_ ( .A(_05957_ ), .B(_05588_ ), .C1(\myexu.pc_jump [22] ), .C2(_05776_ ), .ZN(_05958_ ) );
NAND2_X1 _13768_ ( .A1(\mtvec [22] ), .A2(\myifu.to_reset ), .ZN(_05959_ ) );
AOI21_X1 _13769_ ( .A(fanout_net_4 ), .B1(_05958_ ), .B2(_05959_ ), .ZN(_00277_ ) );
OAI21_X1 _13770_ ( .A(_05587_ ), .B1(_05775_ ), .B2(\myexu.pc_jump [31] ), .ZN(_05960_ ) );
OAI22_X1 _13771_ ( .A1(_05765_ ), .A2(_05766_ ), .B1(\IF_ID_pc [30] ), .B2(_05598_ ), .ZN(_05961_ ) );
NAND2_X1 _13772_ ( .A1(_05598_ ), .A2(\IF_ID_pc [30] ), .ZN(_05962_ ) );
AND2_X1 _13773_ ( .A1(_05961_ ), .A2(_05962_ ), .ZN(_05963_ ) );
XOR2_X1 _13774_ ( .A(_05598_ ), .B(\IF_ID_pc [31] ), .Z(_05964_ ) );
OR2_X1 _13775_ ( .A1(_05963_ ), .A2(_05964_ ), .ZN(_05965_ ) );
AOI21_X1 _13776_ ( .A(_05792_ ), .B1(_05963_ ), .B2(_05964_ ), .ZN(_05966_ ) );
AOI21_X1 _13777_ ( .A(_05960_ ), .B1(_05965_ ), .B2(_05966_ ), .ZN(_05967_ ) );
AND2_X1 _13778_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_05968_ ) );
OR3_X1 _13779_ ( .A1(_05967_ ), .A2(fanout_net_4 ), .A3(_05968_ ), .ZN(_00278_ ) );
OR4_X4 _13780_ ( .A1(\io_master_araddr [23] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [21] ), .A4(\io_master_araddr [22] ), .ZN(_05969_ ) );
OR2_X1 _13781_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [18] ), .ZN(_05970_ ) );
OR4_X4 _13782_ ( .A1(\io_master_araddr [16] ), .A2(_05969_ ), .A3(\io_master_araddr [17] ), .A4(_05970_ ), .ZN(_05971_ ) );
BUF_X2 _13783_ ( .A(_05971_ ), .Z(_05972_ ) );
OR4_X1 _13784_ ( .A1(\io_master_araddr [31] ), .A2(\io_master_araddr [29] ), .A3(\io_master_araddr [30] ), .A4(\io_master_araddr [28] ), .ZN(_05973_ ) );
INV_X1 _13785_ ( .A(_02004_ ), .ZN(\io_master_araddr [26] ) );
NAND2_X1 _13786_ ( .A1(_01990_ ), .A2(\io_master_araddr [25] ), .ZN(_05974_ ) );
OR4_X4 _13787_ ( .A1(\io_master_araddr [24] ), .A2(_05973_ ), .A3(\io_master_araddr [26] ), .A4(_05974_ ), .ZN(_05975_ ) );
BUF_X2 _13788_ ( .A(_05975_ ), .Z(_05976_ ) );
OR3_X4 _13789_ ( .A1(_05972_ ), .A2(_05976_ ), .A3(\myclint.state_r_$_NOT__A_Y ), .ZN(_05977_ ) );
OAI21_X1 _13790_ ( .A(io_master_rvalid ), .B1(_05972_ ), .B2(_05976_ ), .ZN(_05978_ ) );
NAND2_X1 _13791_ ( .A1(_05977_ ), .A2(_05978_ ), .ZN(_05979_ ) );
NOR2_X4 _13792_ ( .A1(_05975_ ), .A2(_05971_ ), .ZN(_05980_ ) );
BUF_X4 _13793_ ( .A(_05980_ ), .Z(_05981_ ) );
BUF_X4 _13794_ ( .A(_05981_ ), .Z(_05982_ ) );
NOR2_X1 _13795_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_05983_ ) );
OR2_X1 _13796_ ( .A1(_05982_ ), .A2(_05983_ ), .ZN(_05984_ ) );
AND3_X2 _13797_ ( .A1(_05979_ ), .A2(_02053_ ), .A3(_05984_ ), .ZN(_05985_ ) );
BUF_X4 _13798_ ( .A(_05981_ ), .Z(_05986_ ) );
NOR2_X1 _13799_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_05987_ ) );
OAI21_X1 _13800_ ( .A(_02053_ ), .B1(_05986_ ), .B2(_05987_ ), .ZN(_05988_ ) );
INV_X1 _13801_ ( .A(\io_master_rid [1] ), .ZN(_05989_ ) );
AND2_X1 _13802_ ( .A1(_05989_ ), .A2(\io_master_rid [0] ), .ZN(_05990_ ) );
NOR2_X1 _13803_ ( .A1(_05986_ ), .A2(_05990_ ), .ZN(_05991_ ) );
NOR3_X1 _13804_ ( .A1(_05972_ ), .A2(_05976_ ), .A3(_05183_ ), .ZN(_05992_ ) );
NOR3_X1 _13805_ ( .A1(_05988_ ), .A2(_05991_ ), .A3(_05992_ ), .ZN(_05993_ ) );
NAND2_X2 _13806_ ( .A1(_05985_ ), .A2(_05993_ ), .ZN(_05994_ ) );
BUF_X2 _13807_ ( .A(_05994_ ), .Z(_05995_ ) );
NOR2_X1 _13808_ ( .A1(_05181_ ), .A2(io_master_rlast ), .ZN(_05996_ ) );
OR2_X1 _13809_ ( .A1(_05995_ ), .A2(_05996_ ), .ZN(_05997_ ) );
INV_X1 _13810_ ( .A(\myifu.tmp_offset [2] ), .ZN(_05998_ ) );
AND3_X1 _13811_ ( .A1(_05997_ ), .A2(_01698_ ), .A3(_05998_ ), .ZN(_00279_ ) );
NOR3_X1 _13812_ ( .A1(fanout_net_4 ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00280_ ) );
AND3_X1 _13813_ ( .A1(_02106_ ), .A2(_05428_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_05999_ ) );
INV_X1 _13814_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_06000_ ) );
MUX2_X1 _13815_ ( .A(_02106_ ), .B(_06000_ ), .S(\myifu.to_reset ), .Z(_06001_ ) );
AOI211_X1 _13816_ ( .A(fanout_net_4 ), .B(_05999_ ), .C1(_06001_ ), .C2(\myifu.state [1] ), .ZN(_00281_ ) );
INV_X1 _13817_ ( .A(\myec.state [0] ), .ZN(_06002_ ) );
NOR2_X1 _13818_ ( .A1(_06002_ ), .A2(\myec.state [1] ), .ZN(_06003_ ) );
INV_X1 _13819_ ( .A(\EX_LS_pc [2] ), .ZN(_06004_ ) );
NOR3_X1 _13820_ ( .A1(_03086_ ), .A2(_06003_ ), .A3(_06004_ ), .ZN(_00282_ ) );
NOR2_X1 _13821_ ( .A1(_03085_ ), .A2(_06003_ ), .ZN(_06005_ ) );
BUF_X2 _13822_ ( .A(_06005_ ), .Z(_06006_ ) );
AND2_X1 _13823_ ( .A1(_06006_ ), .A2(fanout_net_45 ), .ZN(_00283_ ) );
BUF_X4 _13824_ ( .A(_02039_ ), .Z(_06007_ ) );
AOI21_X1 _13825_ ( .A(\LS_WB_waddr_csreg [11] ), .B1(_06007_ ), .B2(\EX_LS_flag [2] ), .ZN(_06008_ ) );
NOR2_X1 _13826_ ( .A1(_02048_ ), .A2(_05191_ ), .ZN(_06009_ ) );
INV_X1 _13827_ ( .A(_06009_ ), .ZN(_06010_ ) );
NOR2_X1 _13828_ ( .A1(_01972_ ), .A2(\EX_LS_flag [1] ), .ZN(_06011_ ) );
OR2_X1 _13829_ ( .A1(_06011_ ), .A2(_02020_ ), .ZN(_06012_ ) );
NOR2_X1 _13830_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_06013_ ) );
AND2_X1 _13831_ ( .A1(_06013_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_06014_ ) );
NOR2_X1 _13832_ ( .A1(_06012_ ), .A2(_06014_ ), .ZN(_06015_ ) );
NAND2_X2 _13833_ ( .A1(_06010_ ), .A2(_06015_ ), .ZN(_06016_ ) );
BUF_X4 _13834_ ( .A(_06016_ ), .Z(_06017_ ) );
INV_X1 _13835_ ( .A(\EX_LS_dest_csreg_mem [11] ), .ZN(_06018_ ) );
BUF_X4 _13836_ ( .A(_02173_ ), .Z(_06019_ ) );
AOI211_X1 _13837_ ( .A(_06008_ ), .B(_06017_ ), .C1(_06018_ ), .C2(_06019_ ), .ZN(_00284_ ) );
BUF_X4 _13838_ ( .A(_02021_ ), .Z(_06020_ ) );
NOR2_X1 _13839_ ( .A1(_06009_ ), .A2(_06014_ ), .ZN(_06021_ ) );
INV_X1 _13840_ ( .A(_06021_ ), .ZN(_06022_ ) );
NAND3_X1 _13841_ ( .A1(_06007_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_06023_ ) );
BUF_X4 _13842_ ( .A(_01972_ ), .Z(_06024_ ) );
NAND2_X1 _13843_ ( .A1(_06024_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06025_ ) );
AOI211_X1 _13844_ ( .A(_06020_ ), .B(_06022_ ), .C1(_06023_ ), .C2(_06025_ ), .ZN(_00285_ ) );
NAND3_X1 _13845_ ( .A1(_06007_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_06026_ ) );
NAND2_X1 _13846_ ( .A1(_06024_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06027_ ) );
AOI211_X1 _13847_ ( .A(_06020_ ), .B(_06022_ ), .C1(_06026_ ), .C2(_06027_ ), .ZN(_00286_ ) );
NAND3_X1 _13848_ ( .A1(_06007_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_06028_ ) );
NAND2_X1 _13849_ ( .A1(_06024_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_06029_ ) );
AOI211_X1 _13850_ ( .A(_06020_ ), .B(_06022_ ), .C1(_06028_ ), .C2(_06029_ ), .ZN(_00287_ ) );
NAND3_X1 _13851_ ( .A1(_06007_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_06030_ ) );
NAND2_X1 _13852_ ( .A1(_06024_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06031_ ) );
AOI211_X1 _13853_ ( .A(_06020_ ), .B(_06022_ ), .C1(_06030_ ), .C2(_06031_ ), .ZN(_00288_ ) );
NAND3_X1 _13854_ ( .A1(_06007_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_06032_ ) );
NAND2_X1 _13855_ ( .A1(_06024_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_06033_ ) );
AOI211_X1 _13856_ ( .A(_06020_ ), .B(_06022_ ), .C1(_06032_ ), .C2(_06033_ ), .ZN(_00289_ ) );
NAND3_X1 _13857_ ( .A1(_06007_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_06034_ ) );
NAND2_X1 _13858_ ( .A1(_06024_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_06035_ ) );
AOI211_X1 _13859_ ( .A(_06020_ ), .B(_06022_ ), .C1(_06034_ ), .C2(_06035_ ), .ZN(_00290_ ) );
NAND3_X1 _13860_ ( .A1(_06007_ ), .A2(fanout_net_6 ), .A3(\EX_LS_flag [2] ), .ZN(_06036_ ) );
NAND2_X1 _13861_ ( .A1(_06024_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_06037_ ) );
AOI211_X1 _13862_ ( .A(_06020_ ), .B(_06022_ ), .C1(_06036_ ), .C2(_06037_ ), .ZN(_00291_ ) );
INV_X1 _13863_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_06038_ ) );
AND4_X1 _13864_ ( .A1(_06038_ ), .A2(_02169_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06039_ ) );
NOR2_X1 _13865_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_06040_ ) );
OAI211_X1 _13866_ ( .A(_06021_ ), .B(_05188_ ), .C1(_06039_ ), .C2(_06040_ ), .ZN(_00292_ ) );
INV_X1 _13867_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_06041_ ) );
AND4_X1 _13868_ ( .A1(_06041_ ), .A2(_02169_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06042_ ) );
NOR2_X1 _13869_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06043_ ) );
OAI211_X1 _13870_ ( .A(_06021_ ), .B(_05188_ ), .C1(_06042_ ), .C2(_06043_ ), .ZN(_00293_ ) );
AND4_X1 _13871_ ( .A1(_04424_ ), .A2(_02169_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06044_ ) );
NOR2_X1 _13872_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06045_ ) );
OAI211_X1 _13873_ ( .A(_06021_ ), .B(_05188_ ), .C1(_06044_ ), .C2(_06045_ ), .ZN(_00294_ ) );
INV_X1 _13874_ ( .A(fanout_net_5 ), .ZN(_06046_ ) );
AND4_X1 _13875_ ( .A1(_06046_ ), .A2(_02169_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06047_ ) );
NOR2_X1 _13876_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_06048_ ) );
OAI211_X1 _13877_ ( .A(_06021_ ), .B(_05188_ ), .C1(_06047_ ), .C2(_06048_ ), .ZN(_00295_ ) );
NOR3_X1 _13878_ ( .A1(_03085_ ), .A2(_06003_ ), .A3(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06049_ ) );
NOR2_X1 _13879_ ( .A1(fanout_net_45 ), .A2(\mylsu.state [1] ), .ZN(_06050_ ) );
NAND2_X1 _13880_ ( .A1(_06049_ ), .A2(_06050_ ), .ZN(_06051_ ) );
BUF_X2 _13881_ ( .A(_01972_ ), .Z(_06052_ ) );
NOR2_X1 _13882_ ( .A1(_02111_ ), .A2(_02113_ ), .ZN(_06053_ ) );
AOI21_X1 _13883_ ( .A(_06052_ ), .B1(_06053_ ), .B2(_02038_ ), .ZN(_06054_ ) );
NOR3_X1 _13884_ ( .A1(_06009_ ), .A2(_06014_ ), .A3(_06054_ ), .ZN(_06055_ ) );
AOI21_X1 _13885_ ( .A(_06051_ ), .B1(_06055_ ), .B2(_02037_ ), .ZN(_00296_ ) );
INV_X1 _13886_ ( .A(_06007_ ), .ZN(_06056_ ) );
AOI21_X1 _13887_ ( .A(_02103_ ), .B1(_06056_ ), .B2(_06054_ ), .ZN(_06057_ ) );
AOI21_X1 _13888_ ( .A(_06051_ ), .B1(_06057_ ), .B2(_06021_ ), .ZN(_00297_ ) );
NAND3_X1 _13889_ ( .A1(_06053_ ), .A2(\EX_LS_flag [2] ), .A3(_02020_ ), .ZN(_06058_ ) );
NOR2_X1 _13890_ ( .A1(_06058_ ), .A2(_06051_ ), .ZN(_00298_ ) );
BUF_X4 _13891_ ( .A(_06010_ ), .Z(_06059_ ) );
AOI21_X1 _13892_ ( .A(_06051_ ), .B1(_06059_ ), .B2(_02037_ ), .ZN(_00299_ ) );
AOI21_X1 _13893_ ( .A(_06051_ ), .B1(_06021_ ), .B2(_06058_ ), .ZN(_00300_ ) );
INV_X1 _13894_ ( .A(_06014_ ), .ZN(_06060_ ) );
AND2_X1 _13895_ ( .A1(_06060_ ), .A2(_06005_ ), .ZN(_06061_ ) );
NOR3_X1 _13896_ ( .A1(_05187_ ), .A2(fanout_net_45 ), .A3(\mylsu.state [1] ), .ZN(_06062_ ) );
OAI211_X1 _13897_ ( .A(_06061_ ), .B(_06062_ ), .C1(_02044_ ), .C2(_02046_ ), .ZN(_06063_ ) );
NOR3_X1 _13898_ ( .A1(_02113_ ), .A2(_06007_ ), .A3(_01972_ ), .ZN(_06064_ ) );
OAI21_X1 _13899_ ( .A(_06064_ ), .B1(_02111_ ), .B2(\EX_LS_flag [1] ), .ZN(_06065_ ) );
NOR2_X1 _13900_ ( .A1(_05186_ ), .A2(_06065_ ), .ZN(_06066_ ) );
OAI211_X1 _13901_ ( .A(_06020_ ), .B(_02036_ ), .C1(_06066_ ), .C2(_02019_ ), .ZN(_06067_ ) );
INV_X1 _13902_ ( .A(_02041_ ), .ZN(_06068_ ) );
AND2_X1 _13903_ ( .A1(_06068_ ), .A2(_06065_ ), .ZN(_06069_ ) );
AOI21_X1 _13904_ ( .A(_06063_ ), .B1(_06067_ ), .B2(_06069_ ), .ZN(_00301_ ) );
INV_X1 _13905_ ( .A(_00283_ ), .ZN(_06070_ ) );
OAI211_X1 _13906_ ( .A(_06006_ ), .B(_06062_ ), .C1(_06019_ ), .C2(_02170_ ), .ZN(_06071_ ) );
OAI21_X1 _13907_ ( .A(_06070_ ), .B1(_02041_ ), .B2(_06071_ ), .ZN(_00302_ ) );
INV_X1 _13908_ ( .A(\mysc.state [2] ), .ZN(_06072_ ) );
NOR2_X1 _13909_ ( .A1(_06072_ ), .A2(fanout_net_4 ), .ZN(_00303_ ) );
AND3_X1 _13910_ ( .A1(_01584_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00093_ ) );
AND2_X1 _13911_ ( .A1(_02056_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _13912_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .ZN(_06073_ ) );
BUF_X2 _13913_ ( .A(_06073_ ), .Z(_06074_ ) );
AND3_X1 _13914_ ( .A1(_02056_ ), .A2(_06074_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00242_ ) );
NAND2_X1 _13915_ ( .A1(_05905_ ), .A2(fanout_net_9 ), .ZN(_06075_ ) );
INV_X1 _13916_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_06076_ ) );
BUF_X4 _13917_ ( .A(_06076_ ), .Z(_06077_ ) );
NOR3_X1 _13918_ ( .A1(_02057_ ), .A2(_06075_ ), .A3(_06077_ ), .ZN(_00243_ ) );
NAND2_X1 _13919_ ( .A1(_05916_ ), .A2(fanout_net_13 ), .ZN(_06078_ ) );
NOR3_X1 _13920_ ( .A1(_02057_ ), .A2(_06078_ ), .A3(_06077_ ), .ZN(_00244_ ) );
BUF_X2 _13921_ ( .A(_02055_ ), .Z(\io_master_arburst [0] ) );
BUF_X2 _13922_ ( .A(_01985_ ), .Z(_06079_ ) );
NOR3_X1 _13923_ ( .A1(_06079_ ), .A2(fanout_net_6 ), .A3(_05187_ ), .ZN(_06080_ ) );
BUF_X4 _13924_ ( .A(_05185_ ), .Z(_06081_ ) );
BUF_X4 _13925_ ( .A(_06081_ ), .Z(_06082_ ) );
INV_X1 _13926_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06083_ ) );
AOI211_X1 _13927_ ( .A(_06080_ ), .B(_06082_ ), .C1(_06083_ ), .C2(_02015_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _13928_ ( .A1(_06079_ ), .A2(fanout_net_5 ), .A3(_05187_ ), .ZN(_06084_ ) );
INV_X1 _13929_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06085_ ) );
AOI211_X1 _13930_ ( .A(_06084_ ), .B(_06082_ ), .C1(_06085_ ), .C2(_02015_ ), .ZN(\io_master_araddr [0] ) );
NOR2_X1 _13931_ ( .A1(_02088_ ), .A2(\mylsu.araddr_tmp [15] ), .ZN(_06086_ ) );
NOR3_X1 _13932_ ( .A1(_06079_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(_02005_ ), .ZN(_06087_ ) );
NOR3_X1 _13933_ ( .A1(_01977_ ), .A2(_06086_ ), .A3(_06087_ ), .ZN(_06088_ ) );
MUX2_X1 _13934_ ( .A(_06088_ ), .B(\IF_ID_pc [15] ), .S(\io_master_arburst [0] ), .Z(\io_master_araddr [15] ) );
MUX2_X1 _13935_ ( .A(\mylsu.araddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_02088_ ), .Z(_06089_ ) );
INV_X1 _13936_ ( .A(_01977_ ), .ZN(_06090_ ) );
AND2_X1 _13937_ ( .A1(_06089_ ), .A2(_06090_ ), .ZN(_06091_ ) );
MUX2_X1 _13938_ ( .A(_06091_ ), .B(\IF_ID_pc [14] ), .S(\io_master_arburst [0] ), .Z(\io_master_araddr [14] ) );
AND2_X1 _13939_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _13940_ ( .A1(_02020_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_04421_ ), .A4(_06052_ ), .ZN(_06092_ ) );
OAI21_X1 _13941_ ( .A(_06092_ ), .B1(_02088_ ), .B2(\mylsu.araddr_tmp [5] ), .ZN(_06093_ ) );
BUF_X4 _13942_ ( .A(_01998_ ), .Z(_06094_ ) );
BUF_X4 _13943_ ( .A(_06094_ ), .Z(_06095_ ) );
OAI22_X1 _13944_ ( .A1(_06082_ ), .A2(_06093_ ), .B1(_05689_ ), .B2(_06095_ ), .ZN(\io_master_araddr [5] ) );
AND4_X1 _13945_ ( .A1(\EX_LS_dest_csreg_mem [4] ), .A2(_02020_ ), .A3(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A4(_06052_ ), .ZN(_06096_ ) );
AOI21_X1 _13946_ ( .A(_06096_ ), .B1(_02015_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_06097_ ) );
OAI22_X1 _13947_ ( .A1(_06082_ ), .A2(_06097_ ), .B1(_05905_ ), .B2(_06095_ ), .ZN(\io_master_araddr [4] ) );
NAND4_X1 _13948_ ( .A1(_02020_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_04426_ ), .A4(_06052_ ), .ZN(_06098_ ) );
OAI21_X1 _13949_ ( .A(_06098_ ), .B1(_02088_ ), .B2(\mylsu.araddr_tmp [3] ), .ZN(_06099_ ) );
OAI22_X1 _13950_ ( .A1(_06082_ ), .A2(_06099_ ), .B1(_05916_ ), .B2(_06095_ ), .ZN(\io_master_araddr [3] ) );
OAI221_X1 _13951_ ( .A(\IF_ID_pc [13] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01988_ ), .C2(_01968_ ), .ZN(_06100_ ) );
OR3_X1 _13952_ ( .A1(_06079_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(_02005_ ), .ZN(_06101_ ) );
OAI211_X1 _13953_ ( .A(_06090_ ), .B(_06101_ ), .C1(\mylsu.araddr_tmp [13] ), .C2(_02088_ ), .ZN(_06102_ ) );
OAI21_X1 _13954_ ( .A(_06100_ ), .B1(\io_master_arburst [0] ), .B2(_06102_ ), .ZN(\io_master_araddr [13] ) );
MUX2_X1 _13955_ ( .A(\mylsu.araddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_02088_ ), .Z(_06103_ ) );
AND2_X1 _13956_ ( .A1(_06103_ ), .A2(_06090_ ), .ZN(_06104_ ) );
MUX2_X1 _13957_ ( .A(_06104_ ), .B(\IF_ID_pc [12] ), .S(\io_master_arburst [0] ), .Z(\io_master_araddr [12] ) );
NOR3_X1 _13958_ ( .A1(_06079_ ), .A2(_06018_ ), .A3(_05187_ ), .ZN(_06105_ ) );
AOI21_X1 _13959_ ( .A(_06105_ ), .B1(_02015_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_06106_ ) );
OAI22_X1 _13960_ ( .A1(_06082_ ), .A2(_06106_ ), .B1(_05724_ ), .B2(_06095_ ), .ZN(\io_master_araddr [11] ) );
OR3_X1 _13961_ ( .A1(_06079_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(_05187_ ), .ZN(_06107_ ) );
OAI21_X1 _13962_ ( .A(_06107_ ), .B1(_02088_ ), .B2(\mylsu.araddr_tmp [10] ), .ZN(_06108_ ) );
OAI22_X1 _13963_ ( .A1(_06082_ ), .A2(_06108_ ), .B1(_05717_ ), .B2(_06095_ ), .ZN(\io_master_araddr [10] ) );
NOR3_X1 _13964_ ( .A1(_06079_ ), .A2(_06038_ ), .A3(_05187_ ), .ZN(_06109_ ) );
AOI21_X1 _13965_ ( .A(_06109_ ), .B1(_02015_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06110_ ) );
OAI22_X1 _13966_ ( .A1(_06082_ ), .A2(_06110_ ), .B1(_05720_ ), .B2(_06095_ ), .ZN(\io_master_araddr [9] ) );
NAND4_X1 _13967_ ( .A1(_02020_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_06041_ ), .A4(_06052_ ), .ZN(_06111_ ) );
OAI21_X1 _13968_ ( .A(_06111_ ), .B1(_02088_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_06112_ ) );
OAI22_X1 _13969_ ( .A1(_06082_ ), .A2(_06112_ ), .B1(_05705_ ), .B2(_06095_ ), .ZN(\io_master_araddr [8] ) );
OAI221_X1 _13970_ ( .A(\IF_ID_pc [7] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01988_ ), .C2(_01968_ ), .ZN(_06113_ ) );
OR3_X1 _13971_ ( .A1(_06079_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(_02005_ ), .ZN(_06114_ ) );
OAI211_X1 _13972_ ( .A(_06090_ ), .B(_06114_ ), .C1(\mylsu.araddr_tmp [7] ), .C2(_02088_ ), .ZN(_06115_ ) );
OAI21_X1 _13973_ ( .A(_06113_ ), .B1(\io_master_arburst [0] ), .B2(_06115_ ), .ZN(\io_master_araddr [7] ) );
NOR3_X1 _13974_ ( .A1(_06079_ ), .A2(_04424_ ), .A3(_05187_ ), .ZN(_06116_ ) );
AOI21_X1 _13975_ ( .A(_06116_ ), .B1(_02015_ ), .B2(\mylsu.araddr_tmp [6] ), .ZN(_06117_ ) );
OAI22_X1 _13976_ ( .A1(_06082_ ), .A2(_06117_ ), .B1(_01955_ ), .B2(_06095_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _13977_ ( .A1(_06079_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(_02005_ ), .ZN(_06118_ ) );
OAI211_X1 _13978_ ( .A(_06090_ ), .B(_06118_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01995_ ), .ZN(_06119_ ) );
CLKBUF_X2 _13979_ ( .A(_06119_ ), .Z(_06120_ ) );
NOR2_X1 _13980_ ( .A1(_01971_ ), .A2(_06120_ ), .ZN(_06121_ ) );
BUF_X4 _13981_ ( .A(_06121_ ), .Z(_06122_ ) );
BUF_X4 _13982_ ( .A(_06122_ ), .Z(_06123_ ) );
BUF_X2 _13983_ ( .A(_06123_ ), .Z(\io_master_araddr [2] ) );
CLKBUF_X2 _13984_ ( .A(_02000_ ), .Z(\io_master_arid [1] ) );
NOR3_X1 _13985_ ( .A1(\io_master_arburst [0] ), .A2(_02026_ ), .A3(_01977_ ), .ZN(\io_master_arsize [2] ) );
INV_X1 _13986_ ( .A(\EX_LS_typ [1] ), .ZN(_06124_ ) );
NOR3_X1 _13987_ ( .A1(\io_master_arburst [0] ), .A2(_06124_ ), .A3(_01977_ ), .ZN(\io_master_arsize [0] ) );
INV_X1 _13988_ ( .A(\EX_LS_typ [2] ), .ZN(_06125_ ) );
OAI22_X1 _13989_ ( .A1(_01969_ ), .A2(_01970_ ), .B1(_06125_ ), .B2(_01977_ ), .ZN(\io_master_arsize [1] ) );
INV_X1 _13990_ ( .A(_05181_ ), .ZN(_06126_ ) );
AND3_X1 _13991_ ( .A1(_06126_ ), .A2(_02051_ ), .A3(_02058_ ), .ZN(io_master_arvalid ) );
AND2_X1 _13992_ ( .A1(_02040_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_06127_ ) );
BUF_X4 _13993_ ( .A(_06127_ ), .Z(_06128_ ) );
BUF_X4 _13994_ ( .A(_06128_ ), .Z(_06129_ ) );
MUX2_X1 _13995_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06129_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _13996_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06129_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _13997_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06129_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _13998_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06129_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _13999_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06129_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _14000_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06129_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _14001_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06129_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _14002_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06129_ ), .Z(\io_master_awaddr [16] ) );
BUF_X4 _14003_ ( .A(_06128_ ), .Z(_06130_ ) );
MUX2_X1 _14004_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06130_ ), .Z(\io_master_awaddr [15] ) );
MUX2_X1 _14005_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06130_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _14006_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06130_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _14007_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06130_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _14008_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06130_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _14009_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06130_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _14010_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06130_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _14011_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06130_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _14012_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06130_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _14013_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06130_ ), .Z(\io_master_awaddr [7] ) );
BUF_X4 _14014_ ( .A(_06128_ ), .Z(_06131_ ) );
MUX2_X1 _14015_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06131_ ), .Z(\io_master_awaddr [6] ) );
MUX2_X1 _14016_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06131_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _14017_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06131_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _14018_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06131_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _14019_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06131_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _14020_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06131_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _14021_ ( .A(\mylsu.awaddr_tmp [1] ), .B(fanout_net_6 ), .S(_06131_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _14022_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_5 ), .S(_06131_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _14023_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06131_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _14024_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06131_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _14025_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06128_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _14026_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06128_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _14027_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06128_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _14028_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06128_ ), .Z(\io_master_awaddr [22] ) );
NOR4_X1 _14029_ ( .A1(_06056_ ), .A2(_02030_ ), .A3(_02042_ ), .A4(_06124_ ), .ZN(\io_master_awsize [0] ) );
NAND2_X1 _14030_ ( .A1(_02043_ ), .A2(_02029_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _14031_ ( .A1(_02037_ ), .A2(_02048_ ), .A3(_06129_ ), .ZN(_06132_ ) );
INV_X1 _14032_ ( .A(\mylsu.state [4] ), .ZN(_06133_ ) );
NAND2_X1 _14033_ ( .A1(_06132_ ), .A2(_06133_ ), .ZN(io_master_awvalid ) );
INV_X1 _14034_ ( .A(\mylsu.state [2] ), .ZN(_06134_ ) );
INV_X1 _14035_ ( .A(\mylsu.state [1] ), .ZN(_06135_ ) );
NAND4_X1 _14036_ ( .A1(_06132_ ), .A2(_06134_ ), .A3(_06133_ ), .A4(_06135_ ), .ZN(io_master_bready ) );
NOR3_X1 _14037_ ( .A1(_01976_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_06136_ ) );
INV_X2 _14038_ ( .A(fanout_net_45 ), .ZN(_06137_ ) );
NAND3_X1 _14039_ ( .A1(_02014_ ), .A2(\io_master_arid [1] ), .A3(_02084_ ), .ZN(_06138_ ) );
NOR2_X1 _14040_ ( .A1(_05989_ ), .A2(\io_master_rid [0] ), .ZN(_06139_ ) );
NAND4_X1 _14041_ ( .A1(_06139_ ), .A2(io_master_rlast ), .A3(_05983_ ), .A4(_05987_ ), .ZN(_06140_ ) );
OAI21_X1 _14042_ ( .A(_06138_ ), .B1(_06081_ ), .B2(_06140_ ), .ZN(_06141_ ) );
AOI21_X1 _14043_ ( .A(_06137_ ), .B1(_05979_ ), .B2(_06141_ ), .ZN(_06142_ ) );
NOR2_X1 _14044_ ( .A1(\io_master_bid [3] ), .A2(\io_master_bid [2] ), .ZN(_06143_ ) );
AND3_X1 _14045_ ( .A1(_06143_ ), .A2(\io_master_bid [1] ), .A3(\io_master_bid [0] ), .ZN(_06144_ ) );
NOR2_X1 _14046_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_06145_ ) );
AND2_X1 _14047_ ( .A1(_06145_ ), .A2(io_master_bvalid ), .ZN(_06146_ ) );
AND2_X1 _14048_ ( .A1(_06144_ ), .A2(_06146_ ), .ZN(_06147_ ) );
INV_X1 _14049_ ( .A(_06147_ ), .ZN(_06148_ ) );
AOI211_X1 _14050_ ( .A(_06136_ ), .B(_06142_ ), .C1(\mylsu.state [1] ), .C2(_06148_ ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _14051_ ( .A(_02089_ ), .B(_02087_ ), .C1(_02014_ ), .C2(_02084_ ), .ZN(io_master_rready ) );
MUX2_X1 _14052_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_5 ), .Z(_06149_ ) );
CLKBUF_X2 _14053_ ( .A(_04420_ ), .Z(_06150_ ) );
AND2_X1 _14054_ ( .A1(_06149_ ), .A2(_06150_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _14055_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_5 ), .Z(_06151_ ) );
AND2_X1 _14056_ ( .A1(_06151_ ), .A2(_06150_ ), .ZN(\io_master_wdata [14] ) );
NOR3_X1 _14057_ ( .A1(_04915_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _14058_ ( .A1(_04934_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [4] ) );
NOR3_X1 _14059_ ( .A1(_04945_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14060_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_06152_ ) );
NOR3_X1 _14061_ ( .A1(_06152_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14062_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06153_ ) );
NOR3_X1 _14063_ ( .A1(_06153_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14064_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06154_ ) );
NOR3_X1 _14065_ ( .A1(_06154_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14066_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_5 ), .Z(_06155_ ) );
AND2_X1 _14067_ ( .A1(_06155_ ), .A2(_06150_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14068_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_5 ), .Z(_06156_ ) );
AND2_X1 _14069_ ( .A1(_06156_ ), .A2(_06150_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14070_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_5 ), .Z(_06157_ ) );
AND2_X1 _14071_ ( .A1(_06157_ ), .A2(_06150_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14072_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_5 ), .Z(_06158_ ) );
AND2_X1 _14073_ ( .A1(_06158_ ), .A2(_06150_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14074_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_5 ), .Z(_06159_ ) );
AND2_X1 _14075_ ( .A1(_06159_ ), .A2(_06150_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14076_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_5 ), .Z(_06160_ ) );
AND2_X1 _14077_ ( .A1(_06160_ ), .A2(_06150_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14078_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06161_ ) );
NOR3_X1 _14079_ ( .A1(_06161_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [7] ) );
NOR3_X1 _14080_ ( .A1(_04896_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14081_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_5 ), .Z(_06162_ ) );
MUX2_X1 _14082_ ( .A(_06162_ ), .B(_06149_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14083_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_5 ), .Z(_06163_ ) );
MUX2_X1 _14084_ ( .A(_06163_ ), .B(_06151_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [30] ) );
MUX2_X1 _14085_ ( .A(_05138_ ), .B(_04733_ ), .S(fanout_net_5 ), .Z(_06164_ ) );
NOR2_X1 _14086_ ( .A1(_04420_ ), .A2(fanout_net_5 ), .ZN(_06165_ ) );
INV_X1 _14087_ ( .A(_06165_ ), .ZN(_06166_ ) );
OAI22_X1 _14088_ ( .A1(_06164_ ), .A2(fanout_net_6 ), .B1(_06166_ ), .B2(_04915_ ), .ZN(\io_master_wdata [21] ) );
MUX2_X1 _14089_ ( .A(_04561_ ), .B(_04749_ ), .S(fanout_net_5 ), .Z(_06167_ ) );
OAI22_X1 _14090_ ( .A1(_06167_ ), .A2(fanout_net_6 ), .B1(_06166_ ), .B2(_04934_ ), .ZN(\io_master_wdata [20] ) );
INV_X1 _14091_ ( .A(\EX_LS_result_csreg_mem [19] ), .ZN(_06168_ ) );
MUX2_X1 _14092_ ( .A(_06168_ ), .B(_04771_ ), .S(fanout_net_5 ), .Z(_06169_ ) );
OAI22_X1 _14093_ ( .A1(_06169_ ), .A2(fanout_net_6 ), .B1(_06166_ ), .B2(_04945_ ), .ZN(\io_master_wdata [19] ) );
INV_X1 _14094_ ( .A(\EX_LS_result_csreg_mem [18] ), .ZN(_06170_ ) );
INV_X1 _14095_ ( .A(\EX_LS_result_csreg_mem [10] ), .ZN(_06171_ ) );
MUX2_X1 _14096_ ( .A(_06170_ ), .B(_06171_ ), .S(fanout_net_5 ), .Z(_06172_ ) );
OAI22_X1 _14097_ ( .A1(_06172_ ), .A2(fanout_net_6 ), .B1(_06166_ ), .B2(_06152_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _14098_ ( .A(_04420_ ), .B1(_06046_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_06173_ ) );
NOR2_X1 _14099_ ( .A1(fanout_net_5 ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_06174_ ) );
OAI22_X1 _14100_ ( .A1(_06166_ ), .A2(_06153_ ), .B1(_06173_ ), .B2(_06174_ ), .ZN(\io_master_wdata [17] ) );
MUX2_X1 _14101_ ( .A(_04664_ ), .B(_04854_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06175_ ) );
OAI22_X1 _14102_ ( .A1(_06175_ ), .A2(fanout_net_6 ), .B1(_06166_ ), .B2(_06154_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14103_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06176_ ) );
MUX2_X1 _14104_ ( .A(_06176_ ), .B(_06155_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14105_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06177_ ) );
MUX2_X1 _14106_ ( .A(_06177_ ), .B(_06156_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14107_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06178_ ) );
MUX2_X1 _14108_ ( .A(_06178_ ), .B(_06157_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14109_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06179_ ) );
MUX2_X1 _14110_ ( .A(_06179_ ), .B(_06158_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14111_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06180_ ) );
MUX2_X1 _14112_ ( .A(_06180_ ), .B(_06159_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14113_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06181_ ) );
MUX2_X1 _14114_ ( .A(_06181_ ), .B(_06160_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [24] ) );
OAI21_X1 _14115_ ( .A(_04420_ ), .B1(_06046_ ), .B2(\EX_LS_result_csreg_mem [15] ), .ZN(_06182_ ) );
NOR2_X1 _14116_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [23] ), .ZN(_06183_ ) );
OAI22_X1 _14117_ ( .A1(_06166_ ), .A2(_06161_ ), .B1(_06182_ ), .B2(_06183_ ), .ZN(\io_master_wdata [23] ) );
MUX2_X1 _14118_ ( .A(_05123_ ), .B(_04708_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06184_ ) );
OAI22_X1 _14119_ ( .A1(_06184_ ), .A2(fanout_net_6 ), .B1(_06166_ ), .B2(_04896_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14120_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06185_ ) );
AND2_X1 _14121_ ( .A1(_06185_ ), .A2(_06150_ ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _14122_ ( .A1(_06046_ ), .A2(_06150_ ), .A3(\EX_LS_typ [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14123_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06186_ ) );
MUX2_X1 _14124_ ( .A(_06186_ ), .B(_06185_ ), .S(fanout_net_6 ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14125_ ( .A1(_06046_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_typ [0] ), .ZN(_06187_ ) );
OAI221_X1 _14126_ ( .A(_06187_ ), .B1(_02025_ ), .B2(_06125_ ), .C1(\EX_LS_dest_csreg_mem [1] ), .C2(_02032_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _14127_ ( .A1(_06132_ ), .A2(_06134_ ), .ZN(io_master_wvalid ) );
MUX2_X1 _14128_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14129_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14130_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14131_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
NAND3_X1 _14132_ ( .A1(_01584_ ), .A2(\LS_WB_waddr_csreg [2] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_06188_ ) );
INV_X1 _14133_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_06189_ ) );
NOR4_X1 _14134_ ( .A1(_06188_ ), .A2(\LS_WB_waddr_csreg [3] ), .A3(\LS_WB_waddr_csreg [1] ), .A4(_06189_ ), .ZN(_06190_ ) );
NOR2_X1 _14135_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06191_ ) );
INV_X1 _14136_ ( .A(_06191_ ), .ZN(_06192_ ) );
NOR3_X1 _14137_ ( .A1(_06192_ ), .A2(\LS_WB_waddr_csreg [7] ), .A3(\LS_WB_waddr_csreg [6] ), .ZN(_06193_ ) );
AND2_X1 _14138_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06194_ ) );
NOR2_X1 _14139_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06195_ ) );
AND2_X1 _14140_ ( .A1(_06194_ ), .A2(_06195_ ), .ZN(_06196_ ) );
AND3_X1 _14141_ ( .A1(_06190_ ), .A2(_06193_ ), .A3(_06196_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ) );
AND2_X1 _14142_ ( .A1(_01583_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(_06197_ ) );
NOR3_X1 _14143_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .A3(\LS_WB_waddr_csreg [7] ), .ZN(_06198_ ) );
AND3_X1 _14144_ ( .A1(_06198_ ), .A2(\LS_WB_waddr_csreg [6] ), .A3(_06191_ ), .ZN(_06199_ ) );
NOR2_X1 _14145_ ( .A1(_06189_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_06200_ ) );
AND4_X1 _14146_ ( .A1(_06197_ ), .A2(_06199_ ), .A3(_06200_ ), .A4(_06196_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ) );
AND4_X1 _14147_ ( .A1(\LS_WB_waddr_csreg [6] ), .A2(_06196_ ), .A3(_06191_ ), .A4(_06198_ ), .ZN(_06201_ ) );
AND4_X1 _14148_ ( .A1(\LS_WB_waddr_csreg [1] ), .A2(_06201_ ), .A3(_06189_ ), .A4(_06197_ ), .ZN(_06202_ ) );
OR2_X1 _14149_ ( .A1(_06202_ ), .A2(_00093_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14150_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .A3(\LS_WB_waddr_csreg [1] ), .A4(\LS_WB_waddr_csreg [0] ), .ZN(_06203_ ) );
AND4_X1 _14151_ ( .A1(_06197_ ), .A2(_06193_ ), .A3(_06196_ ), .A4(_06203_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _14152_ ( .A1(_06053_ ), .A2(exception_quest_IDU ), .ZN(_06204_ ) );
NOR2_X1 _14153_ ( .A1(_02050_ ), .A2(_06204_ ), .ZN(_06205_ ) );
BUF_X4 _14154_ ( .A(_06205_ ), .Z(_06206_ ) );
MUX2_X1 _14155_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14156_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14157_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14158_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14159_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14160_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14161_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14162_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14163_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14164_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_06206_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14165_ ( .A(_06205_ ), .Z(_06207_ ) );
MUX2_X1 _14166_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14167_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14168_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14169_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14170_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14171_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14172_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14173_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14174_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14175_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_06207_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14176_ ( .A(_06205_ ), .Z(_06208_ ) );
MUX2_X1 _14177_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14178_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14179_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14180_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14181_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14182_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14183_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14184_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14185_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14186_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_06208_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14187_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_06205_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14188_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_06205_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
INV_X1 _14189_ ( .A(_02106_ ), .ZN(_06209_ ) );
NOR4_X1 _14190_ ( .A1(_02050_ ), .A2(exception_quest_IDU ), .A3(_06209_ ), .A4(_06204_ ), .ZN(_06210_ ) );
XNOR2_X1 _14191_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06211_ ) );
XNOR2_X1 _14192_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06212_ ) );
XNOR2_X1 _14193_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06213_ ) );
XNOR2_X1 _14194_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06214_ ) );
NAND4_X1 _14195_ ( .A1(_06211_ ), .A2(_06212_ ), .A3(_06213_ ), .A4(_06214_ ), .ZN(_06215_ ) );
XNOR2_X1 _14196_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06216_ ) );
XNOR2_X1 _14197_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06217_ ) );
XNOR2_X1 _14198_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06218_ ) );
XNOR2_X1 _14199_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06219_ ) );
NAND4_X1 _14200_ ( .A1(_06216_ ), .A2(_06217_ ), .A3(_06218_ ), .A4(_06219_ ), .ZN(_06220_ ) );
XNOR2_X1 _14201_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06221_ ) );
XNOR2_X1 _14202_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06222_ ) );
XNOR2_X1 _14203_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06223_ ) );
XNOR2_X1 _14204_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06224_ ) );
NAND4_X1 _14205_ ( .A1(_06221_ ), .A2(_06222_ ), .A3(_06223_ ), .A4(_06224_ ), .ZN(_06225_ ) );
XNOR2_X1 _14206_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06226_ ) );
XNOR2_X1 _14207_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06227_ ) );
XNOR2_X1 _14208_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06228_ ) );
XNOR2_X1 _14209_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06229_ ) );
NAND4_X1 _14210_ ( .A1(_06226_ ), .A2(_06227_ ), .A3(_06228_ ), .A4(_06229_ ), .ZN(_06230_ ) );
NOR4_X1 _14211_ ( .A1(_06215_ ), .A2(_06220_ ), .A3(_06225_ ), .A4(_06230_ ), .ZN(_06231_ ) );
XNOR2_X1 _14212_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06232_ ) );
XNOR2_X1 _14213_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06233_ ) );
XNOR2_X1 _14214_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06234_ ) );
XNOR2_X1 _14215_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06235_ ) );
AND4_X1 _14216_ ( .A1(_06232_ ), .A2(_06233_ ), .A3(_06234_ ), .A4(_06235_ ), .ZN(_06236_ ) );
XNOR2_X1 _14217_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06237_ ) );
XNOR2_X1 _14218_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06238_ ) );
XNOR2_X1 _14219_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06239_ ) );
XNOR2_X1 _14220_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06240_ ) );
AND4_X1 _14221_ ( .A1(_06237_ ), .A2(_06238_ ), .A3(_06239_ ), .A4(_06240_ ), .ZN(_06241_ ) );
XNOR2_X1 _14222_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_06242_ ) );
XNOR2_X1 _14223_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_06243_ ) );
XNOR2_X1 _14224_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_06244_ ) );
XNOR2_X1 _14225_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_06245_ ) );
AND4_X1 _14226_ ( .A1(_06242_ ), .A2(_06243_ ), .A3(_06244_ ), .A4(_06245_ ), .ZN(_06246_ ) );
XNOR2_X1 _14227_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06247_ ) );
XNOR2_X1 _14228_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06248_ ) );
XNOR2_X1 _14229_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06249_ ) );
XNOR2_X1 _14230_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06250_ ) );
AND4_X1 _14231_ ( .A1(_06247_ ), .A2(_06248_ ), .A3(_06249_ ), .A4(_06250_ ), .ZN(_06251_ ) );
AND4_X1 _14232_ ( .A1(_06236_ ), .A2(_06241_ ), .A3(_06246_ ), .A4(_06251_ ), .ZN(_06252_ ) );
NAND3_X1 _14233_ ( .A1(_06231_ ), .A2(excp_written ), .A3(_06252_ ), .ZN(_06253_ ) );
AOI21_X1 _14234_ ( .A(_06210_ ), .B1(_06209_ ), .B2(_06253_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14235_ ( .A1(_04988_ ), .A2(_03033_ ), .ZN(_06254_ ) );
AND2_X1 _14236_ ( .A1(_03029_ ), .A2(_02126_ ), .ZN(_06255_ ) );
BUF_X4 _14237_ ( .A(_06255_ ), .Z(_06256_ ) );
INV_X1 _14238_ ( .A(_06256_ ), .ZN(_06257_ ) );
BUF_X4 _14239_ ( .A(_06257_ ), .Z(_06258_ ) );
BUF_X4 _14240_ ( .A(_06258_ ), .Z(_06259_ ) );
OAI21_X1 _14241_ ( .A(_06254_ ), .B1(_04417_ ), .B2(_06259_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
NOR4_X1 _14242_ ( .A1(_05179_ ), .A2(_02121_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [0] ), .ZN(_06260_ ) );
XNOR2_X1 _14243_ ( .A(_04004_ ), .B(\ID_EX_imm [0] ), .ZN(_06261_ ) );
AOI21_X1 _14244_ ( .A(_06260_ ), .B1(_06261_ ), .B2(_03033_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND2_X1 _14245_ ( .A1(_05480_ ), .A2(\ID_EX_typ [7] ), .ZN(_06262_ ) );
INV_X2 _14246_ ( .A(_06262_ ), .ZN(_06263_ ) );
BUF_X4 _14247_ ( .A(_06263_ ), .Z(_06264_ ) );
AND2_X1 _14248_ ( .A1(_04814_ ), .A2(_06264_ ), .ZN(_06265_ ) );
BUF_X4 _14249_ ( .A(_06257_ ), .Z(_06266_ ) );
MUX2_X1 _14250_ ( .A(\ID_EX_csr [10] ), .B(_06265_ ), .S(_06266_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
NOR4_X1 _14251_ ( .A1(_05179_ ), .A2(_02121_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [9] ), .ZN(_06267_ ) );
AOI21_X1 _14252_ ( .A(_06267_ ), .B1(_04838_ ), .B2(_03033_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR2_X1 _14253_ ( .A1(_04858_ ), .A2(_06262_ ), .ZN(_06268_ ) );
MUX2_X1 _14254_ ( .A(\ID_EX_csr [8] ), .B(_06268_ ), .S(_06266_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _14255_ ( .A1(_04881_ ), .A2(_03033_ ), .ZN(_06269_ ) );
OAI21_X1 _14256_ ( .A(_06269_ ), .B1(_04458_ ), .B2(_06259_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
NOR2_X1 _14257_ ( .A1(_04900_ ), .A2(_03029_ ), .ZN(_06270_ ) );
BUF_X4 _14258_ ( .A(_06256_ ), .Z(_06271_ ) );
BUF_X4 _14259_ ( .A(_06271_ ), .Z(_06272_ ) );
AOI21_X1 _14260_ ( .A(_06270_ ), .B1(_04412_ ), .B2(_06272_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14261_ ( .A1(_04920_ ), .A2(_03033_ ), .ZN(_06273_ ) );
OAI21_X1 _14262_ ( .A(_06273_ ), .B1(_04418_ ), .B2(_06259_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
AND2_X1 _14263_ ( .A1(_04938_ ), .A2(_06263_ ), .ZN(_06274_ ) );
MUX2_X1 _14264_ ( .A(\ID_EX_csr [4] ), .B(_06274_ ), .S(_06266_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _14265_ ( .A1(_04955_ ), .A2(_03032_ ), .ZN(_06275_ ) );
OAI21_X1 _14266_ ( .A(_06275_ ), .B1(_04414_ ), .B2(_06259_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _14267_ ( .A1(_04972_ ), .A2(_03032_ ), .A3(_02792_ ), .ZN(_06276_ ) );
OAI21_X1 _14268_ ( .A(_06276_ ), .B1(_04446_ ), .B2(_06259_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
AND2_X1 _14269_ ( .A1(_04780_ ), .A2(_06263_ ), .ZN(_06277_ ) );
MUX2_X1 _14270_ ( .A(\ID_EX_csr [11] ), .B(_06277_ ), .S(_06266_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
NOR2_X2 _14271_ ( .A1(_04304_ ), .A2(\ID_EX_typ [2] ), .ZN(_06278_ ) );
INV_X1 _14272_ ( .A(_06278_ ), .ZN(_06279_ ) );
AND3_X1 _14273_ ( .A1(_04508_ ), .A2(_05138_ ), .A3(_04502_ ), .ZN(_06280_ ) );
NAND2_X1 _14274_ ( .A1(_05131_ ), .A2(_05132_ ), .ZN(_06281_ ) );
NOR2_X1 _14275_ ( .A1(_05159_ ), .A2(_06281_ ), .ZN(_06282_ ) );
AOI211_X1 _14276_ ( .A(_06279_ ), .B(_06280_ ), .C1(_06282_ ), .C2(_05136_ ), .ZN(_06283_ ) );
AOI22_X1 _14277_ ( .A1(_05140_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02362_ ), .ZN(_06284_ ) );
NAND3_X1 _14278_ ( .A1(_02361_ ), .A2(_02381_ ), .A3(_05027_ ), .ZN(_06285_ ) );
AOI21_X1 _14279_ ( .A(_06283_ ), .B1(_06284_ ), .B2(_06285_ ), .ZN(_06286_ ) );
NOR2_X1 _14280_ ( .A1(_06286_ ), .A2(_06266_ ), .ZN(_06287_ ) );
NOR2_X1 _14281_ ( .A1(_06263_ ), .A2(\ID_EX_pc [21] ), .ZN(_06288_ ) );
BUF_X4 _14282_ ( .A(_06263_ ), .Z(_06289_ ) );
AOI211_X1 _14283_ ( .A(_06256_ ), .B(_06288_ ), .C1(_03447_ ), .C2(_06289_ ), .ZN(_06290_ ) );
OR2_X1 _14284_ ( .A1(_06287_ ), .A2(_06290_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
BUF_X4 _14285_ ( .A(_06256_ ), .Z(_06291_ ) );
BUF_X4 _14286_ ( .A(_06291_ ), .Z(_06292_ ) );
OAI22_X1 _14287_ ( .A1(_04563_ ), .A2(_05195_ ), .B1(_05027_ ), .B2(\ID_EX_imm [20] ), .ZN(_06293_ ) );
AOI21_X1 _14288_ ( .A(_06293_ ), .B1(_05028_ ), .B2(_04251_ ), .ZN(_06294_ ) );
BUF_X4 _14289_ ( .A(_06278_ ), .Z(_06295_ ) );
NAND3_X1 _14290_ ( .A1(_04560_ ), .A2(_06295_ ), .A3(_04562_ ), .ZN(_06296_ ) );
INV_X1 _14291_ ( .A(_06296_ ), .ZN(_06297_ ) );
OAI21_X1 _14292_ ( .A(_06292_ ), .B1(_06294_ ), .B2(_06297_ ), .ZN(_06298_ ) );
BUF_X4 _14293_ ( .A(_06256_ ), .Z(_06299_ ) );
BUF_X4 _14294_ ( .A(_06299_ ), .Z(_06300_ ) );
MUX2_X1 _14295_ ( .A(_05146_ ), .B(_03426_ ), .S(_06289_ ), .Z(_06301_ ) );
OAI21_X1 _14296_ ( .A(_06298_ ), .B1(_06300_ ), .B2(_06301_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND3_X1 _14297_ ( .A1(_04590_ ), .A2(\ID_EX_typ [2] ), .A3(_04593_ ), .ZN(_06302_ ) );
BUF_X2 _14298_ ( .A(_04482_ ), .Z(_06303_ ) );
NAND2_X1 _14299_ ( .A1(_02524_ ), .A2(_06303_ ), .ZN(_06304_ ) );
NAND2_X1 _14300_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [19] ), .ZN(_06305_ ) );
AOI21_X1 _14301_ ( .A(_06302_ ), .B1(_06304_ ), .B2(_06305_ ), .ZN(_06306_ ) );
AOI21_X1 _14302_ ( .A(_06279_ ), .B1(_04590_ ), .B2(_04593_ ), .ZN(_06307_ ) );
OAI21_X1 _14303_ ( .A(_06292_ ), .B1(_06306_ ), .B2(_06307_ ), .ZN(_06308_ ) );
MUX2_X1 _14304_ ( .A(_04576_ ), .B(_03280_ ), .S(_06289_ ), .Z(_06309_ ) );
OAI21_X1 _14305_ ( .A(_06308_ ), .B1(_06300_ ), .B2(_06309_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
AND3_X1 _14306_ ( .A1(_04614_ ), .A2(\ID_EX_typ [2] ), .A3(_04615_ ), .ZN(_06310_ ) );
NAND2_X1 _14307_ ( .A1(_02501_ ), .A2(_06303_ ), .ZN(_06311_ ) );
NAND2_X1 _14308_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [18] ), .ZN(_06312_ ) );
AOI21_X1 _14309_ ( .A(_06310_ ), .B1(_06311_ ), .B2(_06312_ ), .ZN(_06313_ ) );
AOI21_X1 _14310_ ( .A(_06279_ ), .B1(_04614_ ), .B2(_04615_ ), .ZN(_06314_ ) );
OAI21_X1 _14311_ ( .A(_06292_ ), .B1(_06313_ ), .B2(_06314_ ), .ZN(_06315_ ) );
MUX2_X1 _14312_ ( .A(_05175_ ), .B(_03309_ ), .S(_06289_ ), .Z(_06316_ ) );
OAI21_X1 _14313_ ( .A(_06315_ ), .B1(_06300_ ), .B2(_06316_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
OAI22_X1 _14314_ ( .A1(_04645_ ), .A2(_05195_ ), .B1(_05027_ ), .B2(\ID_EX_imm [17] ), .ZN(_06317_ ) );
AOI21_X1 _14315_ ( .A(_06317_ ), .B1(_05028_ ), .B2(_02946_ ), .ZN(_06318_ ) );
INV_X1 _14316_ ( .A(_04644_ ), .ZN(_06319_ ) );
OR2_X1 _14317_ ( .A1(_05159_ ), .A2(_04641_ ), .ZN(_06320_ ) );
OAI211_X1 _14318_ ( .A(_06278_ ), .B(_06319_ ), .C1(_06320_ ), .C2(_04638_ ), .ZN(_06321_ ) );
INV_X1 _14319_ ( .A(_06321_ ), .ZN(_06322_ ) );
OAI21_X1 _14320_ ( .A(_06292_ ), .B1(_06318_ ), .B2(_06322_ ), .ZN(_06323_ ) );
MUX2_X1 _14321_ ( .A(_04627_ ), .B(_03356_ ), .S(_06289_ ), .Z(_06324_ ) );
OAI21_X1 _14322_ ( .A(_06323_ ), .B1(_06300_ ), .B2(_06324_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
OAI22_X1 _14323_ ( .A1(_04666_ ), .A2(_05195_ ), .B1(_05027_ ), .B2(\ID_EX_imm [16] ), .ZN(_06325_ ) );
AOI21_X1 _14324_ ( .A(_06325_ ), .B1(_05028_ ), .B2(_04219_ ), .ZN(_06326_ ) );
NAND3_X1 _14325_ ( .A1(_04663_ ), .A2(_06295_ ), .A3(_04665_ ), .ZN(_06327_ ) );
INV_X1 _14326_ ( .A(_06327_ ), .ZN(_06328_ ) );
OAI21_X1 _14327_ ( .A(_06292_ ), .B1(_06326_ ), .B2(_06328_ ), .ZN(_06329_ ) );
MUX2_X1 _14328_ ( .A(_04650_ ), .B(_03333_ ), .S(_06264_ ), .Z(_06330_ ) );
OAI21_X1 _14329_ ( .A(_06329_ ), .B1(_06300_ ), .B2(_06330_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
OAI211_X1 _14330_ ( .A(_03029_ ), .B(_02126_ ), .C1(_05027_ ), .C2(\ID_EX_imm [15] ), .ZN(_06331_ ) );
AOI21_X1 _14331_ ( .A(_06331_ ), .B1(_04184_ ), .B2(_06303_ ), .ZN(_06332_ ) );
OAI21_X1 _14332_ ( .A(_06332_ ), .B1(_05195_ ), .B2(_04678_ ), .ZN(_06333_ ) );
BUF_X4 _14333_ ( .A(_06278_ ), .Z(_06334_ ) );
BUF_X4 _14334_ ( .A(_06256_ ), .Z(_06335_ ) );
NAND3_X1 _14335_ ( .A1(_04678_ ), .A2(_06334_ ), .A3(_06335_ ), .ZN(_06336_ ) );
MUX2_X1 _14336_ ( .A(_04623_ ), .B(_03771_ ), .S(_06263_ ), .Z(_06337_ ) );
OAI211_X1 _14337_ ( .A(_06333_ ), .B(_06336_ ), .C1(_06272_ ), .C2(_06337_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
BUF_X4 _14338_ ( .A(_06291_ ), .Z(_06338_ ) );
OAI22_X1 _14339_ ( .A1(_04710_ ), .A2(_05195_ ), .B1(_05027_ ), .B2(\ID_EX_imm [14] ), .ZN(_06339_ ) );
AOI21_X1 _14340_ ( .A(_06339_ ), .B1(_05028_ ), .B2(_04166_ ), .ZN(_06340_ ) );
NAND3_X1 _14341_ ( .A1(_04707_ ), .A2(_06295_ ), .A3(_04709_ ), .ZN(_06341_ ) );
INV_X1 _14342_ ( .A(_06341_ ), .ZN(_06342_ ) );
OAI21_X1 _14343_ ( .A(_06338_ ), .B1(_06340_ ), .B2(_06342_ ), .ZN(_06343_ ) );
MUX2_X1 _14344_ ( .A(_04624_ ), .B(_03793_ ), .S(_06264_ ), .Z(_06344_ ) );
OAI21_X1 _14345_ ( .A(_06343_ ), .B1(_06300_ ), .B2(_06344_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
AND2_X1 _14346_ ( .A1(_04729_ ), .A2(_04496_ ), .ZN(_06345_ ) );
NAND3_X1 _14347_ ( .A1(_04554_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_04455_ ), .ZN(_06346_ ) );
AND2_X1 _14348_ ( .A1(_04730_ ), .A2(_06346_ ), .ZN(_06347_ ) );
AOI21_X1 _14349_ ( .A(_04727_ ), .B1(_04502_ ), .B2(_04508_ ), .ZN(_06348_ ) );
NAND3_X1 _14350_ ( .A1(_06345_ ), .A2(_06347_ ), .A3(_06348_ ), .ZN(_06349_ ) );
NAND3_X1 _14351_ ( .A1(_04511_ ), .A2(_04733_ ), .A3(_04513_ ), .ZN(_06350_ ) );
AND2_X1 _14352_ ( .A1(_06349_ ), .A2(_06350_ ), .ZN(_06351_ ) );
OAI22_X1 _14353_ ( .A1(_06351_ ), .A2(_05194_ ), .B1(_05027_ ), .B2(\ID_EX_imm [13] ), .ZN(_06352_ ) );
INV_X1 _14354_ ( .A(_02600_ ), .ZN(_06353_ ) );
AOI21_X1 _14355_ ( .A(_06352_ ), .B1(_05028_ ), .B2(_06353_ ), .ZN(_06354_ ) );
NAND3_X1 _14356_ ( .A1(_06349_ ), .A2(_06295_ ), .A3(_06350_ ), .ZN(_06355_ ) );
INV_X1 _14357_ ( .A(_06355_ ), .ZN(_06356_ ) );
OAI21_X1 _14358_ ( .A(_06338_ ), .B1(_06354_ ), .B2(_06356_ ), .ZN(_06357_ ) );
MUX2_X1 _14359_ ( .A(_04717_ ), .B(_03838_ ), .S(_06264_ ), .Z(_06358_ ) );
OAI21_X1 _14360_ ( .A(_06357_ ), .B1(_06300_ ), .B2(_06358_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AND2_X1 _14361_ ( .A1(_04748_ ), .A2(_04750_ ), .ZN(_06359_ ) );
OAI22_X1 _14362_ ( .A1(_06359_ ), .A2(_05194_ ), .B1(_04482_ ), .B2(\ID_EX_imm [12] ), .ZN(_06360_ ) );
AOI21_X1 _14363_ ( .A(_06360_ ), .B1(_05028_ ), .B2(_04179_ ), .ZN(_06361_ ) );
AND3_X1 _14364_ ( .A1(_04748_ ), .A2(_06278_ ), .A3(_04750_ ), .ZN(_06362_ ) );
OAI21_X1 _14365_ ( .A(_06338_ ), .B1(_06361_ ), .B2(_06362_ ), .ZN(_06363_ ) );
MUX2_X1 _14366_ ( .A(_04715_ ), .B(_03816_ ), .S(_06264_ ), .Z(_06364_ ) );
OAI21_X1 _14367_ ( .A(_06363_ ), .B1(_06300_ ), .B2(_06364_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
BUF_X2 _14368_ ( .A(_04508_ ), .Z(_06365_ ) );
BUF_X2 _14369_ ( .A(_04501_ ), .Z(_06366_ ) );
AND3_X1 _14370_ ( .A1(_06365_ ), .A2(_04430_ ), .A3(_06366_ ), .ZN(_06367_ ) );
NAND2_X1 _14371_ ( .A1(_04470_ ), .A2(_04497_ ), .ZN(_06368_ ) );
NOR2_X1 _14372_ ( .A1(_05159_ ), .A2(_06368_ ), .ZN(_06369_ ) );
AND3_X1 _14373_ ( .A1(_04465_ ), .A2(_04457_ ), .A3(_04477_ ), .ZN(_06370_ ) );
AOI21_X1 _14374_ ( .A(_06367_ ), .B1(_06369_ ), .B2(_06370_ ), .ZN(_06371_ ) );
AOI21_X1 _14375_ ( .A(fanout_net_7 ), .B1(_02197_ ), .B2(_02198_ ), .ZN(_06372_ ) );
AND2_X1 _14376_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [30] ), .ZN(_06373_ ) );
OAI221_X1 _14377_ ( .A(_06271_ ), .B1(_05195_ ), .B2(_06371_ ), .C1(_06372_ ), .C2(_06373_ ), .ZN(_06374_ ) );
AND2_X1 _14378_ ( .A1(_04470_ ), .A2(_04725_ ), .ZN(_06375_ ) );
NAND3_X1 _14379_ ( .A1(_05151_ ), .A2(_06370_ ), .A3(_06375_ ), .ZN(_06376_ ) );
INV_X1 _14380_ ( .A(_06367_ ), .ZN(_06377_ ) );
NAND4_X1 _14381_ ( .A1(_06376_ ), .A2(_06377_ ), .A3(_06295_ ), .A4(_06271_ ), .ZN(_06378_ ) );
AND3_X1 _14382_ ( .A1(_05480_ ), .A2(\ID_EX_pc [30] ), .A3(\ID_EX_typ [7] ), .ZN(_06379_ ) );
BUF_X4 _14383_ ( .A(_06263_ ), .Z(_06380_ ) );
AOI21_X1 _14384_ ( .A(_06379_ ), .B1(_03646_ ), .B2(_06380_ ), .ZN(_06381_ ) );
OAI211_X1 _14385_ ( .A(_06374_ ), .B(_06378_ ), .C1(_06272_ ), .C2(_06381_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
AND3_X1 _14386_ ( .A1(_04511_ ), .A2(_04771_ ), .A3(_04513_ ), .ZN(_06382_ ) );
INV_X1 _14387_ ( .A(_06382_ ), .ZN(_06383_ ) );
AND2_X1 _14388_ ( .A1(_04764_ ), .A2(_04765_ ), .ZN(_06384_ ) );
NAND2_X1 _14389_ ( .A1(_05151_ ), .A2(_06384_ ), .ZN(_06385_ ) );
INV_X1 _14390_ ( .A(_04767_ ), .ZN(_06386_ ) );
NAND3_X1 _14391_ ( .A1(_04473_ ), .A2(\mtvec [11] ), .A3(_04476_ ), .ZN(_06387_ ) );
NAND3_X1 _14392_ ( .A1(_06386_ ), .A2(_04549_ ), .A3(_06387_ ), .ZN(_06388_ ) );
OAI21_X1 _14393_ ( .A(_06383_ ), .B1(_06385_ ), .B2(_06388_ ), .ZN(_06389_ ) );
AOI22_X1 _14394_ ( .A1(_06389_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02695_ ), .ZN(_06390_ ) );
OAI211_X1 _14395_ ( .A(_06390_ ), .B(_06299_ ), .C1(fanout_net_7 ), .C2(_02694_ ), .ZN(_06391_ ) );
NOR4_X1 _14396_ ( .A1(_04767_ ), .A2(_04450_ ), .A3(_04548_ ), .A4(_04768_ ), .ZN(_06392_ ) );
NOR2_X1 _14397_ ( .A1(_05159_ ), .A2(_04766_ ), .ZN(_06393_ ) );
NAND2_X1 _14398_ ( .A1(_06392_ ), .A2(_06393_ ), .ZN(_06394_ ) );
NAND4_X1 _14399_ ( .A1(_06394_ ), .A2(_06334_ ), .A3(_06383_ ), .A4(_06271_ ), .ZN(_06395_ ) );
MUX2_X1 _14400_ ( .A(_03176_ ), .B(_03864_ ), .S(_06263_ ), .Z(_06396_ ) );
OAI211_X1 _14401_ ( .A(_06391_ ), .B(_06395_ ), .C1(_06272_ ), .C2(_06396_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AND3_X1 _14402_ ( .A1(_04809_ ), .A2(\ID_EX_typ [2] ), .A3(_04810_ ), .ZN(_06397_ ) );
NAND2_X1 _14403_ ( .A1(_02718_ ), .A2(_06303_ ), .ZN(_06398_ ) );
NAND2_X1 _14404_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [10] ), .ZN(_06399_ ) );
AOI21_X1 _14405_ ( .A(_06397_ ), .B1(_06398_ ), .B2(_06399_ ), .ZN(_06400_ ) );
AOI21_X1 _14406_ ( .A(_06279_ ), .B1(_04809_ ), .B2(_04810_ ), .ZN(_06401_ ) );
OAI21_X1 _14407_ ( .A(_06338_ ), .B1(_06400_ ), .B2(_06401_ ), .ZN(_06402_ ) );
MUX2_X1 _14408_ ( .A(_05176_ ), .B(_03886_ ), .S(_06264_ ), .Z(_06403_ ) );
OAI21_X1 _14409_ ( .A(_06402_ ), .B1(_06300_ ), .B2(_06403_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
AOI211_X1 _14410_ ( .A(_05194_ ), .B(_04830_ ), .C1(_04724_ ), .C2(_04828_ ), .ZN(_06404_ ) );
NAND2_X1 _14411_ ( .A1(_02670_ ), .A2(_06303_ ), .ZN(_06405_ ) );
NAND2_X1 _14412_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [9] ), .ZN(_06406_ ) );
AOI21_X1 _14413_ ( .A(_06404_ ), .B1(_06405_ ), .B2(_06406_ ), .ZN(_06407_ ) );
AOI21_X1 _14414_ ( .A(_06279_ ), .B1(_04829_ ), .B2(_04831_ ), .ZN(_06408_ ) );
OAI21_X1 _14415_ ( .A(_06338_ ), .B1(_06407_ ), .B2(_06408_ ), .ZN(_06409_ ) );
MUX2_X1 _14416_ ( .A(_05177_ ), .B(_03909_ ), .S(_06264_ ), .Z(_06410_ ) );
OAI21_X1 _14417_ ( .A(_06409_ ), .B1(_06300_ ), .B2(_06410_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
OAI22_X1 _14418_ ( .A1(_04856_ ), .A2(_05194_ ), .B1(_04482_ ), .B2(\ID_EX_imm [8] ), .ZN(_06411_ ) );
INV_X1 _14419_ ( .A(_02647_ ), .ZN(_06412_ ) );
AOI21_X1 _14420_ ( .A(_06411_ ), .B1(_05028_ ), .B2(_06412_ ), .ZN(_06413_ ) );
NAND3_X1 _14421_ ( .A1(_04853_ ), .A2(_06295_ ), .A3(_04855_ ), .ZN(_06414_ ) );
INV_X1 _14422_ ( .A(_06414_ ), .ZN(_06415_ ) );
OAI21_X1 _14423_ ( .A(_06338_ ), .B1(_06413_ ), .B2(_06415_ ), .ZN(_06416_ ) );
MUX2_X1 _14424_ ( .A(_04841_ ), .B(_03931_ ), .S(_06264_ ), .Z(_06417_ ) );
OAI21_X1 _14425_ ( .A(_06416_ ), .B1(_06272_ ), .B2(_06417_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
NAND3_X1 _14426_ ( .A1(_06365_ ), .A2(_06161_ ), .A3(_06366_ ), .ZN(_06418_ ) );
AND2_X1 _14427_ ( .A1(_04867_ ), .A2(_04870_ ), .ZN(_06419_ ) );
NAND3_X1 _14428_ ( .A1(_06419_ ), .A2(_04866_ ), .A3(_04869_ ), .ZN(_06420_ ) );
OAI211_X1 _14429_ ( .A(_06278_ ), .B(_06418_ ), .C1(_06420_ ), .C2(_05159_ ), .ZN(_06421_ ) );
INV_X1 _14430_ ( .A(_06421_ ), .ZN(_06422_ ) );
NOR2_X1 _14431_ ( .A1(_05027_ ), .A2(\ID_EX_imm [7] ), .ZN(_06423_ ) );
AOI21_X1 _14432_ ( .A(_06423_ ), .B1(_04874_ ), .B2(\ID_EX_typ [2] ), .ZN(_06424_ ) );
NAND3_X1 _14433_ ( .A1(_02894_ ), .A2(_02913_ ), .A3(_06303_ ), .ZN(_06425_ ) );
AOI211_X1 _14434_ ( .A(_06258_ ), .B(_06422_ ), .C1(_06424_ ), .C2(_06425_ ), .ZN(_06426_ ) );
MUX2_X1 _14435_ ( .A(_05178_ ), .B(_03672_ ), .S(_06289_ ), .Z(_06427_ ) );
AOI21_X1 _14436_ ( .A(_06426_ ), .B1(_06259_ ), .B2(_06427_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _14437_ ( .A1(_04898_ ), .A2(_05194_ ), .B1(_04482_ ), .B2(\ID_EX_imm [6] ), .ZN(_06428_ ) );
AOI21_X1 _14438_ ( .A(_06428_ ), .B1(_05028_ ), .B2(_02918_ ), .ZN(_06429_ ) );
NAND3_X1 _14439_ ( .A1(_04895_ ), .A2(_06295_ ), .A3(_04897_ ), .ZN(_06430_ ) );
INV_X1 _14440_ ( .A(_06430_ ), .ZN(_06431_ ) );
OAI21_X1 _14441_ ( .A(_06338_ ), .B1(_06429_ ), .B2(_06431_ ), .ZN(_06432_ ) );
MUX2_X1 _14442_ ( .A(_04883_ ), .B(_03702_ ), .S(_06264_ ), .Z(_06433_ ) );
OAI21_X1 _14443_ ( .A(_06432_ ), .B1(_06272_ ), .B2(_06433_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
NAND4_X1 _14444_ ( .A1(_04908_ ), .A2(_04909_ ), .A3(_04912_ ), .A4(_04497_ ), .ZN(_06434_ ) );
NOR3_X1 _14445_ ( .A1(_06434_ ), .A2(_05159_ ), .A3(_04910_ ), .ZN(_06435_ ) );
AND3_X1 _14446_ ( .A1(_04511_ ), .A2(_04915_ ), .A3(_04502_ ), .ZN(_06436_ ) );
NOR2_X1 _14447_ ( .A1(_06435_ ), .A2(_06436_ ), .ZN(_06437_ ) );
OAI22_X1 _14448_ ( .A1(_06437_ ), .A2(_05194_ ), .B1(_04482_ ), .B2(\ID_EX_imm [5] ), .ZN(_06438_ ) );
AOI21_X1 _14449_ ( .A(_06438_ ), .B1(_02923_ ), .B2(_06303_ ), .ZN(_06439_ ) );
AND3_X1 _14450_ ( .A1(_04908_ ), .A2(_04497_ ), .A3(_04912_ ), .ZN(_06440_ ) );
AOI21_X1 _14451_ ( .A(_04910_ ), .B1(_06366_ ), .B2(_06365_ ), .ZN(_06441_ ) );
NAND3_X1 _14452_ ( .A1(_06440_ ), .A2(_06441_ ), .A3(_04909_ ), .ZN(_06442_ ) );
NAND3_X1 _14453_ ( .A1(_06365_ ), .A2(_04915_ ), .A3(_06366_ ), .ZN(_06443_ ) );
NAND3_X1 _14454_ ( .A1(_06442_ ), .A2(_06278_ ), .A3(_06443_ ), .ZN(_06444_ ) );
INV_X1 _14455_ ( .A(_06444_ ), .ZN(_06445_ ) );
OAI21_X1 _14456_ ( .A(_06338_ ), .B1(_06439_ ), .B2(_06445_ ), .ZN(_06446_ ) );
AND4_X1 _14457_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06447_ ) );
AOI21_X1 _14458_ ( .A(_06447_ ), .B1(_03748_ ), .B2(_06380_ ), .ZN(_06448_ ) );
OAI21_X1 _14459_ ( .A(_06446_ ), .B1(_06272_ ), .B2(_06448_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
OAI22_X1 _14460_ ( .A1(_04936_ ), .A2(_05194_ ), .B1(_04482_ ), .B2(\ID_EX_imm [4] ), .ZN(_06449_ ) );
AOI21_X1 _14461_ ( .A(_06449_ ), .B1(_06303_ ), .B2(_04159_ ), .ZN(_06450_ ) );
AND3_X1 _14462_ ( .A1(_04928_ ), .A2(_04497_ ), .A3(_04930_ ), .ZN(_06451_ ) );
AOI21_X1 _14463_ ( .A(_04932_ ), .B1(_06366_ ), .B2(_06365_ ), .ZN(_06452_ ) );
NAND3_X1 _14464_ ( .A1(_06451_ ), .A2(_06452_ ), .A3(_04929_ ), .ZN(_06453_ ) );
NAND3_X1 _14465_ ( .A1(_06365_ ), .A2(_04934_ ), .A3(_06366_ ), .ZN(_06454_ ) );
NAND3_X1 _14466_ ( .A1(_06453_ ), .A2(_06278_ ), .A3(_06454_ ), .ZN(_06455_ ) );
INV_X1 _14467_ ( .A(_06455_ ), .ZN(_06456_ ) );
OAI21_X1 _14468_ ( .A(_06338_ ), .B1(_06450_ ), .B2(_06456_ ), .ZN(_06457_ ) );
MUX2_X1 _14469_ ( .A(_04922_ ), .B(_03726_ ), .S(_06264_ ), .Z(_06458_ ) );
OAI21_X1 _14470_ ( .A(_06457_ ), .B1(_06272_ ), .B2(_06458_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
AND3_X1 _14471_ ( .A1(_04950_ ), .A2(_04497_ ), .A3(_04947_ ), .ZN(_06459_ ) );
AND2_X1 _14472_ ( .A1(_04951_ ), .A2(_04948_ ), .ZN(_06460_ ) );
NAND3_X1 _14473_ ( .A1(_05151_ ), .A2(_06459_ ), .A3(_06460_ ), .ZN(_06461_ ) );
NAND3_X1 _14474_ ( .A1(_06365_ ), .A2(_04945_ ), .A3(_06366_ ), .ZN(_06462_ ) );
NAND2_X1 _14475_ ( .A1(_06461_ ), .A2(_06462_ ), .ZN(_06463_ ) );
AOI22_X1 _14476_ ( .A1(_06463_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02816_ ), .ZN(_06464_ ) );
OAI211_X1 _14477_ ( .A(_06464_ ), .B(_06299_ ), .C1(fanout_net_7 ), .C2(_02815_ ), .ZN(_06465_ ) );
NAND4_X1 _14478_ ( .A1(_06461_ ), .A2(_06334_ ), .A3(_06462_ ), .A4(_06271_ ), .ZN(_06466_ ) );
AND3_X1 _14479_ ( .A1(_05480_ ), .A2(\ID_EX_pc [3] ), .A3(\ID_EX_typ [7] ), .ZN(_06467_ ) );
AOI21_X1 _14480_ ( .A(_06467_ ), .B1(_03978_ ), .B2(_06380_ ), .ZN(_06468_ ) );
OAI211_X1 _14481_ ( .A(_06465_ ), .B(_06466_ ), .C1(_06272_ ), .C2(_06468_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
NAND2_X1 _14482_ ( .A1(_02741_ ), .A2(_04482_ ), .ZN(_06469_ ) );
NAND2_X1 _14483_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [2] ), .ZN(_06470_ ) );
AND2_X1 _14484_ ( .A1(_06469_ ), .A2(_06470_ ), .ZN(_06471_ ) );
OR2_X1 _14485_ ( .A1(_04969_ ), .A2(_06279_ ), .ZN(_06472_ ) );
AOI221_X4 _14486_ ( .A(_06257_ ), .B1(\ID_EX_typ [2] ), .B2(_04969_ ), .C1(_06471_ ), .C2(_06472_ ), .ZN(_06473_ ) );
NOR4_X1 _14487_ ( .A1(_05179_ ), .A2(_02121_ ), .A3(_02126_ ), .A4(\ID_EX_pc [2] ), .ZN(_06474_ ) );
AOI211_X1 _14488_ ( .A(_06256_ ), .B(_06474_ ), .C1(_03956_ ), .C2(_06289_ ), .ZN(_06475_ ) );
OR2_X1 _14489_ ( .A1(_06473_ ), .A2(_06475_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
AOI22_X1 _14490_ ( .A1(_04515_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02993_ ), .ZN(_06476_ ) );
OAI211_X1 _14491_ ( .A(_06476_ ), .B(_06299_ ), .C1(fanout_net_7 ), .C2(_02992_ ), .ZN(_06477_ ) );
NAND4_X1 _14492_ ( .A1(_04510_ ), .A2(_06334_ ), .A3(_04514_ ), .A4(_06271_ ), .ZN(_06478_ ) );
AND3_X1 _14493_ ( .A1(_05480_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_typ [7] ), .ZN(_06479_ ) );
AOI21_X1 _14494_ ( .A(_06479_ ), .B1(_03601_ ), .B2(_06380_ ), .ZN(_06480_ ) );
OAI211_X1 _14495_ ( .A(_06477_ ), .B(_06478_ ), .C1(_06272_ ), .C2(_06480_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
NAND3_X1 _14496_ ( .A1(_06365_ ), .A2(_06153_ ), .A3(_06366_ ), .ZN(_06481_ ) );
AND2_X1 _14497_ ( .A1(_04983_ ), .A2(_04984_ ), .ZN(_06482_ ) );
NAND3_X1 _14498_ ( .A1(_06482_ ), .A2(_04981_ ), .A3(_04982_ ), .ZN(_06483_ ) );
OAI21_X1 _14499_ ( .A(_06481_ ), .B1(_06483_ ), .B2(_05159_ ), .ZN(_06484_ ) );
AOI22_X1 _14500_ ( .A1(_06484_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02765_ ), .ZN(_06485_ ) );
OAI211_X1 _14501_ ( .A(_06485_ ), .B(_06299_ ), .C1(_02764_ ), .C2(fanout_net_7 ), .ZN(_06486_ ) );
AND3_X1 _14502_ ( .A1(_06482_ ), .A2(_04981_ ), .A3(_04982_ ), .ZN(_06487_ ) );
NAND2_X1 _14503_ ( .A1(_06487_ ), .A2(_05151_ ), .ZN(_06488_ ) );
NAND4_X1 _14504_ ( .A1(_06488_ ), .A2(_06334_ ), .A3(_06481_ ), .A4(_06271_ ), .ZN(_06489_ ) );
MUX2_X1 _14505_ ( .A(_04977_ ), .B(_04001_ ), .S(_06289_ ), .Z(_06490_ ) );
BUF_X4 _14506_ ( .A(_06291_ ), .Z(_06491_ ) );
OAI211_X1 _14507_ ( .A(_06486_ ), .B(_06489_ ), .C1(_06490_ ), .C2(_06491_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
NAND3_X1 _14508_ ( .A1(_02768_ ), .A2(_05027_ ), .A3(_02788_ ), .ZN(_06492_ ) );
NAND2_X1 _14509_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [0] ), .ZN(_06493_ ) );
NAND2_X1 _14510_ ( .A1(_06492_ ), .A2(_06493_ ), .ZN(_06494_ ) );
AOI21_X1 _14511_ ( .A(_06279_ ), .B1(_05023_ ), .B2(_05024_ ), .ZN(_06495_ ) );
AND2_X1 _14512_ ( .A1(_05023_ ), .A2(_05024_ ), .ZN(_06496_ ) );
INV_X1 _14513_ ( .A(_06496_ ), .ZN(_06497_ ) );
OAI221_X1 _14514_ ( .A(_06292_ ), .B1(_06494_ ), .B2(_06495_ ), .C1(_05195_ ), .C2(_06497_ ), .ZN(_06498_ ) );
NAND2_X1 _14515_ ( .A1(_04025_ ), .A2(_06380_ ), .ZN(_06499_ ) );
BUF_X4 _14516_ ( .A(_06258_ ), .Z(_06500_ ) );
OAI211_X1 _14517_ ( .A(_06499_ ), .B(_06500_ ), .C1(\ID_EX_pc [0] ), .C2(_06380_ ), .ZN(_06501_ ) );
NAND2_X1 _14518_ ( .A1(_06498_ ), .A2(_06501_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
OR2_X1 _14519_ ( .A1(_04795_ ), .A2(_05195_ ), .ZN(_06502_ ) );
NAND3_X1 _14520_ ( .A1(_02201_ ), .A2(_06303_ ), .A3(_02223_ ), .ZN(_06503_ ) );
OR2_X1 _14521_ ( .A1(_06303_ ), .A2(\ID_EX_imm [28] ), .ZN(_06504_ ) );
NAND4_X1 _14522_ ( .A1(_06502_ ), .A2(_06299_ ), .A3(_06503_ ), .A4(_06504_ ), .ZN(_06505_ ) );
NAND4_X1 _14523_ ( .A1(_04792_ ), .A2(_06334_ ), .A3(_04794_ ), .A4(_06291_ ), .ZN(_06506_ ) );
AND3_X1 _14524_ ( .A1(_05480_ ), .A2(\ID_EX_pc [28] ), .A3(\ID_EX_typ [7] ), .ZN(_06507_ ) );
AOI21_X1 _14525_ ( .A(_06507_ ), .B1(_03579_ ), .B2(_06380_ ), .ZN(_06508_ ) );
OAI211_X1 _14526_ ( .A(_06505_ ), .B(_06506_ ), .C1(_06491_ ), .C2(_06508_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
INV_X1 _14527_ ( .A(_05008_ ), .ZN(_06509_ ) );
AOI22_X1 _14528_ ( .A1(_06509_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02227_ ), .ZN(_06510_ ) );
OAI211_X1 _14529_ ( .A(_06510_ ), .B(_06299_ ), .C1(fanout_net_7 ), .C2(_03478_ ), .ZN(_06511_ ) );
NAND4_X1 _14530_ ( .A1(_05005_ ), .A2(_06334_ ), .A3(_05007_ ), .A4(_06291_ ), .ZN(_06512_ ) );
AND3_X1 _14531_ ( .A1(_05480_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_06513_ ) );
AOI21_X1 _14532_ ( .A(_06513_ ), .B1(_03501_ ), .B2(_06380_ ), .ZN(_06514_ ) );
OAI211_X1 _14533_ ( .A(_06511_ ), .B(_06512_ ), .C1(_06491_ ), .C2(_06514_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
INV_X1 _14534_ ( .A(\EX_LS_result_csreg_mem [26] ), .ZN(_06515_ ) );
NAND3_X1 _14535_ ( .A1(_06365_ ), .A2(_06515_ ), .A3(_06366_ ), .ZN(_06516_ ) );
AND2_X1 _14536_ ( .A1(_05039_ ), .A2(_05040_ ), .ZN(_06517_ ) );
NAND3_X1 _14537_ ( .A1(_06517_ ), .A2(_05037_ ), .A3(_05038_ ), .ZN(_06518_ ) );
OAI21_X1 _14538_ ( .A(_06516_ ), .B1(_06518_ ), .B2(_05159_ ), .ZN(_06519_ ) );
AOI22_X1 _14539_ ( .A1(_06519_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02272_ ), .ZN(_06520_ ) );
OAI211_X1 _14540_ ( .A(_06520_ ), .B(_06299_ ), .C1(_02271_ ), .C2(fanout_net_7 ), .ZN(_06521_ ) );
AND3_X1 _14541_ ( .A1(_06517_ ), .A2(_05037_ ), .A3(_05038_ ), .ZN(_06522_ ) );
NAND2_X1 _14542_ ( .A1(_06522_ ), .A2(_05151_ ), .ZN(_06523_ ) );
NAND4_X1 _14543_ ( .A1(_06523_ ), .A2(_06334_ ), .A3(_06516_ ), .A4(_06291_ ), .ZN(_06524_ ) );
MUX2_X1 _14544_ ( .A(_05031_ ), .B(_04372_ ), .S(_06289_ ), .Z(_06525_ ) );
OAI211_X1 _14545_ ( .A(_06521_ ), .B(_06524_ ), .C1(_06525_ ), .C2(_06491_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
AND2_X1 _14546_ ( .A1(_05060_ ), .A2(_05061_ ), .ZN(_06526_ ) );
AND2_X1 _14547_ ( .A1(_05062_ ), .A2(_05063_ ), .ZN(_06527_ ) );
NAND3_X1 _14548_ ( .A1(_05151_ ), .A2(_06526_ ), .A3(_06527_ ), .ZN(_06528_ ) );
OAI21_X1 _14549_ ( .A(_06528_ ), .B1(\EX_LS_result_csreg_mem [25] ), .B2(_05151_ ), .ZN(_06529_ ) );
AOI22_X1 _14550_ ( .A1(_06529_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02321_ ), .ZN(_06530_ ) );
OAI211_X1 _14551_ ( .A(_06530_ ), .B(_06299_ ), .C1(fanout_net_7 ), .C2(_02320_ ), .ZN(_06531_ ) );
OR2_X1 _14552_ ( .A1(_05151_ ), .A2(\EX_LS_result_csreg_mem [25] ), .ZN(_06532_ ) );
NAND4_X1 _14553_ ( .A1(_06532_ ), .A2(_06334_ ), .A3(_06528_ ), .A4(_06291_ ), .ZN(_06533_ ) );
AND3_X1 _14554_ ( .A1(_05480_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06534_ ) );
AOI21_X1 _14555_ ( .A(_06534_ ), .B1(_03555_ ), .B2(_06380_ ), .ZN(_06535_ ) );
OAI211_X1 _14556_ ( .A(_06531_ ), .B(_06533_ ), .C1(_06491_ ), .C2(_06535_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
INV_X1 _14557_ ( .A(_05079_ ), .ZN(_06536_ ) );
AND4_X1 _14558_ ( .A1(_05075_ ), .A2(_05076_ ), .A3(_06536_ ), .A4(_05077_ ), .ZN(_06537_ ) );
NAND4_X1 _14559_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04588_ ), .A4(_06537_ ), .ZN(_06538_ ) );
NAND3_X1 _14560_ ( .A1(_04429_ ), .A2(_05081_ ), .A3(_04439_ ), .ZN(_06539_ ) );
NAND3_X1 _14561_ ( .A1(_06538_ ), .A2(_06295_ ), .A3(_06539_ ), .ZN(_06540_ ) );
NAND2_X1 _14562_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [24] ), .ZN(_06541_ ) );
NAND2_X1 _14563_ ( .A1(_06540_ ), .A2(_06541_ ), .ZN(_06542_ ) );
AOI21_X1 _14564_ ( .A(fanout_net_7 ), .B1(_02275_ ), .B2(_02295_ ), .ZN(_06543_ ) );
OAI221_X1 _14565_ ( .A(_06292_ ), .B1(_05195_ ), .B2(_05083_ ), .C1(_06542_ ), .C2(_06543_ ), .ZN(_06544_ ) );
NAND4_X1 _14566_ ( .A1(_05049_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06545_ ) );
OAI211_X1 _14567_ ( .A(_06500_ ), .B(_06545_ ), .C1(_03532_ ), .C2(_06262_ ), .ZN(_06546_ ) );
NAND2_X1 _14568_ ( .A1(_06544_ ), .A2(_06546_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
INV_X1 _14569_ ( .A(\EX_LS_result_csreg_mem [23] ), .ZN(_06547_ ) );
NAND3_X1 _14570_ ( .A1(_06365_ ), .A2(_06547_ ), .A3(_06366_ ), .ZN(_06548_ ) );
AND2_X1 _14571_ ( .A1(_05101_ ), .A2(_05102_ ), .ZN(_06549_ ) );
NAND3_X1 _14572_ ( .A1(_06549_ ), .A2(_05099_ ), .A3(_05100_ ), .ZN(_06550_ ) );
OAI21_X1 _14573_ ( .A(_06548_ ), .B1(_06550_ ), .B2(_05159_ ), .ZN(_06551_ ) );
AOI22_X1 _14574_ ( .A1(_06551_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02407_ ), .ZN(_06552_ ) );
OAI211_X1 _14575_ ( .A(_06552_ ), .B(_06271_ ), .C1(_02406_ ), .C2(\ID_EX_typ [0] ), .ZN(_06553_ ) );
AND3_X1 _14576_ ( .A1(_06549_ ), .A2(_05099_ ), .A3(_05100_ ), .ZN(_06554_ ) );
NAND2_X1 _14577_ ( .A1(_06554_ ), .A2(_05151_ ), .ZN(_06555_ ) );
NAND4_X1 _14578_ ( .A1(_06555_ ), .A2(_06334_ ), .A3(_06548_ ), .A4(_06291_ ), .ZN(_06556_ ) );
MUX2_X1 _14579_ ( .A(_03187_ ), .B(_03381_ ), .S(_06289_ ), .Z(_06557_ ) );
OAI211_X1 _14580_ ( .A(_06553_ ), .B(_06556_ ), .C1(_06557_ ), .C2(_06292_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
INV_X1 _14581_ ( .A(_05125_ ), .ZN(_06558_ ) );
AOI22_X1 _14582_ ( .A1(_06558_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02430_ ), .ZN(_06559_ ) );
OAI211_X1 _14583_ ( .A(_06559_ ), .B(_06271_ ), .C1(\ID_EX_typ [0] ), .C2(_02429_ ), .ZN(_06560_ ) );
NAND4_X1 _14584_ ( .A1(_05122_ ), .A2(_06295_ ), .A3(_05124_ ), .A4(_06291_ ), .ZN(_06561_ ) );
MUX2_X1 _14585_ ( .A(_05111_ ), .B(_03403_ ), .S(_06263_ ), .Z(_06562_ ) );
OAI211_X1 _14586_ ( .A(_06560_ ), .B(_06561_ ), .C1(_06491_ ), .C2(_06562_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
INV_X1 _14587_ ( .A(_05161_ ), .ZN(_06563_ ) );
AOI22_X1 _14588_ ( .A1(_06563_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_04274_ ), .ZN(_06564_ ) );
OAI211_X1 _14589_ ( .A(_06564_ ), .B(_06271_ ), .C1(\ID_EX_typ [0] ), .C2(_03025_ ), .ZN(_06565_ ) );
INV_X1 _14590_ ( .A(_05152_ ), .ZN(_06566_ ) );
INV_X1 _14591_ ( .A(_05160_ ), .ZN(_06567_ ) );
NAND4_X1 _14592_ ( .A1(_06566_ ), .A2(_06295_ ), .A3(_06567_ ), .A4(_06291_ ), .ZN(_06568_ ) );
AND3_X1 _14593_ ( .A1(_05480_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06569_ ) );
AOI21_X1 _14594_ ( .A(_06569_ ), .B1(_03624_ ), .B2(_06380_ ), .ZN(_06570_ ) );
OAI211_X1 _14595_ ( .A(_06565_ ), .B(_06568_ ), .C1(_06491_ ), .C2(_06570_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
AND3_X1 _14596_ ( .A1(_04429_ ), .A2(_05138_ ), .A3(_04439_ ), .ZN(_06571_ ) );
INV_X1 _14597_ ( .A(_06571_ ), .ZN(_06572_ ) );
INV_X1 _14598_ ( .A(_04451_ ), .ZN(_06573_ ) );
AND4_X1 _14599_ ( .A1(_05131_ ), .A2(_05134_ ), .A3(_05132_ ), .A4(_05135_ ), .ZN(_06574_ ) );
INV_X1 _14600_ ( .A(_06574_ ), .ZN(_06575_ ) );
OAI211_X1 _14601_ ( .A(_06572_ ), .B(_06299_ ), .C1(_06573_ ), .C2(_06575_ ), .ZN(_06576_ ) );
NOR3_X1 _14602_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_06577_ ) );
AND2_X2 _14603_ ( .A1(\ID_EX_typ [3] ), .A2(\ID_EX_typ [2] ), .ZN(_06578_ ) );
AND2_X1 _14604_ ( .A1(_06577_ ), .A2(_06578_ ), .ZN(_06579_ ) );
BUF_X4 _14605_ ( .A(_06579_ ), .Z(_06580_ ) );
INV_X1 _14606_ ( .A(_06580_ ), .ZN(_06581_ ) );
NOR3_X1 _14607_ ( .A1(_04304_ ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_06582_ ) );
AND2_X2 _14608_ ( .A1(_06582_ ), .A2(_06578_ ), .ZN(_06583_ ) );
INV_X1 _14609_ ( .A(_06583_ ), .ZN(_06584_ ) );
OAI22_X1 _14610_ ( .A1(_05130_ ), .A2(_06581_ ), .B1(_02362_ ), .B2(_06584_ ), .ZN(_06585_ ) );
NAND2_X1 _14611_ ( .A1(_04346_ ), .A2(_03360_ ), .ZN(_06586_ ) );
AND2_X1 _14612_ ( .A1(_06586_ ), .A2(_04354_ ), .ZN(_06587_ ) );
INV_X1 _14613_ ( .A(_03427_ ), .ZN(_06588_ ) );
NOR2_X1 _14614_ ( .A1(_06587_ ), .A2(_06588_ ), .ZN(_06589_ ) );
AOI21_X1 _14615_ ( .A(_06589_ ), .B1(_02358_ ), .B2(_03426_ ), .ZN(_06590_ ) );
XNOR2_X1 _14616_ ( .A(_06590_ ), .B(_03451_ ), .ZN(_06591_ ) );
AND3_X1 _14617_ ( .A1(_03224_ ), .A2(\ID_EX_typ [3] ), .A3(_05194_ ), .ZN(_06592_ ) );
AND2_X1 _14618_ ( .A1(_06592_ ), .A2(_04049_ ), .ZN(_06593_ ) );
BUF_X4 _14619_ ( .A(_06593_ ), .Z(_06594_ ) );
BUF_X4 _14620_ ( .A(_06594_ ), .Z(_06595_ ) );
AOI21_X1 _14621_ ( .A(_06585_ ), .B1(_06591_ ), .B2(_06595_ ), .ZN(_06596_ ) );
NOR2_X1 _14622_ ( .A1(_02126_ ), .A2(\ID_EX_typ [6] ), .ZN(_06597_ ) );
AND2_X1 _14623_ ( .A1(_06597_ ), .A2(_05179_ ), .ZN(_06598_ ) );
INV_X1 _14624_ ( .A(_06598_ ), .ZN(_06599_ ) );
BUF_X4 _14625_ ( .A(_06599_ ), .Z(_06600_ ) );
BUF_X4 _14626_ ( .A(_06600_ ), .Z(_06601_ ) );
OAI21_X1 _14627_ ( .A(_04405_ ), .B1(_06596_ ), .B2(_06601_ ), .ZN(_06602_ ) );
NOR2_X1 _14628_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06603_ ) );
INV_X1 _14629_ ( .A(_06603_ ), .ZN(_06604_ ) );
NOR2_X2 _14630_ ( .A1(_04031_ ), .A2(_06604_ ), .ZN(_06605_ ) );
INV_X1 _14631_ ( .A(_06605_ ), .ZN(_06606_ ) );
BUF_X2 _14632_ ( .A(_06606_ ), .Z(_06607_ ) );
AND2_X1 _14633_ ( .A1(_04222_ ), .A2(_04226_ ), .ZN(_06608_ ) );
AND3_X1 _14634_ ( .A1(_06608_ ), .A2(_04233_ ), .A3(_04215_ ), .ZN(_06609_ ) );
INV_X1 _14635_ ( .A(_06609_ ), .ZN(_06610_ ) );
XNOR2_X1 _14636_ ( .A(_04106_ ), .B(_02670_ ), .ZN(_06611_ ) );
AND2_X1 _14637_ ( .A1(_06611_ ), .A2(_04102_ ), .ZN(_06612_ ) );
INV_X1 _14638_ ( .A(_06612_ ), .ZN(_06613_ ) );
AND2_X1 _14639_ ( .A1(_04126_ ), .A2(_04160_ ), .ZN(_06614_ ) );
AOI21_X1 _14640_ ( .A(_06614_ ), .B1(_02867_ ), .B2(_04125_ ), .ZN(_06615_ ) );
INV_X1 _14641_ ( .A(_04133_ ), .ZN(_06616_ ) );
NOR3_X1 _14642_ ( .A1(_06615_ ), .A2(_04118_ ), .A3(_06616_ ), .ZN(_06617_ ) );
NOR2_X1 _14643_ ( .A1(_04121_ ), .A2(_02918_ ), .ZN(_06618_ ) );
AOI211_X2 _14644_ ( .A(_04115_ ), .B(_06617_ ), .C1(_04117_ ), .C2(_06618_ ), .ZN(_06619_ ) );
BUF_X4 _14645_ ( .A(_04142_ ), .Z(_06620_ ) );
NOR2_X1 _14646_ ( .A1(_06620_ ), .A2(_02793_ ), .ZN(_06621_ ) );
INV_X1 _14647_ ( .A(_06621_ ), .ZN(_06622_ ) );
INV_X1 _14648_ ( .A(_04138_ ), .ZN(_06623_ ) );
NOR2_X1 _14649_ ( .A1(_04148_ ), .A2(_04149_ ), .ZN(_06624_ ) );
INV_X1 _14650_ ( .A(_04004_ ), .ZN(_06625_ ) );
NOR2_X1 _14651_ ( .A1(_04152_ ), .A2(_06625_ ), .ZN(_06626_ ) );
AND2_X1 _14652_ ( .A1(_06624_ ), .A2(_06626_ ), .ZN(_06627_ ) );
NOR2_X1 _14653_ ( .A1(_06627_ ), .A2(_04148_ ), .ZN(_06628_ ) );
INV_X1 _14654_ ( .A(_04143_ ), .ZN(_06629_ ) );
OAI221_X1 _14655_ ( .A(_06622_ ), .B1(_02819_ ), .B2(_06623_ ), .C1(_06628_ ), .C2(_06629_ ), .ZN(_06630_ ) );
BUF_X4 _14656_ ( .A(_04138_ ), .Z(_06631_ ) );
NOR2_X1 _14657_ ( .A1(_06631_ ), .A2(_02815_ ), .ZN(_06632_ ) );
INV_X1 _14658_ ( .A(_06632_ ), .ZN(_06633_ ) );
AND4_X1 _14659_ ( .A1(_04117_ ), .A2(_04126_ ), .A3(_04162_ ), .A4(_04133_ ), .ZN(_06634_ ) );
NAND3_X1 _14660_ ( .A1(_06630_ ), .A2(_06633_ ), .A3(_06634_ ), .ZN(_06635_ ) );
AOI21_X1 _14661_ ( .A(_06613_ ), .B1(_06619_ ), .B2(_06635_ ), .ZN(_06636_ ) );
AND2_X1 _14662_ ( .A1(_04074_ ), .A2(_04070_ ), .ZN(_06637_ ) );
AND2_X1 _14663_ ( .A1(_04091_ ), .A2(_04096_ ), .ZN(_06638_ ) );
AND2_X1 _14664_ ( .A1(_06637_ ), .A2(_06638_ ), .ZN(_06639_ ) );
AND2_X1 _14665_ ( .A1(_04079_ ), .A2(_04086_ ), .ZN(_06640_ ) );
NAND3_X1 _14666_ ( .A1(_06636_ ), .A2(_06639_ ), .A3(_06640_ ), .ZN(_06641_ ) );
NOR2_X1 _14667_ ( .A1(_04101_ ), .A2(_06412_ ), .ZN(_06642_ ) );
AOI21_X1 _14668_ ( .A(_04108_ ), .B1(_06611_ ), .B2(_06642_ ), .ZN(_06643_ ) );
INV_X1 _14669_ ( .A(_04079_ ), .ZN(_06644_ ) );
NOR3_X1 _14670_ ( .A1(_06643_ ), .A2(_06644_ ), .A3(_04174_ ), .ZN(_06645_ ) );
INV_X1 _14671_ ( .A(_02718_ ), .ZN(_06646_ ) );
NOR4_X1 _14672_ ( .A1(_04084_ ), .A2(_04085_ ), .A3(_06646_ ), .A4(_04078_ ), .ZN(_06647_ ) );
NOR3_X1 _14673_ ( .A1(_06645_ ), .A2(_04084_ ), .A3(_06647_ ), .ZN(_06648_ ) );
INV_X1 _14674_ ( .A(_06639_ ), .ZN(_06649_ ) );
NOR2_X1 _14675_ ( .A1(_06648_ ), .A2(_06649_ ), .ZN(_06650_ ) );
NOR2_X1 _14676_ ( .A1(_04073_ ), .A2(_04184_ ), .ZN(_06651_ ) );
NOR2_X1 _14677_ ( .A1(_04090_ ), .A2(_04179_ ), .ZN(_06652_ ) );
NAND2_X1 _14678_ ( .A1(_04096_ ), .A2(_06652_ ), .ZN(_06653_ ) );
OAI21_X1 _14679_ ( .A(_06653_ ), .B1(_06353_ ), .B2(_04095_ ), .ZN(_06654_ ) );
AND2_X1 _14680_ ( .A1(_06654_ ), .A2(_06637_ ), .ZN(_06655_ ) );
NOR2_X1 _14681_ ( .A1(_04069_ ), .A2(_04166_ ), .ZN(_06656_ ) );
INV_X1 _14682_ ( .A(_06656_ ), .ZN(_06657_ ) );
AND2_X1 _14683_ ( .A1(_04073_ ), .A2(_04184_ ), .ZN(_06658_ ) );
NOR3_X1 _14684_ ( .A1(_06657_ ), .A2(_06658_ ), .A3(_06651_ ), .ZN(_06659_ ) );
NOR4_X1 _14685_ ( .A1(_06650_ ), .A2(_06651_ ), .A3(_06655_ ), .A4(_06659_ ), .ZN(_06660_ ) );
AOI21_X1 _14686_ ( .A(_06610_ ), .B1(_06641_ ), .B2(_06660_ ), .ZN(_06661_ ) );
INV_X1 _14687_ ( .A(_06661_ ), .ZN(_06662_ ) );
AOI21_X1 _14688_ ( .A(_04241_ ), .B1(_04226_ ), .B2(_04220_ ), .ZN(_06663_ ) );
INV_X1 _14689_ ( .A(_04215_ ), .ZN(_06664_ ) );
NOR3_X1 _14690_ ( .A1(_06663_ ), .A2(_06664_ ), .A3(_04245_ ), .ZN(_06665_ ) );
INV_X1 _14691_ ( .A(_02501_ ), .ZN(_06666_ ) );
NOR4_X1 _14692_ ( .A1(_04231_ ), .A2(_04232_ ), .A3(_06666_ ), .A4(_04214_ ), .ZN(_06667_ ) );
NOR3_X1 _14693_ ( .A1(_06665_ ), .A2(_04231_ ), .A3(_06667_ ), .ZN(_06668_ ) );
AOI21_X1 _14694_ ( .A(_04204_ ), .B1(_06662_ ), .B2(_06668_ ), .ZN(_06669_ ) );
NOR2_X1 _14695_ ( .A1(_04202_ ), .A2(_04251_ ), .ZN(_06670_ ) );
OR2_X1 _14696_ ( .A1(_06669_ ), .A2(_06670_ ), .ZN(_06671_ ) );
AOI21_X1 _14697_ ( .A(_06607_ ), .B1(_06671_ ), .B2(_04209_ ), .ZN(_06672_ ) );
OAI21_X1 _14698_ ( .A(_06672_ ), .B1(_04209_ ), .B2(_06671_ ), .ZN(_06673_ ) );
AND2_X1 _14699_ ( .A1(_04307_ ), .A2(\ID_EX_typ [2] ), .ZN(_06674_ ) );
BUF_X4 _14700_ ( .A(_06674_ ), .Z(_06675_ ) );
BUF_X4 _14701_ ( .A(_06675_ ), .Z(_06676_ ) );
AND2_X1 _14702_ ( .A1(_04146_ ), .A2(_04152_ ), .ZN(_06677_ ) );
AND2_X1 _14703_ ( .A1(_06677_ ), .A2(_04142_ ), .ZN(_06678_ ) );
AND2_X1 _14704_ ( .A1(_06678_ ), .A2(_06623_ ), .ZN(_06679_ ) );
XNOR2_X1 _14705_ ( .A(_06679_ ), .B(_04130_ ), .ZN(_06680_ ) );
INV_X1 _14706_ ( .A(_06680_ ), .ZN(_06681_ ) );
AND2_X1 _14707_ ( .A1(_06679_ ), .A2(_04130_ ), .ZN(_06682_ ) );
INV_X1 _14708_ ( .A(_04125_ ), .ZN(_06683_ ) );
NOR4_X1 _14709_ ( .A1(_06682_ ), .A2(_04113_ ), .A3(_04121_ ), .A4(_06683_ ), .ZN(_06684_ ) );
AND4_X1 _14710_ ( .A1(_04113_ ), .A2(_04125_ ), .A3(_04130_ ), .A4(_04121_ ), .ZN(_06685_ ) );
NAND3_X1 _14711_ ( .A1(_06678_ ), .A2(_06623_ ), .A3(_06685_ ), .ZN(_06686_ ) );
NAND4_X1 _14712_ ( .A1(_04123_ ), .A2(_04113_ ), .A3(_04121_ ), .A4(_04124_ ), .ZN(_06687_ ) );
NAND2_X1 _14713_ ( .A1(_06686_ ), .A2(_06687_ ), .ZN(_06688_ ) );
NOR2_X1 _14714_ ( .A1(_06684_ ), .A2(_06688_ ), .ZN(_06689_ ) );
NOR2_X1 _14715_ ( .A1(_06689_ ), .A2(_04272_ ), .ZN(_06690_ ) );
AOI22_X1 _14716_ ( .A1(_04105_ ), .A2(_04104_ ), .B1(_04099_ ), .B2(_04100_ ), .ZN(_06691_ ) );
AND2_X1 _14717_ ( .A1(_04106_ ), .A2(_04101_ ), .ZN(_06692_ ) );
MUX2_X1 _14718_ ( .A(_06691_ ), .B(_06692_ ), .S(_06688_ ), .Z(_06693_ ) );
AND2_X1 _14719_ ( .A1(_06690_ ), .A2(_06693_ ), .ZN(_06694_ ) );
AND3_X1 _14720_ ( .A1(_06692_ ), .A2(_04082_ ), .A3(_04078_ ), .ZN(_06695_ ) );
NAND3_X1 _14721_ ( .A1(_06688_ ), .A2(_04073_ ), .A3(_06695_ ), .ZN(_06696_ ) );
NAND3_X1 _14722_ ( .A1(_04069_ ), .A2(_04090_ ), .A3(_04095_ ), .ZN(_06697_ ) );
NAND4_X1 _14723_ ( .A1(_04035_ ), .A2(_04052_ ), .A3(_04045_ ), .A4(_04276_ ), .ZN(_06698_ ) );
NAND4_X1 _14724_ ( .A1(_04214_ ), .A2(_04229_ ), .A3(_04225_ ), .A4(_04055_ ), .ZN(_06699_ ) );
NOR2_X1 _14725_ ( .A1(_06698_ ), .A2(_06699_ ), .ZN(_06700_ ) );
INV_X1 _14726_ ( .A(_04284_ ), .ZN(_06701_ ) );
INV_X1 _14727_ ( .A(_04270_ ), .ZN(_06702_ ) );
AND4_X1 _14728_ ( .A1(_04218_ ), .A2(_06701_ ), .A3(_04295_ ), .A4(_06702_ ), .ZN(_06703_ ) );
NOR2_X1 _14729_ ( .A1(_04252_ ), .A2(_04207_ ), .ZN(_06704_ ) );
AND2_X1 _14730_ ( .A1(_04194_ ), .A2(_04190_ ), .ZN(_06705_ ) );
AND4_X1 _14731_ ( .A1(_06700_ ), .A2(_06703_ ), .A3(_06704_ ), .A4(_06705_ ), .ZN(_06706_ ) );
OR3_X1 _14732_ ( .A1(_06696_ ), .A2(_06697_ ), .A3(_06706_ ), .ZN(_06707_ ) );
AND2_X1 _14733_ ( .A1(_06688_ ), .A2(_06695_ ), .ZN(_06708_ ) );
AOI211_X1 _14734_ ( .A(_04082_ ), .B(_04078_ ), .C1(_06688_ ), .C2(_06692_ ), .ZN(_06709_ ) );
OAI211_X1 _14735_ ( .A(_06694_ ), .B(_06707_ ), .C1(_06708_ ), .C2(_06709_ ), .ZN(_06710_ ) );
NOR4_X1 _14736_ ( .A1(_04073_ ), .A2(_04218_ ), .A3(_04090_ ), .A4(_04095_ ), .ZN(_06711_ ) );
AND4_X1 _14737_ ( .A1(_04256_ ), .A2(_04249_ ), .A3(_04252_ ), .A4(_04207_ ), .ZN(_06712_ ) );
AND4_X1 _14738_ ( .A1(_04167_ ), .A2(_04289_ ), .A3(_04270_ ), .A4(_04284_ ), .ZN(_06713_ ) );
AND3_X1 _14739_ ( .A1(_06711_ ), .A2(_06712_ ), .A3(_06713_ ), .ZN(_06714_ ) );
NOR4_X1 _14740_ ( .A1(_04229_ ), .A2(_04214_ ), .A3(_04225_ ), .A4(_04055_ ), .ZN(_06715_ ) );
NOR4_X1 _14741_ ( .A1(_04035_ ), .A2(_04052_ ), .A3(_04045_ ), .A4(_04276_ ), .ZN(_06716_ ) );
NAND3_X1 _14742_ ( .A1(_06714_ ), .A2(_06715_ ), .A3(_06716_ ), .ZN(_06717_ ) );
AOI21_X1 _14743_ ( .A(_06717_ ), .B1(_06688_ ), .B2(_06695_ ), .ZN(_06718_ ) );
AND4_X1 _14744_ ( .A1(_04072_ ), .A2(_04071_ ), .A3(_04067_ ), .A4(_04068_ ), .ZN(_06719_ ) );
AND4_X1 _14745_ ( .A1(_04090_ ), .A2(_06695_ ), .A3(_04095_ ), .A4(_06719_ ), .ZN(_06720_ ) );
AND2_X1 _14746_ ( .A1(_06688_ ), .A2(_06720_ ), .ZN(_06721_ ) );
NOR2_X1 _14747_ ( .A1(_06718_ ), .A2(_06721_ ), .ZN(_06722_ ) );
NOR2_X1 _14748_ ( .A1(_06710_ ), .A2(_06722_ ), .ZN(_06723_ ) );
BUF_X2 _14749_ ( .A(_06723_ ), .Z(_06724_ ) );
BUF_X2 _14750_ ( .A(_04146_ ), .Z(_06725_ ) );
BUF_X2 _14751_ ( .A(_06725_ ), .Z(_06726_ ) );
BUF_X2 _14752_ ( .A(_06726_ ), .Z(_06727_ ) );
BUF_X4 _14753_ ( .A(_04152_ ), .Z(_06728_ ) );
XNOR2_X1 _14754_ ( .A(_06727_ ), .B(_06728_ ), .ZN(_06729_ ) );
BUF_X4 _14755_ ( .A(_04156_ ), .Z(_06730_ ) );
BUF_X2 _14756_ ( .A(_06730_ ), .Z(_06731_ ) );
OR2_X1 _14757_ ( .A1(_06729_ ), .A2(_06731_ ), .ZN(_06732_ ) );
XNOR2_X1 _14758_ ( .A(_06678_ ), .B(_06631_ ), .ZN(_06733_ ) );
INV_X1 _14759_ ( .A(_06733_ ), .ZN(_06734_ ) );
BUF_X2 _14760_ ( .A(_06734_ ), .Z(_06735_ ) );
BUF_X2 _14761_ ( .A(_06735_ ), .Z(_06736_ ) );
NAND3_X1 _14762_ ( .A1(_06724_ ), .A2(_06732_ ), .A3(_06736_ ), .ZN(_06737_ ) );
NOR4_X1 _14763_ ( .A1(_04214_ ), .A2(_04218_ ), .A3(_04229_ ), .A4(_04225_ ), .ZN(_06738_ ) );
AND4_X1 _14764_ ( .A1(_04249_ ), .A2(_06738_ ), .A3(_04252_ ), .A4(_04207_ ), .ZN(_06739_ ) );
OAI211_X1 _14765_ ( .A(_04256_ ), .B(_06739_ ), .C1(_06696_ ), .C2(_06697_ ), .ZN(_06740_ ) );
AND4_X1 _14766_ ( .A1(_04228_ ), .A2(_04216_ ), .A3(_04227_ ), .A4(_04217_ ), .ZN(_06741_ ) );
AND4_X1 _14767_ ( .A1(_04214_ ), .A2(_06704_ ), .A3(_04225_ ), .A4(_06741_ ), .ZN(_06742_ ) );
AND3_X1 _14768_ ( .A1(_06688_ ), .A2(_06720_ ), .A3(_06742_ ), .ZN(_06743_ ) );
INV_X1 _14769_ ( .A(_06743_ ), .ZN(_06744_ ) );
NAND2_X1 _14770_ ( .A1(_06740_ ), .A2(_06744_ ), .ZN(_06745_ ) );
AND3_X1 _14771_ ( .A1(_06690_ ), .A2(_06693_ ), .A3(_06745_ ), .ZN(_06746_ ) );
NOR2_X1 _14772_ ( .A1(_06744_ ), .A2(_06705_ ), .ZN(_06747_ ) );
INV_X1 _14773_ ( .A(_04095_ ), .ZN(_06748_ ) );
NAND3_X1 _14774_ ( .A1(_04167_ ), .A2(_04185_ ), .A3(_06748_ ), .ZN(_06749_ ) );
OR3_X1 _14775_ ( .A1(_06708_ ), .A2(_04090_ ), .A3(_06749_ ), .ZN(_06750_ ) );
INV_X1 _14776_ ( .A(_06721_ ), .ZN(_06751_ ) );
AOI21_X1 _14777_ ( .A(_06747_ ), .B1(_06750_ ), .B2(_06751_ ), .ZN(_06752_ ) );
OAI211_X1 _14778_ ( .A(_06746_ ), .B(_06752_ ), .C1(_06708_ ), .C2(_06709_ ), .ZN(_06753_ ) );
AND4_X1 _14779_ ( .A1(_04055_ ), .A2(_06701_ ), .A3(_04295_ ), .A4(_04052_ ), .ZN(_06754_ ) );
AND4_X1 _14780_ ( .A1(_04045_ ), .A2(_04035_ ), .A3(_04276_ ), .A4(_06702_ ), .ZN(_06755_ ) );
AND4_X1 _14781_ ( .A1(_06705_ ), .A2(_06743_ ), .A3(_06754_ ), .A4(_06755_ ), .ZN(_06756_ ) );
NAND2_X1 _14782_ ( .A1(_06743_ ), .A2(_06705_ ), .ZN(_06757_ ) );
AND4_X1 _14783_ ( .A1(_04053_ ), .A2(_04287_ ), .A3(_04054_ ), .A4(_04288_ ), .ZN(_06758_ ) );
AND4_X1 _14784_ ( .A1(_04050_ ), .A2(_04282_ ), .A3(_04051_ ), .A4(_04283_ ), .ZN(_06759_ ) );
AND2_X1 _14785_ ( .A1(_06758_ ), .A2(_06759_ ), .ZN(_06760_ ) );
NAND4_X1 _14786_ ( .A1(_06760_ ), .A2(_04043_ ), .A3(_04044_ ), .A4(_04270_ ), .ZN(_06761_ ) );
NOR3_X1 _14787_ ( .A1(_06761_ ), .A2(_04035_ ), .A3(_04276_ ), .ZN(_06762_ ) );
AOI21_X1 _14788_ ( .A(_06756_ ), .B1(_06757_ ), .B2(_06762_ ), .ZN(_06763_ ) );
NOR2_X1 _14789_ ( .A1(_06753_ ), .A2(_06763_ ), .ZN(_06764_ ) );
XNOR2_X1 _14790_ ( .A(_06682_ ), .B(_04125_ ), .ZN(_06765_ ) );
NAND2_X1 _14791_ ( .A1(_06764_ ), .A2(_06765_ ), .ZN(_06766_ ) );
NOR2_X1 _14792_ ( .A1(_06680_ ), .A2(_04125_ ), .ZN(_06767_ ) );
INV_X1 _14793_ ( .A(_06767_ ), .ZN(_06768_ ) );
AOI22_X1 _14794_ ( .A1(_06681_ ), .A2(_06737_ ), .B1(_06766_ ), .B2(_06768_ ), .ZN(_06769_ ) );
BUF_X4 _14795_ ( .A(_04146_ ), .Z(_06770_ ) );
BUF_X4 _14796_ ( .A(_06770_ ), .Z(_06771_ ) );
CLKBUF_X2 _14797_ ( .A(_04150_ ), .Z(_06772_ ) );
BUF_X2 _14798_ ( .A(_04151_ ), .Z(_06773_ ) );
AND3_X1 _14799_ ( .A1(_06772_ ), .A2(_04248_ ), .A3(_06773_ ), .ZN(_06774_ ) );
BUF_X2 _14800_ ( .A(_04150_ ), .Z(_06775_ ) );
BUF_X2 _14801_ ( .A(_06775_ ), .Z(_06776_ ) );
BUF_X2 _14802_ ( .A(_04151_ ), .Z(_06777_ ) );
BUF_X2 _14803_ ( .A(_06777_ ), .Z(_06778_ ) );
AOI21_X1 _14804_ ( .A(_03448_ ), .B1(_06776_ ), .B2(_06778_ ), .ZN(_06779_ ) );
OAI21_X1 _14805_ ( .A(_06771_ ), .B1(_06774_ ), .B2(_06779_ ), .ZN(_06780_ ) );
INV_X1 _14806_ ( .A(_04146_ ), .ZN(_06781_ ) );
BUF_X4 _14807_ ( .A(_06781_ ), .Z(_06782_ ) );
AND3_X1 _14808_ ( .A1(_06772_ ), .A2(_04261_ ), .A3(_06773_ ), .ZN(_06783_ ) );
BUF_X2 _14809_ ( .A(_04150_ ), .Z(_06784_ ) );
BUF_X2 _14810_ ( .A(_06784_ ), .Z(_06785_ ) );
BUF_X2 _14811_ ( .A(_04151_ ), .Z(_06786_ ) );
BUF_X2 _14812_ ( .A(_06786_ ), .Z(_06787_ ) );
AOI21_X1 _14813_ ( .A(_02406_ ), .B1(_06785_ ), .B2(_06787_ ), .ZN(_06788_ ) );
OAI21_X1 _14814_ ( .A(_06782_ ), .B1(_06783_ ), .B2(_06788_ ), .ZN(_06789_ ) );
AOI21_X1 _14815_ ( .A(_06730_ ), .B1(_06780_ ), .B2(_06789_ ), .ZN(_06790_ ) );
BUF_X4 _14816_ ( .A(_06620_ ), .Z(_06791_ ) );
AND3_X1 _14817_ ( .A1(_06776_ ), .A2(_04036_ ), .A3(_06778_ ), .ZN(_06792_ ) );
AOI21_X1 _14818_ ( .A(_02320_ ), .B1(_06776_ ), .B2(_06778_ ), .ZN(_06793_ ) );
OAI21_X1 _14819_ ( .A(_06771_ ), .B1(_06792_ ), .B2(_06793_ ), .ZN(_06794_ ) );
BUF_X4 _14820_ ( .A(_06781_ ), .Z(_06795_ ) );
BUF_X2 _14821_ ( .A(_06795_ ), .Z(_06796_ ) );
AND3_X1 _14822_ ( .A1(_06772_ ), .A2(_04290_ ), .A3(_06773_ ), .ZN(_06797_ ) );
AOI21_X1 _14823_ ( .A(_03478_ ), .B1(_06776_ ), .B2(_06778_ ), .ZN(_06798_ ) );
OAI21_X1 _14824_ ( .A(_06796_ ), .B1(_06797_ ), .B2(_06798_ ), .ZN(_06799_ ) );
AOI21_X1 _14825_ ( .A(_06791_ ), .B1(_06794_ ), .B2(_06799_ ), .ZN(_06800_ ) );
NOR2_X1 _14826_ ( .A1(_06790_ ), .A2(_06800_ ), .ZN(_06801_ ) );
NAND2_X1 _14827_ ( .A1(_06728_ ), .A2(_02992_ ), .ZN(_06802_ ) );
INV_X1 _14828_ ( .A(_02199_ ), .ZN(_06803_ ) );
NAND3_X1 _14829_ ( .A1(_06803_ ), .A2(_06776_ ), .A3(_06778_ ), .ZN(_06804_ ) );
AOI21_X1 _14830_ ( .A(_06782_ ), .B1(_06802_ ), .B2(_06804_ ), .ZN(_06805_ ) );
BUF_X4 _14831_ ( .A(_06782_ ), .Z(_06806_ ) );
AND2_X1 _14832_ ( .A1(_04152_ ), .A2(_03025_ ), .ZN(_06807_ ) );
AOI21_X1 _14833_ ( .A(_06805_ ), .B1(_06806_ ), .B2(_06807_ ), .ZN(_06808_ ) );
BUF_X4 _14834_ ( .A(_06730_ ), .Z(_06809_ ) );
NOR2_X1 _14835_ ( .A1(_06808_ ), .A2(_06809_ ), .ZN(_06810_ ) );
MUX2_X1 _14836_ ( .A(_06801_ ), .B(_06810_ ), .S(_06631_ ), .Z(_06811_ ) );
BUF_X2 _14837_ ( .A(_04130_ ), .Z(_06812_ ) );
BUF_X2 _14838_ ( .A(_06812_ ), .Z(_06813_ ) );
BUF_X2 _14839_ ( .A(_06813_ ), .Z(_06814_ ) );
AND2_X1 _14840_ ( .A1(_06811_ ), .A2(_06814_ ), .ZN(_06815_ ) );
OAI21_X1 _14841_ ( .A(_06676_ ), .B1(_06769_ ), .B2(_06815_ ), .ZN(_06816_ ) );
BUF_X2 _14842_ ( .A(_04388_ ), .Z(_06817_ ) );
INV_X1 _14843_ ( .A(_06812_ ), .ZN(_06818_ ) );
BUF_X4 _14844_ ( .A(_06818_ ), .Z(_06819_ ) );
BUF_X4 _14845_ ( .A(_06819_ ), .Z(_06820_ ) );
BUF_X4 _14846_ ( .A(_06631_ ), .Z(_06821_ ) );
BUF_X4 _14847_ ( .A(_06821_ ), .Z(_06822_ ) );
AND3_X1 _14848_ ( .A1(_06784_ ), .A2(_06412_ ), .A3(_06786_ ), .ZN(_06823_ ) );
AOI21_X1 _14849_ ( .A(_02670_ ), .B1(_06772_ ), .B2(_06773_ ), .ZN(_06824_ ) );
NOR3_X1 _14850_ ( .A1(_06823_ ), .A2(_06796_ ), .A3(_06824_ ), .ZN(_06825_ ) );
BUF_X2 _14851_ ( .A(_04150_ ), .Z(_06826_ ) );
BUF_X2 _14852_ ( .A(_04151_ ), .Z(_06827_ ) );
AND3_X1 _14853_ ( .A1(_06826_ ), .A2(_02918_ ), .A3(_06827_ ), .ZN(_06828_ ) );
AOI21_X1 _14854_ ( .A(_02914_ ), .B1(_06784_ ), .B2(_06786_ ), .ZN(_06829_ ) );
NOR3_X1 _14855_ ( .A1(_06828_ ), .A2(_06829_ ), .A3(_06771_ ), .ZN(_06830_ ) );
NOR2_X1 _14856_ ( .A1(_06825_ ), .A2(_06830_ ), .ZN(_06831_ ) );
BUF_X4 _14857_ ( .A(_06620_ ), .Z(_06832_ ) );
BUF_X4 _14858_ ( .A(_06832_ ), .Z(_06833_ ) );
BUF_X4 _14859_ ( .A(_06833_ ), .Z(_06834_ ) );
NOR2_X1 _14860_ ( .A1(_06831_ ), .A2(_06834_ ), .ZN(_06835_ ) );
AND3_X1 _14861_ ( .A1(_06776_ ), .A2(_04179_ ), .A3(_06778_ ), .ZN(_06836_ ) );
INV_X1 _14862_ ( .A(_06836_ ), .ZN(_06837_ ) );
INV_X1 _14863_ ( .A(_04152_ ), .ZN(_06838_ ) );
OAI211_X1 _14864_ ( .A(_06837_ ), .B(_06727_ ), .C1(_02600_ ), .C2(_06838_ ), .ZN(_06839_ ) );
AOI21_X1 _14865_ ( .A(_02694_ ), .B1(_06772_ ), .B2(_06773_ ), .ZN(_06840_ ) );
INV_X1 _14866_ ( .A(_06840_ ), .ZN(_06841_ ) );
BUF_X4 _14867_ ( .A(_06782_ ), .Z(_06842_ ) );
OAI211_X1 _14868_ ( .A(_06841_ ), .B(_06842_ ), .C1(_02718_ ), .C2(_06728_ ), .ZN(_06843_ ) );
AOI21_X1 _14869_ ( .A(_06731_ ), .B1(_06839_ ), .B2(_06843_ ), .ZN(_06844_ ) );
OAI21_X1 _14870_ ( .A(_06822_ ), .B1(_06835_ ), .B2(_06844_ ), .ZN(_06845_ ) );
BUF_X4 _14871_ ( .A(_06623_ ), .Z(_06846_ ) );
BUF_X4 _14872_ ( .A(_06846_ ), .Z(_06847_ ) );
BUF_X2 _14873_ ( .A(_06847_ ), .Z(_06848_ ) );
AND3_X1 _14874_ ( .A1(_06776_ ), .A2(_04166_ ), .A3(_06778_ ), .ZN(_06849_ ) );
AOI21_X1 _14875_ ( .A(_02553_ ), .B1(_06785_ ), .B2(_06787_ ), .ZN(_06850_ ) );
OR3_X1 _14876_ ( .A1(_06849_ ), .A2(_06850_ ), .A3(_06726_ ), .ZN(_06851_ ) );
AOI21_X1 _14877_ ( .A(_02476_ ), .B1(_06785_ ), .B2(_06787_ ), .ZN(_06852_ ) );
INV_X1 _14878_ ( .A(_06852_ ), .ZN(_06853_ ) );
BUF_X4 _14879_ ( .A(_06770_ ), .Z(_06854_ ) );
OAI211_X1 _14880_ ( .A(_06853_ ), .B(_06854_ ), .C1(_02453_ ), .C2(_06728_ ), .ZN(_06855_ ) );
AOI21_X1 _14881_ ( .A(_06834_ ), .B1(_06851_ ), .B2(_06855_ ), .ZN(_06856_ ) );
AND3_X1 _14882_ ( .A1(_06772_ ), .A2(_04251_ ), .A3(_06773_ ), .ZN(_06857_ ) );
OAI21_X1 _14883_ ( .A(_06727_ ), .B1(_06857_ ), .B2(_06779_ ), .ZN(_06858_ ) );
AND3_X1 _14884_ ( .A1(_06785_ ), .A2(_06666_ ), .A3(_06787_ ), .ZN(_06859_ ) );
AOI21_X1 _14885_ ( .A(_02524_ ), .B1(_06776_ ), .B2(_06778_ ), .ZN(_06860_ ) );
OAI21_X1 _14886_ ( .A(_06842_ ), .B1(_06859_ ), .B2(_06860_ ), .ZN(_06861_ ) );
BUF_X2 _14887_ ( .A(_06832_ ), .Z(_06862_ ) );
AND3_X1 _14888_ ( .A1(_06858_ ), .A2(_06861_ ), .A3(_06862_ ), .ZN(_06863_ ) );
OAI21_X1 _14889_ ( .A(_06848_ ), .B1(_06856_ ), .B2(_06863_ ), .ZN(_06864_ ) );
AOI21_X1 _14890_ ( .A(_06820_ ), .B1(_06845_ ), .B2(_06864_ ), .ZN(_06865_ ) );
BUF_X2 _14891_ ( .A(_06818_ ), .Z(_06866_ ) );
AND3_X1 _14892_ ( .A1(_06625_ ), .A2(_06785_ ), .A3(_06787_ ), .ZN(_06867_ ) );
AOI21_X1 _14893_ ( .A(_02764_ ), .B1(_06776_ ), .B2(_06778_ ), .ZN(_06868_ ) );
NOR3_X1 _14894_ ( .A1(_06867_ ), .A2(_06842_ ), .A3(_06868_ ), .ZN(_06869_ ) );
OR2_X1 _14895_ ( .A1(_06869_ ), .A2(_06862_ ), .ZN(_06870_ ) );
AND3_X1 _14896_ ( .A1(_06826_ ), .A2(_04159_ ), .A3(_06827_ ), .ZN(_06871_ ) );
AOI21_X1 _14897_ ( .A(_02867_ ), .B1(_06826_ ), .B2(_06827_ ), .ZN(_06872_ ) );
OAI21_X1 _14898_ ( .A(_06854_ ), .B1(_06871_ ), .B2(_06872_ ), .ZN(_06873_ ) );
AND3_X1 _14899_ ( .A1(_06776_ ), .A2(_02793_ ), .A3(_06778_ ), .ZN(_06874_ ) );
AOI21_X1 _14900_ ( .A(_02815_ ), .B1(_06785_ ), .B2(_06787_ ), .ZN(_06875_ ) );
OAI21_X1 _14901_ ( .A(_06806_ ), .B1(_06874_ ), .B2(_06875_ ), .ZN(_06876_ ) );
NAND2_X1 _14902_ ( .A1(_06873_ ), .A2(_06876_ ), .ZN(_06877_ ) );
BUF_X4 _14903_ ( .A(_06791_ ), .Z(_06878_ ) );
NAND2_X1 _14904_ ( .A1(_06877_ ), .A2(_06878_ ), .ZN(_06879_ ) );
AND4_X1 _14905_ ( .A1(_06866_ ), .A2(_06870_ ), .A3(_06848_ ), .A4(_06879_ ), .ZN(_06880_ ) );
OAI21_X1 _14906_ ( .A(_06817_ ), .B1(_06865_ ), .B2(_06880_ ), .ZN(_06881_ ) );
OAI21_X1 _14907_ ( .A(_04394_ ), .B1(_04207_ ), .B2(_03448_ ), .ZN(_06882_ ) );
AND2_X1 _14908_ ( .A1(_04392_ ), .A2(\ID_EX_typ [2] ), .ZN(_06883_ ) );
BUF_X2 _14909_ ( .A(_06883_ ), .Z(_06884_ ) );
BUF_X2 _14910_ ( .A(_06884_ ), .Z(_06885_ ) );
NAND3_X1 _14911_ ( .A1(_06811_ ), .A2(_06814_ ), .A3(_06885_ ), .ZN(_06886_ ) );
BUF_X2 _14912_ ( .A(_04308_ ), .Z(_06887_ ) );
AND2_X1 _14913_ ( .A1(_04207_ ), .A2(_03448_ ), .ZN(_06888_ ) );
BUF_X2 _14914_ ( .A(_04031_ ), .Z(_06889_ ) );
BUF_X2 _14915_ ( .A(_06889_ ), .Z(_06890_ ) );
AOI22_X1 _14916_ ( .A1(_04209_ ), .A2(_06887_ ), .B1(_06888_ ), .B2(_06890_ ), .ZN(_06891_ ) );
AND4_X1 _14917_ ( .A1(_06881_ ), .A2(_06882_ ), .A3(_06886_ ), .A4(_06891_ ), .ZN(_06892_ ) );
NAND3_X1 _14918_ ( .A1(_06673_ ), .A2(_06816_ ), .A3(_06892_ ), .ZN(_06893_ ) );
OAI211_X1 _14919_ ( .A(_02123_ ), .B(_06578_ ), .C1(_04392_ ), .C2(_03224_ ), .ZN(_06894_ ) );
NOR2_X1 _14920_ ( .A1(_04407_ ), .A2(\ID_EX_typ [2] ), .ZN(_06895_ ) );
OAI211_X1 _14921_ ( .A(_06895_ ), .B(_04304_ ), .C1(_04049_ ), .C2(_04482_ ), .ZN(_06896_ ) );
AND2_X1 _14922_ ( .A1(_06894_ ), .A2(_06896_ ), .ZN(_06897_ ) );
NOR2_X1 _14923_ ( .A1(_06897_ ), .A2(_06599_ ), .ZN(_06898_ ) );
INV_X2 _14924_ ( .A(_06898_ ), .ZN(_06899_ ) );
BUF_X4 _14925_ ( .A(_06899_ ), .Z(_06900_ ) );
AOI21_X1 _14926_ ( .A(_06602_ ), .B1(_06893_ ), .B2(_06900_ ), .ZN(_06901_ ) );
NAND2_X1 _14927_ ( .A1(_05148_ ), .A2(_05029_ ), .ZN(_06902_ ) );
NAND2_X1 _14928_ ( .A1(_06902_ ), .A2(_06259_ ), .ZN(_06903_ ) );
OAI21_X1 _14929_ ( .A(_06576_ ), .B1(_06901_ ), .B2(_06903_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
INV_X1 _14930_ ( .A(_04558_ ), .ZN(_06904_ ) );
AND4_X1 _14931_ ( .A1(_04550_ ), .A2(_04553_ ), .A3(_04555_ ), .A4(_06904_ ), .ZN(_06905_ ) );
NAND4_X1 _14932_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04588_ ), .A4(_06905_ ), .ZN(_06906_ ) );
BUF_X2 _14933_ ( .A(_04591_ ), .Z(_06907_ ) );
BUF_X2 _14934_ ( .A(_04592_ ), .Z(_06908_ ) );
NAND3_X1 _14935_ ( .A1(_06907_ ), .A2(_04561_ ), .A3(_06908_ ), .ZN(_06909_ ) );
BUF_X4 _14936_ ( .A(_06256_ ), .Z(_06910_ ) );
NAND3_X1 _14937_ ( .A1(_06906_ ), .A2(_06909_ ), .A3(_06910_ ), .ZN(_06911_ ) );
OR2_X1 _14938_ ( .A1(_06587_ ), .A2(_06588_ ), .ZN(_06912_ ) );
NAND3_X1 _14939_ ( .A1(_06586_ ), .A2(_06588_ ), .A3(_04354_ ), .ZN(_06913_ ) );
NAND3_X1 _14940_ ( .A1(_06912_ ), .A2(_06595_ ), .A3(_06913_ ), .ZN(_06914_ ) );
BUF_X2 _14941_ ( .A(_06580_ ), .Z(_06915_ ) );
BUF_X4 _14942_ ( .A(_06583_ ), .Z(_06916_ ) );
AOI22_X1 _14943_ ( .A1(_04545_ ), .A2(_06915_ ), .B1(\ID_EX_imm [20] ), .B2(_06916_ ), .ZN(_06917_ ) );
AOI21_X1 _14944_ ( .A(_06601_ ), .B1(_06914_ ), .B2(_06917_ ), .ZN(_06918_ ) );
CLKBUF_X2 _14945_ ( .A(_04487_ ), .Z(_06919_ ) );
OR2_X1 _14946_ ( .A1(_06918_ ), .A2(_06919_ ), .ZN(_06920_ ) );
AND2_X1 _14947_ ( .A1(_06662_ ), .A2(_06668_ ), .ZN(_06921_ ) );
OAI21_X1 _14948_ ( .A(_06605_ ), .B1(_06921_ ), .B2(_04204_ ), .ZN(_06922_ ) );
AOI21_X1 _14949_ ( .A(_06922_ ), .B1(_04204_ ), .B2(_06921_ ), .ZN(_06923_ ) );
INV_X1 _14950_ ( .A(_06674_ ), .ZN(_06924_ ) );
BUF_X4 _14951_ ( .A(_06924_ ), .Z(_06925_ ) );
BUF_X4 _14952_ ( .A(_06806_ ), .Z(_06926_ ) );
OAI21_X1 _14953_ ( .A(_06833_ ), .B1(_06926_ ), .B2(_06838_ ), .ZN(_06927_ ) );
AND3_X1 _14954_ ( .A1(_06723_ ), .A2(_06735_ ), .A3(_06927_ ), .ZN(_06928_ ) );
AND2_X1 _14955_ ( .A1(_06723_ ), .A2(_06765_ ), .ZN(_06929_ ) );
OAI22_X1 _14956_ ( .A1(_06928_ ), .A2(_06680_ ), .B1(_06929_ ), .B2(_06767_ ), .ZN(_06930_ ) );
AND3_X1 _14957_ ( .A1(_06784_ ), .A2(_02998_ ), .A3(_06786_ ), .ZN(_06931_ ) );
AOI21_X1 _14958_ ( .A(_02224_ ), .B1(_06772_ ), .B2(_06773_ ), .ZN(_06932_ ) );
OAI21_X1 _14959_ ( .A(_06725_ ), .B1(_06931_ ), .B2(_06932_ ), .ZN(_06933_ ) );
AOI21_X1 _14960_ ( .A(_06803_ ), .B1(_06784_ ), .B2(_06786_ ), .ZN(_06934_ ) );
AOI21_X1 _14961_ ( .A(_06934_ ), .B1(_04272_ ), .B2(_06838_ ), .ZN(_06935_ ) );
OAI21_X1 _14962_ ( .A(_06933_ ), .B1(_06935_ ), .B2(_06770_ ), .ZN(_06936_ ) );
BUF_X2 _14963_ ( .A(_06846_ ), .Z(_06937_ ) );
OR3_X1 _14964_ ( .A1(_06936_ ), .A2(_06937_ ), .A3(_06809_ ), .ZN(_06938_ ) );
BUF_X2 _14965_ ( .A(_04156_ ), .Z(_06939_ ) );
AND3_X1 _14966_ ( .A1(_06775_ ), .A2(_04208_ ), .A3(_06777_ ), .ZN(_06940_ ) );
AOI21_X1 _14967_ ( .A(_02358_ ), .B1(_06775_ ), .B2(_06777_ ), .ZN(_06941_ ) );
OR3_X1 _14968_ ( .A1(_06940_ ), .A2(_06781_ ), .A3(_06941_ ), .ZN(_06942_ ) );
AND3_X1 _14969_ ( .A1(_04150_ ), .A2(_04195_ ), .A3(_04151_ ), .ZN(_06943_ ) );
AOI21_X1 _14970_ ( .A(_02429_ ), .B1(_06775_ ), .B2(_06777_ ), .ZN(_06944_ ) );
OR3_X1 _14971_ ( .A1(_06943_ ), .A2(_06944_ ), .A3(_04146_ ), .ZN(_06945_ ) );
AOI21_X1 _14972_ ( .A(_06939_ ), .B1(_06942_ ), .B2(_06945_ ), .ZN(_06946_ ) );
AND3_X1 _14973_ ( .A1(_06784_ ), .A2(_04056_ ), .A3(_06786_ ), .ZN(_06947_ ) );
AOI21_X1 _14974_ ( .A(_02296_ ), .B1(_06784_ ), .B2(_06786_ ), .ZN(_06948_ ) );
OAI21_X1 _14975_ ( .A(_06770_ ), .B1(_06947_ ), .B2(_06948_ ), .ZN(_06949_ ) );
AND3_X1 _14976_ ( .A1(_06784_ ), .A2(_04064_ ), .A3(_06786_ ), .ZN(_06950_ ) );
AOI21_X1 _14977_ ( .A(_02271_ ), .B1(_06784_ ), .B2(_06773_ ), .ZN(_06951_ ) );
OAI21_X1 _14978_ ( .A(_06795_ ), .B1(_06950_ ), .B2(_06951_ ), .ZN(_06952_ ) );
AND3_X1 _14979_ ( .A1(_06949_ ), .A2(_06952_ ), .A3(_06730_ ), .ZN(_06953_ ) );
OAI21_X1 _14980_ ( .A(_06847_ ), .B1(_06946_ ), .B2(_06953_ ), .ZN(_06954_ ) );
NAND2_X1 _14981_ ( .A1(_06938_ ), .A2(_06954_ ), .ZN(_06955_ ) );
NAND2_X1 _14982_ ( .A1(_06955_ ), .A2(_06814_ ), .ZN(_06956_ ) );
AOI21_X1 _14983_ ( .A(_06925_ ), .B1(_06930_ ), .B2(_06956_ ), .ZN(_06957_ ) );
AND3_X1 _14984_ ( .A1(_06955_ ), .A2(_06813_ ), .A3(_06884_ ), .ZN(_06958_ ) );
AOI21_X1 _14985_ ( .A(_06958_ ), .B1(_06670_ ), .B2(_06890_ ), .ZN(_06959_ ) );
AND3_X1 _14986_ ( .A1(_06775_ ), .A2(_04184_ ), .A3(_06777_ ), .ZN(_06960_ ) );
AOI21_X1 _14987_ ( .A(_02453_ ), .B1(_06784_ ), .B2(_06786_ ), .ZN(_06961_ ) );
OR3_X1 _14988_ ( .A1(_06960_ ), .A2(_06782_ ), .A3(_06961_ ), .ZN(_06962_ ) );
AND3_X1 _14989_ ( .A1(_04150_ ), .A2(_06353_ ), .A3(_04151_ ), .ZN(_06963_ ) );
AOI21_X1 _14990_ ( .A(_02575_ ), .B1(_06775_ ), .B2(_06777_ ), .ZN(_06964_ ) );
OR3_X1 _14991_ ( .A1(_06963_ ), .A2(_06964_ ), .A3(_06770_ ), .ZN(_06965_ ) );
AOI21_X1 _14992_ ( .A(_06834_ ), .B1(_06962_ ), .B2(_06965_ ), .ZN(_06966_ ) );
BUF_X4 _14993_ ( .A(_06854_ ), .Z(_06967_ ) );
AND3_X1 _14994_ ( .A1(_06775_ ), .A2(_04230_ ), .A3(_06777_ ), .ZN(_06968_ ) );
OAI21_X1 _14995_ ( .A(_06967_ ), .B1(_06968_ ), .B2(_06941_ ), .ZN(_06969_ ) );
AND3_X1 _14996_ ( .A1(_06826_ ), .A2(_02946_ ), .A3(_06827_ ), .ZN(_06970_ ) );
AOI21_X1 _14997_ ( .A(_02501_ ), .B1(_06826_ ), .B2(_06827_ ), .ZN(_06971_ ) );
OAI21_X1 _14998_ ( .A(_06926_ ), .B1(_06970_ ), .B2(_06971_ ), .ZN(_06972_ ) );
AND3_X1 _14999_ ( .A1(_06969_ ), .A2(_06972_ ), .A3(_06878_ ), .ZN(_06973_ ) );
OAI21_X1 _15000_ ( .A(_06848_ ), .B1(_06966_ ), .B2(_06973_ ), .ZN(_06974_ ) );
AND3_X1 _15001_ ( .A1(_02923_ ), .A2(_06826_ ), .A3(_06827_ ), .ZN(_06975_ ) );
AOI21_X1 _15002_ ( .A(_02890_ ), .B1(_06826_ ), .B2(_06827_ ), .ZN(_06976_ ) );
OAI21_X1 _15003_ ( .A(_06806_ ), .B1(_06975_ ), .B2(_06976_ ), .ZN(_06977_ ) );
AND3_X1 _15004_ ( .A1(_06826_ ), .A2(_04114_ ), .A3(_06827_ ), .ZN(_06978_ ) );
AOI21_X1 _15005_ ( .A(_02647_ ), .B1(_06826_ ), .B2(_06827_ ), .ZN(_06979_ ) );
OAI21_X1 _15006_ ( .A(_06854_ ), .B1(_06978_ ), .B2(_06979_ ), .ZN(_06980_ ) );
NAND2_X1 _15007_ ( .A1(_06977_ ), .A2(_06980_ ), .ZN(_06981_ ) );
BUF_X4 _15008_ ( .A(_06809_ ), .Z(_06982_ ) );
NAND2_X1 _15009_ ( .A1(_06981_ ), .A2(_06982_ ), .ZN(_06983_ ) );
AND3_X1 _15010_ ( .A1(_04150_ ), .A2(_04083_ ), .A3(_04151_ ), .ZN(_06984_ ) );
AOI21_X1 _15011_ ( .A(_02622_ ), .B1(_06775_ ), .B2(_06777_ ), .ZN(_06985_ ) );
OR3_X1 _15012_ ( .A1(_06984_ ), .A2(_06782_ ), .A3(_06985_ ), .ZN(_06986_ ) );
AND3_X1 _15013_ ( .A1(_06775_ ), .A2(_04107_ ), .A3(_06777_ ), .ZN(_06987_ ) );
AOI21_X1 _15014_ ( .A(_02718_ ), .B1(_06775_ ), .B2(_06777_ ), .ZN(_06988_ ) );
OR3_X1 _15015_ ( .A1(_06987_ ), .A2(_06988_ ), .A3(_06770_ ), .ZN(_06989_ ) );
NAND3_X1 _15016_ ( .A1(_06986_ ), .A2(_06989_ ), .A3(_06878_ ), .ZN(_06990_ ) );
BUF_X2 _15017_ ( .A(_06631_ ), .Z(_06991_ ) );
NAND3_X1 _15018_ ( .A1(_06983_ ), .A2(_06990_ ), .A3(_06991_ ), .ZN(_06992_ ) );
AOI21_X1 _15019_ ( .A(_06866_ ), .B1(_06974_ ), .B2(_06992_ ), .ZN(_06993_ ) );
AOI21_X1 _15020_ ( .A(_06625_ ), .B1(_06785_ ), .B2(_06787_ ), .ZN(_06994_ ) );
AND2_X1 _15021_ ( .A1(_06994_ ), .A2(_06727_ ), .ZN(_06995_ ) );
INV_X1 _15022_ ( .A(_06995_ ), .ZN(_06996_ ) );
NOR2_X1 _15023_ ( .A1(_06728_ ), .A2(_02764_ ), .ZN(_06997_ ) );
AOI21_X1 _15024_ ( .A(_02741_ ), .B1(_06772_ ), .B2(_06773_ ), .ZN(_06998_ ) );
OAI21_X1 _15025_ ( .A(_06842_ ), .B1(_06997_ ), .B2(_06998_ ), .ZN(_06999_ ) );
AND3_X1 _15026_ ( .A1(_06772_ ), .A2(_02819_ ), .A3(_06773_ ), .ZN(_07000_ ) );
AOI21_X1 _15027_ ( .A(_02842_ ), .B1(_06826_ ), .B2(_06827_ ), .ZN(_07001_ ) );
OAI21_X1 _15028_ ( .A(_06854_ ), .B1(_07000_ ), .B2(_07001_ ), .ZN(_07002_ ) );
NAND2_X1 _15029_ ( .A1(_06999_ ), .A2(_07002_ ), .ZN(_07003_ ) );
MUX2_X1 _15030_ ( .A(_06996_ ), .B(_07003_ ), .S(_06878_ ), .Z(_07004_ ) );
BUF_X2 _15031_ ( .A(_06812_ ), .Z(_07005_ ) );
BUF_X2 _15032_ ( .A(_07005_ ), .Z(_07006_ ) );
NOR3_X1 _15033_ ( .A1(_07004_ ), .A2(_07006_ ), .A3(_06822_ ), .ZN(_07007_ ) );
OAI21_X1 _15034_ ( .A(_06817_ ), .B1(_06993_ ), .B2(_07007_ ), .ZN(_07008_ ) );
BUF_X4 _15035_ ( .A(_04395_ ), .Z(_07009_ ) );
AOI21_X1 _15036_ ( .A(_07009_ ), .B1(_04202_ ), .B2(_04251_ ), .ZN(_07010_ ) );
AOI21_X1 _15037_ ( .A(_07010_ ), .B1(_04203_ ), .B2(_06887_ ), .ZN(_07011_ ) );
NAND3_X1 _15038_ ( .A1(_06959_ ), .A2(_07008_ ), .A3(_07011_ ), .ZN(_07012_ ) );
OR3_X1 _15039_ ( .A1(_06923_ ), .A2(_06957_ ), .A3(_07012_ ), .ZN(_07013_ ) );
AOI21_X1 _15040_ ( .A(_06920_ ), .B1(_07013_ ), .B2(_06900_ ), .ZN(_07014_ ) );
OAI21_X1 _15041_ ( .A(_06500_ ), .B1(_04540_ ), .B2(_05097_ ), .ZN(_07015_ ) );
OAI21_X1 _15042_ ( .A(_06911_ ), .B1(_07014_ ), .B2(_07015_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OR2_X1 _15043_ ( .A1(_04594_ ), .A2(_06258_ ), .ZN(_07016_ ) );
BUF_X4 _15044_ ( .A(_06600_ ), .Z(_07017_ ) );
INV_X1 _15045_ ( .A(_03334_ ), .ZN(_07018_ ) );
INV_X1 _15046_ ( .A(_03359_ ), .ZN(_07019_ ) );
AOI211_X1 _15047_ ( .A(_07018_ ), .B(_07019_ ), .C1(_04326_ ), .C2(_04344_ ), .ZN(_07020_ ) );
OAI21_X1 _15048_ ( .A(_03310_ ), .B1(_07020_ ), .B2(_04350_ ), .ZN(_07021_ ) );
NAND2_X1 _15049_ ( .A1(_03309_ ), .A2(_02501_ ), .ZN(_07022_ ) );
AND2_X1 _15050_ ( .A1(_07021_ ), .A2(_07022_ ), .ZN(_07023_ ) );
XNOR2_X1 _15051_ ( .A(_07023_ ), .B(_03281_ ), .ZN(_07024_ ) );
NAND2_X1 _15052_ ( .A1(_07024_ ), .A2(_06595_ ), .ZN(_07025_ ) );
AOI22_X1 _15053_ ( .A1(_04573_ ), .A2(_06915_ ), .B1(\ID_EX_imm [19] ), .B2(_06916_ ), .ZN(_07026_ ) );
AOI21_X1 _15054_ ( .A(_07017_ ), .B1(_07025_ ), .B2(_07026_ ), .ZN(_07027_ ) );
OR2_X1 _15055_ ( .A1(_07027_ ), .A2(_06919_ ), .ZN(_07028_ ) );
AND2_X1 _15056_ ( .A1(_06641_ ), .A2(_06660_ ), .ZN(_07029_ ) );
INV_X1 _15057_ ( .A(_04226_ ), .ZN(_07030_ ) );
OR4_X1 _15058_ ( .A1(_04221_ ), .A2(_07029_ ), .A3(_04220_ ), .A4(_07030_ ), .ZN(_07031_ ) );
AOI21_X1 _15059_ ( .A(_06664_ ), .B1(_07031_ ), .B2(_06663_ ), .ZN(_07032_ ) );
NOR2_X1 _15060_ ( .A1(_04214_ ), .A2(_06666_ ), .ZN(_07033_ ) );
OR3_X1 _15061_ ( .A1(_07032_ ), .A2(_04233_ ), .A3(_07033_ ), .ZN(_07034_ ) );
BUF_X4 _15062_ ( .A(_06605_ ), .Z(_07035_ ) );
OAI21_X1 _15063_ ( .A(_04233_ ), .B1(_07032_ ), .B2(_07033_ ), .ZN(_07036_ ) );
NAND3_X1 _15064_ ( .A1(_07034_ ), .A2(_07035_ ), .A3(_07036_ ), .ZN(_07037_ ) );
AND2_X2 _15065_ ( .A1(_06765_ ), .A2(_06680_ ), .ZN(_07038_ ) );
AND2_X1 _15066_ ( .A1(_06764_ ), .A2(_07038_ ), .ZN(_07039_ ) );
NOR3_X1 _15067_ ( .A1(_06783_ ), .A2(_06782_ ), .A3(_06788_ ), .ZN(_07040_ ) );
NOR3_X1 _15068_ ( .A1(_06792_ ), .A2(_06793_ ), .A3(_06726_ ), .ZN(_07041_ ) );
NOR2_X1 _15069_ ( .A1(_07040_ ), .A2(_07041_ ), .ZN(_07042_ ) );
NOR2_X1 _15070_ ( .A1(_07042_ ), .A2(_06791_ ), .ZN(_07043_ ) );
OR3_X1 _15071_ ( .A1(_06857_ ), .A2(_06782_ ), .A3(_06860_ ), .ZN(_07044_ ) );
OR3_X1 _15072_ ( .A1(_06774_ ), .A2(_06779_ ), .A3(_06770_ ), .ZN(_07045_ ) );
AOI21_X1 _15073_ ( .A(_06730_ ), .B1(_07044_ ), .B2(_07045_ ), .ZN(_07046_ ) );
OAI21_X1 _15074_ ( .A(_06937_ ), .B1(_07043_ ), .B2(_07046_ ), .ZN(_07047_ ) );
AND2_X1 _15075_ ( .A1(_06807_ ), .A2(_06725_ ), .ZN(_07048_ ) );
INV_X1 _15076_ ( .A(_07048_ ), .ZN(_07049_ ) );
NOR3_X1 _15077_ ( .A1(_06797_ ), .A2(_06795_ ), .A3(_06798_ ), .ZN(_07050_ ) );
AOI21_X1 _15078_ ( .A(_06770_ ), .B1(_06802_ ), .B2(_06804_ ), .ZN(_07051_ ) );
NOR2_X1 _15079_ ( .A1(_07050_ ), .A2(_07051_ ), .ZN(_07052_ ) );
MUX2_X1 _15080_ ( .A(_07049_ ), .B(_07052_ ), .S(_06791_ ), .Z(_07053_ ) );
OAI21_X1 _15081_ ( .A(_07047_ ), .B1(_06847_ ), .B2(_07053_ ), .ZN(_07054_ ) );
BUF_X2 _15082_ ( .A(_07005_ ), .Z(_07055_ ) );
AND2_X1 _15083_ ( .A1(_07054_ ), .A2(_07055_ ), .ZN(_07056_ ) );
OR2_X1 _15084_ ( .A1(_07039_ ), .A2(_07056_ ), .ZN(_07057_ ) );
BUF_X2 _15085_ ( .A(_06764_ ), .Z(_07058_ ) );
XNOR2_X1 _15086_ ( .A(_06677_ ), .B(_06832_ ), .ZN(_07059_ ) );
AND4_X1 _15087_ ( .A1(_06736_ ), .A2(_07058_ ), .A3(_07059_ ), .A4(_06765_ ), .ZN(_07060_ ) );
OAI21_X1 _15088_ ( .A(_06676_ ), .B1(_07057_ ), .B2(_07060_ ), .ZN(_07061_ ) );
INV_X1 _15089_ ( .A(_06817_ ), .ZN(_07062_ ) );
OAI21_X1 _15090_ ( .A(_06726_ ), .B1(_06874_ ), .B2(_06875_ ), .ZN(_07063_ ) );
AOI21_X1 _15091_ ( .A(_06868_ ), .B1(_06838_ ), .B2(_06625_ ), .ZN(_07064_ ) );
OAI21_X1 _15092_ ( .A(_07063_ ), .B1(_07064_ ), .B2(_06771_ ), .ZN(_07065_ ) );
INV_X1 _15093_ ( .A(_07065_ ), .ZN(_07066_ ) );
NAND3_X1 _15094_ ( .A1(_07066_ ), .A2(_06937_ ), .A3(_06878_ ), .ZN(_07067_ ) );
AOI21_X1 _15095_ ( .A(_07062_ ), .B1(_07067_ ), .B2(_06818_ ), .ZN(_07068_ ) );
OAI21_X1 _15096_ ( .A(_06771_ ), .B1(_06859_ ), .B2(_06860_ ), .ZN(_07069_ ) );
AND3_X1 _15097_ ( .A1(_06785_ ), .A2(_04219_ ), .A3(_06787_ ), .ZN(_07070_ ) );
OAI21_X1 _15098_ ( .A(_06796_ ), .B1(_07070_ ), .B2(_06852_ ), .ZN(_07071_ ) );
AOI21_X1 _15099_ ( .A(_06730_ ), .B1(_07069_ ), .B2(_07071_ ), .ZN(_07072_ ) );
OAI21_X1 _15100_ ( .A(_06726_ ), .B1(_06849_ ), .B2(_06850_ ), .ZN(_07073_ ) );
AOI21_X1 _15101_ ( .A(_02600_ ), .B1(_06785_ ), .B2(_06787_ ), .ZN(_07074_ ) );
OAI21_X1 _15102_ ( .A(_06782_ ), .B1(_06836_ ), .B2(_07074_ ), .ZN(_07075_ ) );
AOI21_X1 _15103_ ( .A(_06832_ ), .B1(_07073_ ), .B2(_07075_ ), .ZN(_07076_ ) );
NOR2_X1 _15104_ ( .A1(_07072_ ), .A2(_07076_ ), .ZN(_07077_ ) );
OR3_X1 _15105_ ( .A1(_06828_ ), .A2(_06781_ ), .A3(_06829_ ), .ZN(_07078_ ) );
OR3_X1 _15106_ ( .A1(_06871_ ), .A2(_06872_ ), .A3(_04146_ ), .ZN(_07079_ ) );
AOI21_X1 _15107_ ( .A(_06832_ ), .B1(_07078_ ), .B2(_07079_ ), .ZN(_07080_ ) );
AND3_X1 _15108_ ( .A1(_06772_ ), .A2(_06646_ ), .A3(_06786_ ), .ZN(_07081_ ) );
OAI21_X1 _15109_ ( .A(_06725_ ), .B1(_07081_ ), .B2(_06840_ ), .ZN(_07082_ ) );
OAI21_X1 _15110_ ( .A(_06795_ ), .B1(_06823_ ), .B2(_06824_ ), .ZN(_07083_ ) );
AND3_X1 _15111_ ( .A1(_07082_ ), .A2(_07083_ ), .A3(_06620_ ), .ZN(_07084_ ) );
OR2_X1 _15112_ ( .A1(_07080_ ), .A2(_07084_ ), .ZN(_07085_ ) );
MUX2_X1 _15113_ ( .A(_07077_ ), .B(_07085_ ), .S(_06631_ ), .Z(_07086_ ) );
OAI21_X1 _15114_ ( .A(_07068_ ), .B1(_07086_ ), .B2(_06819_ ), .ZN(_07087_ ) );
NAND3_X1 _15115_ ( .A1(_07054_ ), .A2(_06813_ ), .A3(_06884_ ), .ZN(_07088_ ) );
OAI211_X1 _15116_ ( .A(_07087_ ), .B(_07088_ ), .C1(_04232_ ), .C2(_07009_ ), .ZN(_07089_ ) );
BUF_X2 _15117_ ( .A(_06887_ ), .Z(_07090_ ) );
AOI221_X4 _15118_ ( .A(_07089_ ), .B1(_04231_ ), .B2(_06890_ ), .C1(_04233_ ), .C2(_07090_ ), .ZN(_07091_ ) );
NAND3_X1 _15119_ ( .A1(_07037_ ), .A2(_07061_ ), .A3(_07091_ ), .ZN(_07092_ ) );
AOI21_X1 _15120_ ( .A(_07028_ ), .B1(_07092_ ), .B2(_06900_ ), .ZN(_07093_ ) );
NAND2_X1 _15121_ ( .A1(_04577_ ), .A2(_05029_ ), .ZN(_07094_ ) );
NAND2_X1 _15122_ ( .A1(_07094_ ), .A2(_06259_ ), .ZN(_07095_ ) );
OAI21_X1 _15123_ ( .A(_07016_ ), .B1(_07093_ ), .B2(_07095_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
OR2_X1 _15124_ ( .A1(_04616_ ), .A2(_06258_ ), .ZN(_07096_ ) );
OR3_X1 _15125_ ( .A1(_07020_ ), .A2(_03310_ ), .A3(_04350_ ), .ZN(_07097_ ) );
NAND3_X1 _15126_ ( .A1(_07097_ ), .A2(_06595_ ), .A3(_07021_ ), .ZN(_07098_ ) );
AOI22_X1 _15127_ ( .A1(_04602_ ), .A2(_06915_ ), .B1(\ID_EX_imm [18] ), .B2(_06916_ ), .ZN(_07099_ ) );
AOI21_X1 _15128_ ( .A(_07017_ ), .B1(_07098_ ), .B2(_07099_ ), .ZN(_07100_ ) );
OR2_X1 _15129_ ( .A1(_07100_ ), .A2(_06919_ ), .ZN(_07101_ ) );
BUF_X4 _15130_ ( .A(_07009_ ), .Z(_07102_ ) );
AOI21_X1 _15131_ ( .A(_07102_ ), .B1(_04214_ ), .B2(_06666_ ), .ZN(_07103_ ) );
AND3_X1 _15132_ ( .A1(_07031_ ), .A2(_06664_ ), .A3(_06663_ ), .ZN(_07104_ ) );
NOR3_X1 _15133_ ( .A1(_07104_ ), .A2(_07032_ ), .A3(_06606_ ), .ZN(_07105_ ) );
NAND3_X1 _15134_ ( .A1(_06935_ ), .A2(_04156_ ), .A3(_06771_ ), .ZN(_07106_ ) );
OAI21_X1 _15135_ ( .A(_06725_ ), .B1(_06950_ ), .B2(_06951_ ), .ZN(_07107_ ) );
OAI21_X1 _15136_ ( .A(_06795_ ), .B1(_06931_ ), .B2(_06932_ ), .ZN(_07108_ ) );
NAND3_X1 _15137_ ( .A1(_07107_ ), .A2(_07108_ ), .A3(_06832_ ), .ZN(_07109_ ) );
AND2_X1 _15138_ ( .A1(_07106_ ), .A2(_07109_ ), .ZN(_07110_ ) );
NOR3_X1 _15139_ ( .A1(_06968_ ), .A2(_06795_ ), .A3(_06971_ ), .ZN(_07111_ ) );
NOR3_X1 _15140_ ( .A1(_06940_ ), .A2(_06941_ ), .A3(_06725_ ), .ZN(_07112_ ) );
NOR3_X1 _15141_ ( .A1(_07111_ ), .A2(_07112_ ), .A3(_04156_ ), .ZN(_07113_ ) );
OAI21_X1 _15142_ ( .A(_06725_ ), .B1(_06943_ ), .B2(_06944_ ), .ZN(_07114_ ) );
OAI21_X1 _15143_ ( .A(_06795_ ), .B1(_06947_ ), .B2(_06948_ ), .ZN(_07115_ ) );
AOI21_X1 _15144_ ( .A(_06620_ ), .B1(_07114_ ), .B2(_07115_ ), .ZN(_07116_ ) );
OR2_X1 _15145_ ( .A1(_07113_ ), .A2(_07116_ ), .ZN(_07117_ ) );
MUX2_X1 _15146_ ( .A(_07110_ ), .B(_07117_ ), .S(_06846_ ), .Z(_07118_ ) );
NOR2_X1 _15147_ ( .A1(_07118_ ), .A2(_06820_ ), .ZN(_07119_ ) );
AOI211_X1 _15148_ ( .A(_07103_ ), .B(_07105_ ), .C1(_06885_ ), .C2(_07119_ ), .ZN(_07120_ ) );
NOR2_X1 _15149_ ( .A1(_06929_ ), .A2(_06767_ ), .ZN(_07121_ ) );
AND3_X1 _15150_ ( .A1(_06764_ ), .A2(_06734_ ), .A3(_07059_ ), .ZN(_07122_ ) );
OAI21_X1 _15151_ ( .A(_07122_ ), .B1(_06926_ ), .B2(_06728_ ), .ZN(_07123_ ) );
AOI21_X1 _15152_ ( .A(_07121_ ), .B1(_07123_ ), .B2(_06681_ ), .ZN(_07124_ ) );
OAI21_X1 _15153_ ( .A(_06676_ ), .B1(_07124_ ), .B2(_07119_ ), .ZN(_07125_ ) );
OAI21_X1 _15154_ ( .A(_06770_ ), .B1(_06997_ ), .B2(_06998_ ), .ZN(_07126_ ) );
OAI21_X1 _15155_ ( .A(_07126_ ), .B1(_06726_ ), .B2(_06994_ ), .ZN(_07127_ ) );
BUF_X2 _15156_ ( .A(_06631_ ), .Z(_07128_ ) );
NOR3_X1 _15157_ ( .A1(_07127_ ), .A2(_07128_ ), .A3(_06731_ ), .ZN(_07129_ ) );
OAI21_X1 _15158_ ( .A(_06817_ ), .B1(_07129_ ), .B2(_07005_ ), .ZN(_07130_ ) );
OR3_X1 _15159_ ( .A1(_06970_ ), .A2(_06796_ ), .A3(_06971_ ), .ZN(_07131_ ) );
OR3_X1 _15160_ ( .A1(_06960_ ), .A2(_06961_ ), .A3(_06726_ ), .ZN(_07132_ ) );
NAND2_X1 _15161_ ( .A1(_07131_ ), .A2(_07132_ ), .ZN(_07133_ ) );
NAND2_X1 _15162_ ( .A1(_07133_ ), .A2(_06878_ ), .ZN(_07134_ ) );
NOR3_X1 _15163_ ( .A1(_06963_ ), .A2(_06806_ ), .A3(_06964_ ), .ZN(_07135_ ) );
NOR3_X1 _15164_ ( .A1(_06984_ ), .A2(_06985_ ), .A3(_06771_ ), .ZN(_07136_ ) );
NOR2_X1 _15165_ ( .A1(_07135_ ), .A2(_07136_ ), .ZN(_07137_ ) );
OAI21_X1 _15166_ ( .A(_07134_ ), .B1(_06834_ ), .B2(_07137_ ), .ZN(_07138_ ) );
BUF_X2 _15167_ ( .A(_06937_ ), .Z(_07139_ ) );
AOI21_X1 _15168_ ( .A(_06819_ ), .B1(_07138_ ), .B2(_07139_ ), .ZN(_07140_ ) );
NOR3_X1 _15169_ ( .A1(_06975_ ), .A2(_06795_ ), .A3(_06976_ ), .ZN(_07141_ ) );
NOR3_X1 _15170_ ( .A1(_07000_ ), .A2(_07001_ ), .A3(_06725_ ), .ZN(_07142_ ) );
OR3_X1 _15171_ ( .A1(_07141_ ), .A2(_07142_ ), .A3(_06862_ ), .ZN(_07143_ ) );
OAI21_X1 _15172_ ( .A(_06854_ ), .B1(_06987_ ), .B2(_06988_ ), .ZN(_07144_ ) );
OAI21_X1 _15173_ ( .A(_06806_ ), .B1(_06978_ ), .B2(_06979_ ), .ZN(_07145_ ) );
NAND2_X1 _15174_ ( .A1(_07144_ ), .A2(_07145_ ), .ZN(_07146_ ) );
NAND2_X1 _15175_ ( .A1(_07146_ ), .A2(_06834_ ), .ZN(_07147_ ) );
NAND3_X1 _15176_ ( .A1(_07143_ ), .A2(_07147_ ), .A3(_06991_ ), .ZN(_07148_ ) );
AOI21_X1 _15177_ ( .A(_07130_ ), .B1(_07140_ ), .B2(_07148_ ), .ZN(_07149_ ) );
AOI221_X4 _15178_ ( .A(_07149_ ), .B1(_07033_ ), .B2(_06889_ ), .C1(_04215_ ), .C2(_06887_ ), .ZN(_07150_ ) );
NAND3_X1 _15179_ ( .A1(_07120_ ), .A2(_07125_ ), .A3(_07150_ ), .ZN(_07151_ ) );
AOI21_X1 _15180_ ( .A(_07101_ ), .B1(_07151_ ), .B2(_06900_ ), .ZN(_07152_ ) );
NAND2_X1 _15181_ ( .A1(_04604_ ), .A2(_05029_ ), .ZN(_07153_ ) );
NAND2_X1 _15182_ ( .A1(_07153_ ), .A2(_06259_ ), .ZN(_07154_ ) );
OAI21_X1 _15183_ ( .A(_07096_ ), .B1(_07152_ ), .B2(_07154_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
INV_X1 _15184_ ( .A(_04641_ ), .ZN(_07155_ ) );
AND4_X1 _15185_ ( .A1(_04634_ ), .A2(_04635_ ), .A3(_04637_ ), .A4(_07155_ ), .ZN(_07156_ ) );
NAND4_X1 _15186_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04588_ ), .A4(_07156_ ), .ZN(_07157_ ) );
NAND3_X1 _15187_ ( .A1(_06907_ ), .A2(_04643_ ), .A3(_06908_ ), .ZN(_07158_ ) );
NAND3_X1 _15188_ ( .A1(_07157_ ), .A2(_07158_ ), .A3(_06910_ ), .ZN(_07159_ ) );
OR2_X1 _15189_ ( .A1(_04345_ ), .A2(_07018_ ), .ZN(_07160_ ) );
AND3_X1 _15190_ ( .A1(_07160_ ), .A2(_04349_ ), .A3(_07019_ ), .ZN(_07161_ ) );
AOI21_X1 _15191_ ( .A(_07019_ ), .B1(_07160_ ), .B2(_04349_ ), .ZN(_07162_ ) );
INV_X1 _15192_ ( .A(_06594_ ), .ZN(_07163_ ) );
BUF_X4 _15193_ ( .A(_07163_ ), .Z(_07164_ ) );
NOR3_X1 _15194_ ( .A1(_07161_ ), .A2(_07162_ ), .A3(_07164_ ), .ZN(_07165_ ) );
OAI22_X1 _15195_ ( .A1(_04631_ ), .A2(_06581_ ), .B1(_02477_ ), .B2(_06584_ ), .ZN(_07166_ ) );
OAI21_X1 _15196_ ( .A(_06598_ ), .B1(_07165_ ), .B2(_07166_ ), .ZN(_07167_ ) );
BUF_X2 _15197_ ( .A(_04404_ ), .Z(_07168_ ) );
NAND2_X1 _15198_ ( .A1(_07167_ ), .A2(_07168_ ), .ZN(_07169_ ) );
NAND4_X1 _15199_ ( .A1(_06724_ ), .A2(_06729_ ), .A3(_06736_ ), .A4(_07059_ ), .ZN(_07170_ ) );
AOI22_X1 _15200_ ( .A1(_06681_ ), .A2(_07170_ ), .B1(_06766_ ), .B2(_06768_ ), .ZN(_07171_ ) );
NAND2_X1 _15201_ ( .A1(_06808_ ), .A2(_06809_ ), .ZN(_07172_ ) );
NAND2_X1 _15202_ ( .A1(_06794_ ), .A2(_06799_ ), .ZN(_07173_ ) );
NAND2_X1 _15203_ ( .A1(_07173_ ), .A2(_06833_ ), .ZN(_07174_ ) );
NAND3_X1 _15204_ ( .A1(_07172_ ), .A2(_07128_ ), .A3(_07174_ ), .ZN(_07175_ ) );
OAI21_X1 _15205_ ( .A(_06771_ ), .B1(_06859_ ), .B2(_06852_ ), .ZN(_07176_ ) );
OAI21_X1 _15206_ ( .A(_06796_ ), .B1(_06857_ ), .B2(_06860_ ), .ZN(_07177_ ) );
AOI21_X1 _15207_ ( .A(_06730_ ), .B1(_07176_ ), .B2(_07177_ ), .ZN(_07178_ ) );
AOI21_X1 _15208_ ( .A(_06832_ ), .B1(_06780_ ), .B2(_06789_ ), .ZN(_07179_ ) );
NOR2_X1 _15209_ ( .A1(_07178_ ), .A2(_07179_ ), .ZN(_07180_ ) );
NAND2_X1 _15210_ ( .A1(_07180_ ), .A2(_06937_ ), .ZN(_07181_ ) );
AOI21_X1 _15211_ ( .A(_06820_ ), .B1(_07175_ ), .B2(_07181_ ), .ZN(_07182_ ) );
OAI21_X1 _15212_ ( .A(_06676_ ), .B1(_07171_ ), .B2(_07182_ ), .ZN(_07183_ ) );
INV_X1 _15213_ ( .A(_04220_ ), .ZN(_07184_ ) );
INV_X1 _15214_ ( .A(_04222_ ), .ZN(_07185_ ) );
OAI211_X1 _15215_ ( .A(_07184_ ), .B(_07030_ ), .C1(_07029_ ), .C2(_07185_ ), .ZN(_07186_ ) );
AOI21_X1 _15216_ ( .A(_07185_ ), .B1(_06641_ ), .B2(_06660_ ), .ZN(_07187_ ) );
OAI21_X1 _15217_ ( .A(_04226_ ), .B1(_07187_ ), .B2(_04220_ ), .ZN(_07188_ ) );
NAND3_X1 _15218_ ( .A1(_07186_ ), .A2(_07035_ ), .A3(_07188_ ), .ZN(_07189_ ) );
AOI21_X1 _15219_ ( .A(_07102_ ), .B1(_04225_ ), .B2(_02946_ ), .ZN(_07190_ ) );
AND3_X1 _15220_ ( .A1(_07064_ ), .A2(_06791_ ), .A3(_06727_ ), .ZN(_07191_ ) );
AND2_X1 _15221_ ( .A1(_07191_ ), .A2(_06847_ ), .ZN(_07192_ ) );
OAI21_X1 _15222_ ( .A(_06817_ ), .B1(_07192_ ), .B2(_07005_ ), .ZN(_07193_ ) );
AOI21_X1 _15223_ ( .A(_06833_ ), .B1(_06839_ ), .B2(_06843_ ), .ZN(_07194_ ) );
AOI21_X1 _15224_ ( .A(_06939_ ), .B1(_06851_ ), .B2(_06855_ ), .ZN(_07195_ ) );
OR2_X1 _15225_ ( .A1(_07194_ ), .A2(_07195_ ), .ZN(_07196_ ) );
AOI21_X1 _15226_ ( .A(_06819_ ), .B1(_07196_ ), .B2(_07139_ ), .ZN(_07197_ ) );
NAND2_X1 _15227_ ( .A1(_06831_ ), .A2(_06862_ ), .ZN(_07198_ ) );
NAND2_X1 _15228_ ( .A1(_06877_ ), .A2(_06809_ ), .ZN(_07199_ ) );
NAND3_X1 _15229_ ( .A1(_07198_ ), .A2(_06991_ ), .A3(_07199_ ), .ZN(_07200_ ) );
AOI21_X1 _15230_ ( .A(_07193_ ), .B1(_07197_ ), .B2(_07200_ ), .ZN(_07201_ ) );
NAND2_X1 _15231_ ( .A1(_07175_ ), .A2(_07181_ ), .ZN(_07202_ ) );
AND3_X1 _15232_ ( .A1(_07202_ ), .A2(_07005_ ), .A3(_06883_ ), .ZN(_07203_ ) );
NOR3_X1 _15233_ ( .A1(_04225_ ), .A2(_02946_ ), .A3(_04032_ ), .ZN(_07204_ ) );
OR3_X1 _15234_ ( .A1(_07201_ ), .A2(_07203_ ), .A3(_07204_ ), .ZN(_07205_ ) );
AOI211_X1 _15235_ ( .A(_07190_ ), .B(_07205_ ), .C1(_04226_ ), .C2(_07090_ ), .ZN(_07206_ ) );
NAND3_X1 _15236_ ( .A1(_07183_ ), .A2(_07189_ ), .A3(_07206_ ), .ZN(_07207_ ) );
AOI21_X1 _15237_ ( .A(_07169_ ), .B1(_07207_ ), .B2(_06900_ ), .ZN(_07208_ ) );
NAND2_X1 _15238_ ( .A1(_04628_ ), .A2(_05029_ ), .ZN(_07209_ ) );
NAND2_X1 _15239_ ( .A1(_07209_ ), .A2(_06259_ ), .ZN(_07210_ ) );
OAI21_X1 _15240_ ( .A(_07159_ ), .B1(_07208_ ), .B2(_07210_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
AND2_X1 _15241_ ( .A1(_04656_ ), .A2(_04655_ ), .ZN(_07211_ ) );
NAND4_X1 _15242_ ( .A1(_04451_ ), .A2(_04588_ ), .A3(_04662_ ), .A4(_07211_ ), .ZN(_07212_ ) );
NAND3_X1 _15243_ ( .A1(_06907_ ), .A2(_04664_ ), .A3(_06908_ ), .ZN(_07213_ ) );
NAND3_X1 _15244_ ( .A1(_07212_ ), .A2(_07213_ ), .A3(_06910_ ), .ZN(_07214_ ) );
AOI21_X1 _15245_ ( .A(_07164_ ), .B1(_04346_ ), .B2(_03334_ ), .ZN(_07215_ ) );
OAI21_X1 _15246_ ( .A(_07215_ ), .B1(_03334_ ), .B2(_04346_ ), .ZN(_07216_ ) );
BUF_X4 _15247_ ( .A(_06580_ ), .Z(_07217_ ) );
AOI22_X1 _15248_ ( .A1(_04652_ ), .A2(_07217_ ), .B1(\ID_EX_imm [16] ), .B2(_06916_ ), .ZN(_07218_ ) );
AOI21_X1 _15249_ ( .A(_07017_ ), .B1(_07216_ ), .B2(_07218_ ), .ZN(_07219_ ) );
OR2_X1 _15250_ ( .A1(_07219_ ), .A2(_06919_ ), .ZN(_07220_ ) );
OAI21_X1 _15251_ ( .A(_06605_ ), .B1(_07029_ ), .B2(_07185_ ), .ZN(_07221_ ) );
AOI21_X1 _15252_ ( .A(_07221_ ), .B1(_07185_ ), .B2(_07029_ ), .ZN(_07222_ ) );
OAI211_X1 _15253_ ( .A(_06724_ ), .B(_06765_ ), .C1(_06820_ ), .C2(_06679_ ), .ZN(_07223_ ) );
OR3_X1 _15254_ ( .A1(_06970_ ), .A2(_06781_ ), .A3(_06961_ ), .ZN(_07224_ ) );
OR3_X1 _15255_ ( .A1(_06968_ ), .A2(_06971_ ), .A3(_04146_ ), .ZN(_07225_ ) );
AOI21_X1 _15256_ ( .A(_04156_ ), .B1(_07224_ ), .B2(_07225_ ), .ZN(_07226_ ) );
AOI21_X1 _15257_ ( .A(_06620_ ), .B1(_06942_ ), .B2(_06945_ ), .ZN(_07227_ ) );
OAI21_X1 _15258_ ( .A(_06846_ ), .B1(_07226_ ), .B2(_07227_ ), .ZN(_07228_ ) );
NAND2_X1 _15259_ ( .A1(_06936_ ), .A2(_06730_ ), .ZN(_07229_ ) );
NAND2_X1 _15260_ ( .A1(_06949_ ), .A2(_06952_ ), .ZN(_07230_ ) );
NAND2_X1 _15261_ ( .A1(_07230_ ), .A2(_06832_ ), .ZN(_07231_ ) );
NAND2_X1 _15262_ ( .A1(_07229_ ), .A2(_07231_ ), .ZN(_07232_ ) );
OAI21_X1 _15263_ ( .A(_07228_ ), .B1(_07232_ ), .B2(_06846_ ), .ZN(_07233_ ) );
NAND2_X1 _15264_ ( .A1(_07233_ ), .A2(_07006_ ), .ZN(_07234_ ) );
AOI21_X1 _15265_ ( .A(_06925_ ), .B1(_07223_ ), .B2(_07234_ ), .ZN(_07235_ ) );
INV_X1 _15266_ ( .A(_06883_ ), .ZN(_07236_ ) );
BUF_X2 _15267_ ( .A(_07236_ ), .Z(_07237_ ) );
OAI22_X1 _15268_ ( .A1(_07234_ ), .A2(_07237_ ), .B1(_04221_ ), .B2(_07009_ ), .ZN(_07238_ ) );
AND3_X1 _15269_ ( .A1(_06994_ ), .A2(_06791_ ), .A3(_06727_ ), .ZN(_07239_ ) );
NAND2_X1 _15270_ ( .A1(_07239_ ), .A2(_06847_ ), .ZN(_07240_ ) );
AOI21_X1 _15271_ ( .A(_07062_ ), .B1(_07240_ ), .B2(_06818_ ), .ZN(_07241_ ) );
AOI21_X1 _15272_ ( .A(_06791_ ), .B1(_06986_ ), .B2(_06989_ ), .ZN(_07242_ ) );
AOI21_X1 _15273_ ( .A(_06939_ ), .B1(_06962_ ), .B2(_06965_ ), .ZN(_07243_ ) );
NOR3_X1 _15274_ ( .A1(_07242_ ), .A2(_07243_ ), .A3(_06631_ ), .ZN(_07244_ ) );
NAND2_X1 _15275_ ( .A1(_07003_ ), .A2(_06731_ ), .ZN(_07245_ ) );
NAND2_X1 _15276_ ( .A1(_06981_ ), .A2(_06862_ ), .ZN(_07246_ ) );
NAND2_X1 _15277_ ( .A1(_07245_ ), .A2(_07246_ ), .ZN(_07247_ ) );
AOI21_X1 _15278_ ( .A(_07244_ ), .B1(_06821_ ), .B2(_07247_ ), .ZN(_07248_ ) );
OAI21_X1 _15279_ ( .A(_07241_ ), .B1(_07248_ ), .B2(_06819_ ), .ZN(_07249_ ) );
BUF_X2 _15280_ ( .A(_04032_ ), .Z(_07250_ ) );
BUF_X4 _15281_ ( .A(_04309_ ), .Z(_07251_ ) );
OAI221_X1 _15282_ ( .A(_07249_ ), .B1(_07184_ ), .B2(_07250_ ), .C1(_07185_ ), .C2(_07251_ ), .ZN(_07252_ ) );
OR2_X1 _15283_ ( .A1(_07238_ ), .A2(_07252_ ), .ZN(_07253_ ) );
OR3_X1 _15284_ ( .A1(_07222_ ), .A2(_07235_ ), .A3(_07253_ ), .ZN(_07254_ ) );
AOI21_X1 _15285_ ( .A(_07220_ ), .B1(_07254_ ), .B2(_06900_ ), .ZN(_07255_ ) );
OAI21_X1 _15286_ ( .A(_06500_ ), .B1(_04651_ ), .B2(_05097_ ), .ZN(_07256_ ) );
OAI21_X1 _15287_ ( .A(_07214_ ), .B1(_07255_ ), .B2(_07256_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
NAND2_X1 _15288_ ( .A1(_04678_ ), .A2(_06292_ ), .ZN(_07257_ ) );
AOI21_X1 _15289_ ( .A(_04319_ ), .B1(_04342_ ), .B2(_03933_ ), .ZN(_07258_ ) );
INV_X1 _15290_ ( .A(_03817_ ), .ZN(_07259_ ) );
INV_X1 _15291_ ( .A(_03841_ ), .ZN(_07260_ ) );
NOR3_X1 _15292_ ( .A1(_07258_ ), .A2(_07259_ ), .A3(_07260_ ), .ZN(_07261_ ) );
OR3_X1 _15293_ ( .A1(_07261_ ), .A2(_03839_ ), .A3(_04321_ ), .ZN(_07262_ ) );
AOI21_X1 _15294_ ( .A(_04323_ ), .B1(_07262_ ), .B2(_03794_ ), .ZN(_07263_ ) );
XNOR2_X1 _15295_ ( .A(_07263_ ), .B(_03772_ ), .ZN(_07264_ ) );
NAND2_X1 _15296_ ( .A1(_07264_ ), .A2(_06595_ ), .ZN(_07265_ ) );
AOI22_X1 _15297_ ( .A1(_04688_ ), .A2(_07217_ ), .B1(\ID_EX_imm [15] ), .B2(_06916_ ), .ZN(_07266_ ) );
AOI21_X1 _15298_ ( .A(_07017_ ), .B1(_07265_ ), .B2(_07266_ ), .ZN(_07267_ ) );
OR2_X1 _15299_ ( .A1(_07267_ ), .A2(_06919_ ), .ZN(_07268_ ) );
AND2_X1 _15300_ ( .A1(_06636_ ), .A2(_06640_ ), .ZN(_07269_ ) );
INV_X1 _15301_ ( .A(_07269_ ), .ZN(_07270_ ) );
AOI211_X1 _15302_ ( .A(_04092_ ), .B(_04097_ ), .C1(_07270_ ), .C2(_06648_ ), .ZN(_07271_ ) );
OAI21_X1 _15303_ ( .A(_04070_ ), .B1(_07271_ ), .B2(_06654_ ), .ZN(_07272_ ) );
AND3_X1 _15304_ ( .A1(_07272_ ), .A2(_04074_ ), .A3(_06657_ ), .ZN(_07273_ ) );
AOI21_X1 _15305_ ( .A(_04074_ ), .B1(_07272_ ), .B2(_06657_ ), .ZN(_07274_ ) );
OAI21_X1 _15306_ ( .A(_07035_ ), .B1(_07273_ ), .B2(_07274_ ), .ZN(_07275_ ) );
NAND4_X1 _15307_ ( .A1(_06724_ ), .A2(_06676_ ), .A3(_06680_ ), .A4(_06765_ ), .ZN(_07276_ ) );
NAND2_X1 _15308_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_07277_ ) );
NAND2_X1 _15309_ ( .A1(_07042_ ), .A2(_06878_ ), .ZN(_07278_ ) );
NAND2_X1 _15310_ ( .A1(_07052_ ), .A2(_06731_ ), .ZN(_07279_ ) );
AND3_X1 _15311_ ( .A1(_07278_ ), .A2(_07279_ ), .A3(_06821_ ), .ZN(_07280_ ) );
BUF_X2 _15312_ ( .A(_06846_ ), .Z(_07281_ ) );
BUF_X2 _15313_ ( .A(_07281_ ), .Z(_07282_ ) );
AOI21_X1 _15314_ ( .A(_06878_ ), .B1(_07044_ ), .B2(_07045_ ), .ZN(_07283_ ) );
OR3_X1 _15315_ ( .A1(_07070_ ), .A2(_06782_ ), .A3(_06850_ ), .ZN(_07284_ ) );
OAI211_X1 _15316_ ( .A(_06853_ ), .B(_06806_ ), .C1(_02501_ ), .C2(_06728_ ), .ZN(_07285_ ) );
AOI21_X1 _15317_ ( .A(_06731_ ), .B1(_07284_ ), .B2(_07285_ ), .ZN(_07286_ ) );
OR2_X1 _15318_ ( .A1(_07283_ ), .A2(_07286_ ), .ZN(_07287_ ) );
AOI211_X1 _15319_ ( .A(_06866_ ), .B(_07280_ ), .C1(_07282_ ), .C2(_07287_ ), .ZN(_07288_ ) );
NAND3_X1 _15320_ ( .A1(_07048_ ), .A2(_06623_ ), .A3(_06832_ ), .ZN(_07289_ ) );
AOI211_X1 _15321_ ( .A(_07277_ ), .B(_07288_ ), .C1(_06820_ ), .C2(_07289_ ), .ZN(_07290_ ) );
NAND3_X1 _15322_ ( .A1(_07078_ ), .A2(_06791_ ), .A3(_07079_ ), .ZN(_07291_ ) );
OAI21_X1 _15323_ ( .A(_07291_ ), .B1(_07066_ ), .B2(_06833_ ), .ZN(_07292_ ) );
NAND2_X1 _15324_ ( .A1(_07292_ ), .A2(_07128_ ), .ZN(_07293_ ) );
AOI21_X1 _15325_ ( .A(_06939_ ), .B1(_07073_ ), .B2(_07075_ ), .ZN(_07294_ ) );
AOI21_X1 _15326_ ( .A(_06833_ ), .B1(_07082_ ), .B2(_07083_ ), .ZN(_07295_ ) );
OAI21_X1 _15327_ ( .A(_06847_ ), .B1(_07294_ ), .B2(_07295_ ), .ZN(_07296_ ) );
AND2_X1 _15328_ ( .A1(_06812_ ), .A2(_04388_ ), .ZN(_07297_ ) );
BUF_X2 _15329_ ( .A(_07297_ ), .Z(_07298_ ) );
AND3_X1 _15330_ ( .A1(_07293_ ), .A2(_07296_ ), .A3(_07298_ ), .ZN(_07299_ ) );
NOR3_X1 _15331_ ( .A1(_06658_ ), .A2(_06651_ ), .A3(_07251_ ), .ZN(_07300_ ) );
NAND3_X1 _15332_ ( .A1(_04185_ ), .A2(_02553_ ), .A3(_06889_ ), .ZN(_07301_ ) );
OAI21_X1 _15333_ ( .A(_07301_ ), .B1(_06658_ ), .B2(_07102_ ), .ZN(_07302_ ) );
NOR4_X1 _15334_ ( .A1(_07290_ ), .A2(_07299_ ), .A3(_07300_ ), .A4(_07302_ ), .ZN(_07303_ ) );
NAND3_X1 _15335_ ( .A1(_07275_ ), .A2(_07276_ ), .A3(_07303_ ), .ZN(_07304_ ) );
AOI21_X1 _15336_ ( .A(_07268_ ), .B1(_07304_ ), .B2(_06900_ ), .ZN(_07305_ ) );
OAI21_X1 _15337_ ( .A(_06500_ ), .B1(_04680_ ), .B2(_05097_ ), .ZN(_07306_ ) );
OAI21_X1 _15338_ ( .A(_07257_ ), .B1(_07305_ ), .B2(_07306_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
AND4_X1 _15339_ ( .A1(_04705_ ), .A2(_04703_ ), .A3(_04701_ ), .A4(_04700_ ), .ZN(_07307_ ) );
NAND4_X1 _15340_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04588_ ), .A4(_07307_ ), .ZN(_07308_ ) );
NAND3_X1 _15341_ ( .A1(_06907_ ), .A2(_04708_ ), .A3(_06908_ ), .ZN(_07309_ ) );
NAND3_X1 _15342_ ( .A1(_07308_ ), .A2(_07309_ ), .A3(_06910_ ), .ZN(_07310_ ) );
AOI21_X1 _15343_ ( .A(_07164_ ), .B1(_07262_ ), .B2(_03794_ ), .ZN(_07311_ ) );
OAI21_X1 _15344_ ( .A(_07311_ ), .B1(_03794_ ), .B2(_07262_ ), .ZN(_07312_ ) );
AOI22_X1 _15345_ ( .A1(_04696_ ), .A2(_07217_ ), .B1(\ID_EX_imm [14] ), .B2(_06916_ ), .ZN(_07313_ ) );
AOI21_X1 _15346_ ( .A(_07017_ ), .B1(_07312_ ), .B2(_07313_ ), .ZN(_07314_ ) );
OR2_X1 _15347_ ( .A1(_07314_ ), .A2(_06919_ ), .ZN(_07315_ ) );
BUF_X4 _15348_ ( .A(_07038_ ), .Z(_07316_ ) );
NAND3_X1 _15349_ ( .A1(_06838_ ), .A2(_06833_ ), .A3(_06967_ ), .ZN(_07317_ ) );
OAI211_X1 _15350_ ( .A(_06724_ ), .B(_07316_ ), .C1(_06735_ ), .C2(_07317_ ), .ZN(_07318_ ) );
AOI21_X1 _15351_ ( .A(_04156_ ), .B1(_07114_ ), .B2(_07115_ ), .ZN(_07319_ ) );
AOI21_X1 _15352_ ( .A(_06620_ ), .B1(_07107_ ), .B2(_07108_ ), .ZN(_07320_ ) );
NOR2_X1 _15353_ ( .A1(_07319_ ), .A2(_07320_ ), .ZN(_07321_ ) );
OAI21_X1 _15354_ ( .A(_06730_ ), .B1(_07111_ ), .B2(_07112_ ), .ZN(_07322_ ) );
OR3_X1 _15355_ ( .A1(_06960_ ), .A2(_06795_ ), .A3(_06964_ ), .ZN(_07323_ ) );
OR3_X1 _15356_ ( .A1(_06970_ ), .A2(_06961_ ), .A3(_06725_ ), .ZN(_07324_ ) );
AND2_X1 _15357_ ( .A1(_07323_ ), .A2(_07324_ ), .ZN(_07325_ ) );
OAI21_X1 _15358_ ( .A(_07322_ ), .B1(_07325_ ), .B2(_06939_ ), .ZN(_07326_ ) );
MUX2_X1 _15359_ ( .A(_07321_ ), .B(_07326_ ), .S(_06937_ ), .Z(_07327_ ) );
AND2_X1 _15360_ ( .A1(_07327_ ), .A2(_06813_ ), .ZN(_07328_ ) );
AND3_X1 _15361_ ( .A1(_06935_ ), .A2(_06620_ ), .A3(_06726_ ), .ZN(_07329_ ) );
AND3_X1 _15362_ ( .A1(_07329_ ), .A2(_06819_ ), .A3(_07139_ ), .ZN(_07330_ ) );
NOR2_X1 _15363_ ( .A1(_07328_ ), .A2(_07330_ ), .ZN(_07331_ ) );
AOI21_X1 _15364_ ( .A(_06924_ ), .B1(_07318_ ), .B2(_07331_ ), .ZN(_07332_ ) );
NOR2_X1 _15365_ ( .A1(_07331_ ), .A2(_07237_ ), .ZN(_07333_ ) );
NOR2_X1 _15366_ ( .A1(_07332_ ), .A2(_07333_ ), .ZN(_07334_ ) );
NOR2_X1 _15367_ ( .A1(_07141_ ), .A2(_07142_ ), .ZN(_07335_ ) );
MUX2_X1 _15368_ ( .A(_07127_ ), .B(_07335_ ), .S(_06832_ ), .Z(_07336_ ) );
BUF_X2 _15369_ ( .A(_06991_ ), .Z(_07337_ ) );
NAND2_X1 _15370_ ( .A1(_07336_ ), .A2(_07337_ ), .ZN(_07338_ ) );
NAND2_X1 _15371_ ( .A1(_07137_ ), .A2(_06862_ ), .ZN(_07339_ ) );
NAND2_X1 _15372_ ( .A1(_07146_ ), .A2(_06809_ ), .ZN(_07340_ ) );
NAND2_X1 _15373_ ( .A1(_07339_ ), .A2(_07340_ ), .ZN(_07341_ ) );
NAND2_X1 _15374_ ( .A1(_07341_ ), .A2(_07282_ ), .ZN(_07342_ ) );
NAND3_X1 _15375_ ( .A1(_07338_ ), .A2(_07298_ ), .A3(_07342_ ), .ZN(_07343_ ) );
AND2_X1 _15376_ ( .A1(_07334_ ), .A2(_07343_ ), .ZN(_07344_ ) );
OR3_X1 _15377_ ( .A1(_07271_ ), .A2(_04070_ ), .A3(_06654_ ), .ZN(_07345_ ) );
NAND3_X1 _15378_ ( .A1(_07345_ ), .A2(_07035_ ), .A3(_07272_ ), .ZN(_07346_ ) );
NAND2_X1 _15379_ ( .A1(_04070_ ), .A2(_07090_ ), .ZN(_07347_ ) );
NAND3_X1 _15380_ ( .A1(_04167_ ), .A2(_02575_ ), .A3(_06890_ ), .ZN(_07348_ ) );
OAI21_X1 _15381_ ( .A(_04394_ ), .B1(_04167_ ), .B2(_02575_ ), .ZN(_07349_ ) );
AND3_X1 _15382_ ( .A1(_07347_ ), .A2(_07348_ ), .A3(_07349_ ), .ZN(_07350_ ) );
NAND3_X1 _15383_ ( .A1(_07344_ ), .A2(_07346_ ), .A3(_07350_ ), .ZN(_07351_ ) );
AOI21_X1 _15384_ ( .A(_07315_ ), .B1(_07351_ ), .B2(_06900_ ), .ZN(_07352_ ) );
NAND2_X1 _15385_ ( .A1(_04698_ ), .A2(_05029_ ), .ZN(_07353_ ) );
NAND2_X1 _15386_ ( .A1(_07353_ ), .A2(_06500_ ), .ZN(_07354_ ) );
OAI21_X1 _15387_ ( .A(_07310_ ), .B1(_07352_ ), .B2(_07354_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
NAND3_X1 _15388_ ( .A1(_04732_ ), .A2(_04734_ ), .A3(_06910_ ), .ZN(_07355_ ) );
NOR2_X1 _15389_ ( .A1(_07258_ ), .A2(_07259_ ), .ZN(_07356_ ) );
AOI21_X1 _15390_ ( .A(_07356_ ), .B1(_02622_ ), .B2(_03816_ ), .ZN(_07357_ ) );
AND2_X1 _15391_ ( .A1(_07357_ ), .A2(_07260_ ), .ZN(_07358_ ) );
OAI21_X1 _15392_ ( .A(_06594_ ), .B1(_07357_ ), .B2(_07260_ ), .ZN(_07359_ ) );
OR2_X1 _15393_ ( .A1(_07358_ ), .A2(_07359_ ), .ZN(_07360_ ) );
BUF_X4 _15394_ ( .A(_06583_ ), .Z(_07361_ ) );
AOI22_X1 _15395_ ( .A1(_04721_ ), .A2(_07217_ ), .B1(\ID_EX_imm [13] ), .B2(_07361_ ), .ZN(_07362_ ) );
AOI21_X1 _15396_ ( .A(_07017_ ), .B1(_07360_ ), .B2(_07362_ ), .ZN(_07363_ ) );
CLKBUF_X2 _15397_ ( .A(_04487_ ), .Z(_07364_ ) );
OR2_X1 _15398_ ( .A1(_07363_ ), .A2(_07364_ ), .ZN(_07365_ ) );
OAI211_X1 _15399_ ( .A(_06723_ ), .B(_07038_ ), .C1(_06732_ ), .C2(_06735_ ), .ZN(_07366_ ) );
NOR2_X1 _15400_ ( .A1(_06801_ ), .A2(_06847_ ), .ZN(_07367_ ) );
NAND3_X1 _15401_ ( .A1(_07176_ ), .A2(_07177_ ), .A3(_06939_ ), .ZN(_07368_ ) );
OAI21_X1 _15402_ ( .A(_06854_ ), .B1(_06849_ ), .B2(_07074_ ), .ZN(_07369_ ) );
OAI21_X1 _15403_ ( .A(_06806_ ), .B1(_07070_ ), .B2(_06850_ ), .ZN(_07370_ ) );
NAND3_X1 _15404_ ( .A1(_07369_ ), .A2(_07370_ ), .A3(_06791_ ), .ZN(_07371_ ) );
AND3_X1 _15405_ ( .A1(_07368_ ), .A2(_07371_ ), .A3(_06937_ ), .ZN(_07372_ ) );
OAI21_X1 _15406_ ( .A(_07005_ ), .B1(_07367_ ), .B2(_07372_ ), .ZN(_07373_ ) );
NOR3_X1 _15407_ ( .A1(_06808_ ), .A2(_06631_ ), .A3(_06809_ ), .ZN(_07374_ ) );
OR2_X1 _15408_ ( .A1(_07374_ ), .A2(_06812_ ), .ZN(_07375_ ) );
NAND2_X1 _15409_ ( .A1(_07373_ ), .A2(_07375_ ), .ZN(_07376_ ) );
AOI21_X1 _15410_ ( .A(_06924_ ), .B1(_07366_ ), .B2(_07376_ ), .ZN(_07377_ ) );
AND3_X1 _15411_ ( .A1(_07373_ ), .A2(_06884_ ), .A3(_07375_ ), .ZN(_07378_ ) );
INV_X1 _15412_ ( .A(_07297_ ), .ZN(_07379_ ) );
OAI21_X1 _15413_ ( .A(_07139_ ), .B1(_06835_ ), .B2(_06844_ ), .ZN(_07380_ ) );
NAND3_X1 _15414_ ( .A1(_06870_ ), .A2(_06879_ ), .A3(_06991_ ), .ZN(_07381_ ) );
AOI21_X1 _15415_ ( .A(_07379_ ), .B1(_07380_ ), .B2(_07381_ ), .ZN(_07382_ ) );
OR3_X1 _15416_ ( .A1(_07377_ ), .A2(_07378_ ), .A3(_07382_ ), .ZN(_07383_ ) );
AOI21_X1 _15417_ ( .A(_04092_ ), .B1(_07270_ ), .B2(_06648_ ), .ZN(_07384_ ) );
OR3_X1 _15418_ ( .A1(_07384_ ), .A2(_06652_ ), .A3(_04097_ ), .ZN(_07385_ ) );
OAI21_X1 _15419_ ( .A(_04097_ ), .B1(_07384_ ), .B2(_06652_ ), .ZN(_07386_ ) );
AOI21_X1 _15420_ ( .A(_06607_ ), .B1(_07385_ ), .B2(_07386_ ), .ZN(_07387_ ) );
NAND2_X1 _15421_ ( .A1(_04096_ ), .A2(_07090_ ), .ZN(_07388_ ) );
NAND3_X1 _15422_ ( .A1(_06748_ ), .A2(_02600_ ), .A3(_06890_ ), .ZN(_07389_ ) );
OAI21_X1 _15423_ ( .A(_04394_ ), .B1(_06748_ ), .B2(_02600_ ), .ZN(_07390_ ) );
NAND3_X1 _15424_ ( .A1(_07388_ ), .A2(_07389_ ), .A3(_07390_ ), .ZN(_07391_ ) );
OR3_X1 _15425_ ( .A1(_07383_ ), .A2(_07387_ ), .A3(_07391_ ), .ZN(_07392_ ) );
AOI21_X1 _15426_ ( .A(_07365_ ), .B1(_07392_ ), .B2(_06900_ ), .ZN(_07393_ ) );
BUF_X4 _15427_ ( .A(_06257_ ), .Z(_07394_ ) );
OAI21_X1 _15428_ ( .A(_07394_ ), .B1(_04718_ ), .B2(_05097_ ), .ZN(_07395_ ) );
OAI21_X1 _15429_ ( .A(_07355_ ), .B1(_07393_ ), .B2(_07395_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _15430_ ( .A1(_04748_ ), .A2(_04750_ ), .A3(_06910_ ), .ZN(_07396_ ) );
AND2_X1 _15431_ ( .A1(_07258_ ), .A2(_07259_ ), .ZN(_07397_ ) );
OR3_X1 _15432_ ( .A1(_07397_ ), .A2(_07356_ ), .A3(_07163_ ), .ZN(_07398_ ) );
AOI22_X1 _15433_ ( .A1(_04740_ ), .A2(_07217_ ), .B1(\ID_EX_imm [12] ), .B2(_07361_ ), .ZN(_07399_ ) );
AOI21_X1 _15434_ ( .A(_07017_ ), .B1(_07398_ ), .B2(_07399_ ), .ZN(_07400_ ) );
OR2_X1 _15435_ ( .A1(_07400_ ), .A2(_07364_ ), .ZN(_07401_ ) );
OAI211_X1 _15436_ ( .A(_06724_ ), .B(_07316_ ), .C1(_06736_ ), .C2(_06927_ ), .ZN(_07402_ ) );
OR3_X1 _15437_ ( .A1(_06936_ ), .A2(_07128_ ), .A3(_06731_ ), .ZN(_07403_ ) );
NAND2_X1 _15438_ ( .A1(_07403_ ), .A2(_06820_ ), .ZN(_07404_ ) );
OAI21_X1 _15439_ ( .A(_07337_ ), .B1(_06946_ ), .B2(_06953_ ), .ZN(_07405_ ) );
OR3_X1 _15440_ ( .A1(_06963_ ), .A2(_06781_ ), .A3(_06985_ ), .ZN(_07406_ ) );
OR3_X1 _15441_ ( .A1(_06960_ ), .A2(_06964_ ), .A3(_04146_ ), .ZN(_07407_ ) );
NAND3_X1 _15442_ ( .A1(_07406_ ), .A2(_07407_ ), .A3(_06834_ ), .ZN(_07408_ ) );
NAND3_X1 _15443_ ( .A1(_07224_ ), .A2(_07225_ ), .A3(_06731_ ), .ZN(_07409_ ) );
NAND3_X1 _15444_ ( .A1(_07408_ ), .A2(_07409_ ), .A3(_06848_ ), .ZN(_07410_ ) );
NAND3_X1 _15445_ ( .A1(_07405_ ), .A2(_07410_ ), .A3(_07055_ ), .ZN(_07411_ ) );
NAND2_X1 _15446_ ( .A1(_07404_ ), .A2(_07411_ ), .ZN(_07412_ ) );
AOI21_X1 _15447_ ( .A(_06925_ ), .B1(_07402_ ), .B2(_07412_ ), .ZN(_07413_ ) );
AND3_X1 _15448_ ( .A1(_07404_ ), .A2(_07411_ ), .A3(_06885_ ), .ZN(_07414_ ) );
NOR2_X1 _15449_ ( .A1(_07413_ ), .A2(_07414_ ), .ZN(_07415_ ) );
AND3_X1 _15450_ ( .A1(_07270_ ), .A2(_04092_ ), .A3(_06648_ ), .ZN(_07416_ ) );
OR3_X1 _15451_ ( .A1(_07416_ ), .A2(_07384_ ), .A3(_06607_ ), .ZN(_07417_ ) );
AOI21_X1 _15452_ ( .A(_06821_ ), .B1(_06983_ ), .B2(_06990_ ), .ZN(_07418_ ) );
AOI21_X1 _15453_ ( .A(_07418_ ), .B1(_06822_ ), .B2(_07004_ ), .ZN(_07419_ ) );
NAND2_X1 _15454_ ( .A1(_07419_ ), .A2(_07298_ ), .ZN(_07420_ ) );
NAND2_X1 _15455_ ( .A1(_04091_ ), .A2(_07090_ ), .ZN(_07421_ ) );
OAI21_X1 _15456_ ( .A(_04394_ ), .B1(_04180_ ), .B2(_02622_ ), .ZN(_07422_ ) );
NAND3_X1 _15457_ ( .A1(_04180_ ), .A2(_02622_ ), .A3(_06890_ ), .ZN(_07423_ ) );
AND4_X1 _15458_ ( .A1(_07420_ ), .A2(_07421_ ), .A3(_07422_ ), .A4(_07423_ ), .ZN(_07424_ ) );
NAND3_X1 _15459_ ( .A1(_07415_ ), .A2(_07417_ ), .A3(_07424_ ), .ZN(_07425_ ) );
AOI21_X1 _15460_ ( .A(_07401_ ), .B1(_07425_ ), .B2(_06900_ ), .ZN(_07426_ ) );
OAI21_X1 _15461_ ( .A(_07394_ ), .B1(_04739_ ), .B2(_05097_ ), .ZN(_07427_ ) );
OAI21_X1 _15462_ ( .A(_07396_ ), .B1(_07426_ ), .B2(_07427_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
NAND3_X1 _15463_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04478_ ), .ZN(_07428_ ) );
INV_X1 _15464_ ( .A(_04440_ ), .ZN(_07429_ ) );
NAND3_X1 _15465_ ( .A1(_07428_ ), .A2(_07429_ ), .A3(_06910_ ), .ZN(_07430_ ) );
OAI21_X1 _15466_ ( .A(_03558_ ), .B1(_04347_ ), .B2(_04366_ ), .ZN(_07431_ ) );
AND2_X1 _15467_ ( .A1(_07431_ ), .A2(_04374_ ), .ZN(_07432_ ) );
INV_X1 _15468_ ( .A(_03580_ ), .ZN(_07433_ ) );
NOR2_X1 _15469_ ( .A1(_07432_ ), .A2(_07433_ ), .ZN(_07434_ ) );
INV_X1 _15470_ ( .A(_07434_ ), .ZN(_07435_ ) );
AOI21_X1 _15471_ ( .A(_04383_ ), .B1(_07435_ ), .B2(_04382_ ), .ZN(_07436_ ) );
AOI21_X1 _15472_ ( .A(_07164_ ), .B1(_07436_ ), .B2(_03647_ ), .ZN(_07437_ ) );
OAI21_X1 _15473_ ( .A(_07437_ ), .B1(_03647_ ), .B2(_07436_ ), .ZN(_07438_ ) );
AOI22_X1 _15474_ ( .A1(_03223_ ), .A2(_06915_ ), .B1(\ID_EX_imm [30] ), .B2(_06916_ ), .ZN(_07439_ ) );
AOI21_X1 _15475_ ( .A(_06601_ ), .B1(_07438_ ), .B2(_07439_ ), .ZN(_07440_ ) );
OR2_X1 _15476_ ( .A1(_07440_ ), .A2(_06919_ ), .ZN(_07441_ ) );
AND4_X1 _15477_ ( .A1(_04046_ ), .A2(_04039_ ), .A3(_04264_ ), .A4(_04259_ ), .ZN(_07442_ ) );
AND2_X1 _15478_ ( .A1(_04209_ ), .A2(_04203_ ), .ZN(_07443_ ) );
AND3_X1 _15479_ ( .A1(_07443_ ), .A2(_04198_ ), .A3(_04191_ ), .ZN(_07444_ ) );
INV_X1 _15480_ ( .A(_07444_ ), .ZN(_07445_ ) );
AOI211_X2 _15481_ ( .A(_06610_ ), .B(_07445_ ), .C1(_06641_ ), .C2(_06660_ ), .ZN(_07446_ ) );
NOR2_X1 _15482_ ( .A1(_06668_ ), .A2(_07445_ ), .ZN(_07447_ ) );
AOI21_X1 _15483_ ( .A(_06888_ ), .B1(_04209_ ), .B2(_06670_ ), .ZN(_07448_ ) );
INV_X1 _15484_ ( .A(_04198_ ), .ZN(_07449_ ) );
INV_X1 _15485_ ( .A(_04191_ ), .ZN(_07450_ ) );
NOR3_X1 _15486_ ( .A1(_07448_ ), .A2(_07449_ ), .A3(_07450_ ), .ZN(_07451_ ) );
NOR4_X1 _15487_ ( .A1(_04196_ ), .A2(_04197_ ), .A3(_04248_ ), .A4(_04190_ ), .ZN(_07452_ ) );
NOR4_X1 _15488_ ( .A1(_07447_ ), .A2(_04196_ ), .A3(_07451_ ), .A4(_07452_ ), .ZN(_07453_ ) );
INV_X1 _15489_ ( .A(_07453_ ), .ZN(_07454_ ) );
OAI21_X1 _15490_ ( .A(_07442_ ), .B1(_07446_ ), .B2(_07454_ ), .ZN(_07455_ ) );
NOR2_X1 _15491_ ( .A1(_04045_ ), .A2(_04064_ ), .ZN(_07456_ ) );
NOR3_X1 _15492_ ( .A1(_04062_ ), .A2(_04037_ ), .A3(_04038_ ), .ZN(_07457_ ) );
AOI21_X1 _15493_ ( .A(_04058_ ), .B1(_04259_ ), .B2(_04262_ ), .ZN(_07458_ ) );
INV_X1 _15494_ ( .A(_07458_ ), .ZN(_07459_ ) );
AOI221_X4 _15495_ ( .A(_07456_ ), .B1(_04046_ ), .B2(_04037_ ), .C1(_07457_ ), .C2(_07459_ ), .ZN(_07460_ ) );
AOI21_X1 _15496_ ( .A(_04292_ ), .B1(_07455_ ), .B2(_07460_ ), .ZN(_07461_ ) );
AND2_X1 _15497_ ( .A1(_04289_ ), .A2(_02224_ ), .ZN(_07462_ ) );
OR3_X2 _15498_ ( .A1(_07461_ ), .A2(_04296_ ), .A3(_07462_ ), .ZN(_07463_ ) );
INV_X1 _15499_ ( .A(_04297_ ), .ZN(_07464_ ) );
AND3_X1 _15500_ ( .A1(_07463_ ), .A2(_07464_ ), .A3(_04271_ ), .ZN(_07465_ ) );
AOI21_X1 _15501_ ( .A(_04271_ ), .B1(_07463_ ), .B2(_07464_ ), .ZN(_07466_ ) );
OR3_X1 _15502_ ( .A1(_07465_ ), .A2(_07466_ ), .A3(_06607_ ), .ZN(_07467_ ) );
OAI211_X1 _15503_ ( .A(_06723_ ), .B(_07317_ ), .C1(_06765_ ), .C2(_06767_ ), .ZN(_07468_ ) );
INV_X1 _15504_ ( .A(_07468_ ), .ZN(_07469_ ) );
AND2_X1 _15505_ ( .A1(_07329_ ), .A2(_06937_ ), .ZN(_07470_ ) );
AND2_X1 _15506_ ( .A1(_07470_ ), .A2(_07005_ ), .ZN(_07471_ ) );
OR2_X1 _15507_ ( .A1(_07469_ ), .A2(_07471_ ), .ZN(_07472_ ) );
NAND3_X1 _15508_ ( .A1(_06764_ ), .A2(_06735_ ), .A3(_06767_ ), .ZN(_07473_ ) );
NAND2_X1 _15509_ ( .A1(_06764_ ), .A2(_07038_ ), .ZN(_07474_ ) );
NAND2_X1 _15510_ ( .A1(_07473_ ), .A2(_07474_ ), .ZN(_07475_ ) );
OAI21_X1 _15511_ ( .A(_06675_ ), .B1(_07472_ ), .B2(_07475_ ), .ZN(_07476_ ) );
NOR2_X1 _15512_ ( .A1(_06812_ ), .A2(_07062_ ), .ZN(_07477_ ) );
NAND3_X1 _15513_ ( .A1(_07338_ ), .A2(_07342_ ), .A3(_07477_ ), .ZN(_07478_ ) );
AND3_X1 _15514_ ( .A1(_07131_ ), .A2(_06809_ ), .A3(_07132_ ), .ZN(_07479_ ) );
OAI21_X1 _15515_ ( .A(_06727_ ), .B1(_06940_ ), .B2(_06944_ ), .ZN(_07480_ ) );
OAI21_X1 _15516_ ( .A(_06842_ ), .B1(_06968_ ), .B2(_06941_ ), .ZN(_07481_ ) );
AOI21_X1 _15517_ ( .A(_06809_ ), .B1(_07480_ ), .B2(_07481_ ), .ZN(_07482_ ) );
OAI21_X1 _15518_ ( .A(_07337_ ), .B1(_07479_ ), .B2(_07482_ ), .ZN(_07483_ ) );
OAI21_X1 _15519_ ( .A(_06967_ ), .B1(_06947_ ), .B2(_06951_ ), .ZN(_07484_ ) );
OAI21_X1 _15520_ ( .A(_06926_ ), .B1(_06943_ ), .B2(_06948_ ), .ZN(_07485_ ) );
NAND3_X1 _15521_ ( .A1(_07484_ ), .A2(_07485_ ), .A3(_06982_ ), .ZN(_07486_ ) );
OAI21_X1 _15522_ ( .A(_06967_ ), .B1(_06934_ ), .B2(_06931_ ), .ZN(_07487_ ) );
NOR2_X1 _15523_ ( .A1(_06950_ ), .A2(_06932_ ), .ZN(_07488_ ) );
OAI21_X1 _15524_ ( .A(_07487_ ), .B1(_07488_ ), .B2(_06967_ ), .ZN(_07489_ ) );
OAI211_X1 _15525_ ( .A(_07282_ ), .B(_07486_ ), .C1(_07489_ ), .C2(_06982_ ), .ZN(_07490_ ) );
NAND3_X1 _15526_ ( .A1(_07483_ ), .A2(_07298_ ), .A3(_07490_ ), .ZN(_07491_ ) );
NAND3_X1 _15527_ ( .A1(_07470_ ), .A2(_07006_ ), .A3(_06884_ ), .ZN(_07492_ ) );
OAI21_X1 _15528_ ( .A(_04394_ ), .B1(_04270_ ), .B2(_06803_ ), .ZN(_07493_ ) );
AND3_X1 _15529_ ( .A1(_06803_ ), .A2(_04269_ ), .A3(_04268_ ), .ZN(_07494_ ) );
AOI22_X1 _15530_ ( .A1(_04271_ ), .A2(_06887_ ), .B1(_07494_ ), .B2(_06889_ ), .ZN(_07495_ ) );
AND3_X1 _15531_ ( .A1(_07492_ ), .A2(_07493_ ), .A3(_07495_ ), .ZN(_07496_ ) );
AND4_X1 _15532_ ( .A1(_07476_ ), .A2(_07478_ ), .A3(_07491_ ), .A4(_07496_ ), .ZN(_07497_ ) );
AOI21_X1 _15533_ ( .A(_06898_ ), .B1(_07467_ ), .B2(_07497_ ), .ZN(_07498_ ) );
OAI22_X1 _15534_ ( .A1(_07441_ ), .A2(_07498_ ), .B1(_07168_ ), .B2(_03104_ ), .ZN(_07499_ ) );
OAI21_X1 _15535_ ( .A(_07430_ ), .B1(_07499_ ), .B2(_06491_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _15536_ ( .A1(_04770_ ), .A2(_04772_ ), .A3(_06335_ ), .ZN(_07500_ ) );
INV_X1 _15537_ ( .A(_03910_ ), .ZN(_07501_ ) );
AND4_X1 _15538_ ( .A1(_02627_ ), .A2(_03911_ ), .A3(_02646_ ), .A4(_03930_ ), .ZN(_07502_ ) );
NOR4_X1 _15539_ ( .A1(_04341_ ), .A2(_07501_ ), .A3(_04310_ ), .A4(_07502_ ), .ZN(_07503_ ) );
OAI21_X1 _15540_ ( .A(_03887_ ), .B1(_07503_ ), .B2(_04313_ ), .ZN(_07504_ ) );
INV_X1 _15541_ ( .A(_04316_ ), .ZN(_07505_ ) );
AND2_X1 _15542_ ( .A1(_07504_ ), .A2(_07505_ ), .ZN(_07506_ ) );
XNOR2_X1 _15543_ ( .A(_07506_ ), .B(_03865_ ), .ZN(_07507_ ) );
NAND2_X1 _15544_ ( .A1(_07507_ ), .A2(_06595_ ), .ZN(_07508_ ) );
AOI22_X1 _15545_ ( .A1(_04761_ ), .A2(_07217_ ), .B1(\ID_EX_imm [11] ), .B2(_07361_ ), .ZN(_07509_ ) );
AOI21_X1 _15546_ ( .A(_07017_ ), .B1(_07508_ ), .B2(_07509_ ), .ZN(_07510_ ) );
OR2_X1 _15547_ ( .A1(_07510_ ), .A2(_07364_ ), .ZN(_07511_ ) );
INV_X1 _15548_ ( .A(_06636_ ), .ZN(_07512_ ) );
AOI21_X1 _15549_ ( .A(_06644_ ), .B1(_07512_ ), .B2(_06643_ ), .ZN(_07513_ ) );
NOR2_X1 _15550_ ( .A1(_04078_ ), .A2(_06646_ ), .ZN(_07514_ ) );
OR3_X1 _15551_ ( .A1(_07513_ ), .A2(_04086_ ), .A3(_07514_ ), .ZN(_07515_ ) );
OAI21_X1 _15552_ ( .A(_04086_ ), .B1(_07513_ ), .B2(_07514_ ), .ZN(_07516_ ) );
AND3_X1 _15553_ ( .A1(_07515_ ), .A2(_06605_ ), .A3(_07516_ ), .ZN(_07517_ ) );
OAI211_X1 _15554_ ( .A(_06724_ ), .B(_07316_ ), .C1(_06736_ ), .C2(_07059_ ), .ZN(_07518_ ) );
OAI21_X1 _15555_ ( .A(_07128_ ), .B1(_07043_ ), .B2(_07046_ ), .ZN(_07519_ ) );
NAND3_X1 _15556_ ( .A1(_07284_ ), .A2(_07285_ ), .A3(_06939_ ), .ZN(_07520_ ) );
OAI21_X1 _15557_ ( .A(_06854_ ), .B1(_06836_ ), .B2(_06840_ ), .ZN(_07521_ ) );
OAI21_X1 _15558_ ( .A(_06796_ ), .B1(_06849_ ), .B2(_07074_ ), .ZN(_07522_ ) );
NAND2_X1 _15559_ ( .A1(_07521_ ), .A2(_07522_ ), .ZN(_07523_ ) );
NAND2_X1 _15560_ ( .A1(_07523_ ), .A2(_06833_ ), .ZN(_07524_ ) );
NAND3_X1 _15561_ ( .A1(_07520_ ), .A2(_07524_ ), .A3(_06937_ ), .ZN(_07525_ ) );
AOI21_X1 _15562_ ( .A(_06818_ ), .B1(_07519_ ), .B2(_07525_ ), .ZN(_07526_ ) );
NOR3_X1 _15563_ ( .A1(_07053_ ), .A2(_06812_ ), .A3(_07128_ ), .ZN(_07527_ ) );
NOR2_X1 _15564_ ( .A1(_07526_ ), .A2(_07527_ ), .ZN(_07528_ ) );
AOI21_X1 _15565_ ( .A(_06925_ ), .B1(_07518_ ), .B2(_07528_ ), .ZN(_07529_ ) );
NOR2_X1 _15566_ ( .A1(_07528_ ), .A2(_07237_ ), .ZN(_07530_ ) );
OAI21_X1 _15567_ ( .A(_07281_ ), .B1(_07080_ ), .B2(_07084_ ), .ZN(_07531_ ) );
NAND3_X1 _15568_ ( .A1(_07066_ ), .A2(_06821_ ), .A3(_06834_ ), .ZN(_07532_ ) );
AOI21_X1 _15569_ ( .A(_07379_ ), .B1(_07531_ ), .B2(_07532_ ), .ZN(_07533_ ) );
NOR3_X1 _15570_ ( .A1(_04084_ ), .A2(_04085_ ), .A3(_07251_ ), .ZN(_07534_ ) );
NAND3_X1 _15571_ ( .A1(_04176_ ), .A2(_02694_ ), .A3(_06889_ ), .ZN(_07535_ ) );
OAI21_X1 _15572_ ( .A(_07535_ ), .B1(_04085_ ), .B2(_04395_ ), .ZN(_07536_ ) );
OR4_X1 _15573_ ( .A1(_07530_ ), .A2(_07533_ ), .A3(_07534_ ), .A4(_07536_ ), .ZN(_07537_ ) );
OR3_X1 _15574_ ( .A1(_07517_ ), .A2(_07529_ ), .A3(_07537_ ), .ZN(_07538_ ) );
BUF_X4 _15575_ ( .A(_06899_ ), .Z(_07539_ ) );
AOI21_X1 _15576_ ( .A(_07511_ ), .B1(_07538_ ), .B2(_07539_ ), .ZN(_07540_ ) );
OAI21_X1 _15577_ ( .A(_07394_ ), .B1(_04755_ ), .B2(_05097_ ), .ZN(_07541_ ) );
OAI21_X1 _15578_ ( .A(_07500_ ), .B1(_07540_ ), .B2(_07541_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OR2_X1 _15579_ ( .A1(_04811_ ), .A2(_06258_ ), .ZN(_07542_ ) );
OR3_X1 _15580_ ( .A1(_07503_ ), .A2(_03887_ ), .A3(_04313_ ), .ZN(_07543_ ) );
NAND3_X1 _15581_ ( .A1(_07543_ ), .A2(_06594_ ), .A3(_07504_ ), .ZN(_07544_ ) );
AOI22_X1 _15582_ ( .A1(_04799_ ), .A2(_07217_ ), .B1(\ID_EX_imm [10] ), .B2(_07361_ ), .ZN(_07545_ ) );
AOI21_X1 _15583_ ( .A(_07017_ ), .B1(_07544_ ), .B2(_07545_ ), .ZN(_07546_ ) );
OR2_X1 _15584_ ( .A1(_07546_ ), .A2(_07364_ ), .ZN(_07547_ ) );
NAND2_X1 _15585_ ( .A1(_07058_ ), .A2(_07059_ ), .ZN(_07548_ ) );
AOI21_X1 _15586_ ( .A(_07548_ ), .B1(_06967_ ), .B2(_06838_ ), .ZN(_07549_ ) );
AND2_X1 _15587_ ( .A1(_07058_ ), .A2(_06735_ ), .ZN(_07550_ ) );
OAI21_X1 _15588_ ( .A(_07316_ ), .B1(_07549_ ), .B2(_07550_ ), .ZN(_07551_ ) );
OAI21_X1 _15589_ ( .A(_06991_ ), .B1(_07113_ ), .B2(_07116_ ), .ZN(_07552_ ) );
AND3_X1 _15590_ ( .A1(_07323_ ), .A2(_07324_ ), .A3(_06939_ ), .ZN(_07553_ ) );
OAI21_X1 _15591_ ( .A(_06771_ ), .B1(_06984_ ), .B2(_06988_ ), .ZN(_07554_ ) );
OAI21_X1 _15592_ ( .A(_06796_ ), .B1(_06963_ ), .B2(_06985_ ), .ZN(_07555_ ) );
AOI21_X1 _15593_ ( .A(_06809_ ), .B1(_07554_ ), .B2(_07555_ ), .ZN(_07556_ ) );
NOR2_X1 _15594_ ( .A1(_07553_ ), .A2(_07556_ ), .ZN(_07557_ ) );
OAI211_X1 _15595_ ( .A(_07006_ ), .B(_07552_ ), .C1(_07557_ ), .C2(_06822_ ), .ZN(_07558_ ) );
AOI21_X1 _15596_ ( .A(_06821_ ), .B1(_07106_ ), .B2(_07109_ ), .ZN(_07559_ ) );
NAND2_X1 _15597_ ( .A1(_07559_ ), .A2(_06866_ ), .ZN(_07560_ ) );
AND2_X1 _15598_ ( .A1(_07558_ ), .A2(_07560_ ), .ZN(_07561_ ) );
AOI21_X1 _15599_ ( .A(_06925_ ), .B1(_07551_ ), .B2(_07561_ ), .ZN(_07562_ ) );
AOI21_X1 _15600_ ( .A(_07237_ ), .B1(_07558_ ), .B2(_07560_ ), .ZN(_07563_ ) );
AND3_X1 _15601_ ( .A1(_07512_ ), .A2(_06644_ ), .A3(_06643_ ), .ZN(_07564_ ) );
OR3_X1 _15602_ ( .A1(_07564_ ), .A2(_07513_ ), .A3(_06606_ ), .ZN(_07565_ ) );
OR3_X1 _15603_ ( .A1(_04078_ ), .A2(_06646_ ), .A3(_07250_ ), .ZN(_07566_ ) );
AOI21_X1 _15604_ ( .A(_07009_ ), .B1(_04078_ ), .B2(_06646_ ), .ZN(_07567_ ) );
AOI21_X1 _15605_ ( .A(_07567_ ), .B1(_04079_ ), .B2(_06887_ ), .ZN(_07568_ ) );
NAND3_X1 _15606_ ( .A1(_07143_ ), .A2(_07147_ ), .A3(_06848_ ), .ZN(_07569_ ) );
OR3_X1 _15607_ ( .A1(_07127_ ), .A2(_07281_ ), .A3(_06982_ ), .ZN(_07570_ ) );
NAND2_X1 _15608_ ( .A1(_07569_ ), .A2(_07570_ ), .ZN(_07571_ ) );
NAND2_X1 _15609_ ( .A1(_07571_ ), .A2(_07298_ ), .ZN(_07572_ ) );
NAND4_X1 _15610_ ( .A1(_07565_ ), .A2(_07566_ ), .A3(_07568_ ), .A4(_07572_ ), .ZN(_07573_ ) );
OR3_X1 _15611_ ( .A1(_07562_ ), .A2(_07563_ ), .A3(_07573_ ), .ZN(_07574_ ) );
AOI21_X1 _15612_ ( .A(_07547_ ), .B1(_07574_ ), .B2(_07539_ ), .ZN(_07575_ ) );
NAND2_X1 _15613_ ( .A1(_04801_ ), .A2(_05029_ ), .ZN(_07576_ ) );
NAND2_X1 _15614_ ( .A1(_07576_ ), .A2(_06500_ ), .ZN(_07577_ ) );
OAI21_X1 _15615_ ( .A(_07542_ ), .B1(_07575_ ), .B2(_07577_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
OR2_X1 _15616_ ( .A1(_04832_ ), .A2(_06258_ ), .ZN(_07578_ ) );
AOI21_X1 _15617_ ( .A(_04310_ ), .B1(_04342_ ), .B2(_03932_ ), .ZN(_07579_ ) );
AOI21_X1 _15618_ ( .A(_07164_ ), .B1(_07579_ ), .B2(_07501_ ), .ZN(_07580_ ) );
OAI21_X1 _15619_ ( .A(_07580_ ), .B1(_07501_ ), .B2(_07579_ ), .ZN(_07581_ ) );
AOI22_X1 _15620_ ( .A1(_04819_ ), .A2(_07217_ ), .B1(\ID_EX_imm [9] ), .B2(_07361_ ), .ZN(_07582_ ) );
AOI21_X1 _15621_ ( .A(_07017_ ), .B1(_07581_ ), .B2(_07582_ ), .ZN(_07583_ ) );
OR2_X1 _15622_ ( .A1(_07583_ ), .A2(_07364_ ), .ZN(_07584_ ) );
NAND2_X1 _15623_ ( .A1(_07058_ ), .A2(_06735_ ), .ZN(_07585_ ) );
NAND3_X1 _15624_ ( .A1(_07058_ ), .A2(_06729_ ), .A3(_07059_ ), .ZN(_07586_ ) );
OAI21_X1 _15625_ ( .A(_07585_ ), .B1(_07586_ ), .B2(_06736_ ), .ZN(_07587_ ) );
NAND2_X1 _15626_ ( .A1(_07587_ ), .A2(_07316_ ), .ZN(_07588_ ) );
OR3_X1 _15627_ ( .A1(_07081_ ), .A2(_06796_ ), .A3(_06824_ ), .ZN(_07589_ ) );
NAND3_X1 _15628_ ( .A1(_06837_ ), .A2(_06842_ ), .A3(_06841_ ), .ZN(_07590_ ) );
AND3_X1 _15629_ ( .A1(_07589_ ), .A2(_06862_ ), .A3(_07590_ ), .ZN(_07591_ ) );
AOI21_X1 _15630_ ( .A(_06862_ ), .B1(_07369_ ), .B2(_07370_ ), .ZN(_07592_ ) );
OAI21_X1 _15631_ ( .A(_07281_ ), .B1(_07591_ ), .B2(_07592_ ), .ZN(_07593_ ) );
OAI211_X1 _15632_ ( .A(_07593_ ), .B(_06813_ ), .C1(_06848_ ), .C2(_07180_ ), .ZN(_07594_ ) );
NAND4_X1 _15633_ ( .A1(_07172_ ), .A2(_06819_ ), .A3(_07139_ ), .A4(_07174_ ), .ZN(_07595_ ) );
AND2_X1 _15634_ ( .A1(_07594_ ), .A2(_07595_ ), .ZN(_07596_ ) );
AOI21_X1 _15635_ ( .A(_06925_ ), .B1(_07588_ ), .B2(_07596_ ), .ZN(_07597_ ) );
AOI21_X1 _15636_ ( .A(_04103_ ), .B1(_06619_ ), .B2(_06635_ ), .ZN(_07598_ ) );
OR3_X1 _15637_ ( .A1(_07598_ ), .A2(_06611_ ), .A3(_06642_ ), .ZN(_07599_ ) );
OAI21_X1 _15638_ ( .A(_06611_ ), .B1(_07598_ ), .B2(_06642_ ), .ZN(_07600_ ) );
AND3_X1 _15639_ ( .A1(_07599_ ), .A2(_06605_ ), .A3(_07600_ ), .ZN(_07601_ ) );
AOI21_X1 _15640_ ( .A(_04395_ ), .B1(_04106_ ), .B2(_04107_ ), .ZN(_07602_ ) );
NAND3_X1 _15641_ ( .A1(_07198_ ), .A2(_06847_ ), .A3(_07199_ ), .ZN(_07603_ ) );
NAND4_X1 _15642_ ( .A1(_07064_ ), .A2(_07128_ ), .A3(_06878_ ), .A4(_06967_ ), .ZN(_07604_ ) );
NAND2_X1 _15643_ ( .A1(_07603_ ), .A2(_07604_ ), .ZN(_07605_ ) );
AOI221_X4 _15644_ ( .A(_07602_ ), .B1(_06611_ ), .B2(_04308_ ), .C1(_07605_ ), .C2(_07297_ ), .ZN(_07606_ ) );
OR3_X1 _15645_ ( .A1(_04106_ ), .A2(_04107_ ), .A3(_07250_ ), .ZN(_07607_ ) );
OAI211_X1 _15646_ ( .A(_07606_ ), .B(_07607_ ), .C1(_07237_ ), .C2(_07596_ ), .ZN(_07608_ ) );
OR3_X1 _15647_ ( .A1(_07597_ ), .A2(_07601_ ), .A3(_07608_ ), .ZN(_07609_ ) );
AOI21_X1 _15648_ ( .A(_07584_ ), .B1(_07609_ ), .B2(_07539_ ), .ZN(_07610_ ) );
NAND2_X1 _15649_ ( .A1(_04821_ ), .A2(_05029_ ), .ZN(_07611_ ) );
NAND2_X1 _15650_ ( .A1(_07611_ ), .A2(_06500_ ), .ZN(_07612_ ) );
OAI21_X1 _15651_ ( .A(_07578_ ), .B1(_07610_ ), .B2(_07612_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
AND4_X1 _15652_ ( .A1(_04851_ ), .A2(_04849_ ), .A3(_04847_ ), .A4(_04846_ ), .ZN(_07613_ ) );
NAND4_X1 _15653_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04588_ ), .A4(_07613_ ), .ZN(_07614_ ) );
NAND3_X1 _15654_ ( .A1(_06907_ ), .A2(_04854_ ), .A3(_06908_ ), .ZN(_07615_ ) );
NAND3_X1 _15655_ ( .A1(_07614_ ), .A2(_07615_ ), .A3(_06335_ ), .ZN(_07616_ ) );
AOI21_X1 _15656_ ( .A(_07164_ ), .B1(_04342_ ), .B2(_03932_ ), .ZN(_07617_ ) );
OAI21_X1 _15657_ ( .A(_07617_ ), .B1(_03932_ ), .B2(_04342_ ), .ZN(_07618_ ) );
AOI22_X1 _15658_ ( .A1(_04843_ ), .A2(_07217_ ), .B1(\ID_EX_imm [8] ), .B2(_07361_ ), .ZN(_07619_ ) );
AOI21_X1 _15659_ ( .A(_06600_ ), .B1(_07618_ ), .B2(_07619_ ), .ZN(_07620_ ) );
OR2_X1 _15660_ ( .A1(_07620_ ), .A2(_07364_ ), .ZN(_07621_ ) );
OAI211_X1 _15661_ ( .A(_07058_ ), .B(_07316_ ), .C1(_07337_ ), .C2(_06678_ ), .ZN(_07622_ ) );
OAI21_X1 _15662_ ( .A(_06820_ ), .B1(_07232_ ), .B2(_07337_ ), .ZN(_07623_ ) );
OAI21_X1 _15663_ ( .A(_06822_ ), .B1(_07226_ ), .B2(_07227_ ), .ZN(_07624_ ) );
AOI21_X1 _15664_ ( .A(_06620_ ), .B1(_07406_ ), .B2(_07407_ ), .ZN(_07625_ ) );
OAI21_X1 _15665_ ( .A(_06725_ ), .B1(_06987_ ), .B2(_06979_ ), .ZN(_07626_ ) );
OAI21_X1 _15666_ ( .A(_06781_ ), .B1(_06984_ ), .B2(_06988_ ), .ZN(_07627_ ) );
AND3_X1 _15667_ ( .A1(_07626_ ), .A2(_07627_ ), .A3(_06620_ ), .ZN(_07628_ ) );
OAI21_X1 _15668_ ( .A(_06848_ ), .B1(_07625_ ), .B2(_07628_ ), .ZN(_07629_ ) );
NAND3_X1 _15669_ ( .A1(_07624_ ), .A2(_07055_ ), .A3(_07629_ ), .ZN(_07630_ ) );
NAND2_X1 _15670_ ( .A1(_07623_ ), .A2(_07630_ ), .ZN(_07631_ ) );
AOI21_X1 _15671_ ( .A(_06925_ ), .B1(_07622_ ), .B2(_07631_ ), .ZN(_07632_ ) );
AND3_X1 _15672_ ( .A1(_07623_ ), .A2(_06885_ ), .A3(_07630_ ), .ZN(_07633_ ) );
NAND2_X1 _15673_ ( .A1(_07247_ ), .A2(_07282_ ), .ZN(_07634_ ) );
OR2_X1 _15674_ ( .A1(_07239_ ), .A2(_06848_ ), .ZN(_07635_ ) );
AND3_X1 _15675_ ( .A1(_07634_ ), .A2(_07298_ ), .A3(_07635_ ), .ZN(_07636_ ) );
NOR3_X1 _15676_ ( .A1(_07632_ ), .A2(_07633_ ), .A3(_07636_ ), .ZN(_07637_ ) );
AND3_X1 _15677_ ( .A1(_06619_ ), .A2(_04103_ ), .A3(_06635_ ), .ZN(_07638_ ) );
OR3_X1 _15678_ ( .A1(_07638_ ), .A2(_07598_ ), .A3(_06607_ ), .ZN(_07639_ ) );
AND2_X1 _15679_ ( .A1(_04102_ ), .A2(_07090_ ), .ZN(_07640_ ) );
NOR3_X1 _15680_ ( .A1(_04101_ ), .A2(_06412_ ), .A3(_07250_ ), .ZN(_07641_ ) );
AOI21_X1 _15681_ ( .A(_07102_ ), .B1(_04101_ ), .B2(_06412_ ), .ZN(_07642_ ) );
NOR3_X1 _15682_ ( .A1(_07640_ ), .A2(_07641_ ), .A3(_07642_ ), .ZN(_07643_ ) );
NAND3_X1 _15683_ ( .A1(_07637_ ), .A2(_07639_ ), .A3(_07643_ ), .ZN(_07644_ ) );
AOI21_X1 _15684_ ( .A(_07621_ ), .B1(_07644_ ), .B2(_07539_ ), .ZN(_07645_ ) );
OAI21_X1 _15685_ ( .A(_07394_ ), .B1(_04842_ ), .B2(_05097_ ), .ZN(_07646_ ) );
OAI21_X1 _15686_ ( .A(_07616_ ), .B1(_07645_ ), .B2(_07646_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
OAI21_X1 _15687_ ( .A(_06338_ ), .B1(_04872_ ), .B2(_04873_ ), .ZN(_07647_ ) );
AND4_X1 _15688_ ( .A1(_04334_ ), .A2(_04333_ ), .A3(_03727_ ), .A4(_03749_ ), .ZN(_07648_ ) );
NOR2_X1 _15689_ ( .A1(_07648_ ), .A2(_04339_ ), .ZN(_07649_ ) );
OR2_X1 _15690_ ( .A1(_07649_ ), .A2(_03703_ ), .ZN(_07650_ ) );
NAND2_X1 _15691_ ( .A1(_02890_ ), .A2(_03702_ ), .ZN(_07651_ ) );
AND3_X1 _15692_ ( .A1(_07650_ ), .A2(_03674_ ), .A3(_07651_ ), .ZN(_07652_ ) );
AOI21_X1 _15693_ ( .A(_03674_ ), .B1(_07650_ ), .B2(_07651_ ), .ZN(_07653_ ) );
OR3_X1 _15694_ ( .A1(_07652_ ), .A2(_07653_ ), .A3(_07163_ ), .ZN(_07654_ ) );
AOI22_X1 _15695_ ( .A1(_04861_ ), .A2(_07217_ ), .B1(\ID_EX_imm [7] ), .B2(_07361_ ), .ZN(_07655_ ) );
AOI21_X1 _15696_ ( .A(_06600_ ), .B1(_07654_ ), .B2(_07655_ ), .ZN(_07656_ ) );
OR2_X1 _15697_ ( .A1(_07656_ ), .A2(_07364_ ), .ZN(_07657_ ) );
NAND4_X1 _15698_ ( .A1(_06929_ ), .A2(_06675_ ), .A3(_06680_ ), .A4(_06736_ ), .ZN(_07658_ ) );
OR3_X1 _15699_ ( .A1(_06823_ ), .A2(_06796_ ), .A3(_06829_ ), .ZN(_07659_ ) );
OR3_X1 _15700_ ( .A1(_07081_ ), .A2(_06824_ ), .A3(_06726_ ), .ZN(_07660_ ) );
NAND2_X1 _15701_ ( .A1(_07659_ ), .A2(_07660_ ), .ZN(_07661_ ) );
BUF_X4 _15702_ ( .A(_06878_ ), .Z(_07662_ ) );
NAND2_X1 _15703_ ( .A1(_07661_ ), .A2(_07662_ ), .ZN(_07663_ ) );
OAI211_X1 _15704_ ( .A(_07663_ ), .B(_07282_ ), .C1(_07662_ ), .C2(_07523_ ), .ZN(_07664_ ) );
OAI211_X1 _15705_ ( .A(_07664_ ), .B(_06814_ ), .C1(_07287_ ), .C2(_07282_ ), .ZN(_07665_ ) );
NAND3_X1 _15706_ ( .A1(_07278_ ), .A2(_07279_ ), .A3(_07281_ ), .ZN(_07666_ ) );
NAND4_X1 _15707_ ( .A1(_06807_ ), .A2(_06821_ ), .A3(_07662_ ), .A4(_06967_ ), .ZN(_07667_ ) );
NAND2_X1 _15708_ ( .A1(_07666_ ), .A2(_07667_ ), .ZN(_07668_ ) );
NAND2_X1 _15709_ ( .A1(_07668_ ), .A2(_06820_ ), .ZN(_07669_ ) );
NAND3_X1 _15710_ ( .A1(_07658_ ), .A2(_07665_ ), .A3(_07669_ ), .ZN(_07670_ ) );
OAI21_X1 _15711_ ( .A(_07670_ ), .B1(_06676_ ), .B2(_06885_ ), .ZN(_07671_ ) );
NAND4_X1 _15712_ ( .A1(_06630_ ), .A2(_04126_ ), .A3(_06633_ ), .A4(_04162_ ), .ZN(_07672_ ) );
NAND2_X1 _15713_ ( .A1(_07672_ ), .A2(_06615_ ), .ZN(_07673_ ) );
NAND2_X1 _15714_ ( .A1(_07673_ ), .A2(_04133_ ), .ZN(_07674_ ) );
INV_X1 _15715_ ( .A(_06618_ ), .ZN(_07675_ ) );
AOI21_X1 _15716_ ( .A(_04117_ ), .B1(_07674_ ), .B2(_07675_ ), .ZN(_07676_ ) );
AOI211_X1 _15717_ ( .A(_04118_ ), .B(_06618_ ), .C1(_07673_ ), .C2(_04133_ ), .ZN(_07677_ ) );
OAI21_X1 _15718_ ( .A(_07035_ ), .B1(_07676_ ), .B2(_07677_ ), .ZN(_07678_ ) );
OR3_X1 _15719_ ( .A1(_04113_ ), .A2(_04114_ ), .A3(_07250_ ), .ZN(_07679_ ) );
OAI21_X1 _15720_ ( .A(_07679_ ), .B1(_04116_ ), .B2(_07102_ ), .ZN(_07680_ ) );
NOR3_X1 _15721_ ( .A1(_07292_ ), .A2(_07337_ ), .A3(_07379_ ), .ZN(_07681_ ) );
AOI211_X1 _15722_ ( .A(_07680_ ), .B(_07681_ ), .C1(_04117_ ), .C2(_07090_ ), .ZN(_07682_ ) );
NAND3_X1 _15723_ ( .A1(_07671_ ), .A2(_07678_ ), .A3(_07682_ ), .ZN(_07683_ ) );
AOI21_X1 _15724_ ( .A(_07657_ ), .B1(_07683_ ), .B2(_07539_ ), .ZN(_07684_ ) );
NAND2_X1 _15725_ ( .A1(_04863_ ), .A2(_05029_ ), .ZN(_07685_ ) );
NAND2_X1 _15726_ ( .A1(_07685_ ), .A2(_06500_ ), .ZN(_07686_ ) );
OAI21_X1 _15727_ ( .A(_07647_ ), .B1(_07684_ ), .B2(_07686_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
NOR2_X1 _15728_ ( .A1(_04884_ ), .A2(_04404_ ), .ZN(_07687_ ) );
NAND4_X1 _15729_ ( .A1(_06723_ ), .A2(_06735_ ), .A3(_07038_ ), .A4(_07317_ ), .ZN(_07688_ ) );
MUX2_X1 _15730_ ( .A(_07329_ ), .B(_07321_ ), .S(_06846_ ), .Z(_07689_ ) );
NAND2_X1 _15731_ ( .A1(_07689_ ), .A2(_06818_ ), .ZN(_07690_ ) );
NAND3_X1 _15732_ ( .A1(_07554_ ), .A2(_07555_ ), .A3(_06730_ ), .ZN(_07691_ ) );
OAI21_X1 _15733_ ( .A(_06854_ ), .B1(_06978_ ), .B2(_06976_ ), .ZN(_07692_ ) );
OAI21_X1 _15734_ ( .A(_06796_ ), .B1(_06987_ ), .B2(_06979_ ), .ZN(_07693_ ) );
NAND2_X1 _15735_ ( .A1(_07692_ ), .A2(_07693_ ), .ZN(_07694_ ) );
OAI211_X1 _15736_ ( .A(_07691_ ), .B(_06846_ ), .C1(_07694_ ), .C2(_06939_ ), .ZN(_07695_ ) );
OAI211_X1 _15737_ ( .A(_06812_ ), .B(_07695_ ), .C1(_07326_ ), .C2(_06937_ ), .ZN(_07696_ ) );
AND2_X1 _15738_ ( .A1(_07690_ ), .A2(_07696_ ), .ZN(_07697_ ) );
AOI21_X1 _15739_ ( .A(_06924_ ), .B1(_07688_ ), .B2(_07697_ ), .ZN(_07698_ ) );
AOI21_X1 _15740_ ( .A(_07237_ ), .B1(_07690_ ), .B2(_07696_ ), .ZN(_07699_ ) );
AOI21_X1 _15741_ ( .A(_07009_ ), .B1(_04121_ ), .B2(_02918_ ), .ZN(_07700_ ) );
OR3_X1 _15742_ ( .A1(_07336_ ), .A2(_06631_ ), .A3(_07379_ ), .ZN(_07701_ ) );
OAI221_X1 _15743_ ( .A(_07701_ ), .B1(_07675_ ), .B2(_04032_ ), .C1(_06616_ ), .C2(_07251_ ), .ZN(_07702_ ) );
OR4_X1 _15744_ ( .A1(_07698_ ), .A2(_07699_ ), .A3(_07700_ ), .A4(_07702_ ), .ZN(_07703_ ) );
NAND3_X1 _15745_ ( .A1(_07672_ ), .A2(_06616_ ), .A3(_06615_ ), .ZN(_07704_ ) );
AND3_X1 _15746_ ( .A1(_07674_ ), .A2(_06605_ ), .A3(_07704_ ), .ZN(_07705_ ) );
OAI21_X1 _15747_ ( .A(_06899_ ), .B1(_07703_ ), .B2(_07705_ ), .ZN(_07706_ ) );
NAND2_X1 _15748_ ( .A1(_07649_ ), .A2(_03703_ ), .ZN(_07707_ ) );
NAND3_X1 _15749_ ( .A1(_07650_ ), .A2(_06594_ ), .A3(_07707_ ), .ZN(_07708_ ) );
AOI22_X1 _15750_ ( .A1(_04886_ ), .A2(_06580_ ), .B1(\ID_EX_imm [6] ), .B2(_06583_ ), .ZN(_07709_ ) );
AOI21_X1 _15751_ ( .A(_06600_ ), .B1(_07708_ ), .B2(_07709_ ), .ZN(_07710_ ) );
NOR2_X1 _15752_ ( .A1(_07710_ ), .A2(_04487_ ), .ZN(_07711_ ) );
AOI21_X1 _15753_ ( .A(_07687_ ), .B1(_07706_ ), .B2(_07711_ ), .ZN(_07712_ ) );
MUX2_X1 _15754_ ( .A(_04898_ ), .B(_07712_ ), .S(_06266_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
AND2_X1 _15755_ ( .A1(_04906_ ), .A2(_04487_ ), .ZN(_07713_ ) );
NAND4_X1 _15756_ ( .A1(_07058_ ), .A2(_06732_ ), .A3(_06736_ ), .A4(_07316_ ), .ZN(_07714_ ) );
AND2_X1 _15757_ ( .A1(_06811_ ), .A2(_06819_ ), .ZN(_07715_ ) );
AOI21_X1 _15758_ ( .A(_06862_ ), .B1(_07589_ ), .B2(_07590_ ), .ZN(_07716_ ) );
NOR3_X1 _15759_ ( .A1(_06828_ ), .A2(_06842_ ), .A3(_06872_ ), .ZN(_07717_ ) );
NOR3_X1 _15760_ ( .A1(_06823_ ), .A2(_06829_ ), .A3(_06727_ ), .ZN(_07718_ ) );
NOR2_X1 _15761_ ( .A1(_07717_ ), .A2(_07718_ ), .ZN(_07719_ ) );
INV_X1 _15762_ ( .A(_07719_ ), .ZN(_07720_ ) );
AOI211_X1 _15763_ ( .A(_06821_ ), .B(_07716_ ), .C1(_07720_ ), .C2(_07662_ ), .ZN(_07721_ ) );
AND3_X1 _15764_ ( .A1(_07368_ ), .A2(_07371_ ), .A3(_07128_ ), .ZN(_07722_ ) );
NOR3_X1 _15765_ ( .A1(_07721_ ), .A2(_06819_ ), .A3(_07722_ ), .ZN(_07723_ ) );
NOR2_X1 _15766_ ( .A1(_07715_ ), .A2(_07723_ ), .ZN(_07724_ ) );
AOI21_X1 _15767_ ( .A(_06925_ ), .B1(_07714_ ), .B2(_07724_ ), .ZN(_07725_ ) );
NAND2_X1 _15768_ ( .A1(_06630_ ), .A2(_06633_ ), .ZN(_07726_ ) );
NOR2_X1 _15769_ ( .A1(_07726_ ), .A2(_04163_ ), .ZN(_07727_ ) );
OR3_X1 _15770_ ( .A1(_07727_ ), .A2(_04126_ ), .A3(_04160_ ), .ZN(_07728_ ) );
OAI21_X1 _15771_ ( .A(_04126_ ), .B1(_07727_ ), .B2(_04160_ ), .ZN(_07729_ ) );
NAND3_X1 _15772_ ( .A1(_07728_ ), .A2(_06605_ ), .A3(_07729_ ), .ZN(_07730_ ) );
OAI21_X1 _15773_ ( .A(_06884_ ), .B1(_07715_ ), .B2(_07723_ ), .ZN(_07731_ ) );
NAND3_X1 _15774_ ( .A1(_04125_ ), .A2(_02867_ ), .A3(_06890_ ), .ZN(_07732_ ) );
AOI21_X1 _15775_ ( .A(_04395_ ), .B1(_06683_ ), .B2(_02923_ ), .ZN(_07733_ ) );
NAND4_X1 _15776_ ( .A1(_06870_ ), .A2(_06879_ ), .A3(_07005_ ), .A4(_07281_ ), .ZN(_07734_ ) );
NOR2_X1 _15777_ ( .A1(_07734_ ), .A2(_07062_ ), .ZN(_07735_ ) );
AOI211_X1 _15778_ ( .A(_07733_ ), .B(_07735_ ), .C1(_04126_ ), .C2(_06887_ ), .ZN(_07736_ ) );
NAND4_X1 _15779_ ( .A1(_07730_ ), .A2(_07731_ ), .A3(_07732_ ), .A4(_07736_ ), .ZN(_07737_ ) );
OAI21_X1 _15780_ ( .A(_06899_ ), .B1(_07725_ ), .B2(_07737_ ), .ZN(_07738_ ) );
AND3_X1 _15781_ ( .A1(_04333_ ), .A2(_04334_ ), .A3(_03727_ ), .ZN(_07739_ ) );
OR3_X1 _15782_ ( .A1(_07739_ ), .A2(_04337_ ), .A3(_03749_ ), .ZN(_07740_ ) );
OAI21_X1 _15783_ ( .A(_03749_ ), .B1(_07739_ ), .B2(_04337_ ), .ZN(_07741_ ) );
NAND3_X1 _15784_ ( .A1(_07740_ ), .A2(_06594_ ), .A3(_07741_ ), .ZN(_07742_ ) );
AOI22_X1 _15785_ ( .A1(_04904_ ), .A2(_06580_ ), .B1(\ID_EX_imm [5] ), .B2(_06583_ ), .ZN(_07743_ ) );
AOI21_X1 _15786_ ( .A(_06600_ ), .B1(_07742_ ), .B2(_07743_ ), .ZN(_07744_ ) );
NOR2_X1 _15787_ ( .A1(_07744_ ), .A2(_04487_ ), .ZN(_07745_ ) );
AOI21_X1 _15788_ ( .A(_07713_ ), .B1(_07738_ ), .B2(_07745_ ), .ZN(_07746_ ) );
MUX2_X1 _15789_ ( .A(_04917_ ), .B(_07746_ ), .S(_06266_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
NOR2_X1 _15790_ ( .A1(_04923_ ), .A2(_04404_ ), .ZN(_07747_ ) );
NAND4_X1 _15791_ ( .A1(_06724_ ), .A2(_06736_ ), .A3(_06927_ ), .A4(_07316_ ), .ZN(_07748_ ) );
OR3_X1 _15792_ ( .A1(_06975_ ), .A2(_06781_ ), .A3(_07001_ ), .ZN(_07749_ ) );
OR3_X1 _15793_ ( .A1(_06978_ ), .A2(_06976_ ), .A3(_04146_ ), .ZN(_07750_ ) );
AOI21_X1 _15794_ ( .A(_06982_ ), .B1(_07749_ ), .B2(_07750_ ), .ZN(_07751_ ) );
AND3_X1 _15795_ ( .A1(_07626_ ), .A2(_07627_ ), .A3(_06731_ ), .ZN(_07752_ ) );
NOR3_X1 _15796_ ( .A1(_07751_ ), .A2(_06991_ ), .A3(_07752_ ), .ZN(_07753_ ) );
AOI21_X1 _15797_ ( .A(_07281_ ), .B1(_07408_ ), .B2(_07409_ ), .ZN(_07754_ ) );
NOR3_X1 _15798_ ( .A1(_07753_ ), .A2(_07754_ ), .A3(_06866_ ), .ZN(_07755_ ) );
AOI21_X1 _15799_ ( .A(_07006_ ), .B1(_06938_ ), .B2(_06954_ ), .ZN(_07756_ ) );
NOR2_X1 _15800_ ( .A1(_07755_ ), .A2(_07756_ ), .ZN(_07757_ ) );
AOI21_X1 _15801_ ( .A(_06925_ ), .B1(_07748_ ), .B2(_07757_ ), .ZN(_07758_ ) );
AOI21_X1 _15802_ ( .A(_06606_ ), .B1(_07726_ ), .B2(_04163_ ), .ZN(_07759_ ) );
OAI21_X1 _15803_ ( .A(_07759_ ), .B1(_04163_ ), .B2(_07726_ ), .ZN(_07760_ ) );
OAI21_X1 _15804_ ( .A(_06884_ ), .B1(_07755_ ), .B2(_07756_ ), .ZN(_07761_ ) );
NOR3_X1 _15805_ ( .A1(_07004_ ), .A2(_06822_ ), .A3(_07379_ ), .ZN(_07762_ ) );
NOR3_X1 _15806_ ( .A1(_04160_ ), .A2(_04161_ ), .A3(_07251_ ), .ZN(_07763_ ) );
NOR3_X1 _15807_ ( .A1(_06813_ ), .A2(_04159_ ), .A3(_04032_ ), .ZN(_07764_ ) );
AOI21_X1 _15808_ ( .A(_04395_ ), .B1(_06813_ ), .B2(_04159_ ), .ZN(_07765_ ) );
NOR4_X1 _15809_ ( .A1(_07762_ ), .A2(_07763_ ), .A3(_07764_ ), .A4(_07765_ ), .ZN(_07766_ ) );
NAND3_X1 _15810_ ( .A1(_07760_ ), .A2(_07761_ ), .A3(_07766_ ), .ZN(_07767_ ) );
OAI21_X1 _15811_ ( .A(_06899_ ), .B1(_07758_ ), .B2(_07767_ ), .ZN(_07768_ ) );
AOI21_X1 _15812_ ( .A(_03727_ ), .B1(_04333_ ), .B2(_04334_ ), .ZN(_07769_ ) );
OR3_X1 _15813_ ( .A1(_07739_ ), .A2(_07769_ ), .A3(_07163_ ), .ZN(_07770_ ) );
AOI22_X1 _15814_ ( .A1(_04925_ ), .A2(_06580_ ), .B1(\ID_EX_imm [4] ), .B2(_06583_ ), .ZN(_07771_ ) );
AOI21_X1 _15815_ ( .A(_06600_ ), .B1(_07770_ ), .B2(_07771_ ), .ZN(_07772_ ) );
NOR2_X1 _15816_ ( .A1(_07772_ ), .A2(_04487_ ), .ZN(_07773_ ) );
AOI21_X1 _15817_ ( .A(_07747_ ), .B1(_07768_ ), .B2(_07773_ ), .ZN(_07774_ ) );
MUX2_X1 _15818_ ( .A(_04936_ ), .B(_07774_ ), .S(_06258_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
NAND3_X1 _15819_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_04952_ ), .ZN(_07775_ ) );
INV_X1 _15820_ ( .A(_04946_ ), .ZN(_07776_ ) );
NAND3_X1 _15821_ ( .A1(_07775_ ), .A2(_07776_ ), .A3(_06335_ ), .ZN(_07777_ ) );
NAND4_X1 _15822_ ( .A1(_07058_ ), .A2(_06736_ ), .A3(_07059_ ), .A4(_07316_ ), .ZN(_07778_ ) );
NAND2_X1 _15823_ ( .A1(_07054_ ), .A2(_06866_ ), .ZN(_07779_ ) );
AOI21_X1 _15824_ ( .A(_06833_ ), .B1(_07659_ ), .B2(_07660_ ), .ZN(_07780_ ) );
NOR2_X1 _15825_ ( .A1(_06871_ ), .A2(_06875_ ), .ZN(_07781_ ) );
NOR2_X1 _15826_ ( .A1(_06828_ ), .A2(_06872_ ), .ZN(_07782_ ) );
MUX2_X1 _15827_ ( .A(_07781_ ), .B(_07782_ ), .S(_06842_ ), .Z(_07783_ ) );
AOI211_X1 _15828_ ( .A(_07128_ ), .B(_07780_ ), .C1(_06834_ ), .C2(_07783_ ), .ZN(_07784_ ) );
AOI21_X1 _15829_ ( .A(_06847_ ), .B1(_07520_ ), .B2(_07524_ ), .ZN(_07785_ ) );
OR3_X1 _15830_ ( .A1(_07784_ ), .A2(_06819_ ), .A3(_07785_ ), .ZN(_07786_ ) );
AND2_X1 _15831_ ( .A1(_07779_ ), .A2(_07786_ ), .ZN(_07787_ ) );
AOI21_X1 _15832_ ( .A(_06925_ ), .B1(_07778_ ), .B2(_07787_ ), .ZN(_07788_ ) );
INV_X1 _15833_ ( .A(_06627_ ), .ZN(_07789_ ) );
INV_X1 _15834_ ( .A(_04148_ ), .ZN(_07790_ ) );
AOI21_X1 _15835_ ( .A(_06629_ ), .B1(_07789_ ), .B2(_07790_ ), .ZN(_07791_ ) );
OAI21_X1 _15836_ ( .A(_04139_ ), .B1(_07791_ ), .B2(_06621_ ), .ZN(_07792_ ) );
AND2_X1 _15837_ ( .A1(_07792_ ), .A2(_06605_ ), .ZN(_07793_ ) );
INV_X1 _15838_ ( .A(_07791_ ), .ZN(_07794_ ) );
AOI21_X1 _15839_ ( .A(_06606_ ), .B1(_07794_ ), .B2(_06622_ ), .ZN(_07795_ ) );
OAI22_X1 _15840_ ( .A1(_07793_ ), .A2(_07090_ ), .B1(_04139_ ), .B2(_07795_ ), .ZN(_07796_ ) );
AND3_X1 _15841_ ( .A1(_06991_ ), .A2(_02815_ ), .A3(_06889_ ), .ZN(_07797_ ) );
NOR2_X1 _15842_ ( .A1(_07067_ ), .A2(_07379_ ), .ZN(_07798_ ) );
AOI211_X1 _15843_ ( .A(_07797_ ), .B(_07798_ ), .C1(_06633_ ), .C2(_04394_ ), .ZN(_07799_ ) );
OAI211_X1 _15844_ ( .A(_07796_ ), .B(_07799_ ), .C1(_07787_ ), .C2(_07237_ ), .ZN(_07800_ ) );
OAI21_X1 _15845_ ( .A(_06899_ ), .B1(_07788_ ), .B2(_07800_ ), .ZN(_07801_ ) );
INV_X1 _15846_ ( .A(_03979_ ), .ZN(_07802_ ) );
AND3_X1 _15847_ ( .A1(_04330_ ), .A2(_07802_ ), .A3(_04332_ ), .ZN(_07803_ ) );
AOI21_X1 _15848_ ( .A(_07802_ ), .B1(_04330_ ), .B2(_04332_ ), .ZN(_07804_ ) );
NOR3_X1 _15849_ ( .A1(_07803_ ), .A2(_07804_ ), .A3(_07164_ ), .ZN(_07805_ ) );
NAND2_X1 _15850_ ( .A1(_04942_ ), .A2(_06915_ ), .ZN(_07806_ ) );
NAND3_X1 _15851_ ( .A1(_06582_ ), .A2(\ID_EX_imm [3] ), .A3(_06578_ ), .ZN(_07807_ ) );
NAND2_X1 _15852_ ( .A1(_07806_ ), .A2(_07807_ ), .ZN(_07808_ ) );
OAI21_X1 _15853_ ( .A(_06598_ ), .B1(_07805_ ), .B2(_07808_ ), .ZN(_07809_ ) );
AND3_X1 _15854_ ( .A1(_07801_ ), .A2(_07168_ ), .A3(_07809_ ), .ZN(_07810_ ) );
OAI21_X1 _15855_ ( .A(_07394_ ), .B1(_04406_ ), .B2(_04940_ ), .ZN(_07811_ ) );
OAI21_X1 _15856_ ( .A(_07777_ ), .B1(_07810_ ), .B2(_07811_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
OR2_X1 _15857_ ( .A1(_04969_ ), .A2(_06258_ ), .ZN(_07812_ ) );
AOI21_X1 _15858_ ( .A(_07164_ ), .B1(_04329_ ), .B2(_03957_ ), .ZN(_07813_ ) );
OAI21_X1 _15859_ ( .A(_07813_ ), .B1(_03957_ ), .B2(_04329_ ), .ZN(_07814_ ) );
AOI22_X1 _15860_ ( .A1(_04958_ ), .A2(_06580_ ), .B1(\ID_EX_imm [2] ), .B2(_07361_ ), .ZN(_07815_ ) );
AOI21_X1 _15861_ ( .A(_06600_ ), .B1(_07814_ ), .B2(_07815_ ), .ZN(_07816_ ) );
OR2_X1 _15862_ ( .A1(_07816_ ), .A2(_07364_ ), .ZN(_07817_ ) );
OR2_X1 _15863_ ( .A1(_07118_ ), .A2(_07005_ ), .ZN(_07818_ ) );
OAI21_X1 _15864_ ( .A(_06842_ ), .B1(_06975_ ), .B2(_07001_ ), .ZN(_07819_ ) );
NOR2_X1 _15865_ ( .A1(_07000_ ), .A2(_06998_ ), .ZN(_07820_ ) );
OAI211_X1 _15866_ ( .A(_07819_ ), .B(_06862_ ), .C1(_06926_ ), .C2(_07820_ ), .ZN(_07821_ ) );
OAI211_X1 _15867_ ( .A(_07821_ ), .B(_06847_ ), .C1(_06834_ ), .C2(_07694_ ), .ZN(_07822_ ) );
OAI211_X1 _15868_ ( .A(_06813_ ), .B(_07822_ ), .C1(_07557_ ), .C2(_07139_ ), .ZN(_07823_ ) );
AOI21_X1 _15869_ ( .A(_07237_ ), .B1(_07818_ ), .B2(_07823_ ), .ZN(_07824_ ) );
OAI211_X1 _15870_ ( .A(_07122_ ), .B(_07316_ ), .C1(_06926_ ), .C2(_06728_ ), .ZN(_07825_ ) );
NAND3_X1 _15871_ ( .A1(_07825_ ), .A2(_07823_ ), .A3(_07818_ ), .ZN(_07826_ ) );
AOI221_X4 _15872_ ( .A(_07824_ ), .B1(_07129_ ), .B2(_07297_ ), .C1(_07826_ ), .C2(_06675_ ), .ZN(_07827_ ) );
AOI21_X1 _15873_ ( .A(_06607_ ), .B1(_06628_ ), .B2(_06629_ ), .ZN(_07828_ ) );
NAND2_X1 _15874_ ( .A1(_07794_ ), .A2(_07828_ ), .ZN(_07829_ ) );
AOI21_X1 _15875_ ( .A(_07009_ ), .B1(_07662_ ), .B2(_02793_ ), .ZN(_07830_ ) );
AOI221_X4 _15876_ ( .A(_07830_ ), .B1(_06621_ ), .B2(_06889_ ), .C1(_04143_ ), .C2(_06887_ ), .ZN(_07831_ ) );
NAND3_X1 _15877_ ( .A1(_07827_ ), .A2(_07829_ ), .A3(_07831_ ), .ZN(_07832_ ) );
AOI21_X1 _15878_ ( .A(_07817_ ), .B1(_07832_ ), .B2(_07539_ ), .ZN(_07833_ ) );
OAI21_X1 _15879_ ( .A(_07394_ ), .B1(_04406_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07834_ ) );
OAI21_X1 _15880_ ( .A(_07812_ ), .B1(_07833_ ), .B2(_07834_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
INV_X1 _15881_ ( .A(_04499_ ), .ZN(_07835_ ) );
AND4_X1 _15882_ ( .A1(_04490_ ), .A2(_04495_ ), .A3(_04492_ ), .A4(_07835_ ), .ZN(_07836_ ) );
NAND3_X1 _15883_ ( .A1(_04724_ ), .A2(_04725_ ), .A3(_07836_ ), .ZN(_07837_ ) );
NAND3_X1 _15884_ ( .A1(_06907_ ), .A2(_04512_ ), .A3(_06908_ ), .ZN(_07838_ ) );
NAND3_X1 _15885_ ( .A1(_07837_ ), .A2(_07838_ ), .A3(_06335_ ), .ZN(_07839_ ) );
OR3_X1 _15886_ ( .A1(_07434_ ), .A2(_04380_ ), .A3(_03602_ ), .ZN(_07840_ ) );
OAI21_X1 _15887_ ( .A(_03602_ ), .B1(_07434_ ), .B2(_04380_ ), .ZN(_07841_ ) );
NAND3_X1 _15888_ ( .A1(_07840_ ), .A2(_06595_ ), .A3(_07841_ ), .ZN(_07842_ ) );
AOI22_X1 _15889_ ( .A1(_04532_ ), .A2(_06915_ ), .B1(\ID_EX_imm [29] ), .B2(_06916_ ), .ZN(_07843_ ) );
AOI21_X1 _15890_ ( .A(_06601_ ), .B1(_07842_ ), .B2(_07843_ ), .ZN(_07844_ ) );
OR2_X1 _15891_ ( .A1(_07844_ ), .A2(_06919_ ), .ZN(_07845_ ) );
OR3_X1 _15892_ ( .A1(_07461_ ), .A2(_04286_ ), .A3(_07462_ ), .ZN(_07846_ ) );
OAI21_X1 _15893_ ( .A(_04286_ ), .B1(_07461_ ), .B2(_07462_ ), .ZN(_07847_ ) );
AOI21_X1 _15894_ ( .A(_06607_ ), .B1(_07846_ ), .B2(_07847_ ), .ZN(_07848_ ) );
OAI21_X1 _15895_ ( .A(_06727_ ), .B1(_06783_ ), .B2(_06793_ ), .ZN(_07849_ ) );
OAI21_X1 _15896_ ( .A(_06842_ ), .B1(_06774_ ), .B2(_06788_ ), .ZN(_07850_ ) );
AND3_X1 _15897_ ( .A1(_07849_ ), .A2(_07850_ ), .A3(_06731_ ), .ZN(_07851_ ) );
AOI21_X1 _15898_ ( .A(_02992_ ), .B1(_06785_ ), .B2(_06787_ ), .ZN(_07852_ ) );
NOR2_X1 _15899_ ( .A1(_06797_ ), .A2(_07852_ ), .ZN(_07853_ ) );
NOR2_X1 _15900_ ( .A1(_06792_ ), .A2(_06798_ ), .ZN(_07854_ ) );
MUX2_X1 _15901_ ( .A(_07853_ ), .B(_07854_ ), .S(_06926_ ), .Z(_07855_ ) );
AOI211_X1 _15902_ ( .A(_06821_ ), .B(_07851_ ), .C1(_07662_ ), .C2(_07855_ ), .ZN(_07856_ ) );
NOR3_X1 _15903_ ( .A1(_06856_ ), .A2(_06863_ ), .A3(_07139_ ), .ZN(_07857_ ) );
OAI21_X1 _15904_ ( .A(_07006_ ), .B1(_07856_ ), .B2(_07857_ ), .ZN(_07858_ ) );
NAND3_X1 _15905_ ( .A1(_07380_ ), .A2(_06866_ ), .A3(_07381_ ), .ZN(_07859_ ) );
AND3_X1 _15906_ ( .A1(_07858_ ), .A2(_06817_ ), .A3(_07859_ ), .ZN(_07860_ ) );
AND3_X1 _15907_ ( .A1(_04284_ ), .A2(_02992_ ), .A3(_06889_ ), .ZN(_07861_ ) );
NAND3_X1 _15908_ ( .A1(_07374_ ), .A2(_07006_ ), .A3(_06884_ ), .ZN(_07862_ ) );
OAI221_X1 _15909_ ( .A(_07862_ ), .B1(_04297_ ), .B2(_07009_ ), .C1(_04286_ ), .C2(_07251_ ), .ZN(_07863_ ) );
NOR4_X1 _15910_ ( .A1(_07848_ ), .A2(_07860_ ), .A3(_07861_ ), .A4(_07863_ ), .ZN(_07864_ ) );
OAI21_X1 _15911_ ( .A(_07058_ ), .B1(_06732_ ), .B2(_06735_ ), .ZN(_07865_ ) );
NOR2_X1 _15912_ ( .A1(_07865_ ), .A2(_06768_ ), .ZN(_07866_ ) );
AND2_X1 _15913_ ( .A1(_07374_ ), .A2(_07006_ ), .ZN(_07867_ ) );
OR3_X1 _15914_ ( .A1(_07866_ ), .A2(_07039_ ), .A3(_07867_ ), .ZN(_07868_ ) );
NAND2_X1 _15915_ ( .A1(_07868_ ), .A2(_06676_ ), .ZN(_07869_ ) );
AOI21_X1 _15916_ ( .A(_06898_ ), .B1(_07864_ ), .B2(_07869_ ), .ZN(_07870_ ) );
OAI22_X1 _15917_ ( .A1(_07845_ ), .A2(_07870_ ), .B1(_07168_ ), .B2(_04528_ ), .ZN(_07871_ ) );
OAI21_X1 _15918_ ( .A(_07839_ ), .B1(_07871_ ), .B2(_06491_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
AND2_X1 _15919_ ( .A1(_04981_ ), .A2(_04983_ ), .ZN(_07872_ ) );
AND2_X1 _15920_ ( .A1(_04982_ ), .A2(_04984_ ), .ZN(_07873_ ) );
AOI22_X1 _15921_ ( .A1(_07872_ ), .A2(_07873_ ), .B1(_06907_ ), .B2(_06908_ ), .ZN(_07874_ ) );
OAI21_X1 _15922_ ( .A(_06910_ ), .B1(_07874_ ), .B2(_04979_ ), .ZN(_07875_ ) );
OAI21_X1 _15923_ ( .A(_06594_ ), .B1(_04003_ ), .B2(_04328_ ), .ZN(_07876_ ) );
AOI21_X1 _15924_ ( .A(_07876_ ), .B1(_04328_ ), .B2(_04003_ ), .ZN(_07877_ ) );
AND2_X1 _15925_ ( .A1(_04975_ ), .A2(_06915_ ), .ZN(_07878_ ) );
AND3_X1 _15926_ ( .A1(_06582_ ), .A2(\ID_EX_imm [1] ), .A3(_06578_ ), .ZN(_07879_ ) );
NOR3_X1 _15927_ ( .A1(_07877_ ), .A2(_07878_ ), .A3(_07879_ ), .ZN(_07880_ ) );
OAI21_X1 _15928_ ( .A(_04405_ ), .B1(_07880_ ), .B2(_06601_ ), .ZN(_07881_ ) );
OAI21_X1 _15929_ ( .A(_06822_ ), .B1(_07591_ ), .B2(_07592_ ), .ZN(_07882_ ) );
NOR2_X1 _15930_ ( .A1(_06874_ ), .A2(_06868_ ), .ZN(_07883_ ) );
MUX2_X1 _15931_ ( .A(_07883_ ), .B(_07781_ ), .S(_06926_ ), .Z(_07884_ ) );
MUX2_X1 _15932_ ( .A(_07884_ ), .B(_07720_ ), .S(_06982_ ), .Z(_07885_ ) );
OAI211_X1 _15933_ ( .A(_07055_ ), .B(_07882_ ), .C1(_07885_ ), .C2(_07337_ ), .ZN(_07886_ ) );
NAND2_X1 _15934_ ( .A1(_07202_ ), .A2(_06820_ ), .ZN(_07887_ ) );
AOI21_X1 _15935_ ( .A(_07237_ ), .B1(_07886_ ), .B2(_07887_ ), .ZN(_07888_ ) );
AND4_X1 _15936_ ( .A1(_07055_ ), .A2(_07191_ ), .A3(_07282_ ), .A4(_06817_ ), .ZN(_07889_ ) );
AND3_X1 _15937_ ( .A1(_06724_ ), .A2(_06735_ ), .A3(_07059_ ), .ZN(_07890_ ) );
NAND4_X1 _15938_ ( .A1(_07890_ ), .A2(_06680_ ), .A3(_06729_ ), .A4(_06765_ ), .ZN(_07891_ ) );
NAND3_X1 _15939_ ( .A1(_07891_ ), .A2(_07886_ ), .A3(_07887_ ), .ZN(_07892_ ) );
AOI211_X1 _15940_ ( .A(_07888_ ), .B(_07889_ ), .C1(_07892_ ), .C2(_06676_ ), .ZN(_07893_ ) );
AOI21_X1 _15941_ ( .A(_06607_ ), .B1(_06624_ ), .B2(_06626_ ), .ZN(_07894_ ) );
OAI21_X1 _15942_ ( .A(_07894_ ), .B1(_06624_ ), .B2(_06626_ ), .ZN(_07895_ ) );
OAI22_X1 _15943_ ( .A1(_07790_ ), .A2(_07250_ ), .B1(_04149_ ), .B2(_07102_ ), .ZN(_07896_ ) );
AOI21_X1 _15944_ ( .A(_07896_ ), .B1(_06624_ ), .B2(_07090_ ), .ZN(_07897_ ) );
NAND3_X1 _15945_ ( .A1(_07893_ ), .A2(_07895_ ), .A3(_07897_ ), .ZN(_07898_ ) );
AOI21_X1 _15946_ ( .A(_07881_ ), .B1(_07898_ ), .B2(_07539_ ), .ZN(_07899_ ) );
OAI21_X1 _15947_ ( .A(_07394_ ), .B1(_04406_ ), .B2(\ID_EX_pc [1] ), .ZN(_07900_ ) );
OAI21_X1 _15948_ ( .A(_07875_ ), .B1(_07899_ ), .B2(_07900_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
AND3_X1 _15949_ ( .A1(_04030_ ), .A2(_06895_ ), .A3(_04049_ ), .ZN(_07901_ ) );
AND4_X1 _15950_ ( .A1(\ID_EX_typ [4] ), .A2(_03224_ ), .A3(\ID_EX_typ [3] ), .A4(_05194_ ), .ZN(_07902_ ) );
OAI21_X1 _15951_ ( .A(_04391_ ), .B1(_07901_ ), .B2(_07902_ ), .ZN(_07903_ ) );
NAND2_X1 _15952_ ( .A1(_04026_ ), .A2(_06594_ ), .ZN(_07904_ ) );
NAND2_X1 _15953_ ( .A1(_07903_ ), .A2(_07904_ ), .ZN(_07905_ ) );
AND3_X1 _15954_ ( .A1(_05013_ ), .A2(_06578_ ), .A3(_06577_ ), .ZN(_07906_ ) );
AND3_X1 _15955_ ( .A1(_06582_ ), .A2(\ID_EX_imm [0] ), .A3(_06578_ ), .ZN(_07907_ ) );
OR2_X1 _15956_ ( .A1(_07906_ ), .A2(_07907_ ), .ZN(_07908_ ) );
OAI21_X1 _15957_ ( .A(_06598_ ), .B1(_07905_ ), .B2(_07908_ ), .ZN(_07909_ ) );
INV_X1 _15958_ ( .A(_04294_ ), .ZN(_07910_ ) );
AOI21_X1 _15959_ ( .A(_04305_ ), .B1(_04276_ ), .B2(_03025_ ), .ZN(_07911_ ) );
NAND3_X1 _15960_ ( .A1(_07910_ ), .A2(_04302_ ), .A3(_07911_ ), .ZN(_07912_ ) );
AND3_X1 _15961_ ( .A1(_06723_ ), .A2(_04125_ ), .A3(_06682_ ), .ZN(_07913_ ) );
NOR2_X1 _15962_ ( .A1(_07233_ ), .A2(_06812_ ), .ZN(_07914_ ) );
AND2_X1 _15963_ ( .A1(_06728_ ), .A2(_06625_ ), .ZN(_07915_ ) );
NOR3_X1 _15964_ ( .A1(_07915_ ), .A2(_06997_ ), .A3(_06795_ ), .ZN(_07916_ ) );
AOI211_X1 _15965_ ( .A(_04156_ ), .B(_07916_ ), .C1(_06806_ ), .C2(_07820_ ), .ZN(_07917_ ) );
AND3_X1 _15966_ ( .A1(_07749_ ), .A2(_04156_ ), .A3(_07750_ ), .ZN(_07918_ ) );
OAI21_X1 _15967_ ( .A(_06846_ ), .B1(_07917_ ), .B2(_07918_ ), .ZN(_07919_ ) );
OR3_X1 _15968_ ( .A1(_07625_ ), .A2(_06846_ ), .A3(_07628_ ), .ZN(_07920_ ) );
AOI21_X1 _15969_ ( .A(_06818_ ), .B1(_07919_ ), .B2(_07920_ ), .ZN(_07921_ ) );
NOR2_X1 _15970_ ( .A1(_07914_ ), .A2(_07921_ ), .ZN(_07922_ ) );
OAI21_X1 _15971_ ( .A(_06675_ ), .B1(_07913_ ), .B2(_07922_ ), .ZN(_07923_ ) );
NAND2_X1 _15972_ ( .A1(_07922_ ), .A2(_06884_ ), .ZN(_07924_ ) );
NAND4_X1 _15973_ ( .A1(_07239_ ), .A2(_06813_ ), .A3(_07139_ ), .A4(_06817_ ), .ZN(_07925_ ) );
NAND4_X1 _15974_ ( .A1(_07912_ ), .A2(_07923_ ), .A3(_07924_ ), .A4(_07925_ ), .ZN(_07926_ ) );
NOR3_X1 _15975_ ( .A1(_07915_ ), .A2(_06626_ ), .A3(_06606_ ), .ZN(_07927_ ) );
OAI21_X1 _15976_ ( .A(_06887_ ), .B1(_06867_ ), .B2(_06994_ ), .ZN(_07928_ ) );
NAND3_X1 _15977_ ( .A1(_06838_ ), .A2(_04004_ ), .A3(_06889_ ), .ZN(_07929_ ) );
OAI211_X1 _15978_ ( .A(_07928_ ), .B(_07929_ ), .C1(_07009_ ), .C2(_07915_ ), .ZN(_07930_ ) );
NOR3_X1 _15979_ ( .A1(_07926_ ), .A2(_07927_ ), .A3(_07930_ ), .ZN(_07931_ ) );
OAI21_X1 _15980_ ( .A(_07909_ ), .B1(_07931_ ), .B2(_06898_ ), .ZN(_07932_ ) );
MUX2_X1 _15981_ ( .A(\ID_EX_pc [0] ), .B(_07932_ ), .S(_04404_ ), .Z(_07933_ ) );
MUX2_X1 _15982_ ( .A(_06497_ ), .B(_07933_ ), .S(_06258_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
NAND3_X1 _15983_ ( .A1(_04792_ ), .A2(_04794_ ), .A3(_06335_ ), .ZN(_07934_ ) );
AND3_X1 _15984_ ( .A1(_06723_ ), .A2(_06733_ ), .A3(_06927_ ), .ZN(_07935_ ) );
OAI21_X1 _15985_ ( .A(_07935_ ), .B1(_06929_ ), .B2(_06767_ ), .ZN(_07936_ ) );
NOR4_X1 _15986_ ( .A1(_06753_ ), .A2(_06733_ ), .A3(_06763_ ), .A4(_06768_ ), .ZN(_07937_ ) );
NOR2_X1 _15987_ ( .A1(_07039_ ), .A2(_07937_ ), .ZN(_07938_ ) );
OAI211_X1 _15988_ ( .A(_07936_ ), .B(_07938_ ), .C1(_06866_ ), .C2(_07403_ ), .ZN(_07939_ ) );
NAND2_X1 _15989_ ( .A1(_07939_ ), .A2(_06675_ ), .ZN(_07940_ ) );
OR3_X1 _15990_ ( .A1(_07403_ ), .A2(_06866_ ), .A3(_07237_ ), .ZN(_07941_ ) );
OAI21_X1 _15991_ ( .A(_06822_ ), .B1(_06966_ ), .B2(_06973_ ), .ZN(_07942_ ) );
NAND2_X1 _15992_ ( .A1(_07488_ ), .A2(_06967_ ), .ZN(_07943_ ) );
OR3_X1 _15993_ ( .A1(_06947_ ), .A2(_06951_ ), .A3(_06727_ ), .ZN(_07944_ ) );
NAND3_X1 _15994_ ( .A1(_07943_ ), .A2(_07944_ ), .A3(_06834_ ), .ZN(_07945_ ) );
OAI21_X1 _15995_ ( .A(_06967_ ), .B1(_06943_ ), .B2(_06948_ ), .ZN(_07946_ ) );
OAI21_X1 _15996_ ( .A(_06926_ ), .B1(_06940_ ), .B2(_06944_ ), .ZN(_07947_ ) );
AND2_X1 _15997_ ( .A1(_07946_ ), .A2(_07947_ ), .ZN(_07948_ ) );
OAI211_X1 _15998_ ( .A(_07945_ ), .B(_07139_ ), .C1(_07662_ ), .C2(_07948_ ), .ZN(_07949_ ) );
AND3_X1 _15999_ ( .A1(_07942_ ), .A2(_07055_ ), .A3(_07949_ ), .ZN(_07950_ ) );
OAI21_X1 _16000_ ( .A(_06817_ ), .B1(_07419_ ), .B2(_07055_ ), .ZN(_07951_ ) );
OAI211_X1 _16001_ ( .A(_07940_ ), .B(_07941_ ), .C1(_07950_ ), .C2(_07951_ ), .ZN(_07952_ ) );
AND2_X1 _16002_ ( .A1(_04291_ ), .A2(_06887_ ), .ZN(_07953_ ) );
AND3_X1 _16003_ ( .A1(_04289_ ), .A2(_02224_ ), .A3(_06890_ ), .ZN(_07954_ ) );
AOI21_X1 _16004_ ( .A(_07102_ ), .B1(_04295_ ), .B2(_04290_ ), .ZN(_07955_ ) );
NOR4_X1 _16005_ ( .A1(_07952_ ), .A2(_07953_ ), .A3(_07954_ ), .A4(_07955_ ), .ZN(_07956_ ) );
AND3_X1 _16006_ ( .A1(_07455_ ), .A2(_04292_ ), .A3(_07460_ ), .ZN(_07957_ ) );
OR3_X1 _16007_ ( .A1(_07957_ ), .A2(_07461_ ), .A3(_06607_ ), .ZN(_07958_ ) );
AOI21_X1 _16008_ ( .A(_06898_ ), .B1(_07956_ ), .B2(_07958_ ), .ZN(_07959_ ) );
NAND3_X1 _16009_ ( .A1(_07431_ ), .A2(_07433_ ), .A3(_04374_ ), .ZN(_07960_ ) );
NAND3_X1 _16010_ ( .A1(_07435_ ), .A2(_06595_ ), .A3(_07960_ ), .ZN(_07961_ ) );
AOI22_X1 _16011_ ( .A1(_04783_ ), .A2(_06915_ ), .B1(\ID_EX_imm [28] ), .B2(_06916_ ), .ZN(_07962_ ) );
AOI21_X1 _16012_ ( .A(_06601_ ), .B1(_07961_ ), .B2(_07962_ ), .ZN(_07963_ ) );
OR2_X1 _16013_ ( .A1(_07963_ ), .A2(_06919_ ), .ZN(_07964_ ) );
OAI22_X1 _16014_ ( .A1(_07959_ ), .A2(_07964_ ), .B1(_07168_ ), .B2(_04782_ ), .ZN(_07965_ ) );
OAI21_X1 _16015_ ( .A(_07934_ ), .B1(_07965_ ), .B2(_06491_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND3_X1 _16016_ ( .A1(_05005_ ), .A2(_05007_ ), .A3(_06335_ ), .ZN(_07966_ ) );
OAI22_X1 _16017_ ( .A1(_04997_ ), .A2(_06581_ ), .B1(_02227_ ), .B2(_06584_ ), .ZN(_07967_ ) );
NOR2_X1 _16018_ ( .A1(_04347_ ), .A2(_04366_ ), .ZN(_07968_ ) );
INV_X1 _16019_ ( .A(_03533_ ), .ZN(_07969_ ) );
NOR2_X1 _16020_ ( .A1(_07968_ ), .A2(_07969_ ), .ZN(_07970_ ) );
NOR3_X1 _16021_ ( .A1(_07970_ ), .A2(_04369_ ), .A3(_04368_ ), .ZN(_07971_ ) );
AOI21_X1 _16022_ ( .A(_07971_ ), .B1(_04056_ ), .B2(_03555_ ), .ZN(_07972_ ) );
AND2_X1 _16023_ ( .A1(_07972_ ), .A2(_03477_ ), .ZN(_07973_ ) );
AOI21_X1 _16024_ ( .A(_07973_ ), .B1(_02271_ ), .B2(_04372_ ), .ZN(_07974_ ) );
NAND2_X1 _16025_ ( .A1(_03500_ ), .A2(_03502_ ), .ZN(_07975_ ) );
OR2_X1 _16026_ ( .A1(_07974_ ), .A2(_07975_ ), .ZN(_07976_ ) );
AOI21_X1 _16027_ ( .A(_07164_ ), .B1(_07974_ ), .B2(_07975_ ), .ZN(_07977_ ) );
AOI21_X1 _16028_ ( .A(_07967_ ), .B1(_07976_ ), .B2(_07977_ ), .ZN(_07978_ ) );
OAI21_X1 _16029_ ( .A(_04405_ ), .B1(_07978_ ), .B2(_06601_ ), .ZN(_07979_ ) );
NOR2_X1 _16030_ ( .A1(_07446_ ), .A2(_07454_ ), .ZN(_07980_ ) );
NOR3_X1 _16031_ ( .A1(_07980_ ), .A2(_04260_ ), .A3(_04265_ ), .ZN(_07981_ ) );
OAI21_X1 _16032_ ( .A(_04039_ ), .B1(_07981_ ), .B2(_07459_ ), .ZN(_07982_ ) );
INV_X1 _16033_ ( .A(_07982_ ), .ZN(_07983_ ) );
OAI21_X1 _16034_ ( .A(_04046_ ), .B1(_07983_ ), .B2(_04037_ ), .ZN(_07984_ ) );
OAI211_X1 _16035_ ( .A(_07982_ ), .B(_04062_ ), .C1(_04036_ ), .C2(_04035_ ), .ZN(_07985_ ) );
NAND3_X1 _16036_ ( .A1(_07984_ ), .A2(_07035_ ), .A3(_07985_ ), .ZN(_07986_ ) );
OAI211_X1 _16037_ ( .A(_07058_ ), .B(_07059_ ), .C1(_06765_ ), .C2(_06767_ ), .ZN(_07987_ ) );
INV_X1 _16038_ ( .A(_07987_ ), .ZN(_07988_ ) );
NOR2_X1 _16039_ ( .A1(_07053_ ), .A2(_06822_ ), .ZN(_07989_ ) );
AND2_X1 _16040_ ( .A1(_07989_ ), .A2(_07055_ ), .ZN(_07990_ ) );
OR2_X1 _16041_ ( .A1(_07988_ ), .A2(_07990_ ), .ZN(_07991_ ) );
OAI21_X1 _16042_ ( .A(_06676_ ), .B1(_07991_ ), .B2(_07475_ ), .ZN(_07992_ ) );
AND2_X1 _16043_ ( .A1(_04045_ ), .A2(_04064_ ), .ZN(_07993_ ) );
OAI22_X1 _16044_ ( .A1(_04062_ ), .A2(_07251_ ), .B1(_07993_ ), .B2(_07009_ ), .ZN(_07994_ ) );
INV_X1 _16045_ ( .A(_07477_ ), .ZN(_07995_ ) );
AOI21_X1 _16046_ ( .A(_07995_ ), .B1(_07531_ ), .B2(_07532_ ), .ZN(_07996_ ) );
AOI211_X1 _16047_ ( .A(_07994_ ), .B(_07996_ ), .C1(_07456_ ), .C2(_06890_ ), .ZN(_07997_ ) );
NAND2_X1 _16048_ ( .A1(_07854_ ), .A2(_06854_ ), .ZN(_07998_ ) );
OR3_X1 _16049_ ( .A1(_06783_ ), .A2(_06793_ ), .A3(_06770_ ), .ZN(_07999_ ) );
NAND2_X1 _16050_ ( .A1(_07998_ ), .A2(_07999_ ), .ZN(_08000_ ) );
NOR3_X1 _16051_ ( .A1(_06774_ ), .A2(_06806_ ), .A3(_06788_ ), .ZN(_08001_ ) );
NOR3_X1 _16052_ ( .A1(_06857_ ), .A2(_06779_ ), .A3(_06771_ ), .ZN(_08002_ ) );
OR2_X1 _16053_ ( .A1(_08001_ ), .A2(_08002_ ), .ZN(_08003_ ) );
MUX2_X1 _16054_ ( .A(_08000_ ), .B(_08003_ ), .S(_06982_ ), .Z(_08004_ ) );
MUX2_X1 _16055_ ( .A(_07077_ ), .B(_08004_ ), .S(_06848_ ), .Z(_08005_ ) );
NAND2_X1 _16056_ ( .A1(_08005_ ), .A2(_07298_ ), .ZN(_08006_ ) );
NAND3_X1 _16057_ ( .A1(_07989_ ), .A2(_06814_ ), .A3(_06885_ ), .ZN(_08007_ ) );
AND3_X1 _16058_ ( .A1(_07997_ ), .A2(_08006_ ), .A3(_08007_ ), .ZN(_08008_ ) );
NAND3_X1 _16059_ ( .A1(_07986_ ), .A2(_07992_ ), .A3(_08008_ ), .ZN(_08009_ ) );
AOI21_X1 _16060_ ( .A(_07979_ ), .B1(_08009_ ), .B2(_07539_ ), .ZN(_08010_ ) );
OAI21_X1 _16061_ ( .A(_07394_ ), .B1(_04992_ ), .B2(_05097_ ), .ZN(_08011_ ) );
OAI21_X1 _16062_ ( .A(_07966_ ), .B1(_08010_ ), .B2(_08011_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
AND2_X1 _16063_ ( .A1(_05037_ ), .A2(_05039_ ), .ZN(_00304_ ) );
AND2_X1 _16064_ ( .A1(_05038_ ), .A2(_05040_ ), .ZN(_00305_ ) );
AOI22_X1 _16065_ ( .A1(_00304_ ), .A2(_00305_ ), .B1(_06907_ ), .B2(_06908_ ), .ZN(_00306_ ) );
AND3_X1 _16066_ ( .A1(_06907_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_06908_ ), .ZN(_00307_ ) );
OAI21_X1 _16067_ ( .A(_06910_ ), .B1(_00306_ ), .B2(_00307_ ), .ZN(_00308_ ) );
AOI21_X1 _16068_ ( .A(_07164_ ), .B1(_07972_ ), .B2(_03477_ ), .ZN(_00309_ ) );
OAI21_X1 _16069_ ( .A(_00309_ ), .B1(_03477_ ), .B2(_07972_ ), .ZN(_00310_ ) );
AOI22_X1 _16070_ ( .A1(_05033_ ), .A2(_06580_ ), .B1(\ID_EX_imm [26] ), .B2(_07361_ ), .ZN(_00311_ ) );
AOI21_X1 _16071_ ( .A(_06600_ ), .B1(_00310_ ), .B2(_00311_ ), .ZN(_00312_ ) );
OR2_X1 _16072_ ( .A1(_00312_ ), .A2(_07364_ ), .ZN(_00313_ ) );
AND2_X1 _16073_ ( .A1(_06723_ ), .A2(_07059_ ), .ZN(_00314_ ) );
OAI21_X1 _16074_ ( .A(_00314_ ), .B1(_06926_ ), .B2(_06728_ ), .ZN(_00315_ ) );
NOR2_X1 _16075_ ( .A1(_00315_ ), .A2(_07121_ ), .ZN(_00316_ ) );
NOR4_X1 _16076_ ( .A1(_06710_ ), .A2(_06733_ ), .A3(_06722_ ), .A4(_06768_ ), .ZN(_00317_ ) );
INV_X1 _16077_ ( .A(_00317_ ), .ZN(_00318_ ) );
NAND2_X1 _16078_ ( .A1(_07559_ ), .A2(_07006_ ), .ZN(_00319_ ) );
INV_X1 _16079_ ( .A(_06929_ ), .ZN(_00320_ ) );
OAI211_X1 _16080_ ( .A(_00318_ ), .B(_00319_ ), .C1(_00320_ ), .C2(_06681_ ), .ZN(_00321_ ) );
OAI21_X1 _16081_ ( .A(_06675_ ), .B1(_00316_ ), .B2(_00321_ ), .ZN(_00322_ ) );
NAND2_X1 _16082_ ( .A1(_07571_ ), .A2(_07477_ ), .ZN(_00323_ ) );
NAND3_X1 _16083_ ( .A1(_07484_ ), .A2(_07485_ ), .A3(_07662_ ), .ZN(_00324_ ) );
NAND3_X1 _16084_ ( .A1(_07480_ ), .A2(_07481_ ), .A3(_06982_ ), .ZN(_00325_ ) );
NAND3_X1 _16085_ ( .A1(_00324_ ), .A2(_00325_ ), .A3(_07282_ ), .ZN(_00326_ ) );
OAI211_X1 _16086_ ( .A(_07298_ ), .B(_00326_ ), .C1(_07138_ ), .C2(_07282_ ), .ZN(_00327_ ) );
NAND3_X1 _16087_ ( .A1(_07559_ ), .A2(_06814_ ), .A3(_06885_ ), .ZN(_00328_ ) );
AND4_X1 _16088_ ( .A1(_00322_ ), .A2(_00323_ ), .A3(_00327_ ), .A4(_00328_ ), .ZN(_00329_ ) );
OR3_X1 _16089_ ( .A1(_07981_ ), .A2(_04039_ ), .A3(_07459_ ), .ZN(_00330_ ) );
NAND3_X1 _16090_ ( .A1(_00330_ ), .A2(_07035_ ), .A3(_07982_ ), .ZN(_00331_ ) );
NOR3_X1 _16091_ ( .A1(_04037_ ), .A2(_04038_ ), .A3(_07251_ ), .ZN(_00332_ ) );
AOI21_X1 _16092_ ( .A(_07102_ ), .B1(_04035_ ), .B2(_04036_ ), .ZN(_00333_ ) );
NOR3_X1 _16093_ ( .A1(_04035_ ), .A2(_04036_ ), .A3(_07250_ ), .ZN(_00334_ ) );
NOR3_X1 _16094_ ( .A1(_00332_ ), .A2(_00333_ ), .A3(_00334_ ), .ZN(_00335_ ) );
NAND3_X1 _16095_ ( .A1(_00329_ ), .A2(_00331_ ), .A3(_00335_ ), .ZN(_00336_ ) );
AOI21_X1 _16096_ ( .A(_00313_ ), .B1(_00336_ ), .B2(_07539_ ), .ZN(_00337_ ) );
OAI21_X1 _16097_ ( .A(_07394_ ), .B1(_05032_ ), .B2(_05097_ ), .ZN(_00338_ ) );
OAI21_X1 _16098_ ( .A(_00308_ ), .B1(_00337_ ), .B2(_00338_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _16099_ ( .A1(_05065_ ), .A2(_06292_ ), .ZN(_00339_ ) );
OR3_X1 _16100_ ( .A1(_07970_ ), .A2(_04369_ ), .A3(_03556_ ), .ZN(_00340_ ) );
OAI21_X1 _16101_ ( .A(_03556_ ), .B1(_07970_ ), .B2(_04369_ ), .ZN(_00341_ ) );
AND3_X1 _16102_ ( .A1(_00340_ ), .A2(_06594_ ), .A3(_00341_ ), .ZN(_00342_ ) );
OAI22_X1 _16103_ ( .A1(_05056_ ), .A2(_06581_ ), .B1(_02321_ ), .B2(_06584_ ), .ZN(_00343_ ) );
OAI21_X1 _16104_ ( .A(_06598_ ), .B1(_00342_ ), .B2(_00343_ ), .ZN(_00344_ ) );
NAND2_X1 _16105_ ( .A1(_00344_ ), .A2(_07168_ ), .ZN(_00345_ ) );
OAI21_X1 _16106_ ( .A(_04264_ ), .B1(_07446_ ), .B2(_07454_ ), .ZN(_00346_ ) );
INV_X1 _16107_ ( .A(_04262_ ), .ZN(_00347_ ) );
AND3_X1 _16108_ ( .A1(_00346_ ), .A2(_04259_ ), .A3(_00347_ ), .ZN(_00348_ ) );
AOI21_X1 _16109_ ( .A(_04259_ ), .B1(_00346_ ), .B2(_00347_ ), .ZN(_00349_ ) );
OAI21_X1 _16110_ ( .A(_07035_ ), .B1(_00348_ ), .B2(_00349_ ), .ZN(_00350_ ) );
NAND3_X1 _16111_ ( .A1(_00314_ ), .A2(_06729_ ), .A3(_06733_ ), .ZN(_00351_ ) );
NOR2_X1 _16112_ ( .A1(_00351_ ), .A2(_07121_ ), .ZN(_00352_ ) );
AND3_X1 _16113_ ( .A1(_07172_ ), .A2(_07281_ ), .A3(_07174_ ), .ZN(_00353_ ) );
AND2_X1 _16114_ ( .A1(_00353_ ), .A2(_07006_ ), .ZN(_00354_ ) );
OR3_X1 _16115_ ( .A1(_07039_ ), .A2(_07937_ ), .A3(_00354_ ), .ZN(_00355_ ) );
OAI21_X1 _16116_ ( .A(_06676_ ), .B1(_00352_ ), .B2(_00355_ ), .ZN(_00356_ ) );
OAI22_X1 _16117_ ( .A1(_04260_ ), .A2(_04309_ ), .B1(_04057_ ), .B2(_04395_ ), .ZN(_00357_ ) );
AOI221_X4 _16118_ ( .A(_00357_ ), .B1(_04058_ ), .B2(_06889_ ), .C1(_07605_ ), .C2(_07477_ ), .ZN(_00358_ ) );
AND2_X1 _16119_ ( .A1(_07196_ ), .A2(_07337_ ), .ZN(_00359_ ) );
AOI21_X1 _16120_ ( .A(_06982_ ), .B1(_07849_ ), .B2(_07850_ ), .ZN(_00360_ ) );
AOI21_X1 _16121_ ( .A(_07662_ ), .B1(_06858_ ), .B2(_06861_ ), .ZN(_00361_ ) );
NOR3_X1 _16122_ ( .A1(_00360_ ), .A2(_00361_ ), .A3(_07337_ ), .ZN(_00362_ ) );
OAI21_X1 _16123_ ( .A(_07298_ ), .B1(_00359_ ), .B2(_00362_ ), .ZN(_00363_ ) );
NAND3_X1 _16124_ ( .A1(_00353_ ), .A2(_06814_ ), .A3(_06885_ ), .ZN(_00364_ ) );
AND3_X1 _16125_ ( .A1(_00358_ ), .A2(_00363_ ), .A3(_00364_ ), .ZN(_00365_ ) );
NAND3_X1 _16126_ ( .A1(_00350_ ), .A2(_00356_ ), .A3(_00365_ ), .ZN(_00366_ ) );
AOI21_X1 _16127_ ( .A(_00345_ ), .B1(_00366_ ), .B2(_07539_ ), .ZN(_00367_ ) );
OAI21_X1 _16128_ ( .A(_07394_ ), .B1(_05052_ ), .B2(_07168_ ), .ZN(_00368_ ) );
OAI21_X1 _16129_ ( .A(_00339_ ), .B1(_00367_ ), .B2(_00368_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND3_X1 _16130_ ( .A1(_06538_ ), .A2(_06539_ ), .A3(_06335_ ), .ZN(_00369_ ) );
OAI21_X1 _16131_ ( .A(_06594_ ), .B1(_07968_ ), .B2(_07969_ ), .ZN(_00370_ ) );
AOI21_X1 _16132_ ( .A(_00370_ ), .B1(_07969_ ), .B2(_07968_ ), .ZN(_00371_ ) );
AND2_X1 _16133_ ( .A1(_05071_ ), .A2(_06915_ ), .ZN(_00372_ ) );
AND3_X1 _16134_ ( .A1(_06582_ ), .A2(\ID_EX_imm [24] ), .A3(_06578_ ), .ZN(_00373_ ) );
NOR3_X1 _16135_ ( .A1(_00371_ ), .A2(_00372_ ), .A3(_00373_ ), .ZN(_00374_ ) );
OAI21_X1 _16136_ ( .A(_04405_ ), .B1(_00374_ ), .B2(_06601_ ), .ZN(_00375_ ) );
OAI211_X1 _16137_ ( .A(_06724_ ), .B(_06767_ ), .C1(_06822_ ), .C2(_06678_ ), .ZN(_00376_ ) );
AND3_X1 _16138_ ( .A1(_07229_ ), .A2(_07281_ ), .A3(_07231_ ), .ZN(_00377_ ) );
NAND2_X1 _16139_ ( .A1(_00377_ ), .A2(_07055_ ), .ZN(_00378_ ) );
NAND3_X1 _16140_ ( .A1(_00376_ ), .A2(_07474_ ), .A3(_00378_ ), .ZN(_00379_ ) );
NAND3_X1 _16141_ ( .A1(_00379_ ), .A2(\ID_EX_typ [2] ), .A3(_04307_ ), .ZN(_00380_ ) );
OR3_X1 _16142_ ( .A1(_07242_ ), .A2(_07243_ ), .A3(_06848_ ), .ZN(_00381_ ) );
AOI21_X1 _16143_ ( .A(_07662_ ), .B1(_06969_ ), .B2(_06972_ ), .ZN(_00382_ ) );
AOI21_X1 _16144_ ( .A(_06982_ ), .B1(_07946_ ), .B2(_07947_ ), .ZN(_00383_ ) );
OAI21_X1 _16145_ ( .A(_07282_ ), .B1(_00382_ ), .B2(_00383_ ), .ZN(_00384_ ) );
NAND3_X1 _16146_ ( .A1(_00381_ ), .A2(_07298_ ), .A3(_00384_ ), .ZN(_00385_ ) );
NAND3_X1 _16147_ ( .A1(_07634_ ), .A2(_07477_ ), .A3(_07635_ ), .ZN(_00386_ ) );
NAND3_X1 _16148_ ( .A1(_00377_ ), .A2(_06814_ ), .A3(_06885_ ), .ZN(_00387_ ) );
AND4_X1 _16149_ ( .A1(_00380_ ), .A2(_00385_ ), .A3(_00386_ ), .A4(_00387_ ), .ZN(_00388_ ) );
AOI21_X1 _16150_ ( .A(_06607_ ), .B1(_07980_ ), .B2(_04265_ ), .ZN(_00389_ ) );
NAND2_X1 _16151_ ( .A1(_00389_ ), .A2(_00346_ ), .ZN(_00390_ ) );
NOR3_X1 _16152_ ( .A1(_04262_ ), .A2(_04263_ ), .A3(_07251_ ), .ZN(_00391_ ) );
NOR3_X1 _16153_ ( .A1(_04052_ ), .A2(_04261_ ), .A3(_07250_ ), .ZN(_00392_ ) );
AOI21_X1 _16154_ ( .A(_07102_ ), .B1(_04052_ ), .B2(_04261_ ), .ZN(_00393_ ) );
NOR3_X1 _16155_ ( .A1(_00391_ ), .A2(_00392_ ), .A3(_00393_ ), .ZN(_00394_ ) );
NAND3_X1 _16156_ ( .A1(_00388_ ), .A2(_00390_ ), .A3(_00394_ ), .ZN(_00395_ ) );
AOI21_X1 _16157_ ( .A(_00375_ ), .B1(_00395_ ), .B2(_06899_ ), .ZN(_00396_ ) );
NAND2_X1 _16158_ ( .A1(_05073_ ), .A2(_06919_ ), .ZN(_00397_ ) );
NAND2_X1 _16159_ ( .A1(_00397_ ), .A2(_06500_ ), .ZN(_00398_ ) );
OAI21_X1 _16160_ ( .A(_00369_ ), .B1(_00396_ ), .B2(_00398_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
AND2_X1 _16161_ ( .A1(_05099_ ), .A2(_05101_ ), .ZN(_00399_ ) );
AND2_X1 _16162_ ( .A1(_05100_ ), .A2(_05102_ ), .ZN(_00400_ ) );
AOI22_X1 _16163_ ( .A1(_00399_ ), .A2(_00400_ ), .B1(_06907_ ), .B2(_06908_ ), .ZN(_00401_ ) );
AND3_X1 _16164_ ( .A1(_04429_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_04439_ ), .ZN(_00402_ ) );
OAI21_X1 _16165_ ( .A(_06910_ ), .B1(_00401_ ), .B2(_00402_ ), .ZN(_00403_ ) );
OAI22_X1 _16166_ ( .A1(_05095_ ), .A2(_06581_ ), .B1(_02407_ ), .B2(_06584_ ), .ZN(_00404_ ) );
AOI21_X1 _16167_ ( .A(_03450_ ), .B1(_06912_ ), .B2(_04359_ ), .ZN(_00405_ ) );
AOI21_X1 _16168_ ( .A(_04362_ ), .B1(_00405_ ), .B2(_03404_ ), .ZN(_00406_ ) );
XNOR2_X1 _16169_ ( .A(_00406_ ), .B(_03382_ ), .ZN(_00407_ ) );
AOI21_X1 _16170_ ( .A(_00404_ ), .B1(_00407_ ), .B2(_06595_ ), .ZN(_00408_ ) );
OAI21_X1 _16171_ ( .A(_04405_ ), .B1(_00408_ ), .B2(_06601_ ), .ZN(_00409_ ) );
OR3_X1 _16172_ ( .A1(_06921_ ), .A2(_04204_ ), .A3(_04210_ ), .ZN(_00410_ ) );
AOI21_X1 _16173_ ( .A(_07450_ ), .B1(_00410_ ), .B2(_07448_ ), .ZN(_00411_ ) );
INV_X1 _16174_ ( .A(_00411_ ), .ZN(_00412_ ) );
NOR2_X1 _16175_ ( .A1(_04190_ ), .A2(_04248_ ), .ZN(_00413_ ) );
INV_X1 _16176_ ( .A(_00413_ ), .ZN(_00414_ ) );
NAND3_X1 _16177_ ( .A1(_00412_ ), .A2(_07449_ ), .A3(_00414_ ), .ZN(_00415_ ) );
OAI21_X1 _16178_ ( .A(_04198_ ), .B1(_00411_ ), .B2(_00413_ ), .ZN(_00416_ ) );
NAND3_X1 _16179_ ( .A1(_00415_ ), .A2(_07035_ ), .A3(_00416_ ), .ZN(_00417_ ) );
NOR3_X1 _16180_ ( .A1(_04196_ ), .A2(_04197_ ), .A3(_07251_ ), .ZN(_00418_ ) );
NOR3_X1 _16181_ ( .A1(_04194_ ), .A2(_04195_ ), .A3(_07250_ ), .ZN(_00419_ ) );
AOI21_X1 _16182_ ( .A(_07102_ ), .B1(_04194_ ), .B2(_04195_ ), .ZN(_00420_ ) );
NOR3_X1 _16183_ ( .A1(_00418_ ), .A2(_00419_ ), .A3(_00420_ ), .ZN(_00421_ ) );
AND2_X1 _16184_ ( .A1(_07668_ ), .A2(_07055_ ), .ZN(_00422_ ) );
OAI21_X1 _16185_ ( .A(_06675_ ), .B1(_07475_ ), .B2(_00422_ ), .ZN(_00423_ ) );
NOR3_X1 _16186_ ( .A1(_08001_ ), .A2(_08002_ ), .A3(_06939_ ), .ZN(_00424_ ) );
AOI21_X1 _16187_ ( .A(_06833_ ), .B1(_07069_ ), .B2(_07071_ ), .ZN(_00425_ ) );
OR3_X1 _16188_ ( .A1(_00424_ ), .A2(_06991_ ), .A3(_00425_ ), .ZN(_00426_ ) );
OR3_X1 _16189_ ( .A1(_07294_ ), .A2(_07295_ ), .A3(_07139_ ), .ZN(_00427_ ) );
NAND3_X1 _16190_ ( .A1(_00426_ ), .A2(_06814_ ), .A3(_00427_ ), .ZN(_00428_ ) );
OAI21_X1 _16191_ ( .A(_06820_ ), .B1(_07292_ ), .B2(_07337_ ), .ZN(_00429_ ) );
NAND3_X1 _16192_ ( .A1(_00428_ ), .A2(_06817_ ), .A3(_00429_ ), .ZN(_00430_ ) );
NAND3_X1 _16193_ ( .A1(_07668_ ), .A2(_06814_ ), .A3(_06885_ ), .ZN(_00431_ ) );
AND3_X1 _16194_ ( .A1(_00423_ ), .A2(_00430_ ), .A3(_00431_ ), .ZN(_00432_ ) );
NAND3_X1 _16195_ ( .A1(_00417_ ), .A2(_00421_ ), .A3(_00432_ ), .ZN(_00433_ ) );
AOI21_X1 _16196_ ( .A(_00409_ ), .B1(_00433_ ), .B2(_06899_ ), .ZN(_00434_ ) );
OAI21_X1 _16197_ ( .A(_06266_ ), .B1(_05088_ ), .B2(_07168_ ), .ZN(_00435_ ) );
OAI21_X1 _16198_ ( .A(_00403_ ), .B1(_00434_ ), .B2(_00435_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _16199_ ( .A1(_05122_ ), .A2(_05124_ ), .A3(_06335_ ), .ZN(_00436_ ) );
AOI21_X1 _16200_ ( .A(_07163_ ), .B1(_00405_ ), .B2(_03404_ ), .ZN(_00437_ ) );
OAI21_X1 _16201_ ( .A(_00437_ ), .B1(_03404_ ), .B2(_00405_ ), .ZN(_00438_ ) );
AOI22_X1 _16202_ ( .A1(_05109_ ), .A2(_06580_ ), .B1(\ID_EX_imm [22] ), .B2(_07361_ ), .ZN(_00439_ ) );
AOI21_X1 _16203_ ( .A(_06600_ ), .B1(_00438_ ), .B2(_00439_ ), .ZN(_00440_ ) );
OR2_X1 _16204_ ( .A1(_00440_ ), .A2(_07364_ ), .ZN(_00441_ ) );
NAND3_X1 _16205_ ( .A1(_00410_ ), .A2(_07450_ ), .A3(_07448_ ), .ZN(_00442_ ) );
NAND3_X1 _16206_ ( .A1(_00412_ ), .A2(_07035_ ), .A3(_00442_ ), .ZN(_00443_ ) );
NAND2_X1 _16207_ ( .A1(_04191_ ), .A2(_07090_ ), .ZN(_00444_ ) );
NAND3_X1 _16208_ ( .A1(_04249_ ), .A2(_02429_ ), .A3(_06890_ ), .ZN(_00445_ ) );
OAI21_X1 _16209_ ( .A(_04394_ ), .B1(_04249_ ), .B2(_02429_ ), .ZN(_00446_ ) );
AND3_X1 _16210_ ( .A1(_00444_ ), .A2(_00445_ ), .A3(_00446_ ), .ZN(_00447_ ) );
OR3_X1 _16211_ ( .A1(_07336_ ), .A2(_07005_ ), .A3(_07128_ ), .ZN(_00448_ ) );
NAND2_X1 _16212_ ( .A1(_07341_ ), .A2(_06821_ ), .ZN(_00449_ ) );
NOR2_X1 _16213_ ( .A1(_07479_ ), .A2(_07482_ ), .ZN(_00450_ ) );
OAI211_X1 _16214_ ( .A(_00449_ ), .B(_06813_ ), .C1(_00450_ ), .C2(_06991_ ), .ZN(_00451_ ) );
AOI21_X1 _16215_ ( .A(_07062_ ), .B1(_00448_ ), .B2(_00451_ ), .ZN(_00452_ ) );
AND2_X1 _16216_ ( .A1(_07689_ ), .A2(_06812_ ), .ZN(_00453_ ) );
AND4_X1 _16217_ ( .A1(_06734_ ), .A2(_06764_ ), .A3(_06767_ ), .A4(_07317_ ), .ZN(_00454_ ) );
OR3_X1 _16218_ ( .A1(_00454_ ), .A2(_07039_ ), .A3(_00453_ ), .ZN(_00455_ ) );
AOI221_X4 _16219_ ( .A(_00452_ ), .B1(_06884_ ), .B2(_00453_ ), .C1(_00455_ ), .C2(_06675_ ), .ZN(_00456_ ) );
NAND3_X1 _16220_ ( .A1(_00443_ ), .A2(_00447_ ), .A3(_00456_ ), .ZN(_00457_ ) );
AOI21_X1 _16221_ ( .A(_00441_ ), .B1(_00457_ ), .B2(_06899_ ), .ZN(_00458_ ) );
OAI21_X1 _16222_ ( .A(_06266_ ), .B1(_05112_ ), .B2(_07168_ ), .ZN(_00459_ ) );
OAI21_X1 _16223_ ( .A(_00436_ ), .B1(_00458_ ), .B2(_00459_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NAND3_X1 _16224_ ( .A1(_06566_ ), .A2(_06567_ ), .A3(_06335_ ), .ZN(_00460_ ) );
AOI22_X1 _16225_ ( .A1(_05169_ ), .A2(_06915_ ), .B1(\ID_EX_imm [31] ), .B2(_06916_ ), .ZN(_00461_ ) );
AOI21_X1 _16226_ ( .A(_04377_ ), .B1(_07436_ ), .B2(_03647_ ), .ZN(_00462_ ) );
XNOR2_X1 _16227_ ( .A(_00462_ ), .B(_03625_ ), .ZN(_00463_ ) );
NAND2_X1 _16228_ ( .A1(_00463_ ), .A2(_06595_ ), .ZN(_00464_ ) );
AOI21_X1 _16229_ ( .A(_06601_ ), .B1(_00461_ ), .B2(_00464_ ), .ZN(_00465_ ) );
OR3_X4 _16230_ ( .A1(_07465_ ), .A2(_04280_ ), .A3(_07494_ ), .ZN(_00466_ ) );
OAI21_X1 _16231_ ( .A(_04280_ ), .B1(_07465_ ), .B2(_07494_ ), .ZN(_00467_ ) );
NAND3_X1 _16232_ ( .A1(_00466_ ), .A2(_06605_ ), .A3(_00467_ ), .ZN(_00468_ ) );
NOR3_X1 _16233_ ( .A1(_07289_ ), .A2(_06818_ ), .A3(_07236_ ), .ZN(_00469_ ) );
AOI221_X4 _16234_ ( .A(_00469_ ), .B1(_04277_ ), .B2(_04394_ ), .C1(_04280_ ), .C2(_04308_ ), .ZN(_00470_ ) );
NAND3_X1 _16235_ ( .A1(_07293_ ), .A2(_07296_ ), .A3(_07477_ ), .ZN(_00471_ ) );
OAI211_X1 _16236_ ( .A(_00470_ ), .B(_00471_ ), .C1(_04278_ ), .C2(_07250_ ), .ZN(_00472_ ) );
NOR2_X1 _16237_ ( .A1(_00424_ ), .A2(_00425_ ), .ZN(_00473_ ) );
OAI21_X1 _16238_ ( .A(_06804_ ), .B1(_06838_ ), .B2(_04272_ ), .ZN(_00474_ ) );
MUX2_X1 _16239_ ( .A(_07853_ ), .B(_00474_ ), .S(_06726_ ), .Z(_00475_ ) );
MUX2_X1 _16240_ ( .A(_08000_ ), .B(_00475_ ), .S(_06791_ ), .Z(_00476_ ) );
MUX2_X1 _16241_ ( .A(_00473_ ), .B(_00476_ ), .S(_07281_ ), .Z(_00477_ ) );
OAI21_X1 _16242_ ( .A(_06766_ ), .B1(_06866_ ), .B2(_07289_ ), .ZN(_00478_ ) );
AOI221_X4 _16243_ ( .A(_00472_ ), .B1(_07297_ ), .B2(_00477_ ), .C1(_00478_ ), .C2(_06675_ ), .ZN(_00479_ ) );
AOI21_X1 _16244_ ( .A(_06898_ ), .B1(_00468_ ), .B2(_00479_ ), .ZN(_00480_ ) );
NOR3_X1 _16245_ ( .A1(_00465_ ), .A2(_05029_ ), .A3(_00480_ ), .ZN(_00481_ ) );
OAI21_X1 _16246_ ( .A(_06266_ ), .B1(_05165_ ), .B2(_07168_ ), .ZN(_00482_ ) );
OAI21_X1 _16247_ ( .A(_00460_ ), .B1(_00481_ ), .B2(_00482_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
NOR4_X1 _16248_ ( .A1(_02116_ ), .A2(fanout_net_4 ), .A3(excp_written ), .A4(EXU_valid_LSU ), .ZN(\myexu.state_$_OR__B_Y_$_ANDNOT__B_Y ) );
AOI21_X1 _16249_ ( .A(_02107_ ), .B1(_02049_ ), .B2(_02114_ ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _16250_ ( .A1(_05507_ ), .A2(IDU_valid_EXU ), .ZN(_00483_ ) );
OAI21_X1 _16251_ ( .A(_00483_ ), .B1(_05439_ ), .B2(_05434_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16252_ ( .A1(_05434_ ), .A2(_05438_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16253_ ( .A1(_05434_ ), .A2(_05438_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16254_ ( .A(_05431_ ), .ZN(_00484_ ) );
NOR4_X1 _16255_ ( .A1(_05438_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_05317_ ), .A4(_00484_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16256_ ( .A1(_05793_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_05317_ ), .A4(_05430_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16257_ ( .A(_06000_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16258_ ( .A(_00483_ ), .B1(_00484_ ), .B2(_05507_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16259_ ( .A1(_05431_ ), .A2(_05507_ ), .B1(_02005_ ), .B2(_02116_ ), .ZN(_00485_ ) );
INV_X1 _16260_ ( .A(loaduse_clear ), .ZN(_00486_ ) );
AOI221_X4 _16261_ ( .A(_00485_ ), .B1(\myidu.state [2] ), .B2(_00486_ ), .C1(_05438_ ), .C2(_06000_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16262_ ( .A(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_00487_ ) );
NAND3_X1 _16263_ ( .A1(_05459_ ), .A2(IDU_valid_EXU ), .A3(_00487_ ), .ZN(_00488_ ) );
NAND3_X1 _16264_ ( .A1(_05459_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_00489_ ) );
NOR2_X1 _16265_ ( .A1(_05482_ ), .A2(_05489_ ), .ZN(_00490_ ) );
OAI21_X1 _16266_ ( .A(_05449_ ), .B1(_05361_ ), .B2(_05547_ ), .ZN(_00491_ ) );
NAND4_X1 _16267_ ( .A1(_05352_ ), .A2(_00491_ ), .A3(_05546_ ), .A4(_05531_ ), .ZN(_00492_ ) );
NOR4_X1 _16268_ ( .A1(_05527_ ), .A2(_05529_ ), .A3(_00492_ ), .A4(_05534_ ), .ZN(_00493_ ) );
INV_X1 _16269_ ( .A(_05272_ ), .ZN(_00494_ ) );
NOR2_X1 _16270_ ( .A1(_00494_ ), .A2(_05512_ ), .ZN(_00495_ ) );
AOI21_X1 _16271_ ( .A(_00490_ ), .B1(_00493_ ), .B2(_00495_ ), .ZN(_00496_ ) );
INV_X1 _16272_ ( .A(_00496_ ), .ZN(_00497_ ) );
OAI21_X1 _16273_ ( .A(_05482_ ), .B1(_05503_ ), .B2(_05216_ ), .ZN(_00498_ ) );
NAND2_X1 _16274_ ( .A1(_00497_ ), .A2(_00498_ ), .ZN(_00499_ ) );
NAND3_X1 _16275_ ( .A1(_05431_ ), .A2(IDU_ready_IFU ), .A3(_05210_ ), .ZN(_00500_ ) );
OAI211_X1 _16276_ ( .A(_00488_ ), .B(_00489_ ), .C1(_00499_ ), .C2(_00500_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16277_ ( .A(_02120_ ), .B(_05459_ ), .C1(_05431_ ), .C2(_05507_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _16278_ ( .A(_05429_ ), .B(_05490_ ), .C1(_05426_ ), .C2(_02117_ ), .ZN(_00501_ ) );
BUF_X4 _16279_ ( .A(_00495_ ), .Z(_00502_ ) );
AOI21_X1 _16280_ ( .A(_00501_ ), .B1(_00493_ ), .B2(_00502_ ), .ZN(_00503_ ) );
OAI211_X1 _16281_ ( .A(_05429_ ), .B(_05482_ ), .C1(_05426_ ), .C2(_02117_ ), .ZN(_00504_ ) );
AOI21_X1 _16282_ ( .A(_00504_ ), .B1(_05505_ ), .B2(_05207_ ), .ZN(_00505_ ) );
OAI211_X1 _16283_ ( .A(IDU_ready_IFU ), .B(_05459_ ), .C1(_00503_ ), .C2(_00505_ ), .ZN(_00506_ ) );
NAND3_X1 _16284_ ( .A1(_05459_ ), .A2(\myidu.state [2] ), .A3(_00486_ ), .ZN(_00507_ ) );
NAND2_X1 _16285_ ( .A1(_00506_ ), .A2(_00507_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
AND4_X1 _16286_ ( .A1(\ID_EX_typ [7] ), .A2(_02121_ ), .A3(_05187_ ), .A4(IDU_valid_EXU ), .ZN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16287_ ( .A1(_05428_ ), .A2(IDU_ready_IFU ), .ZN(_00508_ ) );
NOR2_X1 _16288_ ( .A1(_05428_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00509_ ) );
NOR2_X1 _16289_ ( .A1(\myifu.state [0] ), .A2(\myifu.state [1] ), .ZN(_00510_ ) );
NOR4_X1 _16290_ ( .A1(_00508_ ), .A2(_00509_ ), .A3(fanout_net_4 ), .A4(_00510_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
OR3_X1 _16291_ ( .A1(_01971_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06119_ ), .ZN(_00511_ ) );
OAI211_X1 _16292_ ( .A(_05980_ ), .B(_00511_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06121_ ), .ZN(_00512_ ) );
OAI21_X2 _16293_ ( .A(_00512_ ), .B1(\io_master_rdata [31] ), .B2(_05981_ ), .ZN(_00513_ ) );
NOR2_X1 _16294_ ( .A1(_00513_ ), .A2(_06095_ ), .ZN(\myifu.data_in [31] ) );
CLKBUF_X2 _16295_ ( .A(_05982_ ), .Z(_00514_ ) );
OR2_X1 _16296_ ( .A1(_00514_ ), .A2(\io_master_rdata [30] ), .ZN(_00515_ ) );
BUF_X2 _16297_ ( .A(_05986_ ), .Z(_00516_ ) );
CLKBUF_X2 _16298_ ( .A(_06120_ ), .Z(_00517_ ) );
CLKBUF_X2 _16299_ ( .A(_00517_ ), .Z(_00518_ ) );
OR3_X1 _16300_ ( .A1(_02053_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00519_ ) );
OAI211_X1 _16301_ ( .A(_00516_ ), .B(_00519_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00520_ ) );
AND3_X1 _16302_ ( .A1(_00515_ ), .A2(_00520_ ), .A3(_02055_ ), .ZN(\myifu.data_in [30] ) );
BUF_X4 _16303_ ( .A(_01998_ ), .Z(_00521_ ) );
MUX2_X1 _16304_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06122_ ), .Z(_00522_ ) );
OR3_X1 _16305_ ( .A1(_05972_ ), .A2(_05976_ ), .A3(_00522_ ), .ZN(_00523_ ) );
OAI21_X1 _16306_ ( .A(\io_master_rdata [21] ), .B1(_05972_ ), .B2(_05976_ ), .ZN(_00524_ ) );
AOI21_X1 _16307_ ( .A(_00521_ ), .B1(_00523_ ), .B2(_00524_ ), .ZN(\myifu.data_in [21] ) );
MUX2_X1 _16308_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06122_ ), .Z(_00525_ ) );
OR3_X1 _16309_ ( .A1(_05972_ ), .A2(_05976_ ), .A3(_00525_ ), .ZN(_00526_ ) );
OAI21_X1 _16310_ ( .A(\io_master_rdata [20] ), .B1(_05972_ ), .B2(_05976_ ), .ZN(_00527_ ) );
AOI21_X1 _16311_ ( .A(_01998_ ), .B1(_00526_ ), .B2(_00527_ ), .ZN(\myifu.data_in [20] ) );
OR3_X1 _16312_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00528_ ) );
OAI211_X1 _16313_ ( .A(_05982_ ), .B(_00528_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00529_ ) );
OAI21_X1 _16314_ ( .A(_00529_ ), .B1(\io_master_rdata [19] ), .B2(_05986_ ), .ZN(_00530_ ) );
NOR2_X1 _16315_ ( .A1(_00530_ ), .A2(_06094_ ), .ZN(\myifu.data_in [19] ) );
OR3_X1 _16316_ ( .A1(_01971_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00531_ ) );
OAI211_X1 _16317_ ( .A(_05981_ ), .B(_00531_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06121_ ), .ZN(_00532_ ) );
OAI21_X2 _16318_ ( .A(_00532_ ), .B1(\io_master_rdata [18] ), .B2(_05981_ ), .ZN(_00533_ ) );
NOR2_X1 _16319_ ( .A1(_00533_ ), .A2(_06094_ ), .ZN(\myifu.data_in [18] ) );
OR3_X1 _16320_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00534_ ) );
OAI211_X1 _16321_ ( .A(_05982_ ), .B(_00534_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00535_ ) );
OAI21_X1 _16322_ ( .A(_00535_ ), .B1(\io_master_rdata [17] ), .B2(_05986_ ), .ZN(_00536_ ) );
NOR2_X1 _16323_ ( .A1(_00536_ ), .A2(_00521_ ), .ZN(\myifu.data_in [17] ) );
MUX2_X1 _16324_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06122_ ), .Z(_00537_ ) );
OR3_X1 _16325_ ( .A1(_05972_ ), .A2(_05976_ ), .A3(_00537_ ), .ZN(_00538_ ) );
OAI21_X1 _16326_ ( .A(\io_master_rdata [16] ), .B1(_05972_ ), .B2(_05976_ ), .ZN(_00539_ ) );
AOI21_X1 _16327_ ( .A(_01998_ ), .B1(_00538_ ), .B2(_00539_ ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16328_ ( .A1(_01971_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06119_ ), .ZN(_00540_ ) );
OAI211_X1 _16329_ ( .A(_05980_ ), .B(_00540_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06121_ ), .ZN(_00541_ ) );
OAI21_X2 _16330_ ( .A(_00541_ ), .B1(\io_master_rdata [15] ), .B2(_05981_ ), .ZN(_00542_ ) );
NOR2_X1 _16331_ ( .A1(_00542_ ), .A2(_00521_ ), .ZN(\myifu.data_in [15] ) );
OR2_X1 _16332_ ( .A1(_00514_ ), .A2(\io_master_rdata [14] ), .ZN(_00543_ ) );
OR3_X1 _16333_ ( .A1(_02053_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00544_ ) );
OAI211_X1 _16334_ ( .A(_00516_ ), .B(_00544_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00545_ ) );
AND3_X1 _16335_ ( .A1(_00543_ ), .A2(_00545_ ), .A3(_02055_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16336_ ( .A1(_00514_ ), .A2(\io_master_rdata [13] ), .ZN(_00546_ ) );
OR3_X1 _16337_ ( .A1(_02053_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00547_ ) );
OAI211_X1 _16338_ ( .A(_00516_ ), .B(_00547_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00548_ ) );
AND3_X1 _16339_ ( .A1(_00546_ ), .A2(_00548_ ), .A3(_02055_ ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _16340_ ( .A1(_00516_ ), .A2(\io_master_rdata [12] ), .ZN(_00549_ ) );
OR3_X1 _16341_ ( .A1(_02054_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00550_ ) );
OAI211_X1 _16342_ ( .A(_00516_ ), .B(_00550_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00551_ ) );
AND3_X1 _16343_ ( .A1(_00549_ ), .A2(_00551_ ), .A3(_02055_ ), .ZN(\myifu.data_in [12] ) );
OR2_X1 _16344_ ( .A1(_00514_ ), .A2(\io_master_rdata [29] ), .ZN(_00552_ ) );
OR3_X1 _16345_ ( .A1(_02053_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00553_ ) );
OAI211_X1 _16346_ ( .A(_00516_ ), .B(_00553_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00554_ ) );
AND3_X1 _16347_ ( .A1(_00552_ ), .A2(_00554_ ), .A3(_02055_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16348_ ( .A1(_00514_ ), .A2(\io_master_rdata [11] ), .ZN(_00555_ ) );
OR3_X1 _16349_ ( .A1(_02053_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00556_ ) );
OAI211_X1 _16350_ ( .A(_00514_ ), .B(_00556_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00557_ ) );
AND3_X1 _16351_ ( .A1(_00555_ ), .A2(_00557_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [11] ) );
OR3_X1 _16352_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00558_ ) );
OAI211_X1 _16353_ ( .A(_05982_ ), .B(_00558_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00559_ ) );
OAI21_X1 _16354_ ( .A(_00559_ ), .B1(\io_master_rdata [10] ), .B2(_05986_ ), .ZN(_00560_ ) );
NOR2_X1 _16355_ ( .A1(_00560_ ), .A2(_06094_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16356_ ( .A1(_00514_ ), .A2(\io_master_rdata [9] ), .ZN(_00561_ ) );
OR3_X1 _16357_ ( .A1(_02053_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00562_ ) );
OAI211_X1 _16358_ ( .A(_00514_ ), .B(_00562_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00563_ ) );
AND3_X1 _16359_ ( .A1(_00561_ ), .A2(_00563_ ), .A3(_02055_ ), .ZN(\myifu.data_in [9] ) );
BUF_X2 _16360_ ( .A(_00514_ ), .Z(_00564_ ) );
OR2_X1 _16361_ ( .A1(_00564_ ), .A2(\io_master_rdata [8] ), .ZN(_00565_ ) );
OR3_X1 _16362_ ( .A1(_02054_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00566_ ) );
OAI211_X1 _16363_ ( .A(_00564_ ), .B(_00566_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00567_ ) );
AND3_X1 _16364_ ( .A1(_00565_ ), .A2(_00567_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [8] ) );
OR3_X1 _16365_ ( .A1(_01971_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00568_ ) );
OAI211_X1 _16366_ ( .A(_05981_ ), .B(_00568_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06122_ ), .ZN(_00569_ ) );
OAI21_X1 _16367_ ( .A(_00569_ ), .B1(\io_master_rdata [7] ), .B2(_05981_ ), .ZN(_00570_ ) );
NOR2_X1 _16368_ ( .A1(_00570_ ), .A2(_06094_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16369_ ( .A1(_02054_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00571_ ) );
OAI211_X1 _16370_ ( .A(_00564_ ), .B(_00571_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00572_ ) );
OAI21_X1 _16371_ ( .A(_00572_ ), .B1(\io_master_rdata [6] ), .B2(_00564_ ), .ZN(_00573_ ) );
NOR2_X1 _16372_ ( .A1(_00573_ ), .A2(_06094_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16373_ ( .A1(_02054_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00574_ ) );
OAI211_X1 _16374_ ( .A(_00564_ ), .B(_00574_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00575_ ) );
OAI21_X1 _16375_ ( .A(_00575_ ), .B1(\io_master_rdata [5] ), .B2(_00564_ ), .ZN(_00576_ ) );
NOR2_X1 _16376_ ( .A1(_00576_ ), .A2(_00521_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16377_ ( .A1(_02054_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00577_ ) );
OAI211_X1 _16378_ ( .A(_00564_ ), .B(_00577_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00578_ ) );
OAI21_X1 _16379_ ( .A(_00578_ ), .B1(\io_master_rdata [4] ), .B2(_00564_ ), .ZN(_00579_ ) );
NOR2_X1 _16380_ ( .A1(_00579_ ), .A2(_00521_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16381_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00580_ ) );
OAI211_X1 _16382_ ( .A(_05982_ ), .B(_00580_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06122_ ), .ZN(_00581_ ) );
OAI21_X1 _16383_ ( .A(_00581_ ), .B1(\io_master_rdata [3] ), .B2(_05986_ ), .ZN(_00582_ ) );
NOR2_X1 _16384_ ( .A1(_00582_ ), .A2(_00521_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16385_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00583_ ) );
OAI211_X1 _16386_ ( .A(_05982_ ), .B(_00583_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06122_ ), .ZN(_00584_ ) );
OAI21_X2 _16387_ ( .A(_00584_ ), .B1(\io_master_rdata [2] ), .B2(_05986_ ), .ZN(_00585_ ) );
NOR2_X1 _16388_ ( .A1(_00585_ ), .A2(_00521_ ), .ZN(\myifu.data_in [2] ) );
OR3_X1 _16389_ ( .A1(_02052_ ), .A2(_01638_ ), .A3(_00517_ ), .ZN(_00586_ ) );
OAI211_X1 _16390_ ( .A(_05181_ ), .B(_00586_ ), .C1(_01682_ ), .C2(_06123_ ), .ZN(_00587_ ) );
OAI21_X1 _16391_ ( .A(\io_master_rdata [28] ), .B1(_05972_ ), .B2(_05976_ ), .ZN(_00588_ ) );
AOI21_X1 _16392_ ( .A(_06094_ ), .B1(_00587_ ), .B2(_00588_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16393_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00589_ ) );
OAI211_X1 _16394_ ( .A(_05981_ ), .B(_00589_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06122_ ), .ZN(_00590_ ) );
OAI21_X1 _16395_ ( .A(_00590_ ), .B1(\io_master_rdata [1] ), .B2(_05982_ ), .ZN(_00591_ ) );
NOR2_X1 _16396_ ( .A1(_00591_ ), .A2(_00521_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16397_ ( .A1(_02054_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00518_ ), .ZN(_00592_ ) );
OAI211_X1 _16398_ ( .A(_00516_ ), .B(_00592_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00593_ ) );
OAI21_X1 _16399_ ( .A(_00593_ ), .B1(\io_master_rdata [0] ), .B2(_00564_ ), .ZN(_00594_ ) );
NOR2_X1 _16400_ ( .A1(_00594_ ), .A2(_00521_ ), .ZN(\myifu.data_in [0] ) );
OR3_X1 _16401_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00595_ ) );
OAI211_X1 _16402_ ( .A(_05982_ ), .B(_00595_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06122_ ), .ZN(_00596_ ) );
OAI21_X1 _16403_ ( .A(_00596_ ), .B1(\io_master_rdata [27] ), .B2(_05986_ ), .ZN(_00597_ ) );
NOR2_X1 _16404_ ( .A1(_00597_ ), .A2(_06094_ ), .ZN(\myifu.data_in [27] ) );
OR3_X1 _16405_ ( .A1(_01971_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00598_ ) );
OAI21_X1 _16406_ ( .A(_00598_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06121_ ), .ZN(_00599_ ) );
MUX2_X1 _16407_ ( .A(\io_master_rdata [26] ), .B(_00599_ ), .S(_05181_ ), .Z(_00600_ ) );
AND2_X1 _16408_ ( .A1(_00600_ ), .A2(_02055_ ), .ZN(\myifu.data_in [26] ) );
OR3_X1 _16409_ ( .A1(_02052_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00601_ ) );
OAI211_X1 _16410_ ( .A(_05982_ ), .B(_00601_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06122_ ), .ZN(_00602_ ) );
OAI21_X1 _16411_ ( .A(_00602_ ), .B1(\io_master_rdata [25] ), .B2(_05986_ ), .ZN(_00603_ ) );
NOR2_X1 _16412_ ( .A1(_00603_ ), .A2(_06094_ ), .ZN(\myifu.data_in [25] ) );
OR2_X1 _16413_ ( .A1(_00514_ ), .A2(\io_master_rdata [24] ), .ZN(_00604_ ) );
OR3_X1 _16414_ ( .A1(_02053_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00517_ ), .ZN(_00605_ ) );
OAI211_X1 _16415_ ( .A(_00516_ ), .B(_00605_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06123_ ), .ZN(_00606_ ) );
AND3_X1 _16416_ ( .A1(_00604_ ), .A2(_00606_ ), .A3(_02054_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16417_ ( .A1(_01971_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06120_ ), .ZN(_00607_ ) );
OAI211_X1 _16418_ ( .A(_05980_ ), .B(_00607_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06121_ ), .ZN(_00608_ ) );
OAI21_X2 _16419_ ( .A(_00608_ ), .B1(\io_master_rdata [23] ), .B2(_05981_ ), .ZN(_00609_ ) );
NOR2_X1 _16420_ ( .A1(_00609_ ), .A2(_00521_ ), .ZN(\myifu.data_in [23] ) );
OR2_X1 _16421_ ( .A1(_00516_ ), .A2(\io_master_rdata [22] ), .ZN(_00610_ ) );
OR3_X1 _16422_ ( .A1(_02054_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00518_ ), .ZN(_00611_ ) );
OAI211_X1 _16423_ ( .A(_00516_ ), .B(_00611_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00612_ ) );
AND3_X1 _16424_ ( .A1(_00610_ ), .A2(_00612_ ), .A3(_02054_ ), .ZN(\myifu.data_in [22] ) );
OR2_X1 _16425_ ( .A1(_00242_ ), .A2(_02057_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
OAI21_X1 _16426_ ( .A(_02056_ ), .B1(_06075_ ), .B2(_06077_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
OAI21_X1 _16427_ ( .A(_02056_ ), .B1(_06078_ ), .B2(_06077_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16428_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .ZN(_00613_ ) );
OAI21_X1 _16429_ ( .A(_02056_ ), .B1(_00613_ ), .B2(_06077_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
OAI21_X1 _16430_ ( .A(\IF_ID_inst [16] ), .B1(_05204_ ), .B2(_05206_ ), .ZN(_00614_ ) );
AND2_X1 _16431_ ( .A1(_00495_ ), .A2(_05554_ ), .ZN(_00615_ ) );
AND4_X1 _16432_ ( .A1(_05207_ ), .A2(_05532_ ), .A3(_05460_ ), .A4(_05457_ ), .ZN(_00616_ ) );
NOR4_X1 _16433_ ( .A1(_05527_ ), .A2(_05529_ ), .A3(_05305_ ), .A4(_05534_ ), .ZN(_00617_ ) );
NAND3_X1 _16434_ ( .A1(_00615_ ), .A2(_00616_ ), .A3(_00617_ ), .ZN(_00618_ ) );
AND2_X1 _16435_ ( .A1(_00618_ ), .A2(_05620_ ), .ZN(_00619_ ) );
OAI221_X1 _16436_ ( .A(_00614_ ), .B1(_05291_ ), .B2(_00502_ ), .C1(_00619_ ), .C2(_05214_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
AND3_X1 _16437_ ( .A1(_05594_ ), .A2(_05231_ ), .A3(\IF_ID_inst [31] ), .ZN(_00620_ ) );
INV_X1 _16438_ ( .A(_00620_ ), .ZN(_00621_ ) );
OAI221_X1 _16439_ ( .A(_00621_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_05505_ ), .C1(_00615_ ), .C2(_05209_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
NOR2_X1 _16440_ ( .A1(_05502_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00622_ ) );
NOR2_X1 _16441_ ( .A1(_00495_ ), .A2(_05209_ ), .ZN(_00623_ ) );
NOR2_X2 _16442_ ( .A1(_00622_ ), .A2(_00623_ ), .ZN(_00624_ ) );
BUF_X4 _16443_ ( .A(_00624_ ), .Z(_00625_ ) );
BUF_X4 _16444_ ( .A(_00621_ ), .Z(_00626_ ) );
BUF_X4 _16445_ ( .A(_05554_ ), .Z(_00627_ ) );
OAI211_X1 _16446_ ( .A(_00625_ ), .B(_00626_ ), .C1(_05213_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16447_ ( .A(_00625_ ), .B(_00626_ ), .C1(_05214_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16448_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05217_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
OAI21_X1 _16449_ ( .A(_00625_ ), .B1(_05301_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI21_X1 _16450_ ( .A(_00625_ ), .B1(_05318_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI21_X1 _16451_ ( .A(_00625_ ), .B1(_05319_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI21_X1 _16452_ ( .A(_00625_ ), .B1(_05437_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI21_X1 _16453_ ( .A(_00625_ ), .B1(_05241_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI21_X1 _16454_ ( .A(_00625_ ), .B1(_05329_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI21_X1 _16455_ ( .A(_00625_ ), .B1(_05265_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI21_X1 _16456_ ( .A(_00625_ ), .B1(_05239_ ), .B2(_05310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16457_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05218_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
AOI22_X1 _16458_ ( .A1(_00494_ ), .A2(\IF_ID_inst [31] ), .B1(\IF_ID_inst [7] ), .B2(_05512_ ), .ZN(_00628_ ) );
OAI221_X1 _16459_ ( .A(_00628_ ), .B1(_05217_ ), .B2(_05620_ ), .C1(_05505_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16460_ ( .A(_05649_ ), .ZN(_00629_ ) );
OAI221_X1 _16461_ ( .A(_00629_ ), .B1(_00502_ ), .B2(_05213_ ), .C1(_05505_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
INV_X1 _16462_ ( .A(_05645_ ), .ZN(_00630_ ) );
OAI221_X1 _16463_ ( .A(_00630_ ), .B1(_00502_ ), .B2(_05218_ ), .C1(_05505_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16464_ ( .A(_05700_ ), .ZN(_00631_ ) );
OAI221_X1 _16465_ ( .A(_00631_ ), .B1(_00502_ ), .B2(_05219_ ), .C1(_05505_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
OAI21_X1 _16466_ ( .A(\IF_ID_inst [27] ), .B1(_00494_ ), .B2(_05512_ ), .ZN(_00632_ ) );
OAI221_X1 _16467_ ( .A(_00632_ ), .B1(_05220_ ), .B2(_05620_ ), .C1(_05505_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16468_ ( .A(_05654_ ), .ZN(_00633_ ) );
OAI221_X1 _16469_ ( .A(_00633_ ), .B1(_00502_ ), .B2(_05222_ ), .C1(_05505_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16470_ ( .A(_05658_ ), .ZN(_00634_ ) );
OAI221_X1 _16471_ ( .A(_00634_ ), .B1(_00502_ ), .B2(_05223_ ), .C1(_05505_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16472_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05219_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16473_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05220_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16474_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05222_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16475_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05223_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16476_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05224_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16477_ ( .A(_00624_ ), .B(_00626_ ), .C1(_05225_ ), .C2(_00627_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16478_ ( .A(_00624_ ), .B(_00621_ ), .C1(_05226_ ), .C2(_05554_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16479_ ( .A(\IF_ID_inst [19] ), .B1(_05204_ ), .B2(_05206_ ), .ZN(_00635_ ) );
OAI221_X1 _16480_ ( .A(_00635_ ), .B1(_05245_ ), .B2(_00502_ ), .C1(_00619_ ), .C2(_05224_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16481_ ( .A(\IF_ID_inst [18] ), .B1(_05204_ ), .B2(_05206_ ), .ZN(_00636_ ) );
OAI221_X1 _16482_ ( .A(_00636_ ), .B1(_05246_ ), .B2(_00502_ ), .C1(_00619_ ), .C2(_05225_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16483_ ( .A(\IF_ID_inst [17] ), .B1(_05204_ ), .B2(_05206_ ), .ZN(_00637_ ) );
OAI221_X1 _16484_ ( .A(_00637_ ), .B1(_05247_ ), .B2(_00502_ ), .C1(_00619_ ), .C2(_05226_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OAI21_X1 _16485_ ( .A(\IF_ID_inst [15] ), .B1(_05204_ ), .B2(_05206_ ), .ZN(_00638_ ) );
OAI221_X1 _16486_ ( .A(_00638_ ), .B1(_05240_ ), .B2(_05272_ ), .C1(_00618_ ), .C2(_05217_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AND3_X1 _16487_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00639_ ) );
CLKBUF_X2 _16488_ ( .A(_05902_ ), .Z(_00640_ ) );
AND3_X1 _16489_ ( .A1(_00640_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00641_ ) );
AOI211_X1 _16490_ ( .A(_00639_ ), .B(_00641_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_06074_ ), .ZN(_00642_ ) );
NAND2_X2 _16491_ ( .A1(_06076_ ), .A2(\IF_ID_pc [2] ), .ZN(_00643_ ) );
BUF_X2 _16492_ ( .A(_00643_ ), .Z(_00644_ ) );
NAND2_X2 _16493_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00645_ ) );
BUF_X4 _16494_ ( .A(_00645_ ), .Z(_00646_ ) );
BUF_X4 _16495_ ( .A(_00646_ ), .Z(_00647_ ) );
BUF_X4 _16496_ ( .A(_05914_ ), .Z(_00648_ ) );
BUF_X4 _16497_ ( .A(_00648_ ), .Z(_00649_ ) );
NAND3_X1 _16498_ ( .A1(_00649_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00650_ ) );
NAND4_X1 _16499_ ( .A1(_00642_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_00650_ ), .ZN(_00651_ ) );
NOR2_X1 _16500_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00652_ ) );
BUF_X2 _16501_ ( .A(_00652_ ), .Z(_00653_ ) );
BUF_X4 _16502_ ( .A(_00653_ ), .Z(_00654_ ) );
BUF_X4 _16503_ ( .A(_05903_ ), .Z(_00655_ ) );
NAND3_X1 _16504_ ( .A1(_00655_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00656_ ) );
NAND3_X1 _16505_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00657_ ) );
AND2_X1 _16506_ ( .A1(_00656_ ), .A2(_00657_ ), .ZN(_00658_ ) );
NAND2_X1 _16507_ ( .A1(_00643_ ), .A2(_00645_ ), .ZN(_00659_ ) );
BUF_X4 _16508_ ( .A(_00659_ ), .Z(_00660_ ) );
BUF_X4 _16509_ ( .A(_05914_ ), .Z(_00661_ ) );
BUF_X4 _16510_ ( .A(_00661_ ), .Z(_00662_ ) );
NAND3_X1 _16511_ ( .A1(_00662_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00663_ ) );
BUF_X4 _16512_ ( .A(_05915_ ), .Z(_00664_ ) );
NAND3_X1 _16513_ ( .A1(_05905_ ), .A2(_00664_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00665_ ) );
NAND4_X1 _16514_ ( .A1(_00658_ ), .A2(_00660_ ), .A3(_00663_ ), .A4(_00665_ ), .ZN(_00666_ ) );
NAND3_X1 _16515_ ( .A1(_00651_ ), .A2(_00654_ ), .A3(_00666_ ), .ZN(_00667_ ) );
INV_X1 _16516_ ( .A(\IF_ID_pc [1] ), .ZN(_00668_ ) );
OAI211_X1 _16517_ ( .A(_00668_ ), .B(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .C1(_05408_ ), .C2(\myifu.tmp_offset [2] ), .ZN(_00669_ ) );
NOR2_X1 _16518_ ( .A1(_05998_ ), .A2(\IF_ID_pc [2] ), .ZN(_00670_ ) );
NOR2_X1 _16519_ ( .A1(_00669_ ), .A2(_00670_ ), .ZN(_00671_ ) );
INV_X1 _16520_ ( .A(_00671_ ), .ZN(_00672_ ) );
NOR2_X4 _16521_ ( .A1(_05994_ ), .A2(_00672_ ), .ZN(_00673_ ) );
BUF_X4 _16522_ ( .A(_00673_ ), .Z(_00674_ ) );
OAI21_X1 _16523_ ( .A(\myifu.state [2] ), .B1(_00674_ ), .B2(_05679_ ), .ZN(_00675_ ) );
BUF_X2 _16524_ ( .A(_00672_ ), .Z(_00676_ ) );
NOR3_X1 _16525_ ( .A1(_05995_ ), .A2(\myifu.data_in [8] ), .A3(_00676_ ), .ZN(_00677_ ) );
OAI21_X1 _16526_ ( .A(_00667_ ), .B1(_00675_ ), .B2(_00677_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16527_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00678_ ) );
AND3_X1 _16528_ ( .A1(_00640_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00679_ ) );
BUF_X4 _16529_ ( .A(_06073_ ), .Z(_00680_ ) );
AOI211_X1 _16530_ ( .A(_00678_ ), .B(_00679_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00680_ ), .ZN(_00681_ ) );
NAND3_X1 _16531_ ( .A1(_00649_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00682_ ) );
NAND4_X1 _16532_ ( .A1(_00681_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_00682_ ), .ZN(_00683_ ) );
NAND3_X1 _16533_ ( .A1(_00655_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00684_ ) );
NAND3_X1 _16534_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00685_ ) );
AND2_X1 _16535_ ( .A1(_00684_ ), .A2(_00685_ ), .ZN(_00686_ ) );
NAND3_X1 _16536_ ( .A1(_00662_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00687_ ) );
BUF_X4 _16537_ ( .A(_05902_ ), .Z(_00688_ ) );
BUF_X4 _16538_ ( .A(_00688_ ), .Z(_00689_ ) );
NAND3_X1 _16539_ ( .A1(_00689_ ), .A2(_00664_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00690_ ) );
NAND4_X1 _16540_ ( .A1(_00686_ ), .A2(_00660_ ), .A3(_00687_ ), .A4(_00690_ ), .ZN(_00691_ ) );
NAND3_X1 _16541_ ( .A1(_00683_ ), .A2(_00654_ ), .A3(_00691_ ), .ZN(_00692_ ) );
OAI21_X1 _16542_ ( .A(\myifu.state [2] ), .B1(_00674_ ), .B2(_05335_ ), .ZN(_00693_ ) );
NOR3_X1 _16543_ ( .A1(_05995_ ), .A2(\myifu.data_in [31] ), .A3(_00676_ ), .ZN(_00694_ ) );
OAI21_X1 _16544_ ( .A(_00692_ ), .B1(_00693_ ), .B2(_00694_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
OR3_X1 _16545_ ( .A1(_05995_ ), .A2(\myifu.data_in [30] ), .A3(_00676_ ), .ZN(_00695_ ) );
OAI211_X1 _16546_ ( .A(_00695_ ), .B(\myifu.state [2] ), .C1(_05650_ ), .C2(_00674_ ), .ZN(_00696_ ) );
AND3_X1 _16547_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00697_ ) );
AND3_X1 _16548_ ( .A1(_05904_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00698_ ) );
AOI211_X1 _16549_ ( .A(_00697_ ), .B(_00698_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_06074_ ), .ZN(_00699_ ) );
NAND3_X1 _16550_ ( .A1(_05916_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00700_ ) );
NAND4_X1 _16551_ ( .A1(_00699_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_00700_ ), .ZN(_00701_ ) );
NAND3_X1 _16552_ ( .A1(_00689_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00702_ ) );
NAND3_X1 _16553_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00703_ ) );
AND2_X1 _16554_ ( .A1(_00702_ ), .A2(_00703_ ), .ZN(_00704_ ) );
BUF_X4 _16555_ ( .A(_00659_ ), .Z(_00705_ ) );
BUF_X2 _16556_ ( .A(_00705_ ), .Z(_00706_ ) );
NAND3_X1 _16557_ ( .A1(_05916_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00707_ ) );
NAND3_X1 _16558_ ( .A1(_05905_ ), .A2(_00662_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00708_ ) );
NAND4_X1 _16559_ ( .A1(_00704_ ), .A2(_00706_ ), .A3(_00707_ ), .A4(_00708_ ), .ZN(_00709_ ) );
NAND3_X1 _16560_ ( .A1(_00701_ ), .A2(_00654_ ), .A3(_00709_ ), .ZN(_00710_ ) );
NAND2_X1 _16561_ ( .A1(_00696_ ), .A2(_00710_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
INV_X1 _16562_ ( .A(\myifu.state [2] ), .ZN(_00711_ ) );
BUF_X4 _16563_ ( .A(_00711_ ), .Z(_00712_ ) );
BUF_X2 _16564_ ( .A(_05994_ ), .Z(_00713_ ) );
BUF_X2 _16565_ ( .A(_00672_ ), .Z(_00714_ ) );
NOR3_X1 _16566_ ( .A1(_00713_ ), .A2(\myifu.data_in [21] ), .A3(_00714_ ), .ZN(_00715_ ) );
INV_X1 _16567_ ( .A(_00673_ ), .ZN(_00716_ ) );
BUF_X4 _16568_ ( .A(_00716_ ), .Z(_00717_ ) );
AOI211_X1 _16569_ ( .A(_00712_ ), .B(_00715_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00718_ ) );
AND3_X1 _16570_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00719_ ) );
AND3_X1 _16571_ ( .A1(_05903_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00720_ ) );
AOI211_X1 _16572_ ( .A(_00719_ ), .B(_00720_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_00680_ ), .ZN(_00721_ ) );
BUF_X4 _16573_ ( .A(_00643_ ), .Z(_00722_ ) );
NAND3_X1 _16574_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00723_ ) );
NAND4_X1 _16575_ ( .A1(_00721_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_00723_ ), .ZN(_00724_ ) );
NAND3_X1 _16576_ ( .A1(_00688_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00725_ ) );
NAND3_X1 _16577_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00726_ ) );
AND2_X1 _16578_ ( .A1(_00725_ ), .A2(_00726_ ), .ZN(_00727_ ) );
BUF_X4 _16579_ ( .A(_00659_ ), .Z(_00728_ ) );
NAND3_X1 _16580_ ( .A1(_00661_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00729_ ) );
BUF_X4 _16581_ ( .A(_05903_ ), .Z(_00730_ ) );
NAND3_X1 _16582_ ( .A1(_00730_ ), .A2(_05915_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00731_ ) );
NAND4_X1 _16583_ ( .A1(_00727_ ), .A2(_00728_ ), .A3(_00729_ ), .A4(_00731_ ), .ZN(_00732_ ) );
AND3_X1 _16584_ ( .A1(_00724_ ), .A2(_00653_ ), .A3(_00732_ ), .ZN(_00733_ ) );
OR2_X1 _16585_ ( .A1(_00718_ ), .A2(_00733_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
NOR3_X1 _16586_ ( .A1(_00713_ ), .A2(\myifu.data_in [20] ), .A3(_00714_ ), .ZN(_00734_ ) );
AOI211_X1 _16587_ ( .A(_00712_ ), .B(_00734_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00735_ ) );
AND3_X1 _16588_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00736_ ) );
AND3_X1 _16589_ ( .A1(_05903_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00737_ ) );
AOI211_X1 _16590_ ( .A(_00736_ ), .B(_00737_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_00680_ ), .ZN(_00738_ ) );
NAND3_X1 _16591_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00739_ ) );
NAND4_X1 _16592_ ( .A1(_00738_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_00739_ ), .ZN(_00740_ ) );
NAND3_X1 _16593_ ( .A1(_00688_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00741_ ) );
NAND3_X1 _16594_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00742_ ) );
AND2_X1 _16595_ ( .A1(_00741_ ), .A2(_00742_ ), .ZN(_00743_ ) );
NAND3_X1 _16596_ ( .A1(_00661_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00744_ ) );
NAND3_X1 _16597_ ( .A1(_00730_ ), .A2(_05915_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00745_ ) );
NAND4_X1 _16598_ ( .A1(_00743_ ), .A2(_00728_ ), .A3(_00744_ ), .A4(_00745_ ), .ZN(_00746_ ) );
AND3_X1 _16599_ ( .A1(_00740_ ), .A2(_00653_ ), .A3(_00746_ ), .ZN(_00747_ ) );
OR2_X1 _16600_ ( .A1(_00735_ ), .A2(_00747_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
NOR3_X1 _16601_ ( .A1(_00713_ ), .A2(\myifu.data_in [19] ), .A3(_00714_ ), .ZN(_00748_ ) );
AOI211_X1 _16602_ ( .A(_00712_ ), .B(_00748_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00749_ ) );
AND3_X1 _16603_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00750_ ) );
AND3_X1 _16604_ ( .A1(_05903_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00751_ ) );
AOI211_X1 _16605_ ( .A(_00750_ ), .B(_00751_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_00680_ ), .ZN(_00752_ ) );
NAND3_X1 _16606_ ( .A1(_00648_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00753_ ) );
NAND4_X1 _16607_ ( .A1(_00752_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_00753_ ), .ZN(_00754_ ) );
NAND3_X1 _16608_ ( .A1(_00688_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00755_ ) );
NAND3_X1 _16609_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00756_ ) );
AND2_X1 _16610_ ( .A1(_00755_ ), .A2(_00756_ ), .ZN(_00757_ ) );
NAND3_X1 _16611_ ( .A1(_00661_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00758_ ) );
NAND3_X1 _16612_ ( .A1(_00730_ ), .A2(_05915_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00759_ ) );
NAND4_X1 _16613_ ( .A1(_00757_ ), .A2(_00728_ ), .A3(_00758_ ), .A4(_00759_ ), .ZN(_00760_ ) );
AND3_X1 _16614_ ( .A1(_00754_ ), .A2(_00653_ ), .A3(_00760_ ), .ZN(_00761_ ) );
OR2_X1 _16615_ ( .A1(_00749_ ), .A2(_00761_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
NOR3_X1 _16616_ ( .A1(_00713_ ), .A2(\myifu.data_in [18] ), .A3(_00714_ ), .ZN(_00762_ ) );
AOI211_X1 _16617_ ( .A(_00712_ ), .B(_00762_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00763_ ) );
AND3_X1 _16618_ ( .A1(fanout_net_13 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00764_ ) );
AND3_X1 _16619_ ( .A1(_05903_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00765_ ) );
AOI211_X1 _16620_ ( .A(_00764_ ), .B(_00765_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_00680_ ), .ZN(_00766_ ) );
NAND3_X1 _16621_ ( .A1(_00648_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00767_ ) );
NAND4_X1 _16622_ ( .A1(_00766_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_00767_ ), .ZN(_00768_ ) );
NAND3_X1 _16623_ ( .A1(_00688_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00769_ ) );
NAND3_X1 _16624_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00770_ ) );
AND2_X1 _16625_ ( .A1(_00769_ ), .A2(_00770_ ), .ZN(_00771_ ) );
NAND3_X1 _16626_ ( .A1(_00661_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00772_ ) );
BUF_X4 _16627_ ( .A(_05914_ ), .Z(_00773_ ) );
NAND3_X1 _16628_ ( .A1(_00730_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00774_ ) );
NAND4_X1 _16629_ ( .A1(_00771_ ), .A2(_00728_ ), .A3(_00772_ ), .A4(_00774_ ), .ZN(_00775_ ) );
AND3_X1 _16630_ ( .A1(_00768_ ), .A2(_00653_ ), .A3(_00775_ ), .ZN(_00776_ ) );
OR2_X1 _16631_ ( .A1(_00763_ ), .A2(_00776_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
NOR3_X1 _16632_ ( .A1(_00713_ ), .A2(\myifu.data_in [17] ), .A3(_00714_ ), .ZN(_00777_ ) );
AOI211_X1 _16633_ ( .A(_00712_ ), .B(_00777_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00778_ ) );
AND3_X1 _16634_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00779_ ) );
AND3_X1 _16635_ ( .A1(_05903_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00780_ ) );
BUF_X4 _16636_ ( .A(_06073_ ), .Z(_00781_ ) );
AOI211_X1 _16637_ ( .A(_00779_ ), .B(_00780_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_00781_ ), .ZN(_00782_ ) );
NAND3_X1 _16638_ ( .A1(_00648_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00783_ ) );
NAND4_X1 _16639_ ( .A1(_00782_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_00783_ ), .ZN(_00784_ ) );
NAND3_X1 _16640_ ( .A1(_00688_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00785_ ) );
NAND3_X1 _16641_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00786_ ) );
AND2_X1 _16642_ ( .A1(_00785_ ), .A2(_00786_ ), .ZN(_00787_ ) );
NAND3_X1 _16643_ ( .A1(_00661_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00788_ ) );
NAND3_X1 _16644_ ( .A1(_00730_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00789_ ) );
NAND4_X1 _16645_ ( .A1(_00787_ ), .A2(_00728_ ), .A3(_00788_ ), .A4(_00789_ ), .ZN(_00790_ ) );
AND3_X1 _16646_ ( .A1(_00784_ ), .A2(_00653_ ), .A3(_00790_ ), .ZN(_00791_ ) );
OR2_X1 _16647_ ( .A1(_00778_ ), .A2(_00791_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NOR3_X1 _16648_ ( .A1(_00713_ ), .A2(\myifu.data_in [16] ), .A3(_00714_ ), .ZN(_00792_ ) );
AOI211_X1 _16649_ ( .A(_00712_ ), .B(_00792_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00793_ ) );
NAND3_X1 _16650_ ( .A1(_00688_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00794_ ) );
NAND3_X1 _16651_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00795_ ) );
AND2_X1 _16652_ ( .A1(_00794_ ), .A2(_00795_ ), .ZN(_00796_ ) );
NAND3_X1 _16653_ ( .A1(_00648_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00797_ ) );
NAND3_X1 _16654_ ( .A1(_00655_ ), .A2(_00661_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00798_ ) );
NAND4_X1 _16655_ ( .A1(_00796_ ), .A2(_00660_ ), .A3(_00797_ ), .A4(_00798_ ), .ZN(_00799_ ) );
AND3_X1 _16656_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00800_ ) );
AND3_X1 _16657_ ( .A1(_05902_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00801_ ) );
AOI211_X1 _16658_ ( .A(_00800_ ), .B(_00801_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_06073_ ), .ZN(_00802_ ) );
NAND3_X1 _16659_ ( .A1(_05915_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00803_ ) );
NAND4_X1 _16660_ ( .A1(_00802_ ), .A2(_00643_ ), .A3(_00645_ ), .A4(_00803_ ), .ZN(_00804_ ) );
AND3_X1 _16661_ ( .A1(_00799_ ), .A2(_00653_ ), .A3(_00804_ ), .ZN(_00805_ ) );
OR2_X1 _16662_ ( .A1(_00793_ ), .A2(_00805_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
BUF_X4 _16663_ ( .A(_05994_ ), .Z(_00806_ ) );
NOR3_X1 _16664_ ( .A1(_00806_ ), .A2(\myifu.data_in [15] ), .A3(_00714_ ), .ZN(_00807_ ) );
AOI211_X1 _16665_ ( .A(_00712_ ), .B(_00807_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00808_ ) );
AND3_X1 _16666_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00809_ ) );
CLKBUF_X2 _16667_ ( .A(_05902_ ), .Z(_00810_ ) );
AND3_X1 _16668_ ( .A1(_00810_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00811_ ) );
AOI211_X1 _16669_ ( .A(_00809_ ), .B(_00811_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_00781_ ), .ZN(_00812_ ) );
NAND3_X1 _16670_ ( .A1(_00648_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00813_ ) );
NAND4_X1 _16671_ ( .A1(_00812_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_00813_ ), .ZN(_00814_ ) );
BUF_X4 _16672_ ( .A(_05902_ ), .Z(_00815_ ) );
NAND3_X1 _16673_ ( .A1(_00815_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00816_ ) );
NAND3_X1 _16674_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00817_ ) );
AND2_X1 _16675_ ( .A1(_00816_ ), .A2(_00817_ ), .ZN(_00818_ ) );
BUF_X4 _16676_ ( .A(_05914_ ), .Z(_00819_ ) );
NAND3_X1 _16677_ ( .A1(_00819_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00820_ ) );
NAND3_X1 _16678_ ( .A1(_00730_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00821_ ) );
NAND4_X1 _16679_ ( .A1(_00818_ ), .A2(_00728_ ), .A3(_00820_ ), .A4(_00821_ ), .ZN(_00822_ ) );
AND3_X1 _16680_ ( .A1(_00814_ ), .A2(_00653_ ), .A3(_00822_ ), .ZN(_00823_ ) );
OR2_X1 _16681_ ( .A1(_00808_ ), .A2(_00823_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
NOR3_X1 _16682_ ( .A1(_00806_ ), .A2(\myifu.data_in [14] ), .A3(_00714_ ), .ZN(_00824_ ) );
AOI211_X1 _16683_ ( .A(_00712_ ), .B(_00824_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00825_ ) );
AND3_X1 _16684_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00826_ ) );
AND3_X1 _16685_ ( .A1(_00810_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00827_ ) );
AOI211_X1 _16686_ ( .A(_00826_ ), .B(_00827_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_00781_ ), .ZN(_00828_ ) );
BUF_X4 _16687_ ( .A(_00645_ ), .Z(_00829_ ) );
BUF_X4 _16688_ ( .A(_05914_ ), .Z(_00830_ ) );
NAND3_X1 _16689_ ( .A1(_00830_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00831_ ) );
NAND4_X1 _16690_ ( .A1(_00828_ ), .A2(_00722_ ), .A3(_00829_ ), .A4(_00831_ ), .ZN(_00832_ ) );
CLKBUF_X2 _16691_ ( .A(_00652_ ), .Z(_00833_ ) );
NAND3_X1 _16692_ ( .A1(_00815_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00834_ ) );
NAND3_X1 _16693_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00835_ ) );
AND2_X1 _16694_ ( .A1(_00834_ ), .A2(_00835_ ), .ZN(_00836_ ) );
NAND3_X1 _16695_ ( .A1(_00819_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00837_ ) );
NAND3_X1 _16696_ ( .A1(_00730_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00838_ ) );
NAND4_X1 _16697_ ( .A1(_00836_ ), .A2(_00728_ ), .A3(_00837_ ), .A4(_00838_ ), .ZN(_00839_ ) );
AND3_X1 _16698_ ( .A1(_00832_ ), .A2(_00833_ ), .A3(_00839_ ), .ZN(_00840_ ) );
OR2_X1 _16699_ ( .A1(_00825_ ), .A2(_00840_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
BUF_X4 _16700_ ( .A(_00672_ ), .Z(_00841_ ) );
NOR3_X1 _16701_ ( .A1(_00806_ ), .A2(\myifu.data_in [13] ), .A3(_00841_ ), .ZN(_00842_ ) );
AOI211_X1 _16702_ ( .A(_00712_ ), .B(_00842_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00843_ ) );
AND3_X1 _16703_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00844_ ) );
AND3_X1 _16704_ ( .A1(_00810_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00845_ ) );
AOI211_X1 _16705_ ( .A(_00844_ ), .B(_00845_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_00781_ ), .ZN(_00846_ ) );
BUF_X4 _16706_ ( .A(_00643_ ), .Z(_00847_ ) );
NAND3_X1 _16707_ ( .A1(_00830_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00848_ ) );
NAND4_X1 _16708_ ( .A1(_00846_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_00848_ ), .ZN(_00849_ ) );
NAND3_X1 _16709_ ( .A1(_00815_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00850_ ) );
NAND3_X1 _16710_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00851_ ) );
AND2_X1 _16711_ ( .A1(_00850_ ), .A2(_00851_ ), .ZN(_00852_ ) );
NAND3_X1 _16712_ ( .A1(_00819_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_00853_ ) );
NAND3_X1 _16713_ ( .A1(_00730_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_00854_ ) );
NAND4_X1 _16714_ ( .A1(_00852_ ), .A2(_00728_ ), .A3(_00853_ ), .A4(_00854_ ), .ZN(_00855_ ) );
AND3_X1 _16715_ ( .A1(_00849_ ), .A2(_00833_ ), .A3(_00855_ ), .ZN(_00856_ ) );
OR2_X1 _16716_ ( .A1(_00843_ ), .A2(_00856_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
NOR3_X1 _16717_ ( .A1(_00806_ ), .A2(\myifu.data_in [12] ), .A3(_00841_ ), .ZN(_00857_ ) );
AOI211_X1 _16718_ ( .A(_00712_ ), .B(_00857_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00717_ ), .ZN(_00858_ ) );
AND3_X1 _16719_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_00859_ ) );
AND3_X1 _16720_ ( .A1(_00810_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_00860_ ) );
AOI211_X1 _16721_ ( .A(_00859_ ), .B(_00860_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_00781_ ), .ZN(_00861_ ) );
NAND3_X1 _16722_ ( .A1(_00830_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_00862_ ) );
NAND4_X1 _16723_ ( .A1(_00861_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_00862_ ), .ZN(_00863_ ) );
NAND3_X1 _16724_ ( .A1(_00815_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_00864_ ) );
NAND3_X1 _16725_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_00865_ ) );
AND2_X1 _16726_ ( .A1(_00864_ ), .A2(_00865_ ), .ZN(_00866_ ) );
NAND3_X1 _16727_ ( .A1(_00819_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_00867_ ) );
NAND3_X1 _16728_ ( .A1(_00730_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_00868_ ) );
NAND4_X1 _16729_ ( .A1(_00866_ ), .A2(_00705_ ), .A3(_00867_ ), .A4(_00868_ ), .ZN(_00869_ ) );
AND3_X1 _16730_ ( .A1(_00863_ ), .A2(_00833_ ), .A3(_00869_ ), .ZN(_00870_ ) );
OR2_X1 _16731_ ( .A1(_00858_ ), .A2(_00870_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
OR3_X1 _16732_ ( .A1(_00713_ ), .A2(\myifu.data_in [29] ), .A3(_00676_ ), .ZN(_00871_ ) );
OAI211_X1 _16733_ ( .A(_00871_ ), .B(\myifu.state [2] ), .C1(_05646_ ), .C2(_00674_ ), .ZN(_00872_ ) );
AND3_X1 _16734_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_00873_ ) );
AND3_X1 _16735_ ( .A1(_00640_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_00874_ ) );
AOI211_X1 _16736_ ( .A(_00873_ ), .B(_00874_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_06074_ ), .ZN(_00875_ ) );
NAND3_X1 _16737_ ( .A1(_05916_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_00876_ ) );
NAND4_X1 _16738_ ( .A1(_00875_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_00876_ ), .ZN(_00877_ ) );
NAND3_X1 _16739_ ( .A1(_00689_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_00878_ ) );
NAND3_X1 _16740_ ( .A1(fanout_net_14 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_00879_ ) );
AND2_X1 _16741_ ( .A1(_00878_ ), .A2(_00879_ ), .ZN(_00880_ ) );
NAND3_X1 _16742_ ( .A1(_00649_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_00881_ ) );
NAND3_X1 _16743_ ( .A1(_05905_ ), .A2(_00662_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_00882_ ) );
NAND4_X1 _16744_ ( .A1(_00880_ ), .A2(_00706_ ), .A3(_00881_ ), .A4(_00882_ ), .ZN(_00883_ ) );
NAND3_X1 _16745_ ( .A1(_00877_ ), .A2(_00654_ ), .A3(_00883_ ), .ZN(_00884_ ) );
NAND2_X1 _16746_ ( .A1(_00872_ ), .A2(_00884_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16747_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_00885_ ) );
AND3_X1 _16748_ ( .A1(_00640_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_00886_ ) );
AOI211_X1 _16749_ ( .A(_00885_ ), .B(_00886_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_00680_ ), .ZN(_00887_ ) );
NAND3_X1 _16750_ ( .A1(_00649_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_00888_ ) );
NAND4_X1 _16751_ ( .A1(_00887_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_00888_ ), .ZN(_00889_ ) );
NAND3_X1 _16752_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_00890_ ) );
NAND3_X1 _16753_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_00891_ ) );
AND2_X1 _16754_ ( .A1(_00890_ ), .A2(_00891_ ), .ZN(_00892_ ) );
NAND3_X1 _16755_ ( .A1(_00662_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_00893_ ) );
NAND3_X1 _16756_ ( .A1(_00689_ ), .A2(_00664_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_00894_ ) );
NAND4_X1 _16757_ ( .A1(_00892_ ), .A2(_00660_ ), .A3(_00893_ ), .A4(_00894_ ), .ZN(_00895_ ) );
NAND3_X1 _16758_ ( .A1(_00889_ ), .A2(_00654_ ), .A3(_00895_ ), .ZN(_00896_ ) );
OAI21_X1 _16759_ ( .A(\myifu.state [2] ), .B1(_00674_ ), .B2(_05663_ ), .ZN(_00897_ ) );
NOR3_X1 _16760_ ( .A1(_05995_ ), .A2(\myifu.data_in [11] ), .A3(_00676_ ), .ZN(_00898_ ) );
OAI21_X1 _16761_ ( .A(_00896_ ), .B1(_00897_ ), .B2(_00898_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
OR3_X1 _16762_ ( .A1(_00713_ ), .A2(\myifu.data_in [10] ), .A3(_00676_ ), .ZN(_00899_ ) );
OAI211_X1 _16763_ ( .A(_00899_ ), .B(\myifu.state [2] ), .C1(_05668_ ), .C2(_00674_ ), .ZN(_00900_ ) );
AND3_X1 _16764_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_00901_ ) );
AND3_X1 _16765_ ( .A1(_00640_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_00902_ ) );
AOI211_X1 _16766_ ( .A(_00901_ ), .B(_00902_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_06074_ ), .ZN(_00903_ ) );
NAND3_X1 _16767_ ( .A1(_05916_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_00904_ ) );
NAND4_X1 _16768_ ( .A1(_00903_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_00904_ ), .ZN(_00905_ ) );
NAND3_X1 _16769_ ( .A1(_00689_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_00906_ ) );
NAND3_X1 _16770_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_00907_ ) );
AND2_X1 _16771_ ( .A1(_00906_ ), .A2(_00907_ ), .ZN(_00908_ ) );
NAND3_X1 _16772_ ( .A1(_00649_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_00909_ ) );
NAND3_X1 _16773_ ( .A1(_05905_ ), .A2(_00662_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_00910_ ) );
NAND4_X1 _16774_ ( .A1(_00908_ ), .A2(_00706_ ), .A3(_00909_ ), .A4(_00910_ ), .ZN(_00911_ ) );
NAND3_X1 _16775_ ( .A1(_00905_ ), .A2(_00654_ ), .A3(_00911_ ), .ZN(_00912_ ) );
NAND2_X1 _16776_ ( .A1(_00900_ ), .A2(_00912_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
BUF_X4 _16777_ ( .A(_00711_ ), .Z(_00913_ ) );
NOR3_X1 _16778_ ( .A1(_00806_ ), .A2(\myifu.data_in [9] ), .A3(_00841_ ), .ZN(_00914_ ) );
BUF_X4 _16779_ ( .A(_00716_ ), .Z(_00915_ ) );
AOI211_X1 _16780_ ( .A(_00913_ ), .B(_00914_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .C2(_00915_ ), .ZN(_00916_ ) );
AND3_X1 _16781_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_00917_ ) );
AND3_X1 _16782_ ( .A1(_00810_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_00918_ ) );
AOI211_X1 _16783_ ( .A(_00917_ ), .B(_00918_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_00781_ ), .ZN(_00919_ ) );
NAND3_X1 _16784_ ( .A1(_00830_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_00920_ ) );
NAND4_X1 _16785_ ( .A1(_00919_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_00920_ ), .ZN(_00921_ ) );
NAND3_X1 _16786_ ( .A1(_00815_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_00922_ ) );
NAND3_X1 _16787_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_00923_ ) );
AND2_X1 _16788_ ( .A1(_00922_ ), .A2(_00923_ ), .ZN(_00924_ ) );
NAND3_X1 _16789_ ( .A1(_00819_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_00925_ ) );
NAND3_X1 _16790_ ( .A1(_05904_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_00926_ ) );
NAND4_X1 _16791_ ( .A1(_00924_ ), .A2(_00705_ ), .A3(_00925_ ), .A4(_00926_ ), .ZN(_00927_ ) );
AND3_X1 _16792_ ( .A1(_00921_ ), .A2(_00833_ ), .A3(_00927_ ), .ZN(_00928_ ) );
OR2_X1 _16793_ ( .A1(_00916_ ), .A2(_00928_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
AND3_X1 _16794_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_00929_ ) );
AND3_X1 _16795_ ( .A1(_00640_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_00930_ ) );
AOI211_X1 _16796_ ( .A(_00929_ ), .B(_00930_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_00680_ ), .ZN(_00931_ ) );
NAND3_X1 _16797_ ( .A1(_00649_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_00932_ ) );
NAND4_X1 _16798_ ( .A1(_00931_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_00932_ ), .ZN(_00933_ ) );
NAND3_X1 _16799_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_00934_ ) );
NAND3_X1 _16800_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_00935_ ) );
AND2_X1 _16801_ ( .A1(_00934_ ), .A2(_00935_ ), .ZN(_00936_ ) );
NAND3_X1 _16802_ ( .A1(_00662_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_00937_ ) );
NAND3_X1 _16803_ ( .A1(_00689_ ), .A2(_00664_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_00938_ ) );
NAND4_X1 _16804_ ( .A1(_00936_ ), .A2(_00660_ ), .A3(_00937_ ), .A4(_00938_ ), .ZN(_00939_ ) );
NAND3_X1 _16805_ ( .A1(_00933_ ), .A2(_00654_ ), .A3(_00939_ ), .ZN(_00940_ ) );
OAI21_X1 _16806_ ( .A(\myifu.state [2] ), .B1(_00674_ ), .B2(_05640_ ), .ZN(_00941_ ) );
NOR3_X1 _16807_ ( .A1(_05995_ ), .A2(\myifu.data_in [7] ), .A3(_00676_ ), .ZN(_00942_ ) );
OAI21_X1 _16808_ ( .A(_00940_ ), .B1(_00941_ ), .B2(_00942_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AND3_X1 _16809_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_00943_ ) );
AND3_X1 _16810_ ( .A1(_00640_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_00944_ ) );
AOI211_X1 _16811_ ( .A(_00943_ ), .B(_00944_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00680_ ), .ZN(_00945_ ) );
NAND3_X1 _16812_ ( .A1(_00649_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_00946_ ) );
NAND4_X1 _16813_ ( .A1(_00945_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_00946_ ), .ZN(_00947_ ) );
NAND3_X1 _16814_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_00948_ ) );
NAND3_X1 _16815_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_00949_ ) );
AND2_X1 _16816_ ( .A1(_00948_ ), .A2(_00949_ ), .ZN(_00950_ ) );
NAND3_X1 _16817_ ( .A1(_00664_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_00951_ ) );
NAND3_X1 _16818_ ( .A1(_00689_ ), .A2(_00664_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_00952_ ) );
NAND4_X1 _16819_ ( .A1(_00950_ ), .A2(_00660_ ), .A3(_00951_ ), .A4(_00952_ ), .ZN(_00953_ ) );
NAND3_X1 _16820_ ( .A1(_00947_ ), .A2(_00654_ ), .A3(_00953_ ), .ZN(_00954_ ) );
OAI21_X1 _16821_ ( .A(\myifu.state [2] ), .B1(_00674_ ), .B2(_05302_ ), .ZN(_00955_ ) );
NOR3_X1 _16822_ ( .A1(_05995_ ), .A2(\myifu.data_in [6] ), .A3(_00676_ ), .ZN(_00956_ ) );
OAI21_X1 _16823_ ( .A(_00954_ ), .B1(_00955_ ), .B2(_00956_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
NOR3_X1 _16824_ ( .A1(_00806_ ), .A2(\myifu.data_in [5] ), .A3(_00841_ ), .ZN(_00957_ ) );
AOI211_X1 _16825_ ( .A(_00913_ ), .B(_00957_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_00958_ ) );
AND3_X1 _16826_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_00959_ ) );
AND3_X1 _16827_ ( .A1(_00810_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_00960_ ) );
AOI211_X1 _16828_ ( .A(_00959_ ), .B(_00960_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00781_ ), .ZN(_00961_ ) );
NAND3_X1 _16829_ ( .A1(_00830_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_00962_ ) );
NAND4_X1 _16830_ ( .A1(_00961_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_00962_ ), .ZN(_00963_ ) );
NAND3_X1 _16831_ ( .A1(_00815_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_00964_ ) );
NAND3_X1 _16832_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_00965_ ) );
AND2_X1 _16833_ ( .A1(_00964_ ), .A2(_00965_ ), .ZN(_00966_ ) );
NAND3_X1 _16834_ ( .A1(_00819_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_00967_ ) );
NAND3_X1 _16835_ ( .A1(_05904_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_00968_ ) );
NAND4_X1 _16836_ ( .A1(_00966_ ), .A2(_00705_ ), .A3(_00967_ ), .A4(_00968_ ), .ZN(_00969_ ) );
AND3_X1 _16837_ ( .A1(_00963_ ), .A2(_00833_ ), .A3(_00969_ ), .ZN(_00970_ ) );
OR2_X1 _16838_ ( .A1(_00958_ ), .A2(_00970_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
NOR3_X1 _16839_ ( .A1(_00806_ ), .A2(\myifu.data_in [4] ), .A3(_00841_ ), .ZN(_00971_ ) );
AOI211_X1 _16840_ ( .A(_00913_ ), .B(_00971_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_00972_ ) );
AND3_X1 _16841_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_00973_ ) );
AND3_X1 _16842_ ( .A1(_00810_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_00974_ ) );
AOI211_X1 _16843_ ( .A(_00973_ ), .B(_00974_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00781_ ), .ZN(_00975_ ) );
NAND3_X1 _16844_ ( .A1(_00830_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_00976_ ) );
NAND4_X1 _16845_ ( .A1(_00975_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_00976_ ), .ZN(_00977_ ) );
NAND3_X1 _16846_ ( .A1(_00815_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_00978_ ) );
NAND3_X1 _16847_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_00979_ ) );
AND2_X1 _16848_ ( .A1(_00978_ ), .A2(_00979_ ), .ZN(_00980_ ) );
NAND3_X1 _16849_ ( .A1(_00819_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_00981_ ) );
NAND3_X1 _16850_ ( .A1(_05904_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_00982_ ) );
NAND4_X1 _16851_ ( .A1(_00980_ ), .A2(_00705_ ), .A3(_00981_ ), .A4(_00982_ ), .ZN(_00983_ ) );
AND3_X1 _16852_ ( .A1(_00977_ ), .A2(_00833_ ), .A3(_00983_ ), .ZN(_00984_ ) );
OR2_X1 _16853_ ( .A1(_00972_ ), .A2(_00984_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
NOR3_X1 _16854_ ( .A1(_00806_ ), .A2(\myifu.data_in [3] ), .A3(_00841_ ), .ZN(_00985_ ) );
AOI211_X1 _16855_ ( .A(_00913_ ), .B(_00985_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_00986_ ) );
AND3_X1 _16856_ ( .A1(fanout_net_15 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_00987_ ) );
AND3_X1 _16857_ ( .A1(_00810_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_00988_ ) );
AOI211_X1 _16858_ ( .A(_00987_ ), .B(_00988_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00781_ ), .ZN(_00989_ ) );
NAND3_X1 _16859_ ( .A1(_00830_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_00990_ ) );
NAND4_X1 _16860_ ( .A1(_00989_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_00990_ ), .ZN(_00991_ ) );
NAND3_X1 _16861_ ( .A1(_00815_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_00992_ ) );
NAND3_X1 _16862_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_00993_ ) );
AND2_X1 _16863_ ( .A1(_00992_ ), .A2(_00993_ ), .ZN(_00994_ ) );
NAND3_X1 _16864_ ( .A1(_00819_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_00995_ ) );
NAND3_X1 _16865_ ( .A1(_05904_ ), .A2(_00773_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_00996_ ) );
NAND4_X1 _16866_ ( .A1(_00994_ ), .A2(_00705_ ), .A3(_00995_ ), .A4(_00996_ ), .ZN(_00997_ ) );
AND3_X1 _16867_ ( .A1(_00991_ ), .A2(_00833_ ), .A3(_00997_ ), .ZN(_00998_ ) );
OR2_X1 _16868_ ( .A1(_00986_ ), .A2(_00998_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
NOR3_X1 _16869_ ( .A1(_00806_ ), .A2(\myifu.data_in [2] ), .A3(_00841_ ), .ZN(_00999_ ) );
AOI211_X1 _16870_ ( .A(_00913_ ), .B(_00999_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_01000_ ) );
AND3_X1 _16871_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_01001_ ) );
AND3_X1 _16872_ ( .A1(_00810_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_01002_ ) );
AOI211_X1 _16873_ ( .A(_01001_ ), .B(_01002_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_00781_ ), .ZN(_01003_ ) );
NAND3_X1 _16874_ ( .A1(_00830_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_01004_ ) );
NAND4_X1 _16875_ ( .A1(_01003_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_01004_ ), .ZN(_01005_ ) );
NAND3_X1 _16876_ ( .A1(_00815_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_01006_ ) );
NAND3_X1 _16877_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_01007_ ) );
AND2_X1 _16878_ ( .A1(_01006_ ), .A2(_01007_ ), .ZN(_01008_ ) );
NAND3_X1 _16879_ ( .A1(_00819_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_01009_ ) );
NAND3_X1 _16880_ ( .A1(_05904_ ), .A2(_05914_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_01010_ ) );
NAND4_X1 _16881_ ( .A1(_01008_ ), .A2(_00705_ ), .A3(_01009_ ), .A4(_01010_ ), .ZN(_01011_ ) );
AND3_X1 _16882_ ( .A1(_01005_ ), .A2(_00833_ ), .A3(_01011_ ), .ZN(_01012_ ) );
OR2_X1 _16883_ ( .A1(_01000_ ), .A2(_01012_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
NOR3_X1 _16884_ ( .A1(_00806_ ), .A2(\myifu.data_in [1] ), .A3(_00841_ ), .ZN(_01013_ ) );
AOI211_X1 _16885_ ( .A(_00913_ ), .B(_01013_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_01014_ ) );
AND3_X1 _16886_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01015_ ) );
AND3_X1 _16887_ ( .A1(_00810_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01016_ ) );
AOI211_X1 _16888_ ( .A(_01015_ ), .B(_01016_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_06073_ ), .ZN(_01017_ ) );
NAND3_X1 _16889_ ( .A1(_00830_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01018_ ) );
NAND4_X1 _16890_ ( .A1(_01017_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_01018_ ), .ZN(_01019_ ) );
NAND3_X1 _16891_ ( .A1(_00815_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01020_ ) );
NAND3_X1 _16892_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01021_ ) );
AND2_X1 _16893_ ( .A1(_01020_ ), .A2(_01021_ ), .ZN(_01022_ ) );
NAND3_X1 _16894_ ( .A1(_00819_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01023_ ) );
NAND3_X1 _16895_ ( .A1(_05904_ ), .A2(_05914_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01024_ ) );
NAND4_X1 _16896_ ( .A1(_01022_ ), .A2(_00705_ ), .A3(_01023_ ), .A4(_01024_ ), .ZN(_01025_ ) );
AND3_X1 _16897_ ( .A1(_01019_ ), .A2(_00833_ ), .A3(_01025_ ), .ZN(_01026_ ) );
OR2_X1 _16898_ ( .A1(_01014_ ), .A2(_01026_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
OR3_X1 _16899_ ( .A1(_00713_ ), .A2(\myifu.data_in [28] ), .A3(_00714_ ), .ZN(_01027_ ) );
OAI211_X1 _16900_ ( .A(_01027_ ), .B(\myifu.state [2] ), .C1(_05701_ ), .C2(_00673_ ), .ZN(_01028_ ) );
AND3_X1 _16901_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01029_ ) );
AND3_X1 _16902_ ( .A1(_00640_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01030_ ) );
AOI211_X1 _16903_ ( .A(_01029_ ), .B(_01030_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_06074_ ), .ZN(_01031_ ) );
NAND3_X1 _16904_ ( .A1(_05916_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01032_ ) );
NAND4_X1 _16905_ ( .A1(_01031_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_01032_ ), .ZN(_01033_ ) );
NAND3_X1 _16906_ ( .A1(_00689_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01034_ ) );
NAND3_X1 _16907_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01035_ ) );
AND2_X1 _16908_ ( .A1(_01034_ ), .A2(_01035_ ), .ZN(_01036_ ) );
NAND3_X1 _16909_ ( .A1(_00649_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01037_ ) );
NAND3_X1 _16910_ ( .A1(_05905_ ), .A2(_00662_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01038_ ) );
NAND4_X1 _16911_ ( .A1(_01036_ ), .A2(_00660_ ), .A3(_01037_ ), .A4(_01038_ ), .ZN(_01039_ ) );
NAND3_X1 _16912_ ( .A1(_01033_ ), .A2(_00654_ ), .A3(_01039_ ), .ZN(_01040_ ) );
NAND2_X1 _16913_ ( .A1(_01028_ ), .A2(_01040_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
NOR3_X1 _16914_ ( .A1(_05994_ ), .A2(\myifu.data_in [0] ), .A3(_00841_ ), .ZN(_01041_ ) );
AOI211_X1 _16915_ ( .A(_00913_ ), .B(_01041_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_01042_ ) );
AND3_X1 _16916_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01043_ ) );
AND3_X1 _16917_ ( .A1(_05902_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01044_ ) );
AOI211_X1 _16918_ ( .A(_01043_ ), .B(_01044_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_06073_ ), .ZN(_01045_ ) );
NAND3_X1 _16919_ ( .A1(_00830_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01046_ ) );
NAND4_X1 _16920_ ( .A1(_01045_ ), .A2(_00847_ ), .A3(_00829_ ), .A4(_01046_ ), .ZN(_01047_ ) );
NAND3_X1 _16921_ ( .A1(_05903_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01048_ ) );
NAND3_X1 _16922_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01049_ ) );
AND2_X1 _16923_ ( .A1(_01048_ ), .A2(_01049_ ), .ZN(_01050_ ) );
NAND3_X1 _16924_ ( .A1(_05915_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01051_ ) );
NAND3_X1 _16925_ ( .A1(_05904_ ), .A2(_05914_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01052_ ) );
NAND4_X1 _16926_ ( .A1(_01050_ ), .A2(_00705_ ), .A3(_01051_ ), .A4(_01052_ ), .ZN(_01053_ ) );
AND3_X1 _16927_ ( .A1(_01047_ ), .A2(_00833_ ), .A3(_01053_ ), .ZN(_01054_ ) );
OR2_X1 _16928_ ( .A1(_01042_ ), .A2(_01054_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
AND3_X1 _16929_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01055_ ) );
AND3_X1 _16930_ ( .A1(_00640_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01056_ ) );
AOI211_X1 _16931_ ( .A(_01055_ ), .B(_01056_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00680_ ), .ZN(_01057_ ) );
NAND3_X1 _16932_ ( .A1(_00649_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01058_ ) );
NAND4_X1 _16933_ ( .A1(_01057_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_01058_ ), .ZN(_01059_ ) );
NAND3_X1 _16934_ ( .A1(_00655_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01060_ ) );
NAND3_X1 _16935_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01061_ ) );
AND2_X1 _16936_ ( .A1(_01060_ ), .A2(_01061_ ), .ZN(_01062_ ) );
NAND3_X1 _16937_ ( .A1(_00664_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01063_ ) );
NAND3_X1 _16938_ ( .A1(_00689_ ), .A2(_00664_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01064_ ) );
NAND4_X1 _16939_ ( .A1(_01062_ ), .A2(_00660_ ), .A3(_01063_ ), .A4(_01064_ ), .ZN(_01065_ ) );
NAND3_X1 _16940_ ( .A1(_01059_ ), .A2(_00653_ ), .A3(_01065_ ), .ZN(_01066_ ) );
OAI21_X1 _16941_ ( .A(\myifu.state [2] ), .B1(_00674_ ), .B2(_05692_ ), .ZN(_01067_ ) );
NOR3_X1 _16942_ ( .A1(_05995_ ), .A2(\myifu.data_in [27] ), .A3(_00676_ ), .ZN(_01068_ ) );
OAI21_X1 _16943_ ( .A(_01066_ ), .B1(_01067_ ), .B2(_01068_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
OR3_X1 _16944_ ( .A1(_00713_ ), .A2(\myifu.data_in [26] ), .A3(_00714_ ), .ZN(_01069_ ) );
OAI211_X1 _16945_ ( .A(_01069_ ), .B(\myifu.state [2] ), .C1(_05655_ ), .C2(_00673_ ), .ZN(_01070_ ) );
AND3_X1 _16946_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01071_ ) );
AND3_X1 _16947_ ( .A1(_00640_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01072_ ) );
AOI211_X1 _16948_ ( .A(_01071_ ), .B(_01072_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_06074_ ), .ZN(_01073_ ) );
NAND3_X1 _16949_ ( .A1(_05916_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01074_ ) );
NAND4_X1 _16950_ ( .A1(_01073_ ), .A2(_00644_ ), .A3(_00647_ ), .A4(_01074_ ), .ZN(_01075_ ) );
NAND3_X1 _16951_ ( .A1(_00655_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01076_ ) );
NAND3_X1 _16952_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01077_ ) );
AND2_X1 _16953_ ( .A1(_01076_ ), .A2(_01077_ ), .ZN(_01078_ ) );
NAND3_X1 _16954_ ( .A1(_00649_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01079_ ) );
NAND3_X1 _16955_ ( .A1(_05905_ ), .A2(_00662_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01080_ ) );
NAND4_X1 _16956_ ( .A1(_01078_ ), .A2(_00660_ ), .A3(_01079_ ), .A4(_01080_ ), .ZN(_01081_ ) );
NAND3_X1 _16957_ ( .A1(_01075_ ), .A2(_00654_ ), .A3(_01081_ ), .ZN(_01082_ ) );
NAND2_X1 _16958_ ( .A1(_01070_ ), .A2(_01082_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
AND3_X1 _16959_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01083_ ) );
AND3_X1 _16960_ ( .A1(_00688_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01084_ ) );
AOI211_X1 _16961_ ( .A(_01083_ ), .B(_01084_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00680_ ), .ZN(_01085_ ) );
NAND3_X1 _16962_ ( .A1(_00662_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01086_ ) );
NAND4_X1 _16963_ ( .A1(_01085_ ), .A2(_00722_ ), .A3(_00646_ ), .A4(_01086_ ), .ZN(_01087_ ) );
NAND3_X1 _16964_ ( .A1(_00655_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01088_ ) );
NAND3_X1 _16965_ ( .A1(fanout_net_16 ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01089_ ) );
AND2_X1 _16966_ ( .A1(_01088_ ), .A2(_01089_ ), .ZN(_01090_ ) );
NAND3_X1 _16967_ ( .A1(_00664_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01091_ ) );
NAND3_X1 _16968_ ( .A1(_00689_ ), .A2(_00664_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01092_ ) );
NAND4_X1 _16969_ ( .A1(_01090_ ), .A2(_00660_ ), .A3(_01091_ ), .A4(_01092_ ), .ZN(_01093_ ) );
NAND3_X1 _16970_ ( .A1(_01087_ ), .A2(_00653_ ), .A3(_01093_ ), .ZN(_01094_ ) );
OAI21_X1 _16971_ ( .A(\myifu.state [2] ), .B1(_00674_ ), .B2(_05659_ ), .ZN(_01095_ ) );
NOR3_X1 _16972_ ( .A1(_05995_ ), .A2(\myifu.data_in [25] ), .A3(_00676_ ), .ZN(_01096_ ) );
OAI21_X1 _16973_ ( .A(_01094_ ), .B1(_01095_ ), .B2(_01096_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
NOR3_X1 _16974_ ( .A1(_05994_ ), .A2(\myifu.data_in [24] ), .A3(_00841_ ), .ZN(_01097_ ) );
AOI211_X1 _16975_ ( .A(_00913_ ), .B(_01097_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_01098_ ) );
AND3_X1 _16976_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01099_ ) );
AND3_X1 _16977_ ( .A1(_05902_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01100_ ) );
AOI211_X1 _16978_ ( .A(_01099_ ), .B(_01100_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_06073_ ), .ZN(_01101_ ) );
NAND3_X1 _16979_ ( .A1(_00661_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01102_ ) );
NAND4_X1 _16980_ ( .A1(_01101_ ), .A2(_00847_ ), .A3(_00645_ ), .A4(_01102_ ), .ZN(_01103_ ) );
NAND3_X1 _16981_ ( .A1(_05903_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01104_ ) );
NAND3_X1 _16982_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01105_ ) );
AND2_X1 _16983_ ( .A1(_01104_ ), .A2(_01105_ ), .ZN(_01106_ ) );
NAND3_X1 _16984_ ( .A1(_05915_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01107_ ) );
NAND3_X1 _16985_ ( .A1(_05904_ ), .A2(_05914_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01108_ ) );
NAND4_X1 _16986_ ( .A1(_01106_ ), .A2(_00705_ ), .A3(_01107_ ), .A4(_01108_ ), .ZN(_01109_ ) );
AND3_X1 _16987_ ( .A1(_01103_ ), .A2(_00652_ ), .A3(_01109_ ), .ZN(_01110_ ) );
OR2_X1 _16988_ ( .A1(_01098_ ), .A2(_01110_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
NOR3_X1 _16989_ ( .A1(_05994_ ), .A2(\myifu.data_in [23] ), .A3(_00672_ ), .ZN(_01111_ ) );
AOI211_X1 _16990_ ( .A(_00913_ ), .B(_01111_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00915_ ), .ZN(_01112_ ) );
NAND3_X1 _16991_ ( .A1(_00688_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01113_ ) );
NAND3_X1 _16992_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01114_ ) );
AND2_X1 _16993_ ( .A1(_01113_ ), .A2(_01114_ ), .ZN(_01115_ ) );
NAND3_X1 _16994_ ( .A1(_00648_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01116_ ) );
NAND3_X1 _16995_ ( .A1(_00655_ ), .A2(_00661_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01117_ ) );
NAND4_X1 _16996_ ( .A1(_01115_ ), .A2(_00728_ ), .A3(_01116_ ), .A4(_01117_ ), .ZN(_01118_ ) );
AND3_X1 _16997_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01119_ ) );
AND3_X1 _16998_ ( .A1(_05902_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01120_ ) );
AOI211_X1 _16999_ ( .A(_01119_ ), .B(_01120_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_06073_ ), .ZN(_01121_ ) );
NAND3_X1 _17000_ ( .A1(_05915_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01122_ ) );
NAND4_X1 _17001_ ( .A1(_01121_ ), .A2(_00643_ ), .A3(_00645_ ), .A4(_01122_ ), .ZN(_01123_ ) );
AND3_X1 _17002_ ( .A1(_01118_ ), .A2(_00652_ ), .A3(_01123_ ), .ZN(_01124_ ) );
OR2_X1 _17003_ ( .A1(_01112_ ), .A2(_01124_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
NOR3_X1 _17004_ ( .A1(_05994_ ), .A2(\myifu.data_in [22] ), .A3(_00672_ ), .ZN(_01125_ ) );
AOI211_X1 _17005_ ( .A(_00913_ ), .B(_01125_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .C2(_00915_ ), .ZN(_01126_ ) );
NAND3_X1 _17006_ ( .A1(_00688_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01127_ ) );
NAND3_X1 _17007_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01128_ ) );
AND2_X1 _17008_ ( .A1(_01127_ ), .A2(_01128_ ), .ZN(_01129_ ) );
NAND3_X1 _17009_ ( .A1(_00648_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01130_ ) );
NAND3_X1 _17010_ ( .A1(_00730_ ), .A2(_00661_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01131_ ) );
NAND4_X1 _17011_ ( .A1(_01129_ ), .A2(_00728_ ), .A3(_01130_ ), .A4(_01131_ ), .ZN(_01132_ ) );
AND3_X1 _17012_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01133_ ) );
AND3_X1 _17013_ ( .A1(_05902_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01134_ ) );
AOI211_X1 _17014_ ( .A(_01133_ ), .B(_01134_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_06073_ ), .ZN(_01135_ ) );
NAND3_X1 _17015_ ( .A1(_05915_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01136_ ) );
NAND4_X1 _17016_ ( .A1(_01135_ ), .A2(_00643_ ), .A3(_00645_ ), .A4(_01136_ ), .ZN(_01137_ ) );
AND3_X1 _17017_ ( .A1(_01132_ ), .A2(_00652_ ), .A3(_01137_ ), .ZN(_01138_ ) );
OR2_X1 _17018_ ( .A1(_01126_ ), .A2(_01138_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI211_X1 _17019_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_05428_ ), .C1(_05781_ ), .C2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
AND3_X1 _17020_ ( .A1(_05985_ ), .A2(\myifu.state [2] ), .A3(_05993_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _17021_ ( .A(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .B1(io_master_rlast ), .B2(_00564_ ), .ZN(_01139_ ) );
INV_X1 _17022_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01140_ ) );
AND4_X1 _17023_ ( .A1(_01140_ ), .A2(_01898_ ), .A3(\myifu.state [0] ), .A4(_01964_ ), .ZN(_01141_ ) );
NOR2_X1 _17024_ ( .A1(_01141_ ), .A2(_00508_ ), .ZN(_01142_ ) );
AOI21_X1 _17025_ ( .A(fanout_net_4 ), .B1(_01139_ ), .B2(_01142_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _17026_ ( .A(_01140_ ), .B(_01988_ ), .C1(_05182_ ), .C2(_06095_ ), .ZN(_01143_ ) );
NAND2_X1 _17027_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01144_ ) );
NAND4_X1 _17028_ ( .A1(_01143_ ), .A2(_01585_ ), .A3(_05906_ ), .A4(_01144_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _17029_ ( .A(_01584_ ), .B(\myifu.state [2] ), .C1(_05995_ ), .C2(_05996_ ), .ZN(_01145_ ) );
NOR2_X1 _17030_ ( .A1(_05182_ ), .A2(_06094_ ), .ZN(_01146_ ) );
NAND3_X1 _17031_ ( .A1(_01146_ ), .A2(_01988_ ), .A3(_02056_ ), .ZN(_01147_ ) );
NAND2_X1 _17032_ ( .A1(_01145_ ), .A2(_01147_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
NOR4_X1 _17033_ ( .A1(_00706_ ), .A2(_02057_ ), .A3(_06077_ ), .A4(_06078_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NOR4_X1 _17034_ ( .A1(_00706_ ), .A2(_02057_ ), .A3(_06077_ ), .A4(_00613_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _17035_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00706_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17036_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(_05916_ ), .A4(_00706_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _17037_ ( .A1(_00706_ ), .A2(_02057_ ), .A3(_06076_ ), .A4(_06075_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17038_ ( .A1(_05905_ ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00706_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
AND3_X1 _17039_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06074_ ), .A3(_00706_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17040_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06074_ ), .A3(_00644_ ), .A4(_00647_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
NOR3_X1 _17041_ ( .A1(_02057_ ), .A2(_06075_ ), .A3(_06077_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
NOR3_X1 _17042_ ( .A1(_02057_ ), .A2(_06078_ ), .A3(_06077_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
NOR3_X1 _17043_ ( .A1(_02057_ ), .A2(_06077_ ), .A3(_00613_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
AND3_X1 _17044_ ( .A1(_02056_ ), .A2(_06074_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
NOR2_X1 _17045_ ( .A1(_01146_ ), .A2(_01966_ ), .ZN(_01148_ ) );
AND2_X1 _17046_ ( .A1(_01965_ ), .A2(\myifu.state [0] ), .ZN(_01149_ ) );
OAI21_X1 _17047_ ( .A(\myifu.state [1] ), .B1(_05507_ ), .B2(_05587_ ), .ZN(_01150_ ) );
NAND2_X1 _17048_ ( .A1(_00510_ ), .A2(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01151_ ) );
NAND3_X1 _17049_ ( .A1(_01150_ ), .A2(_01151_ ), .A3(_01144_ ), .ZN(_01152_ ) );
OR3_X1 _17050_ ( .A1(_01148_ ), .A2(_01149_ ), .A3(_01152_ ), .ZN(_01153_ ) );
AOI21_X1 _17051_ ( .A(_01153_ ), .B1(_05997_ ), .B2(_01968_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17052_ ( .A1(_05793_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_05430_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _17053_ ( .A1(_05253_ ), .A2(_05255_ ), .A3(_05257_ ), .A4(_05260_ ), .ZN(_01154_ ) );
AND2_X1 _17054_ ( .A1(_05294_ ), .A2(_01154_ ), .ZN(_01155_ ) );
INV_X1 _17055_ ( .A(_01155_ ), .ZN(_01156_ ) );
AOI211_X1 _17056_ ( .A(_05507_ ), .B(_00484_ ), .C1(_05208_ ), .C2(_01156_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
NOR3_X1 _17057_ ( .A1(_01988_ ), .A2(fanout_net_4 ), .A3(_01152_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _17058_ ( .A(_06137_ ), .B(_05187_ ), .S(\mylsu.state [0] ), .Z(_01157_ ) );
NOR2_X1 _17059_ ( .A1(_06142_ ), .A2(_01157_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17060_ ( .A(_06006_ ), .ZN(_01158_ ) );
NOR3_X1 _17061_ ( .A1(_06142_ ), .A2(_01158_ ), .A3(_01157_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
AND2_X1 _17062_ ( .A1(_06020_ ), .A2(_00487_ ), .ZN(_01159_ ) );
AND3_X1 _17063_ ( .A1(_05186_ ), .A2(\mylsu.state [0] ), .A3(_01159_ ), .ZN(_01160_ ) );
NAND3_X1 _17064_ ( .A1(_01160_ ), .A2(_02037_ ), .A3(_06061_ ), .ZN(_01161_ ) );
AND2_X1 _17065_ ( .A1(_05979_ ), .A2(_06141_ ), .ZN(_01162_ ) );
OAI21_X1 _17066_ ( .A(_01161_ ), .B1(_01162_ ), .B2(_06070_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND3_X1 _17067_ ( .A1(_06006_ ), .A2(\mylsu.state [0] ), .A3(_00487_ ), .ZN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
INV_X1 _17068_ ( .A(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .ZN(_01163_ ) );
NOR2_X1 _17069_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01164_ ) );
NOR4_X1 _17070_ ( .A1(_02105_ ), .A2(_05191_ ), .A3(_01163_ ), .A4(_01164_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OR3_X1 _17071_ ( .A1(_01158_ ), .A2(_06134_ ), .A3(io_master_wready ), .ZN(_01165_ ) );
AND2_X1 _17072_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01166_ ) );
NOR2_X1 _17073_ ( .A1(_06014_ ), .A2(_01166_ ), .ZN(_01167_ ) );
BUF_X2 _17074_ ( .A(_02040_ ), .Z(_01168_ ) );
AND4_X1 _17075_ ( .A1(io_master_awready ), .A2(_01167_ ), .A3(_01168_ ), .A4(_06049_ ), .ZN(_01169_ ) );
NAND2_X1 _17076_ ( .A1(_01169_ ), .A2(\mylsu.state [0] ), .ZN(_01170_ ) );
OAI21_X1 _17077_ ( .A(_01165_ ), .B1(_02105_ ), .B2(_01170_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
BUF_X2 _17078_ ( .A(_02040_ ), .Z(_01171_ ) );
NAND4_X1 _17079_ ( .A1(_06060_ ), .A2(_01171_ ), .A3(EXU_valid_LSU ), .A4(_01166_ ), .ZN(_01172_ ) );
NOR4_X1 _17080_ ( .A1(_02041_ ), .A2(_02047_ ), .A3(_01158_ ), .A4(_01172_ ), .ZN(_01173_ ) );
NAND2_X1 _17081_ ( .A1(_01173_ ), .A2(\mylsu.state [0] ), .ZN(_01174_ ) );
NAND3_X1 _17082_ ( .A1(_06006_ ), .A2(\mylsu.state [4] ), .A3(io_master_awready ), .ZN(_01175_ ) );
NAND3_X1 _17083_ ( .A1(_06006_ ), .A2(\mylsu.state [2] ), .A3(io_master_wready ), .ZN(_01176_ ) );
NAND3_X1 _17084_ ( .A1(_06148_ ), .A2(\mylsu.state [1] ), .A3(_06006_ ), .ZN(_01177_ ) );
NAND4_X1 _17085_ ( .A1(_01174_ ), .A2(_01175_ ), .A3(_01176_ ), .A4(_01177_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
NOR4_X1 _17086_ ( .A1(_06124_ ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .A4(\EX_LS_typ [0] ), .ZN(_01178_ ) );
NAND4_X1 _17087_ ( .A1(_02021_ ), .A2(_01178_ ), .A3(\EX_LS_dest_csreg_mem [0] ), .A4(_02034_ ), .ZN(_01179_ ) );
NAND4_X1 _17088_ ( .A1(_02035_ ), .A2(_02026_ ), .A3(\EX_LS_typ [2] ), .A4(_02027_ ), .ZN(_01180_ ) );
OAI21_X1 _17089_ ( .A(_01179_ ), .B1(_02024_ ), .B2(_01180_ ), .ZN(_01181_ ) );
NAND3_X1 _17090_ ( .A1(_02019_ ), .A2(_06020_ ), .A3(_06005_ ), .ZN(_01182_ ) );
AND4_X1 _17091_ ( .A1(\EX_LS_typ [1] ), .A2(_02035_ ), .A3(\EX_LS_typ [0] ), .A4(_02029_ ), .ZN(_01183_ ) );
AOI211_X1 _17092_ ( .A(_01181_ ), .B(_01182_ ), .C1(\EX_LS_dest_csreg_mem [0] ), .C2(_01183_ ), .ZN(_01184_ ) );
AND3_X1 _17093_ ( .A1(_01184_ ), .A2(\mylsu.state [0] ), .A3(_01159_ ), .ZN(_01185_ ) );
NOR3_X1 _17094_ ( .A1(_05186_ ), .A2(_02005_ ), .A3(_05188_ ), .ZN(_01186_ ) );
AND4_X1 _17095_ ( .A1(\mylsu.state [0] ), .A2(_01186_ ), .A3(_02037_ ), .A4(_06061_ ), .ZN(_01187_ ) );
AOI22_X1 _17096_ ( .A1(_02039_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .B1(_02020_ ), .B2(_01972_ ), .ZN(_01188_ ) );
AND4_X1 _17097_ ( .A1(_00487_ ), .A2(_06060_ ), .A3(_01188_ ), .A4(_06006_ ), .ZN(_01189_ ) );
AOI211_X1 _17098_ ( .A(_01185_ ), .B(_01187_ ), .C1(\mylsu.state [0] ), .C2(_01189_ ), .ZN(_01190_ ) );
NAND3_X1 _17099_ ( .A1(_05979_ ), .A2(_00283_ ), .A3(_06141_ ), .ZN(_01191_ ) );
AND4_X1 _17100_ ( .A1(_01171_ ), .A2(_01167_ ), .A3(_06049_ ), .A4(_01164_ ), .ZN(_01192_ ) );
NAND3_X1 _17101_ ( .A1(_02048_ ), .A2(\mylsu.state [0] ), .A3(_01192_ ), .ZN(_01193_ ) );
AND3_X1 _17102_ ( .A1(_06005_ ), .A2(_00487_ ), .A3(_02021_ ), .ZN(_01194_ ) );
NAND4_X1 _17103_ ( .A1(_01194_ ), .A2(_02033_ ), .A3(_02034_ ), .A4(_02021_ ), .ZN(_01195_ ) );
NAND4_X1 _17104_ ( .A1(_02019_ ), .A2(_06061_ ), .A3(EXU_valid_LSU ), .A4(_02040_ ), .ZN(_01196_ ) );
OAI21_X1 _17105_ ( .A(_01195_ ), .B1(_01196_ ), .B2(_02047_ ), .ZN(_01197_ ) );
NAND2_X1 _17106_ ( .A1(_01197_ ), .A2(\mylsu.state [0] ), .ZN(_01198_ ) );
NAND2_X1 _17107_ ( .A1(_01198_ ), .A2(_06006_ ), .ZN(_01199_ ) );
NAND3_X1 _17108_ ( .A1(_02047_ ), .A2(_02040_ ), .A3(_06006_ ), .ZN(_01200_ ) );
NAND3_X1 _17109_ ( .A1(_01200_ ), .A2(EXU_valid_LSU ), .A3(_06060_ ), .ZN(_01201_ ) );
AOI221_X4 _17110_ ( .A(_01199_ ), .B1(\mylsu.state [1] ), .B2(_06147_ ), .C1(\mylsu.state [0] ), .C2(_01201_ ), .ZN(_01202_ ) );
NAND4_X1 _17111_ ( .A1(_01190_ ), .A2(_01191_ ), .A3(_01193_ ), .A4(_01202_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND4_X1 _17112_ ( .A1(_02048_ ), .A2(io_master_wready ), .A3(_06129_ ), .A4(_01167_ ), .ZN(_01203_ ) );
AOI211_X1 _17113_ ( .A(io_master_awready ), .B(_01158_ ), .C1(_01203_ ), .C2(_06133_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
BUF_X4 _17114_ ( .A(_06015_ ), .Z(_01204_ ) );
BUF_X4 _17115_ ( .A(_01204_ ), .Z(_01205_ ) );
AOI21_X1 _17116_ ( .A(\EX_LS_pc [21] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01206_ ) );
BUF_X4 _17117_ ( .A(_02174_ ), .Z(_01207_ ) );
OAI21_X1 _17118_ ( .A(_01204_ ), .B1(_01207_ ), .B2(_05138_ ), .ZN(_01208_ ) );
BUF_X4 _17119_ ( .A(_02174_ ), .Z(_01209_ ) );
AOI221_X4 _17120_ ( .A(_01208_ ), .B1(\LS_WB_wdata_csreg [21] ), .B2(_01209_ ), .C1(_02105_ ), .C2(_01168_ ), .ZN(_01210_ ) );
NOR2_X1 _17121_ ( .A1(_01206_ ), .A2(_01210_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _17122_ ( .A(\LS_WB_wdata_csreg [20] ), .B(\EX_LS_result_csreg_mem [20] ), .S(_02173_ ), .Z(_01211_ ) );
MUX2_X1 _17123_ ( .A(_01211_ ), .B(\EX_LS_pc [20] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
OAI22_X1 _17124_ ( .A1(_06019_ ), .A2(_02095_ ), .B1(_06024_ ), .B2(_06168_ ), .ZN(_01212_ ) );
MUX2_X1 _17125_ ( .A(_01212_ ), .B(\EX_LS_pc [19] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
OAI22_X1 _17126_ ( .A1(_06019_ ), .A2(_02096_ ), .B1(_06024_ ), .B2(_06170_ ), .ZN(_01213_ ) );
MUX2_X1 _17127_ ( .A(_01213_ ), .B(\EX_LS_pc [18] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
OAI22_X1 _17128_ ( .A1(_06019_ ), .A2(_02097_ ), .B1(_06024_ ), .B2(_04643_ ), .ZN(_01214_ ) );
MUX2_X1 _17129_ ( .A(_01214_ ), .B(\EX_LS_pc [17] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _17130_ ( .A(\EX_LS_pc [16] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01215_ ) );
OAI21_X1 _17131_ ( .A(_01204_ ), .B1(_01207_ ), .B2(_04664_ ), .ZN(_01216_ ) );
AOI221_X4 _17132_ ( .A(_01216_ ), .B1(\LS_WB_wdata_csreg [16] ), .B2(_01209_ ), .C1(_02105_ ), .C2(_01168_ ), .ZN(_01217_ ) );
NOR2_X1 _17133_ ( .A1(_01215_ ), .A2(_01217_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
AOI221_X4 _17134_ ( .A(_06016_ ), .B1(\LS_WB_wdata_csreg [15] ), .B2(_01209_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [15] ), .ZN(_01218_ ) );
BUF_X4 _17135_ ( .A(_06010_ ), .Z(_01219_ ) );
BUF_X4 _17136_ ( .A(_01204_ ), .Z(_01220_ ) );
AOI21_X1 _17137_ ( .A(\EX_LS_pc [15] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01221_ ) );
NOR2_X1 _17138_ ( .A1(_01218_ ), .A2(_01221_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _17139_ ( .A(\EX_LS_pc [14] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01222_ ) );
OAI21_X1 _17140_ ( .A(_01204_ ), .B1(_01207_ ), .B2(_04708_ ), .ZN(_01223_ ) );
AOI221_X4 _17141_ ( .A(_01223_ ), .B1(\LS_WB_wdata_csreg [14] ), .B2(_01209_ ), .C1(_02105_ ), .C2(_01168_ ), .ZN(_01224_ ) );
NOR2_X1 _17142_ ( .A1(_01222_ ), .A2(_01224_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
AOI21_X1 _17143_ ( .A(\EX_LS_pc [13] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01225_ ) );
OAI21_X1 _17144_ ( .A(_01204_ ), .B1(_01207_ ), .B2(_04733_ ), .ZN(_01226_ ) );
AOI221_X4 _17145_ ( .A(_01226_ ), .B1(\LS_WB_wdata_csreg [13] ), .B2(_01209_ ), .C1(_02105_ ), .C2(_01168_ ), .ZN(_01227_ ) );
NOR2_X1 _17146_ ( .A1(_01225_ ), .A2(_01227_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
OAI22_X1 _17147_ ( .A1(_06019_ ), .A2(_02098_ ), .B1(_06052_ ), .B2(_04749_ ), .ZN(_01228_ ) );
MUX2_X1 _17148_ ( .A(_01228_ ), .B(\EX_LS_pc [12] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _17149_ ( .A(\EX_LS_pc [30] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01229_ ) );
OAI21_X1 _17150_ ( .A(_01204_ ), .B1(_01207_ ), .B2(_04430_ ), .ZN(_01230_ ) );
BUF_X4 _17151_ ( .A(_02174_ ), .Z(_01231_ ) );
AOI221_X4 _17152_ ( .A(_01230_ ), .B1(\LS_WB_wdata_csreg [30] ), .B2(_01231_ ), .C1(_02105_ ), .C2(_01168_ ), .ZN(_01232_ ) );
NOR2_X1 _17153_ ( .A1(_01229_ ), .A2(_01232_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
AOI21_X1 _17154_ ( .A(\EX_LS_pc [11] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01233_ ) );
OAI21_X1 _17155_ ( .A(_01204_ ), .B1(_01207_ ), .B2(_04771_ ), .ZN(_01234_ ) );
AOI221_X4 _17156_ ( .A(_01234_ ), .B1(\LS_WB_wdata_csreg [11] ), .B2(_01231_ ), .C1(_02105_ ), .C2(_01168_ ), .ZN(_01235_ ) );
NOR2_X1 _17157_ ( .A1(_01233_ ), .A2(_01235_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _17158_ ( .A(\EX_LS_pc [10] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01236_ ) );
BUF_X4 _17159_ ( .A(_06015_ ), .Z(_01237_ ) );
OAI21_X1 _17160_ ( .A(_01237_ ), .B1(_01207_ ), .B2(_06171_ ), .ZN(_01238_ ) );
AOI221_X4 _17161_ ( .A(_01238_ ), .B1(\LS_WB_wdata_csreg [10] ), .B2(_01231_ ), .C1(_02105_ ), .C2(_01168_ ), .ZN(_01239_ ) );
NOR2_X1 _17162_ ( .A1(_01236_ ), .A2(_01239_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
AOI221_X4 _17163_ ( .A(_06016_ ), .B1(\LS_WB_wdata_csreg [9] ), .B2(_01209_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [9] ), .ZN(_01240_ ) );
AOI21_X1 _17164_ ( .A(\EX_LS_pc [9] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01241_ ) );
NOR2_X1 _17165_ ( .A1(_01240_ ), .A2(_01241_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
OAI22_X1 _17166_ ( .A1(_06019_ ), .A2(_02100_ ), .B1(_06052_ ), .B2(_04854_ ), .ZN(_01242_ ) );
MUX2_X1 _17167_ ( .A(_01242_ ), .B(\EX_LS_pc [8] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
OAI22_X1 _17168_ ( .A1(_06019_ ), .A2(_02101_ ), .B1(_06052_ ), .B2(_06161_ ), .ZN(_01243_ ) );
MUX2_X1 _17169_ ( .A(_01243_ ), .B(\EX_LS_pc [7] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _17170_ ( .A1(_06019_ ), .A2(_02102_ ), .B1(_06052_ ), .B2(_04896_ ), .ZN(_01244_ ) );
MUX2_X1 _17171_ ( .A(_01244_ ), .B(\EX_LS_pc [6] ), .S(_06017_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
AOI21_X1 _17172_ ( .A(\EX_LS_pc [5] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01245_ ) );
BUF_X4 _17173_ ( .A(_02174_ ), .Z(_01246_ ) );
OAI21_X1 _17174_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_04915_ ), .ZN(_01247_ ) );
BUF_X2 _17175_ ( .A(_02104_ ), .Z(_01248_ ) );
AOI221_X4 _17176_ ( .A(_01247_ ), .B1(\LS_WB_wdata_csreg [5] ), .B2(_01231_ ), .C1(_01248_ ), .C2(_01168_ ), .ZN(_01249_ ) );
NOR2_X1 _17177_ ( .A1(_01245_ ), .A2(_01249_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
AOI21_X1 _17178_ ( .A(\EX_LS_pc [4] ), .B1(_06059_ ), .B2(_01205_ ), .ZN(_01250_ ) );
OAI21_X1 _17179_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_04934_ ), .ZN(_01251_ ) );
AOI221_X4 _17180_ ( .A(_01251_ ), .B1(\LS_WB_wdata_csreg [4] ), .B2(_01231_ ), .C1(_01248_ ), .C2(_01168_ ), .ZN(_01252_ ) );
NOR2_X1 _17181_ ( .A1(_01250_ ), .A2(_01252_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
AOI221_X4 _17182_ ( .A(_06016_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [3] ), .C1(\LS_WB_wdata_csreg [3] ), .C2(_01209_ ), .ZN(_01253_ ) );
AOI21_X1 _17183_ ( .A(\EX_LS_pc [3] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01254_ ) );
NOR2_X1 _17184_ ( .A1(_01253_ ), .A2(_01254_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
OAI21_X1 _17185_ ( .A(_06015_ ), .B1(_01246_ ), .B2(_06152_ ), .ZN(_01255_ ) );
AOI221_X4 _17186_ ( .A(_01255_ ), .B1(\LS_WB_wdata_csreg [2] ), .B2(_01207_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01256_ ) );
AOI21_X1 _17187_ ( .A(_01256_ ), .B1(_06004_ ), .B2(_06017_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
AOI21_X1 _17188_ ( .A(\EX_LS_pc [29] ), .B1(_01219_ ), .B2(_01205_ ), .ZN(_01257_ ) );
OAI21_X1 _17189_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_04512_ ), .ZN(_01258_ ) );
AOI221_X4 _17190_ ( .A(_01258_ ), .B1(\LS_WB_wdata_csreg [29] ), .B2(_01231_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01259_ ) );
NOR2_X1 _17191_ ( .A1(_01257_ ), .A2(_01259_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
AOI221_X4 _17192_ ( .A(_06016_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [1] ), .C1(\LS_WB_wdata_csreg [1] ), .C2(_01209_ ), .ZN(_01260_ ) );
AOI21_X1 _17193_ ( .A(\EX_LS_pc [1] ), .B1(_06010_ ), .B2(_01220_ ), .ZN(_01261_ ) );
NOR2_X1 _17194_ ( .A1(_01260_ ), .A2(_01261_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI21_X1 _17195_ ( .A(\EX_LS_pc [0] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01262_ ) );
OAI21_X1 _17196_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_06154_ ), .ZN(_01263_ ) );
AOI221_X4 _17197_ ( .A(_01263_ ), .B1(\LS_WB_wdata_csreg [0] ), .B2(_01231_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01264_ ) );
NOR2_X1 _17198_ ( .A1(_01262_ ), .A2(_01264_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
AOI21_X1 _17199_ ( .A(\EX_LS_pc [28] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01265_ ) );
OAI21_X1 _17200_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_04793_ ), .ZN(_01266_ ) );
AOI221_X4 _17201_ ( .A(_01266_ ), .B1(\LS_WB_wdata_csreg [28] ), .B2(_01231_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01267_ ) );
NOR2_X1 _17202_ ( .A1(_01265_ ), .A2(_01267_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _17203_ ( .A(\EX_LS_pc [27] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01268_ ) );
OAI21_X1 _17204_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_05006_ ), .ZN(_01269_ ) );
AOI221_X4 _17205_ ( .A(_01269_ ), .B1(\LS_WB_wdata_csreg [27] ), .B2(_01231_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01270_ ) );
NOR2_X1 _17206_ ( .A1(_01268_ ), .A2(_01270_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI21_X1 _17207_ ( .A(\EX_LS_pc [26] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01271_ ) );
OAI21_X1 _17208_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_06515_ ), .ZN(_01272_ ) );
AOI221_X4 _17209_ ( .A(_01272_ ), .B1(\LS_WB_wdata_csreg [26] ), .B2(_01231_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01273_ ) );
NOR2_X1 _17210_ ( .A1(_01271_ ), .A2(_01273_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI221_X4 _17211_ ( .A(_06016_ ), .B1(\LS_WB_wdata_csreg [25] ), .B2(_01209_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [25] ), .ZN(_01274_ ) );
AOI21_X1 _17212_ ( .A(\EX_LS_pc [25] ), .B1(_06010_ ), .B2(_01204_ ), .ZN(_01275_ ) );
NOR2_X1 _17213_ ( .A1(_01274_ ), .A2(_01275_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _17214_ ( .A(\EX_LS_pc [24] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01276_ ) );
OAI21_X1 _17215_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_05081_ ), .ZN(_01277_ ) );
AOI221_X4 _17216_ ( .A(_01277_ ), .B1(\LS_WB_wdata_csreg [24] ), .B2(_01207_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01278_ ) );
NOR2_X1 _17217_ ( .A1(_01276_ ), .A2(_01278_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
OAI22_X1 _17218_ ( .A1(_06019_ ), .A2(_02094_ ), .B1(_06052_ ), .B2(_06547_ ), .ZN(_01279_ ) );
MUX2_X1 _17219_ ( .A(_01279_ ), .B(\EX_LS_pc [23] ), .S(_06016_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
AOI21_X1 _17220_ ( .A(\EX_LS_pc [22] ), .B1(_01219_ ), .B2(_01220_ ), .ZN(_01280_ ) );
OAI21_X1 _17221_ ( .A(_01237_ ), .B1(_01246_ ), .B2(_05123_ ), .ZN(_01281_ ) );
AOI221_X4 _17222_ ( .A(_01281_ ), .B1(\LS_WB_wdata_csreg [22] ), .B2(_01207_ ), .C1(_01248_ ), .C2(_01171_ ), .ZN(_01282_ ) );
NOR2_X1 _17223_ ( .A1(_01280_ ), .A2(_01282_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
AOI221_X4 _17224_ ( .A(_06016_ ), .B1(\LS_WB_wdata_csreg [31] ), .B2(_01209_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [31] ), .ZN(_01283_ ) );
AOI21_X1 _17225_ ( .A(\EX_LS_pc [31] ), .B1(_06010_ ), .B2(_01204_ ), .ZN(_01284_ ) );
NOR2_X1 _17226_ ( .A1(_01283_ ), .A2(_01284_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17227_ ( .A1(_00570_ ), .A2(_05184_ ), .ZN(_01285_ ) );
NOR2_X1 _17228_ ( .A1(_06083_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01286_ ) );
INV_X1 _17229_ ( .A(_01286_ ), .ZN(_01287_ ) );
OR3_X1 _17230_ ( .A1(_00609_ ), .A2(_05183_ ), .A3(_01287_ ), .ZN(_01288_ ) );
NOR2_X1 _17231_ ( .A1(_06085_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01289_ ) );
INV_X1 _17232_ ( .A(_01289_ ), .ZN(_01290_ ) );
OR3_X1 _17233_ ( .A1(_00542_ ), .A2(_05183_ ), .A3(_01290_ ), .ZN(_01291_ ) );
XOR2_X1 _17234_ ( .A(\mylsu.araddr_tmp [0] ), .B(\mylsu.araddr_tmp [1] ), .Z(_01292_ ) );
OR3_X1 _17235_ ( .A1(_00513_ ), .A2(_05183_ ), .A3(_01292_ ), .ZN(_01293_ ) );
NAND3_X1 _17236_ ( .A1(_01288_ ), .A2(_01291_ ), .A3(_01293_ ), .ZN(_01294_ ) );
NOR2_X2 _17237_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01295_ ) );
INV_X1 _17238_ ( .A(_01295_ ), .ZN(_01296_ ) );
MUX2_X2 _17239_ ( .A(_01285_ ), .B(_01294_ ), .S(_01296_ ), .Z(_01297_ ) );
INV_X1 _17240_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01298_ ) );
NAND2_X1 _17241_ ( .A1(_01298_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01299_ ) );
NOR2_X1 _17242_ ( .A1(_01299_ ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01300_ ) );
BUF_X4 _17243_ ( .A(_01300_ ), .Z(_01301_ ) );
AND2_X4 _17244_ ( .A1(_01297_ ), .A2(_01301_ ), .ZN(_01302_ ) );
INV_X4 _17245_ ( .A(_01302_ ), .ZN(_01303_ ) );
BUF_X8 _17246_ ( .A(_01303_ ), .Z(_01304_ ) );
NOR2_X1 _17247_ ( .A1(_00513_ ), .A2(_05183_ ), .ZN(_01305_ ) );
NOR2_X1 _17248_ ( .A1(_00542_ ), .A2(_05183_ ), .ZN(_01306_ ) );
MUX2_X1 _17249_ ( .A(_01305_ ), .B(_01306_ ), .S(_01295_ ), .Z(_01307_ ) );
AND2_X1 _17250_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01308_ ) );
AND2_X2 _17251_ ( .A1(_01308_ ), .A2(_01298_ ), .ZN(_01309_ ) );
INV_X1 _17252_ ( .A(_01309_ ), .ZN(_01310_ ) );
NOR2_X1 _17253_ ( .A1(_01307_ ), .A2(_01310_ ), .ZN(_01311_ ) );
OR2_X1 _17254_ ( .A1(_01298_ ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01312_ ) );
NOR2_X1 _17255_ ( .A1(_01312_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01313_ ) );
NOR2_X1 _17256_ ( .A1(_01313_ ), .A2(_01300_ ), .ZN(_01314_ ) );
INV_X1 _17257_ ( .A(_01314_ ), .ZN(_01315_ ) );
NOR2_X1 _17258_ ( .A1(_01311_ ), .A2(_01315_ ), .ZN(_01316_ ) );
BUF_X4 _17259_ ( .A(_01316_ ), .Z(_01317_ ) );
AND2_X1 _17260_ ( .A1(_01308_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01318_ ) );
BUF_X2 _17261_ ( .A(_01318_ ), .Z(_01319_ ) );
AOI211_X1 _17262_ ( .A(_05185_ ), .B(_01319_ ), .C1(_00523_ ), .C2(_00524_ ), .ZN(_01320_ ) );
OR2_X1 _17263_ ( .A1(_01320_ ), .A2(_01309_ ), .ZN(_01321_ ) );
NAND2_X1 _17264_ ( .A1(_01317_ ), .A2(_01321_ ), .ZN(_01322_ ) );
NAND2_X1 _17265_ ( .A1(_01304_ ), .A2(_01322_ ), .ZN(_01323_ ) );
MUX2_X1 _17266_ ( .A(\EX_LS_result_reg [21] ), .B(_01323_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
AOI211_X1 _17267_ ( .A(_05185_ ), .B(_01319_ ), .C1(_00526_ ), .C2(_00527_ ), .ZN(_01324_ ) );
OR2_X1 _17268_ ( .A1(_01324_ ), .A2(_01309_ ), .ZN(_01325_ ) );
NAND2_X1 _17269_ ( .A1(_01317_ ), .A2(_01325_ ), .ZN(_01326_ ) );
NAND2_X1 _17270_ ( .A1(_01304_ ), .A2(_01326_ ), .ZN(_01327_ ) );
MUX2_X1 _17271_ ( .A(\EX_LS_result_reg [20] ), .B(_01327_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
OR2_X1 _17272_ ( .A1(_00530_ ), .A2(_06081_ ), .ZN(_01328_ ) );
OAI21_X1 _17273_ ( .A(_01310_ ), .B1(_01328_ ), .B2(_01319_ ), .ZN(_01329_ ) );
NAND2_X1 _17274_ ( .A1(_01317_ ), .A2(_01329_ ), .ZN(_01330_ ) );
NAND2_X1 _17275_ ( .A1(_01304_ ), .A2(_01330_ ), .ZN(_01331_ ) );
MUX2_X1 _17276_ ( .A(\EX_LS_result_reg [19] ), .B(_01331_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
OR2_X1 _17277_ ( .A1(_00533_ ), .A2(_05183_ ), .ZN(_01332_ ) );
OAI21_X1 _17278_ ( .A(_01310_ ), .B1(_01332_ ), .B2(_01319_ ), .ZN(_01333_ ) );
NAND2_X1 _17279_ ( .A1(_01317_ ), .A2(_01333_ ), .ZN(_01334_ ) );
NAND2_X1 _17280_ ( .A1(_01304_ ), .A2(_01334_ ), .ZN(_01335_ ) );
MUX2_X1 _17281_ ( .A(\EX_LS_result_reg [18] ), .B(_01335_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
OR2_X1 _17282_ ( .A1(_00536_ ), .A2(_05185_ ), .ZN(_01336_ ) );
OAI21_X1 _17283_ ( .A(_01310_ ), .B1(_01336_ ), .B2(_01319_ ), .ZN(_01337_ ) );
NAND2_X1 _17284_ ( .A1(_01317_ ), .A2(_01337_ ), .ZN(_01338_ ) );
NAND2_X1 _17285_ ( .A1(_01304_ ), .A2(_01338_ ), .ZN(_01339_ ) );
MUX2_X1 _17286_ ( .A(\EX_LS_result_reg [17] ), .B(_01339_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
AOI211_X1 _17287_ ( .A(_05185_ ), .B(_01319_ ), .C1(_00538_ ), .C2(_00539_ ), .ZN(_01340_ ) );
OR2_X1 _17288_ ( .A1(_01340_ ), .A2(_01309_ ), .ZN(_01341_ ) );
NAND2_X1 _17289_ ( .A1(_01317_ ), .A2(_01341_ ), .ZN(_01342_ ) );
NAND2_X1 _17290_ ( .A1(_01304_ ), .A2(_01342_ ), .ZN(_01343_ ) );
MUX2_X1 _17291_ ( .A(\EX_LS_result_reg [16] ), .B(_01343_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
BUF_X2 _17292_ ( .A(_01308_ ), .Z(_01344_ ) );
NOR4_X1 _17293_ ( .A1(_00542_ ), .A2(_06081_ ), .A3(_01344_ ), .A4(_01315_ ), .ZN(_01345_ ) );
AND2_X1 _17294_ ( .A1(_01307_ ), .A2(_01344_ ), .ZN(_01346_ ) );
OR3_X1 _17295_ ( .A1(_01302_ ), .A2(_01345_ ), .A3(_01346_ ), .ZN(_01347_ ) );
MUX2_X1 _17296_ ( .A(\EX_LS_result_reg [15] ), .B(_01347_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
AND2_X2 _17297_ ( .A1(_01296_ ), .A2(_01308_ ), .ZN(_01348_ ) );
NOR3_X1 _17298_ ( .A1(_01348_ ), .A2(_01313_ ), .A3(_01301_ ), .ZN(_01349_ ) );
AND2_X1 _17299_ ( .A1(_02000_ ), .A2(_01349_ ), .ZN(_01350_ ) );
NAND3_X1 _17300_ ( .A1(_00543_ ), .A2(_00545_ ), .A3(_01350_ ), .ZN(_01351_ ) );
NAND4_X1 _17301_ ( .A1(_00515_ ), .A2(_00520_ ), .A3(\io_master_arid [1] ), .A4(_01348_ ), .ZN(_01352_ ) );
NAND3_X1 _17302_ ( .A1(_01303_ ), .A2(_01351_ ), .A3(_01352_ ), .ZN(_01353_ ) );
MUX2_X1 _17303_ ( .A(\EX_LS_result_reg [14] ), .B(_01353_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
NAND3_X1 _17304_ ( .A1(_00546_ ), .A2(_00548_ ), .A3(_01350_ ), .ZN(_01354_ ) );
NAND4_X1 _17305_ ( .A1(_00552_ ), .A2(_00554_ ), .A3(\io_master_arid [1] ), .A4(_01348_ ), .ZN(_01355_ ) );
NAND3_X1 _17306_ ( .A1(_01303_ ), .A2(_01354_ ), .A3(_01355_ ), .ZN(_01356_ ) );
MUX2_X1 _17307_ ( .A(\EX_LS_result_reg [13] ), .B(_01356_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
AND2_X1 _17308_ ( .A1(_00587_ ), .A2(_00588_ ), .ZN(_01357_ ) );
NOR2_X1 _17309_ ( .A1(_01357_ ), .A2(_05185_ ), .ZN(_01358_ ) );
AND2_X1 _17310_ ( .A1(_01358_ ), .A2(_01348_ ), .ZN(_01359_ ) );
AND3_X1 _17311_ ( .A1(_00549_ ), .A2(_00551_ ), .A3(_01350_ ), .ZN(_01360_ ) );
OR3_X1 _17312_ ( .A1(_01302_ ), .A2(_01359_ ), .A3(_01360_ ), .ZN(_01361_ ) );
MUX2_X1 _17313_ ( .A(\EX_LS_result_reg [12] ), .B(_01361_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
BUF_X4 _17314_ ( .A(_01309_ ), .Z(_01362_ ) );
NAND2_X1 _17315_ ( .A1(_01344_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01363_ ) );
AND4_X1 _17316_ ( .A1(\io_master_arid [1] ), .A2(_00515_ ), .A3(_00520_ ), .A4(_01363_ ), .ZN(_01364_ ) );
OAI21_X1 _17317_ ( .A(_01317_ ), .B1(_01362_ ), .B2(_01364_ ), .ZN(_01365_ ) );
NAND2_X1 _17318_ ( .A1(_01304_ ), .A2(_01365_ ), .ZN(_01366_ ) );
MUX2_X1 _17319_ ( .A(\EX_LS_result_reg [30] ), .B(_01366_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17320_ ( .A1(_00555_ ), .A2(_00557_ ), .A3(_01350_ ), .ZN(_01367_ ) );
NOR2_X1 _17321_ ( .A1(_00597_ ), .A2(_05185_ ), .ZN(_01368_ ) );
AND2_X1 _17322_ ( .A1(_01368_ ), .A2(_01348_ ), .ZN(_01369_ ) );
OR3_X1 _17323_ ( .A1(_01302_ ), .A2(_01367_ ), .A3(_01369_ ), .ZN(_01370_ ) );
MUX2_X1 _17324_ ( .A(\EX_LS_result_reg [11] ), .B(_01370_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
NOR2_X1 _17325_ ( .A1(_00560_ ), .A2(_05185_ ), .ZN(_01371_ ) );
OAI21_X1 _17326_ ( .A(_01314_ ), .B1(_01371_ ), .B2(_01348_ ), .ZN(_01372_ ) );
AND2_X1 _17327_ ( .A1(_00600_ ), .A2(_02000_ ), .ZN(_01373_ ) );
INV_X1 _17328_ ( .A(_01373_ ), .ZN(_01374_ ) );
AOI21_X1 _17329_ ( .A(_01372_ ), .B1(_01348_ ), .B2(_01374_ ), .ZN(_01375_ ) );
OR2_X1 _17330_ ( .A1(_01302_ ), .A2(_01375_ ), .ZN(_01376_ ) );
MUX2_X1 _17331_ ( .A(\EX_LS_result_reg [10] ), .B(_01376_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17332_ ( .A1(_00561_ ), .A2(_00563_ ), .A3(_01350_ ), .ZN(_01377_ ) );
NOR2_X1 _17333_ ( .A1(_00603_ ), .A2(_05185_ ), .ZN(_01378_ ) );
AND2_X1 _17334_ ( .A1(_01378_ ), .A2(_01348_ ), .ZN(_01379_ ) );
OR3_X1 _17335_ ( .A1(_01302_ ), .A2(_01377_ ), .A3(_01379_ ), .ZN(_01380_ ) );
MUX2_X1 _17336_ ( .A(\EX_LS_result_reg [9] ), .B(_01380_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _17337_ ( .A1(_00565_ ), .A2(_00567_ ), .A3(_01350_ ), .ZN(_01381_ ) );
NAND4_X1 _17338_ ( .A1(_00604_ ), .A2(_00606_ ), .A3(\io_master_arid [1] ), .A4(_01348_ ), .ZN(_01382_ ) );
NAND3_X1 _17339_ ( .A1(_01303_ ), .A2(_01381_ ), .A3(_01382_ ), .ZN(_01383_ ) );
MUX2_X1 _17340_ ( .A(\EX_LS_result_reg [8] ), .B(_01383_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
NOR2_X1 _17341_ ( .A1(_00609_ ), .A2(_05184_ ), .ZN(_01384_ ) );
MUX2_X1 _17342_ ( .A(_01285_ ), .B(_01384_ ), .S(_01348_ ), .Z(_01385_ ) );
MUX2_X2 _17343_ ( .A(_01385_ ), .B(_01297_ ), .S(_01313_ ), .Z(_01386_ ) );
MUX2_X1 _17344_ ( .A(_01386_ ), .B(_01297_ ), .S(_01301_ ), .Z(_01387_ ) );
MUX2_X1 _17345_ ( .A(\EX_LS_result_reg [7] ), .B(_01387_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _17346_ ( .A1(_06137_ ), .A2(\EX_LS_result_reg [6] ), .ZN(_01388_ ) );
NOR3_X1 _17347_ ( .A1(_01313_ ), .A2(_01301_ ), .A3(_01344_ ), .ZN(_01389_ ) );
NOR2_X1 _17348_ ( .A1(_01389_ ), .A2(_01295_ ), .ZN(_01390_ ) );
INV_X1 _17349_ ( .A(_01390_ ), .ZN(_01391_ ) );
AOI211_X1 _17350_ ( .A(_06137_ ), .B(_06081_ ), .C1(_00573_ ), .C2(_01391_ ), .ZN(_01392_ ) );
NAND2_X1 _17351_ ( .A1(_00610_ ), .A2(_00612_ ), .ZN(_01393_ ) );
NOR2_X1 _17352_ ( .A1(_01314_ ), .A2(_06085_ ), .ZN(_01394_ ) );
INV_X1 _17353_ ( .A(_01394_ ), .ZN(_01395_ ) );
AND2_X1 _17354_ ( .A1(_01395_ ), .A2(_01390_ ), .ZN(_01396_ ) );
NAND2_X1 _17355_ ( .A1(_01393_ ), .A2(_01396_ ), .ZN(_01397_ ) );
NAND2_X1 _17356_ ( .A1(_01392_ ), .A2(_01397_ ), .ZN(_01398_ ) );
NAND3_X1 _17357_ ( .A1(_00515_ ), .A2(_00520_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01399_ ) );
NAND3_X1 _17358_ ( .A1(_00543_ ), .A2(_00545_ ), .A3(_06083_ ), .ZN(_01400_ ) );
AND3_X1 _17359_ ( .A1(_01399_ ), .A2(_01400_ ), .A3(_01394_ ), .ZN(_01401_ ) );
OAI21_X1 _17360_ ( .A(_01388_ ), .B1(_01398_ ), .B2(_01401_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _17361_ ( .A1(_06137_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01402_ ) );
NAND2_X1 _17362_ ( .A1(_00576_ ), .A2(_01391_ ), .ZN(_01403_ ) );
AND2_X1 _17363_ ( .A1(\io_master_arid [1] ), .A2(fanout_net_45 ), .ZN(_01404_ ) );
NAND3_X1 _17364_ ( .A1(_00523_ ), .A2(_00524_ ), .A3(_01396_ ), .ZN(_01405_ ) );
NAND3_X1 _17365_ ( .A1(_01403_ ), .A2(_01404_ ), .A3(_01405_ ), .ZN(_01406_ ) );
NAND3_X1 _17366_ ( .A1(_00552_ ), .A2(_00554_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01407_ ) );
NAND3_X1 _17367_ ( .A1(_00546_ ), .A2(_00548_ ), .A3(_06083_ ), .ZN(_01408_ ) );
AND3_X1 _17368_ ( .A1(_01407_ ), .A2(_01408_ ), .A3(_01394_ ), .ZN(_01409_ ) );
OAI21_X1 _17369_ ( .A(_01402_ ), .B1(_01406_ ), .B2(_01409_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
NAND2_X1 _17370_ ( .A1(_06137_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_01410_ ) );
AND3_X1 _17371_ ( .A1(_00549_ ), .A2(_00551_ ), .A3(_06083_ ), .ZN(_01411_ ) );
AOI21_X1 _17372_ ( .A(_06083_ ), .B1(_00587_ ), .B2(_00588_ ), .ZN(_01412_ ) );
NOR3_X1 _17373_ ( .A1(_01411_ ), .A2(_01395_ ), .A3(_01412_ ), .ZN(_01413_ ) );
NAND2_X1 _17374_ ( .A1(_00579_ ), .A2(_01391_ ), .ZN(_01414_ ) );
NAND3_X1 _17375_ ( .A1(_00526_ ), .A2(_00527_ ), .A3(_01396_ ), .ZN(_01415_ ) );
NAND3_X1 _17376_ ( .A1(_01414_ ), .A2(_01404_ ), .A3(_01415_ ), .ZN(_01416_ ) );
OAI21_X1 _17377_ ( .A(_01410_ ), .B1(_01413_ ), .B2(_01416_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
BUF_X2 _17378_ ( .A(_05184_ ), .Z(_01417_ ) );
NOR3_X1 _17379_ ( .A1(_00530_ ), .A2(_01417_ ), .A3(_01287_ ), .ZN(_01418_ ) );
NOR3_X1 _17380_ ( .A1(_00597_ ), .A2(_05184_ ), .A3(_01286_ ), .ZN(_01419_ ) );
OAI21_X1 _17381_ ( .A(_01290_ ), .B1(_01418_ ), .B2(_01419_ ), .ZN(_01420_ ) );
NAND4_X1 _17382_ ( .A1(_00555_ ), .A2(_00557_ ), .A3(_02000_ ), .A4(_01289_ ), .ZN(_01421_ ) );
AOI21_X1 _17383_ ( .A(_01295_ ), .B1(_01420_ ), .B2(_01421_ ), .ZN(_01422_ ) );
NOR3_X1 _17384_ ( .A1(_00582_ ), .A2(_05184_ ), .A3(_01296_ ), .ZN(_01423_ ) );
OAI21_X1 _17385_ ( .A(_01301_ ), .B1(_01422_ ), .B2(_01423_ ), .ZN(_01424_ ) );
NOR3_X1 _17386_ ( .A1(_00530_ ), .A2(_01417_ ), .A3(_01295_ ), .ZN(_01425_ ) );
OAI21_X1 _17387_ ( .A(_01319_ ), .B1(_01425_ ), .B2(_01423_ ), .ZN(_01426_ ) );
OR3_X1 _17388_ ( .A1(_00582_ ), .A2(_01417_ ), .A3(_01319_ ), .ZN(_01427_ ) );
AOI21_X1 _17389_ ( .A(_01309_ ), .B1(_01426_ ), .B2(_01427_ ), .ZN(_01428_ ) );
INV_X1 _17390_ ( .A(_01425_ ), .ZN(_01429_ ) );
INV_X1 _17391_ ( .A(_01423_ ), .ZN(_01430_ ) );
AOI21_X1 _17392_ ( .A(_01310_ ), .B1(_01429_ ), .B2(_01430_ ), .ZN(_01431_ ) );
OAI22_X1 _17393_ ( .A1(_01428_ ), .A2(_01431_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01312_ ), .ZN(_01432_ ) );
OAI21_X1 _17394_ ( .A(_01313_ ), .B1(_01422_ ), .B2(_01423_ ), .ZN(_01433_ ) );
AND2_X1 _17395_ ( .A1(_01432_ ), .A2(_01433_ ), .ZN(_01434_ ) );
OAI21_X1 _17396_ ( .A(_01424_ ), .B1(_01434_ ), .B2(_01301_ ), .ZN(_01435_ ) );
MUX2_X1 _17397_ ( .A(\EX_LS_result_reg [3] ), .B(_01435_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
MUX2_X1 _17398_ ( .A(_01332_ ), .B(_01374_ ), .S(_01287_ ), .Z(_01436_ ) );
OR2_X2 _17399_ ( .A1(_01436_ ), .A2(_01289_ ), .ZN(_01437_ ) );
OR3_X1 _17400_ ( .A1(_00560_ ), .A2(_01417_ ), .A3(_01290_ ), .ZN(_01438_ ) );
AOI21_X2 _17401_ ( .A(_01295_ ), .B1(_01437_ ), .B2(_01438_ ), .ZN(_01439_ ) );
NOR3_X1 _17402_ ( .A1(_00585_ ), .A2(_05184_ ), .A3(_01296_ ), .ZN(_01440_ ) );
OAI21_X1 _17403_ ( .A(_01301_ ), .B1(_01439_ ), .B2(_01440_ ), .ZN(_01441_ ) );
OAI21_X1 _17404_ ( .A(_01313_ ), .B1(_01439_ ), .B2(_01440_ ), .ZN(_01442_ ) );
NOR3_X1 _17405_ ( .A1(_00533_ ), .A2(_01417_ ), .A3(_01295_ ), .ZN(_01443_ ) );
OAI21_X1 _17406_ ( .A(_01319_ ), .B1(_01443_ ), .B2(_01440_ ), .ZN(_01444_ ) );
OR3_X1 _17407_ ( .A1(_00585_ ), .A2(_01417_ ), .A3(_01318_ ), .ZN(_01445_ ) );
AOI21_X1 _17408_ ( .A(_01309_ ), .B1(_01444_ ), .B2(_01445_ ), .ZN(_01446_ ) );
OR3_X1 _17409_ ( .A1(_00533_ ), .A2(_01417_ ), .A3(_01295_ ), .ZN(_01447_ ) );
OR3_X1 _17410_ ( .A1(_00585_ ), .A2(_05184_ ), .A3(_01296_ ), .ZN(_01448_ ) );
AOI21_X1 _17411_ ( .A(_01310_ ), .B1(_01447_ ), .B2(_01448_ ), .ZN(_01449_ ) );
OAI22_X1 _17412_ ( .A1(_01446_ ), .A2(_01449_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01312_ ), .ZN(_01450_ ) );
AND2_X1 _17413_ ( .A1(_01442_ ), .A2(_01450_ ), .ZN(_01451_ ) );
OAI21_X1 _17414_ ( .A(_01441_ ), .B1(_01451_ ), .B2(_01301_ ), .ZN(_01452_ ) );
MUX2_X1 _17415_ ( .A(\EX_LS_result_reg [2] ), .B(_01452_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
AND4_X1 _17416_ ( .A1(\io_master_arid [1] ), .A2(_00552_ ), .A3(_00554_ ), .A4(_01363_ ), .ZN(_01453_ ) );
OAI21_X1 _17417_ ( .A(_01317_ ), .B1(_01362_ ), .B2(_01453_ ), .ZN(_01454_ ) );
NAND2_X1 _17418_ ( .A1(_01304_ ), .A2(_01454_ ), .ZN(_01455_ ) );
MUX2_X1 _17419_ ( .A(\EX_LS_result_reg [29] ), .B(_01455_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
NOR3_X1 _17420_ ( .A1(_00536_ ), .A2(_01417_ ), .A3(_01287_ ), .ZN(_01456_ ) );
NOR3_X1 _17421_ ( .A1(_00603_ ), .A2(_05184_ ), .A3(_01286_ ), .ZN(_01457_ ) );
OAI21_X1 _17422_ ( .A(_01290_ ), .B1(_01456_ ), .B2(_01457_ ), .ZN(_01458_ ) );
NAND4_X1 _17423_ ( .A1(_00561_ ), .A2(_00563_ ), .A3(_02000_ ), .A4(_01289_ ), .ZN(_01459_ ) );
AOI21_X1 _17424_ ( .A(_01295_ ), .B1(_01458_ ), .B2(_01459_ ), .ZN(_01460_ ) );
NOR3_X1 _17425_ ( .A1(_00591_ ), .A2(_05184_ ), .A3(_01296_ ), .ZN(_01461_ ) );
OAI21_X1 _17426_ ( .A(_01301_ ), .B1(_01460_ ), .B2(_01461_ ), .ZN(_01462_ ) );
NOR3_X1 _17427_ ( .A1(_00536_ ), .A2(_01417_ ), .A3(_01295_ ), .ZN(_01463_ ) );
OAI21_X1 _17428_ ( .A(_01319_ ), .B1(_01463_ ), .B2(_01461_ ), .ZN(_01464_ ) );
OR3_X1 _17429_ ( .A1(_00591_ ), .A2(_01417_ ), .A3(_01318_ ), .ZN(_01465_ ) );
AOI21_X1 _17430_ ( .A(_01309_ ), .B1(_01464_ ), .B2(_01465_ ), .ZN(_01466_ ) );
INV_X1 _17431_ ( .A(_01463_ ), .ZN(_01467_ ) );
INV_X1 _17432_ ( .A(_01461_ ), .ZN(_01468_ ) );
AOI21_X1 _17433_ ( .A(_01310_ ), .B1(_01467_ ), .B2(_01468_ ), .ZN(_01469_ ) );
OAI22_X1 _17434_ ( .A1(_01466_ ), .A2(_01469_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01312_ ), .ZN(_01470_ ) );
OAI21_X1 _17435_ ( .A(_01313_ ), .B1(_01460_ ), .B2(_01461_ ), .ZN(_01471_ ) );
AND2_X1 _17436_ ( .A1(_01470_ ), .A2(_01471_ ), .ZN(_01472_ ) );
OAI21_X1 _17437_ ( .A(_01462_ ), .B1(_01472_ ), .B2(_01301_ ), .ZN(_01473_ ) );
MUX2_X1 _17438_ ( .A(\EX_LS_result_reg [1] ), .B(_01473_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
NAND2_X1 _17439_ ( .A1(_06137_ ), .A2(\EX_LS_result_reg [0] ), .ZN(_01474_ ) );
NAND2_X1 _17440_ ( .A1(_00594_ ), .A2(_01391_ ), .ZN(_01475_ ) );
NAND3_X1 _17441_ ( .A1(_00538_ ), .A2(_00539_ ), .A3(_01396_ ), .ZN(_01476_ ) );
NAND3_X1 _17442_ ( .A1(_01475_ ), .A2(_01404_ ), .A3(_01476_ ), .ZN(_01477_ ) );
NAND3_X1 _17443_ ( .A1(_00604_ ), .A2(_00606_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01478_ ) );
NAND3_X1 _17444_ ( .A1(_00565_ ), .A2(_00567_ ), .A3(_06083_ ), .ZN(_01479_ ) );
AND3_X1 _17445_ ( .A1(_01478_ ), .A2(_01479_ ), .A3(_01394_ ), .ZN(_01480_ ) );
OAI21_X1 _17446_ ( .A(_01474_ ), .B1(_01477_ ), .B2(_01480_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
AOI211_X1 _17447_ ( .A(_06081_ ), .B(_01344_ ), .C1(_00587_ ), .C2(_00588_ ), .ZN(_01481_ ) );
OAI21_X1 _17448_ ( .A(_01316_ ), .B1(_01362_ ), .B2(_01481_ ), .ZN(_01482_ ) );
NAND2_X1 _17449_ ( .A1(_01304_ ), .A2(_01482_ ), .ZN(_01483_ ) );
MUX2_X1 _17450_ ( .A(\EX_LS_result_reg [28] ), .B(_01483_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
NOR2_X1 _17451_ ( .A1(_01302_ ), .A2(_06137_ ), .ZN(_01484_ ) );
NOR3_X1 _17452_ ( .A1(_00597_ ), .A2(_06081_ ), .A3(_01344_ ), .ZN(_01485_ ) );
OAI21_X1 _17453_ ( .A(_01317_ ), .B1(_01362_ ), .B2(_01485_ ), .ZN(_01486_ ) );
AOI22_X1 _17454_ ( .A1(_01484_ ), .A2(_01486_ ), .B1(_06137_ ), .B2(_03479_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
NOR2_X1 _17455_ ( .A1(_01374_ ), .A2(_01344_ ), .ZN(_01487_ ) );
OAI21_X1 _17456_ ( .A(_01316_ ), .B1(_01362_ ), .B2(_01487_ ), .ZN(_01488_ ) );
NAND2_X1 _17457_ ( .A1(_01304_ ), .A2(_01488_ ), .ZN(_01489_ ) );
MUX2_X1 _17458_ ( .A(\EX_LS_result_reg [26] ), .B(_01489_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
NOR3_X1 _17459_ ( .A1(_00603_ ), .A2(_06081_ ), .A3(_01344_ ), .ZN(_01490_ ) );
OAI21_X1 _17460_ ( .A(_01317_ ), .B1(_01362_ ), .B2(_01490_ ), .ZN(_01491_ ) );
AOI22_X1 _17461_ ( .A1(_01484_ ), .A2(_01491_ ), .B1(_06137_ ), .B2(_03553_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
AND4_X1 _17462_ ( .A1(\io_master_arid [1] ), .A2(_00604_ ), .A3(_00606_ ), .A4(_01363_ ), .ZN(_01492_ ) );
OAI21_X1 _17463_ ( .A(_01316_ ), .B1(_01362_ ), .B2(_01492_ ), .ZN(_01493_ ) );
NAND2_X1 _17464_ ( .A1(_01303_ ), .A2(_01493_ ), .ZN(_01494_ ) );
MUX2_X1 _17465_ ( .A(\EX_LS_result_reg [24] ), .B(_01494_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _17466_ ( .A1(_00609_ ), .A2(_06081_ ), .A3(_01344_ ), .ZN(_01495_ ) );
OAI21_X1 _17467_ ( .A(_01316_ ), .B1(_01362_ ), .B2(_01495_ ), .ZN(_01496_ ) );
NAND2_X1 _17468_ ( .A1(_01303_ ), .A2(_01496_ ), .ZN(_01497_ ) );
MUX2_X1 _17469_ ( .A(\EX_LS_result_reg [23] ), .B(_01497_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
AND4_X1 _17470_ ( .A1(\io_master_arid [1] ), .A2(_00610_ ), .A3(_00612_ ), .A4(_01363_ ), .ZN(_01498_ ) );
OAI21_X1 _17471_ ( .A(_01316_ ), .B1(_01362_ ), .B2(_01498_ ), .ZN(_01499_ ) );
NAND2_X1 _17472_ ( .A1(_01303_ ), .A2(_01499_ ), .ZN(_01500_ ) );
MUX2_X1 _17473_ ( .A(\EX_LS_result_reg [22] ), .B(_01500_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
NOR3_X1 _17474_ ( .A1(_00513_ ), .A2(_06081_ ), .A3(_01344_ ), .ZN(_01501_ ) );
OAI21_X1 _17475_ ( .A(_01316_ ), .B1(_01362_ ), .B2(_01501_ ), .ZN(_01502_ ) );
NAND2_X1 _17476_ ( .A1(_01303_ ), .A2(_01502_ ), .ZN(_01503_ ) );
MUX2_X1 _17477_ ( .A(\EX_LS_result_reg [31] ), .B(_01503_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17478_ ( .A1(\LS_WB_waddr_reg [1] ), .A2(\LS_WB_waddr_reg [0] ), .ZN(_01504_ ) );
INV_X1 _17479_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01505_ ) );
INV_X1 _17480_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01506_ ) );
NAND3_X1 _17481_ ( .A1(_01504_ ), .A2(_01505_ ), .A3(_01506_ ), .ZN(_01507_ ) );
AND2_X1 _17482_ ( .A1(_01583_ ), .A2(LS_WB_wen_reg ), .ZN(_01508_ ) );
NAND2_X1 _17483_ ( .A1(_01507_ ), .A2(_01508_ ), .ZN(_01509_ ) );
BUF_X4 _17484_ ( .A(_01509_ ), .Z(_01510_ ) );
INV_X1 _17485_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01511_ ) );
INV_X1 _17486_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01512_ ) );
AOI21_X1 _17487_ ( .A(_01510_ ), .B1(_01511_ ), .B2(_01512_ ), .ZN(_01513_ ) );
NOR2_X1 _17488_ ( .A1(_01509_ ), .A2(_01505_ ), .ZN(_01514_ ) );
NOR4_X1 _17489_ ( .A1(_01513_ ), .A2(_01514_ ), .A3(_01506_ ), .A4(_01510_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _17490_ ( .A1(_01510_ ), .A2(_01506_ ), .ZN(_01515_ ) );
NOR2_X1 _17491_ ( .A1(_01510_ ), .A2(_01512_ ), .ZN(_01516_ ) );
AND4_X1 _17492_ ( .A1(_01505_ ), .A2(_01515_ ), .A3(_01516_ ), .A4(_01511_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
NOR2_X1 _17493_ ( .A1(_01509_ ), .A2(_01511_ ), .ZN(_01517_ ) );
AND4_X1 _17494_ ( .A1(_01506_ ), .A2(_01514_ ), .A3(_01517_ ), .A4(_01512_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
AND4_X1 _17495_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(_01515_ ), .A3(_01517_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
CLKBUF_X1 _17496_ ( .A(fanout_net_4 ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
AOI21_X1 _17497_ ( .A(_01510_ ), .B1(_01505_ ), .B2(_01506_ ), .ZN(_01518_ ) );
NOR4_X1 _17498_ ( .A1(_01518_ ), .A2(_01517_ ), .A3(_01512_ ), .A4(_01510_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17499_ ( .A1(_01518_ ), .A2(_01516_ ), .A3(_01511_ ), .A4(_01510_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17500_ ( .A1(_01505_ ), .A2(_01515_ ), .A3(_01517_ ), .A4(_01512_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17501_ ( .A1(_01505_ ), .A2(_01515_ ), .A3(_01517_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _17502_ ( .A1(_01513_ ), .A2(_01515_ ), .A3(_01505_ ), .A4(_01510_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
NOR4_X1 _17503_ ( .A1(_01513_ ), .A2(_01505_ ), .A3(_01506_ ), .A4(_01510_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17504_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01514_ ), .A3(_01516_ ), .A4(_01511_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17505_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01514_ ), .A3(_01517_ ), .A4(_01512_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17506_ ( .A1(_01506_ ), .A2(_01514_ ), .A3(_01517_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17507_ ( .A1(_01506_ ), .A2(_01514_ ), .A3(_01516_ ), .A4(_01511_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17508_ ( .A1(_01518_ ), .A2(_01511_ ), .A3(_01512_ ), .A4(_01510_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17509_ ( .A1(_01969_ ), .A2(_01585_ ), .A3(_01977_ ), .ZN(_01519_ ) );
NAND2_X1 _17510_ ( .A1(_01519_ ), .A2(_01585_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17511_ ( .A(fanout_net_4 ), .B(_01969_ ), .C1(_01970_ ), .C2(_06090_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17512_ ( .A(_01507_ ), .Z(_01520_ ) );
CLKBUF_X2 _17513_ ( .A(_01508_ ), .Z(_01521_ ) );
AND3_X1 _17514_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17515_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17516_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17517_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17518_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17519_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17520_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17521_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17522_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17523_ ( .A1(_01520_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01521_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17524_ ( .A(_01507_ ), .Z(_01522_ ) );
CLKBUF_X2 _17525_ ( .A(_01508_ ), .Z(_01523_ ) );
AND3_X1 _17526_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17527_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17528_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17529_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17530_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17531_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17532_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17533_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17534_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17535_ ( .A1(_01522_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01523_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17536_ ( .A(_01507_ ), .Z(_01524_ ) );
CLKBUF_X2 _17537_ ( .A(_01508_ ), .Z(_01525_ ) );
AND3_X1 _17538_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17539_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17540_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17541_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17542_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17543_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17544_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17545_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17546_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17547_ ( .A1(_01524_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01525_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17548_ ( .A1(_01507_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01508_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17549_ ( .A1(_01507_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01508_ ), .ZN(\myreg.Reg[2]_$_DFFE_PP__Q_D ) );
AND3_X1 _17550_ ( .A1(_01585_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17551_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01526_ ) );
AND2_X1 _17552_ ( .A1(_01526_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01527_ ) );
INV_X1 _17553_ ( .A(_01527_ ), .ZN(_01528_ ) );
NOR2_X1 _17554_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01529_ ) );
OAI211_X1 _17555_ ( .A(_01584_ ), .B(\mysc.state [0] ), .C1(_01528_ ), .C2(_01529_ ), .ZN(_01530_ ) );
INV_X1 _17556_ ( .A(_01530_ ), .ZN(_01531_ ) );
OR3_X1 _17557_ ( .A1(_01531_ ), .A2(fanout_net_4 ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17558_ ( .A1(_01528_ ), .A2(reset ), .A3(_01529_ ), .ZN(_01532_ ) );
NAND2_X1 _17559_ ( .A1(_01532_ ), .A2(\mysc.state [0] ), .ZN(_01533_ ) );
OR3_X1 _17560_ ( .A1(_06072_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01534_ ) );
NAND2_X1 _17561_ ( .A1(_01533_ ), .A2(_01534_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17562_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_08012_ ) );
CLKGATE_X1 _17563_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_08013_ ) );
CLKGATE_X1 _17564_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08014_ ) );
CLKGATE_X1 _17565_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08015_ ) );
CLKGATE_X1 _17566_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08016_ ) );
CLKGATE_X1 _17567_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08017_ ) );
CLKGATE_X1 _17568_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_08018_ ) );
CLKGATE_X1 _17569_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_08019_ ) );
CLKGATE_X1 _17570_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_08020_ ) );
CLKGATE_X1 _17571_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_08021_ ) );
CLKGATE_X1 _17572_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_08022_ ) );
CLKGATE_X1 _17573_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08023_ ) );
CLKGATE_X1 _17574_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08024_ ) );
CLKGATE_X1 _17575_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08025_ ) );
CLKGATE_X1 _17576_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_08026_ ) );
CLKGATE_X1 _17577_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_08027_ ) );
CLKGATE_X1 _17578_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_08028_ ) );
CLKGATE_X1 _17579_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08029_ ) );
CLKGATE_X1 _17580_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_08030_ ) );
CLKGATE_X1 _17581_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ), .GCK(_08031_ ) );
CLKGATE_X1 _17582_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .GCK(_08032_ ) );
CLKGATE_X1 _17583_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08033_ ) );
CLKGATE_X1 _17584_ ( .CK(clock ), .E(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_08034_ ) );
CLKGATE_X1 _17585_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_08035_ ) );
CLKGATE_X1 _17586_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_08036_ ) );
CLKGATE_X1 _17587_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_08037_ ) );
CLKGATE_X1 _17588_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_08038_ ) );
CLKGATE_X1 _17589_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_08039_ ) );
CLKGATE_X1 _17590_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_08040_ ) );
CLKGATE_X1 _17591_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_08041_ ) );
CLKGATE_X1 _17592_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_08042_ ) );
CLKGATE_X1 _17593_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_08043_ ) );
CLKGATE_X1 _17594_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_08044_ ) );
CLKGATE_X1 _17595_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_08045_ ) );
CLKGATE_X1 _17596_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_08046_ ) );
CLKGATE_X1 _17597_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08047_ ) );
CLKGATE_X1 _17598_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08048_ ) );
CLKGATE_X1 _17599_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08049_ ) );
CLKGATE_X1 _17600_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08050_ ) );
CLKGATE_X1 _17601_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08051_ ) );
CLKGATE_X1 _17602_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08052_ ) );
CLKGATE_X1 _17603_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08053_ ) );
CLKGATE_X1 _17604_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08054_ ) );
CLKGATE_X1 _17605_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08055_ ) );
CLKGATE_X1 _17606_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08056_ ) );
CLKGATE_X1 _17607_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_08057_ ) );
CLKGATE_X1 _17608_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08058_ ) );
CLKGATE_X1 _17609_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08059_ ) );
CLKGATE_X1 _17610_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08060_ ) );
CLKGATE_X1 _17611_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08061_ ) );
CLKGATE_X1 _17612_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08062_ ) );
CLKGATE_X1 _17613_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_08063_ ) );
CLKGATE_X1 _17614_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08064_ ) );
CLKGATE_X1 _17615_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08065_ ) );
CLKGATE_X1 _17616_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08066_ ) );
CLKGATE_X1 _17617_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08067_ ) );
CLKGATE_X1 _17618_ ( .CK(clock ), .E(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08068_ ) );
CLKGATE_X1 _17619_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_08069_ ) );
CLKGATE_X1 _17620_ ( .CK(clock ), .E(\myexu.state_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_08070_ ) );
CLKGATE_X1 _17621_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08071_ ) );
CLKGATE_X1 _17622_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08072_ ) );
CLKGATE_X1 _17623_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08073_ ) );
CLKGATE_X1 _17624_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ), .GCK(_08074_ ) );
CLKGATE_X1 _17625_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ), .GCK(_08075_ ) );
CLKGATE_X1 _17626_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08076_ ) );
LOGIC1_X1 _17627_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17628_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08307_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08308_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08309_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08310_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08311_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08312_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08313_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08314_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08315_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08316_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08317_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08318_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08319_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08320_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08321_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08322_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08323_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08324_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08325_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08326_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08327_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08328_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08329_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08330_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08331_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08332_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08333_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08334_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08335_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08336_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08337_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08076_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08338_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08075_ ), .Q(\mtvec [31] ), .QN(_08339_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08075_ ), .Q(\mtvec [30] ), .QN(_08340_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08075_ ), .Q(\mtvec [21] ), .QN(_08341_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08075_ ), .Q(\mtvec [20] ), .QN(_08342_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08075_ ), .Q(\mtvec [19] ), .QN(_08343_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08075_ ), .Q(\mtvec [18] ), .QN(_08344_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08075_ ), .Q(\mtvec [17] ), .QN(_08345_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08075_ ), .Q(\mtvec [16] ), .QN(_08346_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08075_ ), .Q(\mtvec [15] ), .QN(_08347_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08075_ ), .Q(\mtvec [14] ), .QN(_08348_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08075_ ), .Q(\mtvec [13] ), .QN(_08349_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08075_ ), .Q(\mtvec [12] ), .QN(_08350_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08075_ ), .Q(\mtvec [29] ), .QN(_08351_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08075_ ), .Q(\mtvec [11] ), .QN(_08352_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08075_ ), .Q(\mtvec [10] ), .QN(_08353_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08075_ ), .Q(\mtvec [9] ), .QN(_08354_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08075_ ), .Q(\mtvec [8] ), .QN(_08355_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08075_ ), .Q(\mtvec [7] ), .QN(_08356_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08075_ ), .Q(\mtvec [6] ), .QN(_08357_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08075_ ), .Q(\mtvec [5] ), .QN(_08358_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08075_ ), .Q(\mtvec [4] ), .QN(_08359_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08075_ ), .Q(\mtvec [3] ), .QN(_08360_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08075_ ), .Q(\mtvec [2] ), .QN(_08361_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08075_ ), .Q(\mtvec [28] ), .QN(_08362_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08075_ ), .Q(\mtvec [1] ), .QN(_08363_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08075_ ), .Q(\mtvec [0] ), .QN(_08364_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08075_ ), .Q(\mtvec [27] ), .QN(_08365_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08075_ ), .Q(\mtvec [26] ), .QN(_08366_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08075_ ), .Q(\mtvec [25] ), .QN(_08367_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08075_ ), .Q(\mtvec [24] ), .QN(_08368_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08075_ ), .Q(\mtvec [23] ), .QN(_08369_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08075_ ), .Q(\mtvec [22] ), .QN(_08370_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08074_ ), .Q(\mepc [31] ), .QN(_08371_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08074_ ), .Q(\mepc [30] ), .QN(_08372_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08074_ ), .Q(\mepc [21] ), .QN(_08373_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08074_ ), .Q(\mepc [20] ), .QN(_08374_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08074_ ), .Q(\mepc [19] ), .QN(_08375_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08074_ ), .Q(\mepc [18] ), .QN(_08376_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08074_ ), .Q(\mepc [17] ), .QN(_08377_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08074_ ), .Q(\mepc [16] ), .QN(_08378_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08074_ ), .Q(\mepc [15] ), .QN(_08379_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08074_ ), .Q(\mepc [14] ), .QN(_08380_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08074_ ), .Q(\mepc [13] ), .QN(_08381_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08074_ ), .Q(\mepc [12] ), .QN(_08382_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08074_ ), .Q(\mepc [29] ), .QN(_08383_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08074_ ), .Q(\mepc [11] ), .QN(_08384_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08074_ ), .Q(\mepc [10] ), .QN(_08385_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08074_ ), .Q(\mepc [9] ), .QN(_08386_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08074_ ), .Q(\mepc [8] ), .QN(_08387_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08074_ ), .Q(\mepc [7] ), .QN(_08388_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08074_ ), .Q(\mepc [6] ), .QN(_08389_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08074_ ), .Q(\mepc [5] ), .QN(_08390_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08074_ ), .Q(\mepc [4] ), .QN(_08391_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08074_ ), .Q(\mepc [3] ), .QN(_08392_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08074_ ), .Q(\mepc [2] ), .QN(_08393_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08074_ ), .Q(\mepc [28] ), .QN(_08394_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08074_ ), .Q(\mepc [1] ), .QN(_08395_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08074_ ), .Q(\mepc [0] ), .QN(_08396_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08074_ ), .Q(\mepc [27] ), .QN(_08397_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08074_ ), .Q(\mepc [26] ), .QN(_08398_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08074_ ), .Q(\mepc [25] ), .QN(_08399_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08074_ ), .Q(\mepc [24] ), .QN(_08400_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08074_ ), .Q(\mepc [23] ), .QN(_08401_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08074_ ), .Q(\mepc [22] ), .QN(_08402_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08403_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08404_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08405_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08306_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08305_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08304_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08303_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08302_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08301_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08300_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08299_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08298_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08297_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08296_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08295_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08294_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08293_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08292_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08291_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08290_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08289_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08288_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08287_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08286_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08285_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00086_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08284_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00087_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08283_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00088_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08282_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00089_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08281_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00090_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08280_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00091_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08279_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00092_ ), .CK(_08073_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08406_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PN0__Q ( .D(_00093_ ), .CK(clock ), .Q(excp_written ), .QN(_08407_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08278_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08408_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08409_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08410_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08411_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08412_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08413_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08414_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08415_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08416_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08417_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08418_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08419_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08420_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08421_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08422_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08423_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08424_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08425_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08426_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08427_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08428_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08429_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08430_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08431_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08432_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08433_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08434_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08435_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08436_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08437_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08072_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08277_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00094_ ), .CK(_08071_ ), .Q(\myec.state [1] ), .QN(_08276_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00095_ ), .CK(_08071_ ), .Q(\myec.state [0] ), .QN(_08438_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PP0__Q ( .D(_00096_ ), .CK(clock ), .Q(check_quest ), .QN(_08439_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08275_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08440_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08441_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08442_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08443_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08444_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08445_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08446_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08447_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08448_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08449_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08274_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00097_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08273_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00098_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08272_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00099_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08271_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00100_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08270_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00101_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08269_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00102_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08268_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00103_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08267_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00104_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08266_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00105_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08265_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00106_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08264_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00107_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08263_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00108_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08262_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00109_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08261_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00110_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08260_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00111_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08259_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00112_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08258_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00113_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08257_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00114_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08256_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00115_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08255_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00116_ ), .CK(_08070_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08254_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q ( .D(_00117_ ), .CK(_08069_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08253_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_1 ( .D(_00118_ ), .CK(_08069_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08252_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_2 ( .D(_00119_ ), .CK(_08069_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08251_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_3 ( .D(_00120_ ), .CK(_08069_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08250_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_4 ( .D(_00121_ ), .CK(_08069_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08249_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q ( .D(_00122_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [30] ), .QN(_08248_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_1 ( .D(_00123_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [29] ), .QN(_08247_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_10 ( .D(_00124_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [20] ), .QN(_08246_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_11 ( .D(_00125_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [19] ), .QN(_08245_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_12 ( .D(_00126_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [18] ), .QN(_08244_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_13 ( .D(_00127_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [17] ), .QN(_08243_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_14 ( .D(_00128_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [16] ), .QN(_08242_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_15 ( .D(_00129_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [15] ), .QN(_08241_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_16 ( .D(_00130_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [14] ), .QN(_08240_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_17 ( .D(_00131_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [13] ), .QN(_08239_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_18 ( .D(_00132_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [12] ), .QN(_08238_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_19 ( .D(_00133_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [11] ), .QN(_08237_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_2 ( .D(_00134_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [28] ), .QN(_08236_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_20 ( .D(_00135_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [10] ), .QN(_08235_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_21 ( .D(_00136_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [9] ), .QN(_08234_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_22 ( .D(_00137_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [8] ), .QN(_08233_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_23 ( .D(_00138_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [7] ), .QN(_08232_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_24 ( .D(_00139_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [6] ), .QN(_08231_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_25 ( .D(_00140_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [5] ), .QN(_08230_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_26 ( .D(_00141_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [4] ), .QN(_08229_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_27 ( .D(_00142_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [3] ), .QN(_08228_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_28 ( .D(_00143_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [2] ), .QN(_08227_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_29 ( .D(_00144_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [1] ), .QN(_08226_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_3 ( .D(_00145_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [27] ), .QN(_08225_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_30 ( .D(_00146_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [0] ), .QN(_08224_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_4 ( .D(_00147_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [26] ), .QN(_08223_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_5 ( .D(_00148_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [25] ), .QN(_08222_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_6 ( .D(_00149_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [24] ), .QN(_08221_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_7 ( .D(_00150_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [23] ), .QN(_08220_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_8 ( .D(_00151_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [22] ), .QN(_08219_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_9 ( .D(_00152_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [21] ), .QN(_08218_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP1P__Q ( .D(_00153_ ), .CK(_08068_ ), .Q(\myexu.pc_jump [31] ), .QN(_08217_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q ( .D(_00154_ ), .CK(_08069_ ), .Q(\EX_LS_pc [31] ), .QN(_08216_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_1 ( .D(_00155_ ), .CK(_08069_ ), .Q(\EX_LS_pc [30] ), .QN(_08215_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_10 ( .D(_00156_ ), .CK(_08069_ ), .Q(\EX_LS_pc [21] ), .QN(_08214_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_11 ( .D(_00157_ ), .CK(_08069_ ), .Q(\EX_LS_pc [20] ), .QN(_08213_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_12 ( .D(_00158_ ), .CK(_08069_ ), .Q(\EX_LS_pc [19] ), .QN(_08212_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_13 ( .D(_00159_ ), .CK(_08069_ ), .Q(\EX_LS_pc [18] ), .QN(_08211_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_14 ( .D(_00160_ ), .CK(_08069_ ), .Q(\EX_LS_pc [17] ), .QN(_08210_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_15 ( .D(_00161_ ), .CK(_08069_ ), .Q(\EX_LS_pc [16] ), .QN(_08209_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_16 ( .D(_00162_ ), .CK(_08069_ ), .Q(\EX_LS_pc [15] ), .QN(_08208_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_17 ( .D(_00163_ ), .CK(_08069_ ), .Q(\EX_LS_pc [14] ), .QN(_08207_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_18 ( .D(_00164_ ), .CK(_08069_ ), .Q(\EX_LS_pc [13] ), .QN(_08206_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_19 ( .D(_00165_ ), .CK(_08069_ ), .Q(\EX_LS_pc [12] ), .QN(_08205_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_2 ( .D(_00166_ ), .CK(_08069_ ), .Q(\EX_LS_pc [29] ), .QN(_08204_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_20 ( .D(_00167_ ), .CK(_08069_ ), .Q(\EX_LS_pc [11] ), .QN(_08203_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_21 ( .D(_00168_ ), .CK(_08069_ ), .Q(\EX_LS_pc [10] ), .QN(_08202_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_22 ( .D(_00169_ ), .CK(_08069_ ), .Q(\EX_LS_pc [9] ), .QN(_08201_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_23 ( .D(_00170_ ), .CK(_08069_ ), .Q(\EX_LS_pc [8] ), .QN(_08200_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_24 ( .D(_00171_ ), .CK(_08069_ ), .Q(\EX_LS_pc [7] ), .QN(_08199_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_25 ( .D(_00172_ ), .CK(_08069_ ), .Q(\EX_LS_pc [6] ), .QN(_08198_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_26 ( .D(_00173_ ), .CK(_08069_ ), .Q(\EX_LS_pc [5] ), .QN(_08197_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_27 ( .D(_00174_ ), .CK(_08069_ ), .Q(\EX_LS_pc [4] ), .QN(_08196_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_28 ( .D(_00175_ ), .CK(_08069_ ), .Q(\EX_LS_pc [3] ), .QN(_08195_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_29 ( .D(_00176_ ), .CK(_08069_ ), .Q(\EX_LS_pc [2] ), .QN(_08194_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_3 ( .D(_00177_ ), .CK(_08069_ ), .Q(\EX_LS_pc [28] ), .QN(_08193_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_30 ( .D(_00178_ ), .CK(_08069_ ), .Q(\EX_LS_pc [1] ), .QN(_08192_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_31 ( .D(_00179_ ), .CK(_08069_ ), .Q(\EX_LS_pc [0] ), .QN(_08191_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_4 ( .D(_00180_ ), .CK(_08069_ ), .Q(\EX_LS_pc [27] ), .QN(_08190_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_5 ( .D(_00181_ ), .CK(_08069_ ), .Q(\EX_LS_pc [26] ), .QN(_08189_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_6 ( .D(_00182_ ), .CK(_08069_ ), .Q(\EX_LS_pc [25] ), .QN(_08188_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_7 ( .D(_00183_ ), .CK(_08069_ ), .Q(\EX_LS_pc [24] ), .QN(_08187_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_8 ( .D(_00184_ ), .CK(_08069_ ), .Q(\EX_LS_pc [23] ), .QN(_08186_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_9 ( .D(_00185_ ), .CK(_08069_ ), .Q(\EX_LS_pc [22] ), .QN(_08450_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08451_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08452_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08453_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08454_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08455_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08456_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08457_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08458_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08459_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08460_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08461_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08462_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08463_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08464_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08465_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08466_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08467_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08468_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08469_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08470_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08471_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08472_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08473_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08474_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08475_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08476_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08477_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08478_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08479_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08480_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08481_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08070_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08482_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08070_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PP0__Q ( .D(_00187_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q ( .D(_00186_ ), .CK(_08069_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_1 ( .D(_00188_ ), .CK(_08069_ ), .Q(\EX_LS_flag [1] ), .QN(_08185_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_2 ( .D(_00189_ ), .CK(_08069_ ), .Q(\EX_LS_flag [0] ), .QN(_08184_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_3 ( .D(_00190_ ), .CK(_08069_ ), .Q(\EX_LS_typ [4] ), .QN(_08183_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_4 ( .D(_00191_ ), .CK(_08069_ ), .Q(\EX_LS_typ [3] ), .QN(_08182_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_5 ( .D(_00192_ ), .CK(_08069_ ), .Q(\EX_LS_typ [2] ), .QN(_08181_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_6 ( .D(_00193_ ), .CK(_08069_ ), .Q(\EX_LS_typ [1] ), .QN(_08180_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_7 ( .D(_00194_ ), .CK(_08069_ ), .Q(\EX_LS_typ [0] ), .QN(_08179_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00195_ ), .CK(_08067_ ), .Q(\ID_EX_csr [11] ), .QN(_08178_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00196_ ), .CK(_08067_ ), .Q(\ID_EX_csr [10] ), .QN(_08177_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00197_ ), .CK(_08067_ ), .Q(\ID_EX_csr [1] ), .QN(_08176_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00198_ ), .CK(_08067_ ), .Q(\ID_EX_csr [0] ), .QN(_08175_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00199_ ), .CK(_08067_ ), .Q(\ID_EX_csr [9] ), .QN(_08174_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00200_ ), .CK(_08067_ ), .Q(\ID_EX_csr [8] ), .QN(_08173_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00201_ ), .CK(_08067_ ), .Q(\ID_EX_csr [7] ), .QN(_08172_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00202_ ), .CK(_08067_ ), .Q(\ID_EX_csr [6] ), .QN(_08171_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00203_ ), .CK(_08067_ ), .Q(\ID_EX_csr [5] ), .QN(_08170_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00204_ ), .CK(_08067_ ), .Q(\ID_EX_csr [4] ), .QN(_08169_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00205_ ), .CK(_08067_ ), .Q(\ID_EX_csr [3] ), .QN(_08168_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00206_ ), .CK(_08067_ ), .Q(\ID_EX_csr [2] ), .QN(_08167_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00207_ ), .CK(_08066_ ), .Q(exception_quest_IDU ), .QN(_08166_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00208_ ), .CK(_08065_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08064_ ), .Q(\ID_EX_imm [31] ), .QN(_08483_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08064_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08064_ ), .Q(\ID_EX_imm [21] ), .QN(_08484_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08064_ ), .Q(\ID_EX_imm [20] ), .QN(_08485_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08064_ ), .Q(\ID_EX_imm [19] ), .QN(_08486_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08064_ ), .Q(\ID_EX_imm [18] ), .QN(_08487_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08064_ ), .Q(\ID_EX_imm [17] ), .QN(_08488_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08064_ ), .Q(\ID_EX_imm [16] ), .QN(_08489_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08064_ ), .Q(\ID_EX_imm [15] ), .QN(_08490_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08064_ ), .Q(\ID_EX_imm [14] ), .QN(_08491_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08064_ ), .Q(\ID_EX_imm [13] ), .QN(_08492_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08064_ ), .Q(\ID_EX_imm [12] ), .QN(_08493_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08064_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08064_ ), .Q(\ID_EX_imm [11] ), .QN(_08494_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08064_ ), .Q(\ID_EX_imm [10] ), .QN(_08495_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08064_ ), .Q(\ID_EX_imm [9] ), .QN(_08496_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08064_ ), .Q(\ID_EX_imm [8] ), .QN(_08497_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08064_ ), .Q(\ID_EX_imm [7] ), .QN(_08498_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08064_ ), .Q(\ID_EX_imm [6] ), .QN(_08499_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08064_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08064_ ), .Q(\ID_EX_imm [4] ), .QN(_08500_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08064_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08064_ ), .Q(\ID_EX_imm [2] ), .QN(_08501_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08064_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08064_ ), .Q(\ID_EX_imm [1] ), .QN(_08502_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08064_ ), .Q(\ID_EX_imm [0] ), .QN(_08503_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08064_ ), .Q(\ID_EX_imm [27] ), .QN(_08504_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08064_ ), .Q(\ID_EX_imm [26] ), .QN(_08505_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08064_ ), .Q(\ID_EX_imm [25] ), .QN(_08506_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08064_ ), .Q(\ID_EX_imm [24] ), .QN(_08507_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08064_ ), .Q(\ID_EX_imm [23] ), .QN(_08508_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08064_ ), .Q(\ID_EX_imm [22] ), .QN(_08509_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08063_ ), .Q(\ID_EX_pc [31] ), .QN(_08510_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08063_ ), .Q(\ID_EX_pc [30] ), .QN(_08511_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08063_ ), .Q(\ID_EX_pc [21] ), .QN(_08512_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08063_ ), .Q(\ID_EX_pc [20] ), .QN(_08513_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08063_ ), .Q(\ID_EX_pc [19] ), .QN(_08514_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08063_ ), .Q(\ID_EX_pc [18] ), .QN(_08515_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08063_ ), .Q(\ID_EX_pc [17] ), .QN(_08516_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08063_ ), .Q(\ID_EX_pc [16] ), .QN(_08517_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08063_ ), .Q(\ID_EX_pc [15] ), .QN(_08518_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08063_ ), .Q(\ID_EX_pc [14] ), .QN(_08519_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08063_ ), .Q(\ID_EX_pc [13] ), .QN(_08520_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08063_ ), .Q(\ID_EX_pc [12] ), .QN(_08521_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08063_ ), .Q(\ID_EX_pc [29] ), .QN(_08522_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08063_ ), .Q(\ID_EX_pc [11] ), .QN(_08523_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08063_ ), .Q(\ID_EX_pc [10] ), .QN(_08524_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08063_ ), .Q(\ID_EX_pc [9] ), .QN(_08525_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08063_ ), .Q(\ID_EX_pc [8] ), .QN(_08526_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08063_ ), .Q(\ID_EX_pc [7] ), .QN(_08527_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08063_ ), .Q(\ID_EX_pc [6] ), .QN(_08528_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08063_ ), .Q(\ID_EX_pc [5] ), .QN(_08529_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08063_ ), .Q(\ID_EX_pc [4] ), .QN(_08530_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08063_ ), .Q(\ID_EX_pc [3] ), .QN(_08531_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08063_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08063_ ), .Q(\ID_EX_pc [28] ), .QN(_08532_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08063_ ), .Q(\ID_EX_pc [1] ), .QN(_08533_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08063_ ), .Q(\ID_EX_pc [0] ), .QN(_08534_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08063_ ), .Q(\ID_EX_pc [27] ), .QN(_08535_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08063_ ), .Q(\ID_EX_pc [26] ), .QN(_08536_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08063_ ), .Q(\ID_EX_pc [25] ), .QN(_08537_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08063_ ), .Q(\ID_EX_pc [24] ), .QN(_08538_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08063_ ), .Q(\ID_EX_pc [23] ), .QN(_08539_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08063_ ), .Q(\ID_EX_pc [22] ), .QN(_08165_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00209_ ), .CK(_08062_ ), .Q(\ID_EX_rd [4] ), .QN(_08164_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00210_ ), .CK(_08062_ ), .Q(\ID_EX_rd [3] ), .QN(_08163_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00211_ ), .CK(_08062_ ), .Q(\ID_EX_rd [2] ), .QN(_08162_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00212_ ), .CK(_08062_ ), .Q(\ID_EX_rd [1] ), .QN(_08161_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00213_ ), .CK(_08062_ ), .Q(\ID_EX_rd [0] ), .QN(_08160_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00214_ ), .CK(_08061_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08159_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00215_ ), .CK(_08061_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08158_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00217_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08156_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00216_ ), .CK(_08061_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08157_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00219_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08154_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00218_ ), .CK(_08061_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08155_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00221_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08152_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00220_ ), .CK(_08061_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08153_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00223_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08150_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00222_ ), .CK(_08060_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08151_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00224_ ), .CK(_08060_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08149_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00226_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08147_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00225_ ), .CK(_08060_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08148_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00228_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08145_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00227_ ), .CK(_08060_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08146_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00230_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08143_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00229_ ), .CK(_08060_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08144_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00232_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08141_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_08059_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08142_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00233_ ), .CK(_08058_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08140_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08541_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00234_ ), .CK(_08057_ ), .Q(\ID_EX_typ [7] ), .QN(_08540_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00235_ ), .CK(_08057_ ), .Q(\ID_EX_typ [6] ), .QN(_08139_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00236_ ), .CK(_08057_ ), .Q(\ID_EX_typ [5] ), .QN(_08138_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00237_ ), .CK(_08057_ ), .Q(\ID_EX_typ [4] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00238_ ), .CK(_08057_ ), .Q(\ID_EX_typ [3] ), .QN(_08137_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00239_ ), .CK(_08057_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00240_ ), .CK(_08057_ ), .Q(\ID_EX_typ [1] ), .QN(_08136_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00241_ ), .CK(_08057_ ), .Q(\ID_EX_typ [0] ), .QN(_08542_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08056_ ), .Q(check_assert ), .QN(_08543_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08055_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08055_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08055_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08055_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08055_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08055_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08055_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08055_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08055_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08055_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08055_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08055_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08055_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08055_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08055_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08055_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08055_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08055_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08055_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08055_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08055_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08055_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08055_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08055_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08055_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08055_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08055_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08055_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08055_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08055_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08055_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08055_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08544_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08545_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08546_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08547_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08548_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08549_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08550_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08551_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08552_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08553_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08554_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08555_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08556_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08557_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08558_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08559_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08560_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08561_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08562_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08563_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08564_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08565_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08566_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08567_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08054_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08053_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08052_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08051_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08050_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08049_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08048_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08047_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08046_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08045_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08855_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08856_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08857_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08858_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08859_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08860_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08861_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08862_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08863_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08864_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08865_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08866_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08867_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08868_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08869_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08870_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08871_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08872_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08873_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08874_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08875_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08876_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08877_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08878_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08879_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08044_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08880_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08881_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08882_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08883_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08884_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08885_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08886_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08887_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08888_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08889_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08890_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08891_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08892_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08893_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08894_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08895_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08896_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08897_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08898_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08899_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08900_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08901_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08902_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08903_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08904_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08905_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08906_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08043_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08135_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00242_ ), .CK(_08042_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08134_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00243_ ), .CK(_08041_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08133_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00244_ ), .CK(_08040_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08907_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_08039_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08132_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_08038_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_08037_ ), .Q(\IF_ID_pc [30] ), .QN(_08131_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00247_ ), .CK(_08037_ ), .Q(\IF_ID_pc [21] ), .QN(_08130_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00248_ ), .CK(_08037_ ), .Q(\IF_ID_pc [20] ), .QN(_08129_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00249_ ), .CK(_08037_ ), .Q(\IF_ID_pc [19] ), .QN(_08128_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00250_ ), .CK(_08037_ ), .Q(\IF_ID_pc [18] ), .QN(_08127_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00251_ ), .CK(_08037_ ), .Q(\IF_ID_pc [17] ), .QN(_08126_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00252_ ), .CK(_08037_ ), .Q(\IF_ID_pc [16] ), .QN(_08125_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00253_ ), .CK(_08037_ ), .Q(\IF_ID_pc [15] ), .QN(_08124_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00254_ ), .CK(_08037_ ), .Q(\IF_ID_pc [14] ), .QN(_08123_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00255_ ), .CK(_08037_ ), .Q(\IF_ID_pc [13] ), .QN(_08122_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00256_ ), .CK(_08037_ ), .Q(\IF_ID_pc [12] ), .QN(_08121_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00257_ ), .CK(_08037_ ), .Q(\IF_ID_pc [29] ), .QN(_08120_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00258_ ), .CK(_08037_ ), .Q(\IF_ID_pc [11] ), .QN(_08119_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00259_ ), .CK(_08037_ ), .Q(\IF_ID_pc [10] ), .QN(_08118_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00260_ ), .CK(_08037_ ), .Q(\IF_ID_pc [9] ), .QN(_08117_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00261_ ), .CK(_08037_ ), .Q(\IF_ID_pc [8] ), .QN(_08116_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00262_ ), .CK(_08037_ ), .Q(\IF_ID_pc [7] ), .QN(_08115_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00263_ ), .CK(_08037_ ), .Q(\IF_ID_pc [6] ), .QN(_08114_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00264_ ), .CK(_08037_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00265_ ), .CK(_08037_ ), .Q(\IF_ID_pc [4] ), .QN(_08113_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00267_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08112_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00266_ ), .CK(_08037_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00269_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08110_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00268_ ), .CK(_08037_ ), .Q(\IF_ID_pc [2] ), .QN(_08111_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00270_ ), .CK(_08037_ ), .Q(\IF_ID_pc [28] ), .QN(_08109_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00271_ ), .CK(_08037_ ), .Q(\IF_ID_pc [1] ), .QN(_08108_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00272_ ), .CK(_08037_ ), .Q(\IF_ID_pc [27] ), .QN(_08107_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00273_ ), .CK(_08037_ ), .Q(\IF_ID_pc [26] ), .QN(_08106_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00274_ ), .CK(_08037_ ), .Q(\IF_ID_pc [25] ), .QN(_08105_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00275_ ), .CK(_08037_ ), .Q(\IF_ID_pc [24] ), .QN(_08104_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00276_ ), .CK(_08037_ ), .Q(\IF_ID_pc [23] ), .QN(_08103_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00277_ ), .CK(_08037_ ), .Q(\IF_ID_pc [22] ), .QN(_08102_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00278_ ), .CK(_08037_ ), .Q(\IF_ID_pc [31] ), .QN(_08101_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08909_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08100_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00279_ ), .CK(_08036_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08908_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00281_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00280_ ), .CK(_08035_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08099_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08910_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08911_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08912_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08913_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08914_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08915_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08916_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08917_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08918_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08919_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08920_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08921_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08922_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08923_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08924_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08925_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08926_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08927_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08928_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08929_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08930_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08931_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08932_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08933_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08934_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08935_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08936_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08937_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08938_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08939_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08940_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08034_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08941_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08942_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08943_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08944_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08945_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08946_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08947_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08948_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08949_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08950_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08951_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08952_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08953_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08954_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08955_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08956_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08957_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08958_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08959_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08960_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08961_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08962_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08963_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08964_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08965_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08966_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08967_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08968_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08969_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08970_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08971_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08972_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08033_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08098_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PP0P__Q ( .D(_00282_ ), .CK(_08032_ ), .Q(LS_WB_pc ), .QN(_08097_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PP0P__Q ( .D(_00283_ ), .CK(_08031_ ), .Q(\mylsu.previous_load_done ), .QN(_08973_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08974_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08975_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08976_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(_08977_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_08034_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_08034_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08978_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_08034_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08096_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00284_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08095_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00285_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08094_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00286_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08093_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00287_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08092_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00288_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08091_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00289_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08090_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00290_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08089_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00291_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08088_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00292_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08087_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00293_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08086_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00294_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08085_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00295_ ), .CK(_08034_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08979_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_08034_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08980_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_08034_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08981_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_08034_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08982_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_08034_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08983_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08984_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08985_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08986_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08987_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08988_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08989_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08990_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08991_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08992_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08993_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08994_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08995_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08996_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08997_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08998_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08999_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_09000_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_09001_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_09002_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_09003_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_09004_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_09005_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_09006_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_09007_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_09008_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_09009_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_09010_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_09011_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_09012_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_09013_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_09014_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_08034_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_09015_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_09016_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_09017_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_09018_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_09019_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_09020_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_09021_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_09022_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_09023_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_09024_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_09025_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_09026_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_09027_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_09028_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_09029_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_09030_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_09031_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_09032_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_09033_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_09034_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_09035_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_09036_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_09037_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_09038_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_09039_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_09040_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_09041_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_09042_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_09043_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_09044_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_09045_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_09046_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_08030_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08084_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q ( .D(_00296_ ), .CK(_08029_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_08083_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_1 ( .D(_00297_ ), .CK(_08029_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08082_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_2 ( .D(_00298_ ), .CK(_08029_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08081_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_3 ( .D(_00299_ ), .CK(_08029_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08080_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_4 ( .D(_00300_ ), .CK(_08029_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08079_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_5 ( .D(_00301_ ), .CK(_08029_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08078_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PP0P__Q ( .D(_00302_ ), .CK(_08029_ ), .Q(LS_WB_wen_reg ), .QN(_09047_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_09048_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_09049_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08028_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08027_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08026_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08025_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08024_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08023_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08022_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08021_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08020_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08019_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08018_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08017_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08016_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08015_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08014_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_1_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_10_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_11_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_12_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_13_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_14_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_15_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_16_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_17_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_18_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_19_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_2_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_20_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_21_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_22_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_23_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_24_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_25_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_26_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_27_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_28_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_29_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_3_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_30_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_31_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_4_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_5_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_6_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_7_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_8_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[2]_$_DFFE_PP__Q_9_D ), .CK(_08013_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00303_ ), .CK(_08012_ ), .Q(loaduse_clear ), .QN(_09050_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_09051_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_09052_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08077_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(excp_written ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(\myifu.to_reset ), .Z(fanout_net_44 ) );
BUF_X8 fanout_buf_45 ( .A(\mylsu.state [3] ), .Z(fanout_net_45 ) );

endmodule
