//Generate the verilog at 2025-09-29T16:42:59 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[0]_$_DFFE_PP__Q_E ;
wire \mycsreg.CSReg[1]_$_DFFE_PP__Q_E ;
wire \mycsreg.CSReg[2]_$_DFFE_PP__Q_E ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_E ;
wire \mycsreg.excp_written_$_SDFFE_PP0P__Q_E ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ;
wire \myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[4]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[5]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[6]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data[7]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.tag[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[3]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

AND3_X4 _09025_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01510_ ) );
AND3_X4 _09026_ ( .A1(_01510_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01511_ ) );
AND3_X4 _09027_ ( .A1(_01511_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01512_ ) );
AND2_X2 _09028_ ( .A1(_01512_ ), .A2(\myclint.mtime [7] ), .ZN(_01513_ ) );
AND4_X1 _09029_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01514_ ) );
AND2_X1 _09030_ ( .A1(\myclint.mtime [10] ), .A2(\myclint.mtime [11] ), .ZN(_01515_ ) );
AND4_X1 _09031_ ( .A1(\myclint.mtime [8] ), .A2(_01514_ ), .A3(\myclint.mtime [9] ), .A4(_01515_ ), .ZN(_01516_ ) );
NAND2_X1 _09032_ ( .A1(_01513_ ), .A2(_01516_ ), .ZN(_01517_ ) );
AND2_X1 _09033_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_01518_ ) );
AND3_X1 _09034_ ( .A1(_01518_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01519_ ) );
AND4_X1 _09035_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01520_ ) );
AND2_X1 _09036_ ( .A1(_01519_ ), .A2(_01520_ ), .ZN(_01521_ ) );
AND2_X1 _09037_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01522_ ) );
AND2_X1 _09038_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01523_ ) );
AND2_X1 _09039_ ( .A1(\myclint.mtime [26] ), .A2(\myclint.mtime [27] ), .ZN(_01524_ ) );
AND3_X1 _09040_ ( .A1(_01524_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_01525_ ) );
NAND4_X1 _09041_ ( .A1(_01521_ ), .A2(_01522_ ), .A3(_01523_ ), .A4(_01525_ ), .ZN(_01526_ ) );
NOR2_X1 _09042_ ( .A1(_01517_ ), .A2(_01526_ ), .ZN(_01527_ ) );
AND2_X1 _09043_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01528_ ) );
AND3_X1 _09044_ ( .A1(_01528_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01529_ ) );
AND2_X1 _09045_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [39] ), .ZN(_01530_ ) );
AND2_X1 _09046_ ( .A1(\myclint.mtime [36] ), .A2(\myclint.mtime [37] ), .ZN(_01531_ ) );
AND3_X1 _09047_ ( .A1(_01529_ ), .A2(_01530_ ), .A3(_01531_ ), .ZN(_01532_ ) );
AND2_X1 _09048_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01533_ ) );
AND3_X1 _09049_ ( .A1(_01533_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01534_ ) );
AND2_X2 _09050_ ( .A1(\myclint.mtime [42] ), .A2(\myclint.mtime [43] ), .ZN(_01535_ ) );
AND3_X1 _09051_ ( .A1(_01535_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01536_ ) );
AND3_X1 _09052_ ( .A1(_01532_ ), .A2(_01534_ ), .A3(_01536_ ), .ZN(_01537_ ) );
AND2_X1 _09053_ ( .A1(_01527_ ), .A2(_01537_ ), .ZN(_01538_ ) );
AND2_X1 _09054_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01539_ ) );
AND2_X1 _09055_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01540_ ) );
AND2_X1 _09056_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01541_ ) );
AND2_X1 _09057_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01542_ ) );
AND4_X1 _09058_ ( .A1(_01539_ ), .A2(_01540_ ), .A3(_01541_ ), .A4(_01542_ ), .ZN(_01543_ ) );
AND2_X1 _09059_ ( .A1(_01538_ ), .A2(_01543_ ), .ZN(_01544_ ) );
AND4_X1 _09060_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01545_ ) );
AND2_X1 _09061_ ( .A1(_01544_ ), .A2(_01545_ ), .ZN(_01546_ ) );
AND3_X1 _09062_ ( .A1(_01546_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01547_ ) );
INV_X1 _09063_ ( .A(_01547_ ), .ZN(_01548_ ) );
OR3_X1 _09064_ ( .A1(_01548_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [63] ), .ZN(_01549_ ) );
OAI21_X1 _09065_ ( .A(\myclint.mtime [63] ), .B1(_01548_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01550_ ) );
AOI21_X1 _09066_ ( .A(fanout_net_1 ), .B1(_01549_ ), .B2(_01550_ ), .ZN(_00000_ ) );
XNOR2_X1 _09067_ ( .A(_01547_ ), .B(\myclint.mtime [62] ), .ZN(_01551_ ) );
NOR2_X1 _09068_ ( .A1(_01551_ ), .A2(fanout_net_1 ), .ZN(_00001_ ) );
AND2_X1 _09069_ ( .A1(_01541_ ), .A2(_01542_ ), .ZN(_01552_ ) );
AND2_X1 _09070_ ( .A1(_01538_ ), .A2(_01552_ ), .ZN(_01553_ ) );
INV_X1 _09071_ ( .A(_01553_ ), .ZN(_01554_ ) );
OR3_X1 _09072_ ( .A1(_01554_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [53] ), .ZN(_01555_ ) );
OAI21_X1 _09073_ ( .A(\myclint.mtime [53] ), .B1(_01554_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01556_ ) );
AOI21_X1 _09074_ ( .A(fanout_net_1 ), .B1(_01555_ ), .B2(_01556_ ), .ZN(_00002_ ) );
XNOR2_X1 _09075_ ( .A(_01553_ ), .B(\myclint.mtime [52] ), .ZN(_01557_ ) );
NOR2_X1 _09076_ ( .A1(_01557_ ), .A2(fanout_net_1 ), .ZN(_00003_ ) );
INV_X1 _09077_ ( .A(fanout_net_1 ), .ZN(_01558_ ) );
BUF_X4 _09078_ ( .A(_01558_ ), .Z(_01559_ ) );
BUF_X4 _09079_ ( .A(_01559_ ), .Z(_01560_ ) );
AND3_X4 _09080_ ( .A1(_01512_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01561_ ) );
AND3_X2 _09081_ ( .A1(_01561_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01562_ ) );
AND3_X4 _09082_ ( .A1(_01562_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01563_ ) );
AND3_X2 _09083_ ( .A1(_01563_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01564_ ) );
AND3_X4 _09084_ ( .A1(_01564_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01565_ ) );
AND3_X4 _09085_ ( .A1(_01565_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01566_ ) );
AND3_X4 _09086_ ( .A1(_01566_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01567_ ) );
AND3_X4 _09087_ ( .A1(_01567_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01568_ ) );
AND3_X4 _09088_ ( .A1(_01568_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01569_ ) );
AND3_X4 _09089_ ( .A1(_01569_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01570_ ) );
AND2_X4 _09090_ ( .A1(_01570_ ), .A2(\myclint.mtime [27] ), .ZN(_01571_ ) );
AND4_X1 _09091_ ( .A1(\myclint.mtime [33] ), .A2(_01571_ ), .A3(_01522_ ), .A4(_01523_ ), .ZN(_01572_ ) );
AND3_X2 _09092_ ( .A1(_01572_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01573_ ) );
AND2_X1 _09093_ ( .A1(_01573_ ), .A2(\myclint.mtime [35] ), .ZN(_01574_ ) );
AND3_X1 _09094_ ( .A1(_01574_ ), .A2(_01530_ ), .A3(_01531_ ), .ZN(_01575_ ) );
AND2_X2 _09095_ ( .A1(_01575_ ), .A2(\myclint.mtime [40] ), .ZN(_01576_ ) );
AND2_X2 _09096_ ( .A1(_01576_ ), .A2(\myclint.mtime [41] ), .ZN(_01577_ ) );
AND2_X2 _09097_ ( .A1(_01577_ ), .A2(_01535_ ), .ZN(_01578_ ) );
NAND2_X1 _09098_ ( .A1(_01578_ ), .A2(_01534_ ), .ZN(_01579_ ) );
INV_X1 _09099_ ( .A(_01542_ ), .ZN(_01580_ ) );
NOR3_X1 _09100_ ( .A1(_01579_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01580_ ), .ZN(_01581_ ) );
OAI21_X1 _09101_ ( .A(_01560_ ), .B1(_01581_ ), .B2(\myclint.mtime [51] ), .ZN(_01582_ ) );
AND2_X1 _09102_ ( .A1(_01571_ ), .A2(_01523_ ), .ZN(_01583_ ) );
AND3_X1 _09103_ ( .A1(_01583_ ), .A2(_01528_ ), .A3(_01522_ ), .ZN(_01584_ ) );
AND2_X2 _09104_ ( .A1(_01584_ ), .A2(\myclint.mtime [34] ), .ZN(_01585_ ) );
AND2_X1 _09105_ ( .A1(_01585_ ), .A2(\myclint.mtime [35] ), .ZN(_01586_ ) );
AND3_X1 _09106_ ( .A1(_01586_ ), .A2(_01530_ ), .A3(_01531_ ), .ZN(_01587_ ) );
AND2_X1 _09107_ ( .A1(_01587_ ), .A2(\myclint.mtime [40] ), .ZN(_01588_ ) );
AND2_X2 _09108_ ( .A1(_01588_ ), .A2(\myclint.mtime [41] ), .ZN(_01589_ ) );
AND2_X1 _09109_ ( .A1(_01589_ ), .A2(_01535_ ), .ZN(_01590_ ) );
AND2_X1 _09110_ ( .A1(_01590_ ), .A2(_01534_ ), .ZN(_01591_ ) );
INV_X1 _09111_ ( .A(_01591_ ), .ZN(_01592_ ) );
NOR3_X1 _09112_ ( .A1(_01592_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01580_ ), .ZN(_01593_ ) );
AOI21_X1 _09113_ ( .A(_01582_ ), .B1(_01593_ ), .B2(\myclint.mtime [51] ), .ZN(_00004_ ) );
INV_X1 _09114_ ( .A(_01527_ ), .ZN(_01594_ ) );
INV_X1 _09115_ ( .A(_01537_ ), .ZN(_01595_ ) );
OR4_X1 _09116_ ( .A1(\myclint.mtime [50] ), .A2(_01594_ ), .A3(_01580_ ), .A4(_01595_ ), .ZN(_01596_ ) );
AND3_X1 _09117_ ( .A1(_01527_ ), .A2(_01542_ ), .A3(_01537_ ), .ZN(_01597_ ) );
INV_X1 _09118_ ( .A(_01597_ ), .ZN(_01598_ ) );
NAND2_X1 _09119_ ( .A1(_01598_ ), .A2(\myclint.mtime [50] ), .ZN(_01599_ ) );
AOI21_X1 _09120_ ( .A(fanout_net_1 ), .B1(_01596_ ), .B2(_01599_ ), .ZN(_00005_ ) );
INV_X1 _09121_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01600_ ) );
AND4_X1 _09122_ ( .A1(\myclint.mtime [49] ), .A2(_01590_ ), .A3(_01600_ ), .A4(_01534_ ), .ZN(_01601_ ) );
BUF_X4 _09123_ ( .A(_01559_ ), .Z(_01602_ ) );
AND3_X1 _09124_ ( .A1(_01578_ ), .A2(_01600_ ), .A3(_01534_ ), .ZN(_01603_ ) );
OAI21_X1 _09125_ ( .A(_01602_ ), .B1(_01603_ ), .B2(\myclint.mtime [49] ), .ZN(_01604_ ) );
NOR2_X1 _09126_ ( .A1(_01601_ ), .A2(_01604_ ), .ZN(_00006_ ) );
OAI21_X1 _09127_ ( .A(\myclint.mtime [48] ), .B1(_01594_ ), .B2(_01595_ ), .ZN(_01605_ ) );
OR4_X1 _09128_ ( .A1(\myclint.mtime [48] ), .A2(_01517_ ), .A3(_01595_ ), .A4(_01526_ ), .ZN(_01606_ ) );
AOI21_X1 _09129_ ( .A(fanout_net_1 ), .B1(_01605_ ), .B2(_01606_ ), .ZN(_00007_ ) );
NAND3_X1 _09130_ ( .A1(_01577_ ), .A2(_01533_ ), .A3(_01535_ ), .ZN(_01607_ ) );
NOR2_X1 _09131_ ( .A1(_01607_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01608_ ) );
OAI21_X1 _09132_ ( .A(_01560_ ), .B1(_01608_ ), .B2(\myclint.mtime [47] ), .ZN(_01609_ ) );
NAND3_X1 _09133_ ( .A1(_01589_ ), .A2(\myclint.mtime [44] ), .A3(_01535_ ), .ZN(_01610_ ) );
INV_X1 _09134_ ( .A(\myclint.mtime [45] ), .ZN(_01611_ ) );
NOR3_X1 _09135_ ( .A1(_01610_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01611_ ), .ZN(_01612_ ) );
AOI21_X1 _09136_ ( .A(_01609_ ), .B1(_01612_ ), .B2(\myclint.mtime [47] ), .ZN(_00008_ ) );
AND2_X1 _09137_ ( .A1(_01527_ ), .A2(_01532_ ), .ZN(_01613_ ) );
AND3_X1 _09138_ ( .A1(_01613_ ), .A2(_01533_ ), .A3(_01536_ ), .ZN(_01614_ ) );
XNOR2_X1 _09139_ ( .A(_01614_ ), .B(\myclint.mtime [46] ), .ZN(_01615_ ) );
NOR2_X1 _09140_ ( .A1(_01615_ ), .A2(fanout_net_1 ), .ZN(_00009_ ) );
INV_X1 _09141_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01616_ ) );
NAND3_X1 _09142_ ( .A1(_01577_ ), .A2(_01616_ ), .A3(_01535_ ), .ZN(_01617_ ) );
AOI21_X1 _09143_ ( .A(fanout_net_1 ), .B1(_01617_ ), .B2(_01611_ ), .ZN(_01618_ ) );
NAND4_X1 _09144_ ( .A1(_01589_ ), .A2(\myclint.mtime [45] ), .A3(_01616_ ), .A4(_01535_ ), .ZN(_01619_ ) );
AND2_X1 _09145_ ( .A1(_01618_ ), .A2(_01619_ ), .ZN(_00010_ ) );
AND2_X1 _09146_ ( .A1(_01613_ ), .A2(_01536_ ), .ZN(_01620_ ) );
XNOR2_X1 _09147_ ( .A(_01620_ ), .B(\myclint.mtime [44] ), .ZN(_01621_ ) );
NOR2_X1 _09148_ ( .A1(_01621_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
INV_X1 _09149_ ( .A(_01546_ ), .ZN(_01622_ ) );
OR3_X1 _09150_ ( .A1(_01622_ ), .A2(\myclint.mtime [61] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01623_ ) );
OAI21_X1 _09151_ ( .A(\myclint.mtime [61] ), .B1(_01622_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01624_ ) );
AOI21_X1 _09152_ ( .A(fanout_net_1 ), .B1(_01623_ ), .B2(_01624_ ), .ZN(_00012_ ) );
INV_X1 _09153_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01625_ ) );
AND4_X1 _09154_ ( .A1(_01625_ ), .A2(_01588_ ), .A3(\myclint.mtime [41] ), .A4(\myclint.mtime [43] ), .ZN(_01626_ ) );
AND3_X1 _09155_ ( .A1(_01576_ ), .A2(_01625_ ), .A3(\myclint.mtime [41] ), .ZN(_01627_ ) );
OAI21_X1 _09156_ ( .A(_01602_ ), .B1(_01627_ ), .B2(\myclint.mtime [43] ), .ZN(_01628_ ) );
NOR2_X1 _09157_ ( .A1(_01626_ ), .A2(_01628_ ), .ZN(_00013_ ) );
AND3_X1 _09158_ ( .A1(_01613_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01629_ ) );
XNOR2_X1 _09159_ ( .A(_01629_ ), .B(\myclint.mtime [42] ), .ZN(_01630_ ) );
NOR2_X1 _09160_ ( .A1(_01630_ ), .A2(fanout_net_1 ), .ZN(_00014_ ) );
BUF_X4 _09161_ ( .A(_01559_ ), .Z(_01631_ ) );
INV_X1 _09162_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01632_ ) );
AND2_X1 _09163_ ( .A1(_01575_ ), .A2(_01632_ ), .ZN(_01633_ ) );
OAI21_X1 _09164_ ( .A(_01631_ ), .B1(_01633_ ), .B2(\myclint.mtime [41] ), .ZN(_01634_ ) );
AND3_X1 _09165_ ( .A1(_01587_ ), .A2(\myclint.mtime [41] ), .A3(_01632_ ), .ZN(_01635_ ) );
NOR2_X1 _09166_ ( .A1(_01634_ ), .A2(_01635_ ), .ZN(_00015_ ) );
XNOR2_X1 _09167_ ( .A(_01613_ ), .B(\myclint.mtime [40] ), .ZN(_01636_ ) );
NOR2_X1 _09168_ ( .A1(_01636_ ), .A2(fanout_net_1 ), .ZN(_00016_ ) );
NAND3_X1 _09169_ ( .A1(_01527_ ), .A2(_01531_ ), .A3(_01529_ ), .ZN(_01637_ ) );
OR3_X1 _09170_ ( .A1(_01637_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [39] ), .ZN(_01638_ ) );
OAI21_X1 _09171_ ( .A(\myclint.mtime [39] ), .B1(_01637_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01639_ ) );
AOI21_X1 _09172_ ( .A(fanout_net_1 ), .B1(_01638_ ), .B2(_01639_ ), .ZN(_00017_ ) );
OR2_X1 _09173_ ( .A1(_01637_ ), .A2(\myclint.mtime [38] ), .ZN(_01640_ ) );
NAND2_X1 _09174_ ( .A1(_01637_ ), .A2(\myclint.mtime [38] ), .ZN(_01641_ ) );
AOI21_X1 _09175_ ( .A(fanout_net_1 ), .B1(_01640_ ), .B2(_01641_ ), .ZN(_00018_ ) );
INV_X1 _09176_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01642_ ) );
AND4_X1 _09177_ ( .A1(\myclint.mtime [37] ), .A2(_01585_ ), .A3(_01642_ ), .A4(\myclint.mtime [35] ), .ZN(_01643_ ) );
AND3_X1 _09178_ ( .A1(_01573_ ), .A2(_01642_ ), .A3(\myclint.mtime [35] ), .ZN(_01644_ ) );
OAI21_X1 _09179_ ( .A(_01602_ ), .B1(_01644_ ), .B2(\myclint.mtime [37] ), .ZN(_01645_ ) );
NOR2_X1 _09180_ ( .A1(_01643_ ), .A2(_01645_ ), .ZN(_00019_ ) );
AND2_X1 _09181_ ( .A1(_01527_ ), .A2(_01529_ ), .ZN(_01646_ ) );
XNOR2_X1 _09182_ ( .A(_01646_ ), .B(\myclint.mtime [36] ), .ZN(_01647_ ) );
NOR2_X1 _09183_ ( .A1(_01647_ ), .A2(fanout_net_1 ), .ZN(_00020_ ) );
AND2_X1 _09184_ ( .A1(_01513_ ), .A2(_01516_ ), .ZN(_01648_ ) );
AND4_X1 _09185_ ( .A1(_01522_ ), .A2(_01521_ ), .A3(_01523_ ), .A4(_01525_ ), .ZN(_01649_ ) );
NAND3_X1 _09186_ ( .A1(_01648_ ), .A2(_01528_ ), .A3(_01649_ ), .ZN(_01650_ ) );
OR3_X1 _09187_ ( .A1(_01650_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [35] ), .ZN(_01651_ ) );
OAI21_X1 _09188_ ( .A(\myclint.mtime [35] ), .B1(_01650_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01652_ ) );
AOI21_X1 _09189_ ( .A(fanout_net_1 ), .B1(_01651_ ), .B2(_01652_ ), .ZN(_00021_ ) );
NAND4_X1 _09190_ ( .A1(_01571_ ), .A2(\myclint.mtime [33] ), .A3(_01522_ ), .A4(_01523_ ), .ZN(_01653_ ) );
INV_X1 _09191_ ( .A(\myclint.mtime [32] ), .ZN(_01654_ ) );
NOR2_X1 _09192_ ( .A1(_01653_ ), .A2(_01654_ ), .ZN(_01655_ ) );
OAI21_X1 _09193_ ( .A(_01631_ ), .B1(_01655_ ), .B2(\myclint.mtime [34] ), .ZN(_01656_ ) );
NOR2_X1 _09194_ ( .A1(_01656_ ), .A2(_01573_ ), .ZN(_00022_ ) );
XNOR2_X1 _09195_ ( .A(_01546_ ), .B(\myclint.mtime [60] ), .ZN(_01657_ ) );
NOR2_X1 _09196_ ( .A1(_01657_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
INV_X1 _09197_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01658_ ) );
AND3_X1 _09198_ ( .A1(_01583_ ), .A2(_01658_ ), .A3(_01522_ ), .ZN(_01659_ ) );
AND2_X1 _09199_ ( .A1(_01659_ ), .A2(\myclint.mtime [33] ), .ZN(_01660_ ) );
OAI21_X1 _09200_ ( .A(_01560_ ), .B1(_01659_ ), .B2(\myclint.mtime [33] ), .ZN(_01661_ ) );
NOR2_X1 _09201_ ( .A1(_01660_ ), .A2(_01661_ ), .ZN(_00024_ ) );
OAI21_X1 _09202_ ( .A(\myclint.mtime [32] ), .B1(_01517_ ), .B2(_01526_ ), .ZN(_01662_ ) );
NAND4_X1 _09203_ ( .A1(_01649_ ), .A2(_01513_ ), .A3(_01654_ ), .A4(_01516_ ), .ZN(_01663_ ) );
AOI21_X1 _09204_ ( .A(fanout_net_1 ), .B1(_01662_ ), .B2(_01663_ ), .ZN(_00025_ ) );
AND2_X1 _09205_ ( .A1(_01648_ ), .A2(_01521_ ), .ZN(_01664_ ) );
NAND3_X1 _09206_ ( .A1(_01664_ ), .A2(_01523_ ), .A3(_01525_ ), .ZN(_01665_ ) );
OR3_X1 _09207_ ( .A1(_01665_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [31] ), .ZN(_01666_ ) );
OAI21_X1 _09208_ ( .A(\myclint.mtime [31] ), .B1(_01665_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01667_ ) );
AOI21_X1 _09209_ ( .A(fanout_net_1 ), .B1(_01666_ ), .B2(_01667_ ), .ZN(_00026_ ) );
OR2_X1 _09210_ ( .A1(_01665_ ), .A2(\myclint.mtime [30] ), .ZN(_01668_ ) );
NAND2_X1 _09211_ ( .A1(_01665_ ), .A2(\myclint.mtime [30] ), .ZN(_01669_ ) );
AOI21_X1 _09212_ ( .A(fanout_net_1 ), .B1(_01668_ ), .B2(_01669_ ), .ZN(_00027_ ) );
INV_X1 _09213_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01670_ ) );
AND3_X1 _09214_ ( .A1(_01570_ ), .A2(_01670_ ), .A3(\myclint.mtime [27] ), .ZN(_01671_ ) );
AND2_X1 _09215_ ( .A1(_01671_ ), .A2(\myclint.mtime [29] ), .ZN(_01672_ ) );
OAI21_X1 _09216_ ( .A(_01560_ ), .B1(_01671_ ), .B2(\myclint.mtime [29] ), .ZN(_01673_ ) );
NOR2_X1 _09217_ ( .A1(_01672_ ), .A2(_01673_ ), .ZN(_00028_ ) );
NAND2_X1 _09218_ ( .A1(_01664_ ), .A2(_01525_ ), .ZN(_01674_ ) );
OR2_X1 _09219_ ( .A1(_01674_ ), .A2(\myclint.mtime [28] ), .ZN(_01675_ ) );
NAND2_X1 _09220_ ( .A1(_01674_ ), .A2(\myclint.mtime [28] ), .ZN(_01676_ ) );
AOI21_X1 _09221_ ( .A(fanout_net_1 ), .B1(_01675_ ), .B2(_01676_ ), .ZN(_00029_ ) );
INV_X1 _09222_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01677_ ) );
AND3_X1 _09223_ ( .A1(_01569_ ), .A2(_01677_ ), .A3(\myclint.mtime [25] ), .ZN(_01678_ ) );
AND2_X1 _09224_ ( .A1(_01678_ ), .A2(\myclint.mtime [27] ), .ZN(_01679_ ) );
OAI21_X1 _09225_ ( .A(_01560_ ), .B1(_01678_ ), .B2(\myclint.mtime [27] ), .ZN(_01680_ ) );
NOR2_X1 _09226_ ( .A1(_01679_ ), .A2(_01680_ ), .ZN(_00030_ ) );
AND2_X1 _09227_ ( .A1(_01569_ ), .A2(\myclint.mtime [25] ), .ZN(_01681_ ) );
OAI21_X1 _09228_ ( .A(_01631_ ), .B1(_01681_ ), .B2(\myclint.mtime [26] ), .ZN(_01682_ ) );
NOR2_X1 _09229_ ( .A1(_01682_ ), .A2(_01570_ ), .ZN(_00031_ ) );
INV_X1 _09230_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01683_ ) );
AND3_X1 _09231_ ( .A1(_01568_ ), .A2(_01683_ ), .A3(\myclint.mtime [23] ), .ZN(_01684_ ) );
AND2_X1 _09232_ ( .A1(_01684_ ), .A2(\myclint.mtime [25] ), .ZN(_01685_ ) );
OAI21_X1 _09233_ ( .A(_01560_ ), .B1(_01684_ ), .B2(\myclint.mtime [25] ), .ZN(_01686_ ) );
NOR2_X1 _09234_ ( .A1(_01685_ ), .A2(_01686_ ), .ZN(_00032_ ) );
AND2_X1 _09235_ ( .A1(_01568_ ), .A2(\myclint.mtime [23] ), .ZN(_01687_ ) );
OAI21_X1 _09236_ ( .A(_01631_ ), .B1(_01687_ ), .B2(\myclint.mtime [24] ), .ZN(_01688_ ) );
NOR2_X1 _09237_ ( .A1(_01688_ ), .A2(_01569_ ), .ZN(_00033_ ) );
NOR2_X1 _09238_ ( .A1(_01579_ ), .A2(_01580_ ), .ZN(_01689_ ) );
AND2_X1 _09239_ ( .A1(_01689_ ), .A2(_01541_ ), .ZN(_01690_ ) );
AND2_X1 _09240_ ( .A1(_01690_ ), .A2(_01540_ ), .ZN(_01691_ ) );
AND2_X1 _09241_ ( .A1(_01691_ ), .A2(_01539_ ), .ZN(_01692_ ) );
INV_X1 _09242_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01693_ ) );
AND2_X1 _09243_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01694_ ) );
AND3_X1 _09244_ ( .A1(_01692_ ), .A2(_01693_ ), .A3(_01694_ ), .ZN(_01695_ ) );
OAI21_X1 _09245_ ( .A(_01560_ ), .B1(_01695_ ), .B2(\myclint.mtime [59] ), .ZN(_01696_ ) );
AND2_X2 _09246_ ( .A1(_01591_ ), .A2(_01542_ ), .ZN(_01697_ ) );
AND2_X1 _09247_ ( .A1(_01697_ ), .A2(_01541_ ), .ZN(_01698_ ) );
AND2_X1 _09248_ ( .A1(_01698_ ), .A2(_01540_ ), .ZN(_01699_ ) );
AND2_X1 _09249_ ( .A1(_01699_ ), .A2(_01539_ ), .ZN(_01700_ ) );
AND3_X1 _09250_ ( .A1(_01700_ ), .A2(_01693_ ), .A3(_01694_ ), .ZN(_01701_ ) );
AOI21_X1 _09251_ ( .A(_01696_ ), .B1(_01701_ ), .B2(\myclint.mtime [59] ), .ZN(_00034_ ) );
AND2_X1 _09252_ ( .A1(_01648_ ), .A2(_01519_ ), .ZN(_01702_ ) );
NAND3_X1 _09253_ ( .A1(_01702_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01703_ ) );
OR3_X1 _09254_ ( .A1(_01703_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01704_ ) );
OAI21_X1 _09255_ ( .A(\myclint.mtime [23] ), .B1(_01703_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01705_ ) );
AOI21_X1 _09256_ ( .A(fanout_net_1 ), .B1(_01704_ ), .B2(_01705_ ), .ZN(_00035_ ) );
AND2_X1 _09257_ ( .A1(_01567_ ), .A2(\myclint.mtime [21] ), .ZN(_01706_ ) );
OAI21_X1 _09258_ ( .A(_01631_ ), .B1(_01706_ ), .B2(\myclint.mtime [22] ), .ZN(_01707_ ) );
NOR2_X1 _09259_ ( .A1(_01707_ ), .A2(_01568_ ), .ZN(_00036_ ) );
INV_X1 _09260_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01708_ ) );
AND3_X1 _09261_ ( .A1(_01566_ ), .A2(_01708_ ), .A3(\myclint.mtime [19] ), .ZN(_01709_ ) );
AND2_X1 _09262_ ( .A1(_01709_ ), .A2(\myclint.mtime [21] ), .ZN(_01710_ ) );
OAI21_X1 _09263_ ( .A(_01560_ ), .B1(_01709_ ), .B2(\myclint.mtime [21] ), .ZN(_01711_ ) );
NOR2_X1 _09264_ ( .A1(_01710_ ), .A2(_01711_ ), .ZN(_00037_ ) );
AND2_X1 _09265_ ( .A1(_01566_ ), .A2(\myclint.mtime [19] ), .ZN(_01712_ ) );
OAI21_X1 _09266_ ( .A(_01631_ ), .B1(_01712_ ), .B2(\myclint.mtime [20] ), .ZN(_01713_ ) );
NOR2_X1 _09267_ ( .A1(_01713_ ), .A2(_01567_ ), .ZN(_00038_ ) );
NAND3_X1 _09268_ ( .A1(_01648_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01714_ ) );
OR3_X1 _09269_ ( .A1(_01714_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01715_ ) );
OAI21_X1 _09270_ ( .A(\myclint.mtime [19] ), .B1(_01714_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01716_ ) );
AOI21_X1 _09271_ ( .A(fanout_net_1 ), .B1(_01715_ ), .B2(_01716_ ), .ZN(_00039_ ) );
AND2_X1 _09272_ ( .A1(_01565_ ), .A2(\myclint.mtime [17] ), .ZN(_01717_ ) );
OAI21_X1 _09273_ ( .A(_01631_ ), .B1(_01717_ ), .B2(\myclint.mtime [18] ), .ZN(_01718_ ) );
NOR2_X1 _09274_ ( .A1(_01718_ ), .A2(_01566_ ), .ZN(_00040_ ) );
INV_X1 _09275_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01719_ ) );
AND3_X1 _09276_ ( .A1(_01564_ ), .A2(_01719_ ), .A3(\myclint.mtime [15] ), .ZN(_01720_ ) );
AND2_X1 _09277_ ( .A1(_01720_ ), .A2(\myclint.mtime [17] ), .ZN(_01721_ ) );
OAI21_X1 _09278_ ( .A(_01560_ ), .B1(_01720_ ), .B2(\myclint.mtime [17] ), .ZN(_01722_ ) );
NOR2_X1 _09279_ ( .A1(_01721_ ), .A2(_01722_ ), .ZN(_00041_ ) );
AND2_X1 _09280_ ( .A1(_01564_ ), .A2(\myclint.mtime [15] ), .ZN(_01723_ ) );
OAI21_X1 _09281_ ( .A(_01602_ ), .B1(_01723_ ), .B2(\myclint.mtime [16] ), .ZN(_01724_ ) );
NOR2_X1 _09282_ ( .A1(_01724_ ), .A2(_01565_ ), .ZN(_00042_ ) );
AND3_X1 _09283_ ( .A1(_01515_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01725_ ) );
AND2_X1 _09284_ ( .A1(_01513_ ), .A2(_01725_ ), .ZN(_01726_ ) );
NAND3_X1 _09285_ ( .A1(_01726_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01727_ ) );
OR3_X1 _09286_ ( .A1(_01727_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01728_ ) );
OAI21_X1 _09287_ ( .A(\myclint.mtime [15] ), .B1(_01727_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01729_ ) );
AOI21_X1 _09288_ ( .A(fanout_net_1 ), .B1(_01728_ ), .B2(_01729_ ), .ZN(_00043_ ) );
AND2_X1 _09289_ ( .A1(_01563_ ), .A2(\myclint.mtime [13] ), .ZN(_01730_ ) );
OAI21_X1 _09290_ ( .A(_01602_ ), .B1(_01730_ ), .B2(\myclint.mtime [14] ), .ZN(_01731_ ) );
NOR2_X1 _09291_ ( .A1(_01731_ ), .A2(_01564_ ), .ZN(_00044_ ) );
NAND3_X1 _09292_ ( .A1(_01538_ ), .A2(_01694_ ), .A3(_01543_ ), .ZN(_01732_ ) );
OR2_X1 _09293_ ( .A1(_01732_ ), .A2(\myclint.mtime [58] ), .ZN(_01733_ ) );
NAND2_X1 _09294_ ( .A1(_01732_ ), .A2(\myclint.mtime [58] ), .ZN(_01734_ ) );
AOI21_X1 _09295_ ( .A(fanout_net_1 ), .B1(_01733_ ), .B2(_01734_ ), .ZN(_00045_ ) );
INV_X1 _09296_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01735_ ) );
AND3_X1 _09297_ ( .A1(_01562_ ), .A2(_01735_ ), .A3(\myclint.mtime [11] ), .ZN(_01736_ ) );
AND2_X1 _09298_ ( .A1(_01736_ ), .A2(\myclint.mtime [13] ), .ZN(_01737_ ) );
OAI21_X1 _09299_ ( .A(_01560_ ), .B1(_01736_ ), .B2(\myclint.mtime [13] ), .ZN(_01738_ ) );
NOR2_X1 _09300_ ( .A1(_01737_ ), .A2(_01738_ ), .ZN(_00046_ ) );
XNOR2_X1 _09301_ ( .A(_01726_ ), .B(\myclint.mtime [12] ), .ZN(_01739_ ) );
NOR2_X1 _09302_ ( .A1(_01739_ ), .A2(fanout_net_1 ), .ZN(_00047_ ) );
NAND3_X1 _09303_ ( .A1(_01513_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01740_ ) );
OR3_X1 _09304_ ( .A1(_01740_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_01741_ ) );
OAI21_X1 _09305_ ( .A(\myclint.mtime [11] ), .B1(_01740_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01742_ ) );
AOI21_X1 _09306_ ( .A(fanout_net_1 ), .B1(_01741_ ), .B2(_01742_ ), .ZN(_00048_ ) );
AOI21_X1 _09307_ ( .A(\myclint.mtime [10] ), .B1(_01561_ ), .B2(\myclint.mtime [9] ), .ZN(_01743_ ) );
NOR3_X1 _09308_ ( .A1(_01562_ ), .A2(_01743_ ), .A3(fanout_net_1 ), .ZN(_00049_ ) );
INV_X1 _09309_ ( .A(_01513_ ), .ZN(_01744_ ) );
OR3_X1 _09310_ ( .A1(_01744_ ), .A2(\myclint.mtime [9] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01745_ ) );
OAI21_X1 _09311_ ( .A(\myclint.mtime [9] ), .B1(_01744_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01746_ ) );
AOI21_X1 _09312_ ( .A(fanout_net_1 ), .B1(_01745_ ), .B2(_01746_ ), .ZN(_00050_ ) );
OAI21_X1 _09313_ ( .A(_01602_ ), .B1(_01513_ ), .B2(\myclint.mtime [8] ), .ZN(_01747_ ) );
NOR2_X1 _09314_ ( .A1(_01747_ ), .A2(_01561_ ), .ZN(_00051_ ) );
AND2_X1 _09315_ ( .A1(_01511_ ), .A2(\myclint.mtime [5] ), .ZN(_01748_ ) );
INV_X1 _09316_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01749_ ) );
AND3_X1 _09317_ ( .A1(_01748_ ), .A2(_01749_ ), .A3(\myclint.mtime [7] ), .ZN(_01750_ ) );
AOI21_X1 _09318_ ( .A(\myclint.mtime [7] ), .B1(_01748_ ), .B2(_01749_ ), .ZN(_01751_ ) );
NOR3_X1 _09319_ ( .A1(_01750_ ), .A2(_01751_ ), .A3(fanout_net_2 ), .ZN(_00052_ ) );
OAI21_X1 _09320_ ( .A(_01602_ ), .B1(_01748_ ), .B2(\myclint.mtime [6] ), .ZN(_01752_ ) );
NOR2_X1 _09321_ ( .A1(_01752_ ), .A2(_01512_ ), .ZN(_00053_ ) );
AND2_X1 _09322_ ( .A1(_01510_ ), .A2(\myclint.mtime [3] ), .ZN(_01753_ ) );
INV_X1 _09323_ ( .A(_01753_ ), .ZN(_01754_ ) );
OR3_X1 _09324_ ( .A1(_01754_ ), .A2(\myclint.mtime [5] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01755_ ) );
OAI21_X1 _09325_ ( .A(\myclint.mtime [5] ), .B1(_01754_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01756_ ) );
AOI21_X1 _09326_ ( .A(fanout_net_2 ), .B1(_01755_ ), .B2(_01756_ ), .ZN(_00054_ ) );
OAI21_X1 _09327_ ( .A(_01602_ ), .B1(_01753_ ), .B2(\myclint.mtime [4] ), .ZN(_01757_ ) );
NOR2_X1 _09328_ ( .A1(_01757_ ), .A2(_01511_ ), .ZN(_00055_ ) );
INV_X1 _09329_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01758_ ) );
AND3_X1 _09330_ ( .A1(_01691_ ), .A2(_01758_ ), .A3(_01539_ ), .ZN(_01759_ ) );
OAI21_X1 _09331_ ( .A(_01559_ ), .B1(_01759_ ), .B2(\myclint.mtime [57] ), .ZN(_01760_ ) );
AND3_X1 _09332_ ( .A1(_01699_ ), .A2(_01758_ ), .A3(_01539_ ), .ZN(_01761_ ) );
AOI21_X1 _09333_ ( .A(_01760_ ), .B1(_01761_ ), .B2(\myclint.mtime [57] ), .ZN(_00056_ ) );
AND2_X1 _09334_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01762_ ) );
INV_X1 _09335_ ( .A(_01762_ ), .ZN(_01763_ ) );
OR3_X1 _09336_ ( .A1(_01763_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01764_ ) );
OAI21_X1 _09337_ ( .A(\myclint.mtime [3] ), .B1(_01763_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01765_ ) );
AOI21_X1 _09338_ ( .A(fanout_net_2 ), .B1(_01764_ ), .B2(_01765_ ), .ZN(_00057_ ) );
AOI21_X1 _09339_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01766_ ) );
NOR3_X1 _09340_ ( .A1(_01510_ ), .A2(_01766_ ), .A3(fanout_net_2 ), .ZN(_00058_ ) );
NOR2_X1 _09341_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01767_ ) );
NOR3_X1 _09342_ ( .A1(_01762_ ), .A2(_01767_ ), .A3(fanout_net_2 ), .ZN(_00059_ ) );
INV_X1 _09343_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_01768_ ) );
NOR2_X1 _09344_ ( .A1(_01768_ ), .A2(fanout_net_2 ), .ZN(_00060_ ) );
XNOR2_X1 _09345_ ( .A(_01544_ ), .B(\myclint.mtime [56] ), .ZN(_01769_ ) );
NOR2_X1 _09346_ ( .A1(_01769_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
NAND3_X1 _09347_ ( .A1(_01538_ ), .A2(_01540_ ), .A3(_01552_ ), .ZN(_01770_ ) );
OR3_X1 _09348_ ( .A1(_01770_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01771_ ) );
OAI21_X1 _09349_ ( .A(\myclint.mtime [55] ), .B1(_01770_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01772_ ) );
AOI21_X1 _09350_ ( .A(fanout_net_2 ), .B1(_01771_ ), .B2(_01772_ ), .ZN(_00062_ ) );
OR2_X1 _09351_ ( .A1(_01770_ ), .A2(\myclint.mtime [54] ), .ZN(_01773_ ) );
NAND2_X1 _09352_ ( .A1(_01770_ ), .A2(\myclint.mtime [54] ), .ZN(_01774_ ) );
AOI21_X1 _09353_ ( .A(fanout_net_2 ), .B1(_01773_ ), .B2(_01774_ ), .ZN(_00063_ ) );
INV_X32 _09354_ ( .A(fanout_net_41 ), .ZN(_01775_ ) );
BUF_X32 _09355_ ( .A(_01775_ ), .Z(_01776_ ) );
OR2_X2 _09356_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[1][10] ), .ZN(_01777_ ) );
INV_X16 _09357_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01778_ ) );
BUF_X4 _09358_ ( .A(_01778_ ), .Z(_01779_ ) );
OAI211_X1 _09359_ ( .A(_01777_ ), .B(_01779_ ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[0][10] ), .ZN(_01780_ ) );
OR2_X2 _09360_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[3][10] ), .ZN(_01781_ ) );
OAI211_X2 _09361_ ( .A(_01781_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[2][10] ), .ZN(_01782_ ) );
NAND2_X1 _09362_ ( .A1(_01780_ ), .A2(_01782_ ), .ZN(_01783_ ) );
XNOR2_X1 _09363_ ( .A(_01783_ ), .B(\IF_ID_pc [15] ), .ZN(_01784_ ) );
INV_X1 _09364_ ( .A(\IF_ID_pc [23] ), .ZN(_01785_ ) );
MUX2_X1 _09365_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(fanout_net_41 ), .Z(_01786_ ) );
MUX2_X1 _09366_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(fanout_net_41 ), .Z(_01787_ ) );
MUX2_X2 _09367_ ( .A(_01786_ ), .B(_01787_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01788_ ) );
INV_X1 _09368_ ( .A(\IF_ID_pc [7] ), .ZN(_01789_ ) );
MUX2_X1 _09369_ ( .A(\myifu.myicache.tag[2][2] ), .B(\myifu.myicache.tag[3][2] ), .S(fanout_net_41 ), .Z(_01790_ ) );
OR2_X1 _09370_ ( .A1(_01790_ ), .A2(_01779_ ), .ZN(_01791_ ) );
MUX2_X1 _09371_ ( .A(\myifu.myicache.tag[0][2] ), .B(\myifu.myicache.tag[1][2] ), .S(fanout_net_41 ), .Z(_01792_ ) );
OR2_X1 _09372_ ( .A1(_01792_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01793_ ) );
AND2_X1 _09373_ ( .A1(_01791_ ), .A2(_01793_ ), .ZN(_01794_ ) );
OAI221_X1 _09374_ ( .A(_01784_ ), .B1(_01785_ ), .B2(_01788_ ), .C1(_01789_ ), .C2(_01794_ ), .ZN(_01795_ ) );
OR2_X4 _09375_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[1][22] ), .ZN(_01796_ ) );
OAI211_X4 _09376_ ( .A(_01796_ ), .B(_01778_ ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[0][22] ), .ZN(_01797_ ) );
OR2_X1 _09377_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[3][22] ), .ZN(_01798_ ) );
OAI211_X2 _09378_ ( .A(_01798_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[2][22] ), .ZN(_01799_ ) );
AOI21_X2 _09379_ ( .A(\IF_ID_pc [27] ), .B1(_01797_ ), .B2(_01799_ ), .ZN(_01800_ ) );
INV_X1 _09380_ ( .A(\IF_ID_pc [29] ), .ZN(_01801_ ) );
MUX2_X1 _09381_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(fanout_net_41 ), .Z(_01802_ ) );
MUX2_X1 _09382_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(fanout_net_41 ), .Z(_01803_ ) );
MUX2_X2 _09383_ ( .A(_01802_ ), .B(_01803_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01804_ ) );
AOI21_X2 _09384_ ( .A(_01800_ ), .B1(_01801_ ), .B2(_01804_ ), .ZN(_01805_ ) );
INV_X1 _09385_ ( .A(\IF_ID_pc [21] ), .ZN(_01806_ ) );
MUX2_X1 _09386_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(fanout_net_41 ), .Z(_01807_ ) );
MUX2_X1 _09387_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(fanout_net_41 ), .Z(_01808_ ) );
MUX2_X2 _09388_ ( .A(_01807_ ), .B(_01808_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01809_ ) );
INV_X1 _09389_ ( .A(\IF_ID_pc [8] ), .ZN(_01810_ ) );
MUX2_X1 _09390_ ( .A(\myifu.myicache.tag[0][3] ), .B(\myifu.myicache.tag[1][3] ), .S(fanout_net_41 ), .Z(_01811_ ) );
MUX2_X1 _09391_ ( .A(\myifu.myicache.tag[2][3] ), .B(\myifu.myicache.tag[3][3] ), .S(fanout_net_41 ), .Z(_01812_ ) );
MUX2_X2 _09392_ ( .A(_01811_ ), .B(_01812_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01813_ ) );
OAI221_X1 _09393_ ( .A(_01805_ ), .B1(_01806_ ), .B2(_01809_ ), .C1(_01810_ ), .C2(_01813_ ), .ZN(_01814_ ) );
MUX2_X1 _09394_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(fanout_net_41 ), .Z(_01815_ ) );
MUX2_X1 _09395_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_41 ), .Z(_01816_ ) );
MUX2_X2 _09396_ ( .A(_01815_ ), .B(_01816_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01817_ ) );
XNOR2_X2 _09397_ ( .A(_01817_ ), .B(\IF_ID_pc [25] ), .ZN(_01818_ ) );
BUF_X16 _09398_ ( .A(_01775_ ), .Z(_01819_ ) );
OR2_X2 _09399_ ( .A1(_01819_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01820_ ) );
OAI211_X1 _09400_ ( .A(_01820_ ), .B(_01779_ ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01821_ ) );
OR2_X2 _09401_ ( .A1(_01819_ ), .A2(\myifu.myicache.tag[3][12] ), .ZN(_01822_ ) );
OAI211_X1 _09402_ ( .A(_01822_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[2][12] ), .ZN(_01823_ ) );
INV_X1 _09403_ ( .A(\IF_ID_pc [17] ), .ZN(_01824_ ) );
AND3_X1 _09404_ ( .A1(_01821_ ), .A2(_01823_ ), .A3(_01824_ ), .ZN(_01825_ ) );
AOI21_X1 _09405_ ( .A(_01824_ ), .B1(_01821_ ), .B2(_01823_ ), .ZN(_01826_ ) );
OAI21_X1 _09406_ ( .A(_01818_ ), .B1(_01825_ ), .B2(_01826_ ), .ZN(_01827_ ) );
NAND2_X1 _09407_ ( .A1(_01809_ ), .A2(_01806_ ), .ZN(_01828_ ) );
MUX2_X1 _09408_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(fanout_net_41 ), .Z(_01829_ ) );
MUX2_X1 _09409_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(fanout_net_41 ), .Z(_01830_ ) );
MUX2_X2 _09410_ ( .A(_01829_ ), .B(_01830_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01831_ ) );
INV_X1 _09411_ ( .A(\IF_ID_pc [12] ), .ZN(_01832_ ) );
NAND2_X1 _09412_ ( .A1(_01831_ ), .A2(_01832_ ), .ZN(_01833_ ) );
OR2_X4 _09413_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[3][13] ), .ZN(_01834_ ) );
OAI211_X4 _09414_ ( .A(_01834_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[2][13] ), .ZN(_01835_ ) );
OR2_X1 _09415_ ( .A1(fanout_net_41 ), .A2(\myifu.myicache.tag[0][13] ), .ZN(_01836_ ) );
OAI211_X1 _09416_ ( .A(_01836_ ), .B(_01778_ ), .C1(_01819_ ), .C2(\myifu.myicache.tag[1][13] ), .ZN(_01837_ ) );
NAND3_X1 _09417_ ( .A1(_01835_ ), .A2(\IF_ID_pc [18] ), .A3(_01837_ ), .ZN(_01838_ ) );
NAND3_X1 _09418_ ( .A1(_01797_ ), .A2(_01799_ ), .A3(\IF_ID_pc [27] ), .ZN(_01839_ ) );
NAND4_X2 _09419_ ( .A1(_01828_ ), .A2(_01833_ ), .A3(_01838_ ), .A4(_01839_ ), .ZN(_01840_ ) );
NOR4_X1 _09420_ ( .A1(_01795_ ), .A2(_01814_ ), .A3(_01827_ ), .A4(_01840_ ), .ZN(_01841_ ) );
MUX2_X1 _09421_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(fanout_net_41 ), .Z(_01842_ ) );
MUX2_X1 _09422_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(fanout_net_41 ), .Z(_01843_ ) );
MUX2_X2 _09423_ ( .A(_01842_ ), .B(_01843_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01844_ ) );
INV_X2 _09424_ ( .A(_01844_ ), .ZN(_01845_ ) );
AOI22_X1 _09425_ ( .A1(_01845_ ), .A2(\IF_ID_pc [14] ), .B1(_01785_ ), .B2(_01788_ ), .ZN(_01846_ ) );
INV_X1 _09426_ ( .A(\IF_ID_pc [31] ), .ZN(_01847_ ) );
MUX2_X1 _09427_ ( .A(\myifu.myicache.tag[0][26] ), .B(\myifu.myicache.tag[1][26] ), .S(fanout_net_41 ), .Z(_01848_ ) );
MUX2_X1 _09428_ ( .A(\myifu.myicache.tag[2][26] ), .B(\myifu.myicache.tag[3][26] ), .S(fanout_net_41 ), .Z(_01849_ ) );
MUX2_X2 _09429_ ( .A(_01848_ ), .B(_01849_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01850_ ) );
OR2_X4 _09430_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[1][0] ), .ZN(_01851_ ) );
OAI211_X1 _09431_ ( .A(_01851_ ), .B(_01778_ ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[0][0] ), .ZN(_01852_ ) );
OR2_X4 _09432_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[3][0] ), .ZN(_01853_ ) );
OAI211_X1 _09433_ ( .A(_01853_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myifu.myicache.tag[2][0] ), .ZN(_01854_ ) );
NAND2_X1 _09434_ ( .A1(_01852_ ), .A2(_01854_ ), .ZN(_01855_ ) );
OAI221_X1 _09435_ ( .A(_01846_ ), .B1(_01847_ ), .B2(_01850_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .C2(_01855_ ), .ZN(_01856_ ) );
AOI21_X2 _09436_ ( .A(\IF_ID_pc [18] ), .B1(_01835_ ), .B2(_01837_ ), .ZN(_01857_ ) );
AOI21_X1 _09437_ ( .A(_01857_ ), .B1(_01847_ ), .B2(_01850_ ), .ZN(_01858_ ) );
INV_X1 _09438_ ( .A(\IF_ID_pc [16] ), .ZN(_01859_ ) );
MUX2_X1 _09439_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_41 ), .Z(_01860_ ) );
MUX2_X1 _09440_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01861_ ) );
MUX2_X2 _09441_ ( .A(_01860_ ), .B(_01861_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01862_ ) );
INV_X1 _09442_ ( .A(\IF_ID_pc [10] ), .ZN(_01863_ ) );
OR2_X2 _09443_ ( .A1(_01819_ ), .A2(\myifu.myicache.tag[1][5] ), .ZN(_01864_ ) );
OAI211_X1 _09444_ ( .A(_01864_ ), .B(_01779_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][5] ), .ZN(_01865_ ) );
OR2_X4 _09445_ ( .A1(_01819_ ), .A2(\myifu.myicache.tag[3][5] ), .ZN(_01866_ ) );
OAI211_X1 _09446_ ( .A(_01866_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][5] ), .ZN(_01867_ ) );
NAND2_X1 _09447_ ( .A1(_01865_ ), .A2(_01867_ ), .ZN(_01868_ ) );
OAI221_X1 _09448_ ( .A(_01858_ ), .B1(_01859_ ), .B2(_01862_ ), .C1(_01863_ ), .C2(_01868_ ), .ZN(_01869_ ) );
INV_X1 _09449_ ( .A(\IF_ID_pc [9] ), .ZN(_01870_ ) );
OR2_X4 _09450_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[1][4] ), .ZN(_01871_ ) );
OAI211_X2 _09451_ ( .A(_01871_ ), .B(_01779_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][4] ), .ZN(_01872_ ) );
OR2_X4 _09452_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[3][4] ), .ZN(_01873_ ) );
OAI211_X4 _09453_ ( .A(_01873_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][4] ), .ZN(_01874_ ) );
NAND2_X2 _09454_ ( .A1(_01872_ ), .A2(_01874_ ), .ZN(_01875_ ) );
AOI22_X1 _09455_ ( .A1(_01870_ ), .A2(_01875_ ), .B1(_01855_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01876_ ) );
NAND3_X1 _09456_ ( .A1(_01791_ ), .A2(_01793_ ), .A3(_01789_ ), .ZN(_01877_ ) );
OAI211_X1 _09457_ ( .A(_01876_ ), .B(_01877_ ), .C1(_01870_ ), .C2(_01875_ ), .ZN(_01878_ ) );
NAND2_X1 _09458_ ( .A1(_01862_ ), .A2(_01859_ ), .ZN(_01879_ ) );
NAND2_X1 _09459_ ( .A1(_01868_ ), .A2(_01863_ ), .ZN(_01880_ ) );
OAI211_X1 _09460_ ( .A(_01879_ ), .B(_01880_ ), .C1(_01801_ ), .C2(_01804_ ), .ZN(_01881_ ) );
NOR4_X1 _09461_ ( .A1(_01856_ ), .A2(_01869_ ), .A3(_01878_ ), .A4(_01881_ ), .ZN(_01882_ ) );
AND2_X1 _09462_ ( .A1(_01841_ ), .A2(_01882_ ), .ZN(_01883_ ) );
MUX2_X1 _09463_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01884_ ) );
MUX2_X1 _09464_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01885_ ) );
MUX2_X1 _09465_ ( .A(_01884_ ), .B(_01885_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01886_ ) );
MUX2_X1 _09466_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01887_ ) );
MUX2_X1 _09467_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01888_ ) );
MUX2_X2 _09468_ ( .A(_01887_ ), .B(_01888_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01889_ ) );
INV_X1 _09469_ ( .A(\IF_ID_pc [20] ), .ZN(_01890_ ) );
OR2_X1 _09470_ ( .A1(_01889_ ), .A2(_01890_ ), .ZN(_01891_ ) );
MUX2_X1 _09471_ ( .A(\myifu.myicache.tag[2][21] ), .B(\myifu.myicache.tag[3][21] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01892_ ) );
NOR2_X1 _09472_ ( .A1(_01892_ ), .A2(_01779_ ), .ZN(_01893_ ) );
MUX2_X1 _09473_ ( .A(\myifu.myicache.tag[0][21] ), .B(\myifu.myicache.tag[1][21] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01894_ ) );
NOR2_X1 _09474_ ( .A1(_01894_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01895_ ) );
OAI21_X1 _09475_ ( .A(\IF_ID_pc [26] ), .B1(_01893_ ), .B2(_01895_ ), .ZN(_01896_ ) );
NAND2_X1 _09476_ ( .A1(_01813_ ), .A2(_01810_ ), .ZN(_01897_ ) );
AND4_X2 _09477_ ( .A1(_01886_ ), .A2(_01891_ ), .A3(_01896_ ), .A4(_01897_ ), .ZN(_01898_ ) );
OR2_X1 _09478_ ( .A1(_01819_ ), .A2(\myifu.myicache.tag[1][19] ), .ZN(_01899_ ) );
OAI211_X1 _09479_ ( .A(_01899_ ), .B(_01779_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][19] ), .ZN(_01900_ ) );
OR2_X1 _09480_ ( .A1(_01819_ ), .A2(\myifu.myicache.tag[3][19] ), .ZN(_01901_ ) );
OAI211_X1 _09481_ ( .A(_01901_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][19] ), .ZN(_01902_ ) );
INV_X1 _09482_ ( .A(\IF_ID_pc [24] ), .ZN(_01903_ ) );
AND3_X1 _09483_ ( .A1(_01900_ ), .A2(_01902_ ), .A3(_01903_ ), .ZN(_01904_ ) );
AOI21_X1 _09484_ ( .A(_01903_ ), .B1(_01900_ ), .B2(_01902_ ), .ZN(_01905_ ) );
OR2_X1 _09485_ ( .A1(_01819_ ), .A2(\myifu.myicache.tag[3][1] ), .ZN(_01906_ ) );
OAI211_X1 _09486_ ( .A(_01906_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][1] ), .ZN(_01907_ ) );
INV_X1 _09487_ ( .A(\IF_ID_pc [6] ), .ZN(_01908_ ) );
OR2_X1 _09488_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_01909_ ) );
OAI211_X1 _09489_ ( .A(_01909_ ), .B(_01779_ ), .C1(_01819_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_01910_ ) );
AND3_X1 _09490_ ( .A1(_01907_ ), .A2(_01908_ ), .A3(_01910_ ), .ZN(_01911_ ) );
AOI21_X1 _09491_ ( .A(_01908_ ), .B1(_01907_ ), .B2(_01910_ ), .ZN(_01912_ ) );
OAI221_X2 _09492_ ( .A(_01898_ ), .B1(_01904_ ), .B2(_01905_ ), .C1(_01911_ ), .C2(_01912_ ), .ZN(_01913_ ) );
OR2_X4 _09493_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_01914_ ) );
OAI211_X1 _09494_ ( .A(_01914_ ), .B(_01779_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_01915_ ) );
OR2_X1 _09495_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][25] ), .ZN(_01916_ ) );
OAI211_X1 _09496_ ( .A(_01916_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01819_ ), .C2(\myifu.myicache.tag[3][25] ), .ZN(_01917_ ) );
AND3_X1 _09497_ ( .A1(_01915_ ), .A2(_01917_ ), .A3(\IF_ID_pc [30] ), .ZN(_01918_ ) );
OR2_X4 _09498_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_01919_ ) );
OAI211_X2 _09499_ ( .A(_01919_ ), .B(_01778_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_01920_ ) );
OR2_X4 _09500_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[3][6] ), .ZN(_01921_ ) );
OAI211_X2 _09501_ ( .A(_01921_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][6] ), .ZN(_01922_ ) );
INV_X1 _09502_ ( .A(\IF_ID_pc [11] ), .ZN(_01923_ ) );
AND3_X1 _09503_ ( .A1(_01920_ ), .A2(_01922_ ), .A3(_01923_ ), .ZN(_01924_ ) );
AOI21_X1 _09504_ ( .A(_01923_ ), .B1(_01920_ ), .B2(_01922_ ), .ZN(_01925_ ) );
OR2_X4 _09505_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[3][23] ), .ZN(_01926_ ) );
OAI211_X2 _09506_ ( .A(_01926_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][23] ), .ZN(_01927_ ) );
INV_X1 _09507_ ( .A(\IF_ID_pc [28] ), .ZN(_01928_ ) );
OR2_X4 _09508_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][23] ), .ZN(_01929_ ) );
OAI211_X2 _09509_ ( .A(_01929_ ), .B(_01778_ ), .C1(_01776_ ), .C2(\myifu.myicache.tag[1][23] ), .ZN(_01930_ ) );
AND3_X1 _09510_ ( .A1(_01927_ ), .A2(_01928_ ), .A3(_01930_ ), .ZN(_01931_ ) );
AOI21_X1 _09511_ ( .A(_01928_ ), .B1(_01927_ ), .B2(_01930_ ), .ZN(_01932_ ) );
OAI22_X1 _09512_ ( .A1(_01924_ ), .A2(_01925_ ), .B1(_01931_ ), .B2(_01932_ ), .ZN(_01933_ ) );
OR2_X4 _09513_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[1][14] ), .ZN(_01934_ ) );
OAI211_X2 _09514_ ( .A(_01934_ ), .B(_01778_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][14] ), .ZN(_01935_ ) );
OR2_X4 _09515_ ( .A1(_01775_ ), .A2(\myifu.myicache.tag[3][14] ), .ZN(_01936_ ) );
OAI211_X2 _09516_ ( .A(_01936_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][14] ), .ZN(_01937_ ) );
NAND2_X1 _09517_ ( .A1(_01935_ ), .A2(_01937_ ), .ZN(_01938_ ) );
INV_X1 _09518_ ( .A(\IF_ID_pc [19] ), .ZN(_01939_ ) );
XNOR2_X1 _09519_ ( .A(_01938_ ), .B(_01939_ ), .ZN(_01940_ ) );
AOI21_X1 _09520_ ( .A(\IF_ID_pc [30] ), .B1(_01915_ ), .B2(_01917_ ), .ZN(_01941_ ) );
OR4_X4 _09521_ ( .A1(_01918_ ), .A2(_01933_ ), .A3(_01940_ ), .A4(_01941_ ), .ZN(_01942_ ) );
OR2_X4 _09522_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[1][17] ), .ZN(_01943_ ) );
OAI211_X1 _09523_ ( .A(_01943_ ), .B(_01779_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][17] ), .ZN(_01944_ ) );
OR2_X4 _09524_ ( .A1(_01776_ ), .A2(\myifu.myicache.tag[3][17] ), .ZN(_01945_ ) );
OAI211_X2 _09525_ ( .A(_01945_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][17] ), .ZN(_01946_ ) );
NAND2_X1 _09526_ ( .A1(_01944_ ), .A2(_01946_ ), .ZN(_01947_ ) );
XNOR2_X1 _09527_ ( .A(_01947_ ), .B(\IF_ID_pc [22] ), .ZN(_01948_ ) );
INV_X1 _09528_ ( .A(\IF_ID_pc [13] ), .ZN(_01949_ ) );
MUX2_X1 _09529_ ( .A(\myifu.myicache.tag[2][8] ), .B(\myifu.myicache.tag[3][8] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01950_ ) );
OR2_X2 _09530_ ( .A1(_01950_ ), .A2(_01778_ ), .ZN(_01951_ ) );
MUX2_X2 _09531_ ( .A(\myifu.myicache.tag[0][8] ), .B(\myifu.myicache.tag[1][8] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01952_ ) );
OAI21_X2 _09532_ ( .A(_01951_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01952_ ), .ZN(_01953_ ) );
INV_X1 _09533_ ( .A(_01953_ ), .ZN(_01954_ ) );
OAI221_X4 _09534_ ( .A(_01948_ ), .B1(\IF_ID_pc [14] ), .B2(_01845_ ), .C1(_01949_ ), .C2(_01954_ ), .ZN(_01955_ ) );
NOR3_X1 _09535_ ( .A1(_01893_ ), .A2(_01895_ ), .A3(\IF_ID_pc [26] ), .ZN(_01956_ ) );
AOI21_X1 _09536_ ( .A(_01956_ ), .B1(_01954_ ), .B2(_01949_ ), .ZN(_01957_ ) );
NAND2_X1 _09537_ ( .A1(_01889_ ), .A2(_01890_ ), .ZN(_01958_ ) );
OAI211_X1 _09538_ ( .A(_01957_ ), .B(_01958_ ), .C1(_01832_ ), .C2(_01831_ ), .ZN(_01959_ ) );
NOR4_X4 _09539_ ( .A1(_01913_ ), .A2(_01942_ ), .A3(_01955_ ), .A4(_01959_ ), .ZN(_01960_ ) );
NAND2_X2 _09540_ ( .A1(_01883_ ), .A2(_01960_ ), .ZN(_01961_ ) );
AND2_X4 _09541_ ( .A1(_01961_ ), .A2(\myifu.state [0] ), .ZN(_01962_ ) );
INV_X2 _09542_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01963_ ) );
NOR2_X4 _09543_ ( .A1(_01962_ ), .A2(_01963_ ), .ZN(_01964_ ) );
NOR2_X1 _09544_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01965_ ) );
NOR2_X4 _09545_ ( .A1(_01964_ ), .A2(_01965_ ), .ZN(_01966_ ) );
INV_X1 _09546_ ( .A(\EX_LS_flag [2] ), .ZN(_01967_ ) );
NAND4_X1 _09547_ ( .A1(_01967_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(EXU_valid_LSU ), .ZN(_01968_ ) );
NOR2_X1 _09548_ ( .A1(_01968_ ), .A2(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01969_ ) );
INV_X1 _09549_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01970_ ) );
NOR2_X1 _09550_ ( .A1(_01969_ ), .A2(_01970_ ), .ZN(_01971_ ) );
NOR2_X4 _09551_ ( .A1(_01966_ ), .A2(_01971_ ), .ZN(_01972_ ) );
BUF_X4 _09552_ ( .A(_01972_ ), .Z(_01973_ ) );
CLKBUF_X2 _09553_ ( .A(_01968_ ), .Z(_01974_ ) );
CLKBUF_X2 _09554_ ( .A(_01974_ ), .Z(_01975_ ) );
OR3_X1 _09555_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01976_ ) );
BUF_X4 _09556_ ( .A(_01969_ ), .Z(_01977_ ) );
BUF_X4 _09557_ ( .A(_01977_ ), .Z(_01978_ ) );
OAI211_X1 _09558_ ( .A(_01973_ ), .B(_01976_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01978_ ), .ZN(_01979_ ) );
INV_X1 _09559_ ( .A(\IF_ID_pc [22] ), .ZN(_01980_ ) );
INV_X8 _09560_ ( .A(_01966_ ), .ZN(_01981_ ) );
BUF_X8 _09561_ ( .A(_01981_ ), .Z(_01982_ ) );
OAI21_X1 _09562_ ( .A(_01979_ ), .B1(_01980_ ), .B2(_01982_ ), .ZN(\io_master_araddr [22] ) );
OR3_X1 _09563_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01983_ ) );
OAI211_X1 _09564_ ( .A(_01973_ ), .B(_01983_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01978_ ), .ZN(_01984_ ) );
OAI21_X1 _09565_ ( .A(_01984_ ), .B1(_01824_ ), .B2(_01982_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09566_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01985_ ) );
OAI211_X1 _09567_ ( .A(_01973_ ), .B(_01985_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01977_ ), .ZN(_01986_ ) );
OAI21_X1 _09568_ ( .A(_01986_ ), .B1(_01785_ ), .B2(_01982_ ), .ZN(\io_master_araddr [23] ) );
OR3_X1 _09569_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01987_ ) );
OAI211_X1 _09570_ ( .A(_01973_ ), .B(_01987_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01978_ ), .ZN(_01988_ ) );
OAI21_X1 _09571_ ( .A(_01988_ ), .B1(_01939_ ), .B2(_01982_ ), .ZN(\io_master_araddr [19] ) );
OR4_X1 _09572_ ( .A1(\io_master_araddr [22] ), .A2(\io_master_araddr [17] ), .A3(\io_master_araddr [23] ), .A4(\io_master_araddr [19] ), .ZN(_01989_ ) );
OR3_X1 _09573_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01990_ ) );
OAI211_X1 _09574_ ( .A(_01973_ ), .B(_01990_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01977_ ), .ZN(_01991_ ) );
OAI21_X1 _09575_ ( .A(_01991_ ), .B1(_01859_ ), .B2(_01981_ ), .ZN(\io_master_araddr [16] ) );
OR3_X1 _09576_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01992_ ) );
OAI211_X1 _09577_ ( .A(_01972_ ), .B(_01992_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01969_ ), .ZN(_01993_ ) );
OAI21_X1 _09578_ ( .A(_01993_ ), .B1(_01801_ ), .B2(_01981_ ), .ZN(\io_master_araddr [29] ) );
OR3_X1 _09579_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01994_ ) );
OAI211_X1 _09580_ ( .A(_01972_ ), .B(_01994_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01977_ ), .ZN(_01995_ ) );
OAI221_X1 _09581_ ( .A(\IF_ID_pc [26] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01962_ ), .C2(_01963_ ), .ZN(_01996_ ) );
AND2_X1 _09582_ ( .A1(_01995_ ), .A2(_01996_ ), .ZN(_01997_ ) );
INV_X1 _09583_ ( .A(EXU_valid_LSU ), .ZN(_01998_ ) );
NOR2_X1 _09584_ ( .A1(_01998_ ), .A2(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01999_ ) );
INV_X1 _09585_ ( .A(\EX_LS_dest_csreg_mem [25] ), .ZN(_02000_ ) );
AND2_X4 _09586_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02001_ ) );
NAND4_X1 _09587_ ( .A1(_01999_ ), .A2(_02000_ ), .A3(_02001_ ), .A4(_01967_ ), .ZN(_02002_ ) );
OAI211_X2 _09588_ ( .A(_01972_ ), .B(_02002_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_01977_ ), .ZN(_02003_ ) );
INV_X1 _09589_ ( .A(\IF_ID_pc [25] ), .ZN(_02004_ ) );
OAI21_X2 _09590_ ( .A(_02003_ ), .B1(_02004_ ), .B2(_01981_ ), .ZN(\io_master_araddr [25] ) );
NAND2_X1 _09591_ ( .A1(_01997_ ), .A2(\io_master_araddr [25] ), .ZN(_02005_ ) );
OR4_X2 _09592_ ( .A1(_01989_ ), .A2(\io_master_araddr [16] ), .A3(\io_master_araddr [29] ), .A4(_02005_ ), .ZN(_02006_ ) );
OR3_X1 _09593_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02007_ ) );
OAI211_X1 _09594_ ( .A(_01972_ ), .B(_02007_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01977_ ), .ZN(_02008_ ) );
OAI221_X1 _09595_ ( .A(\IF_ID_pc [27] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01962_ ), .C2(_01963_ ), .ZN(_02009_ ) );
AND2_X1 _09596_ ( .A1(_02008_ ), .A2(_02009_ ), .ZN(_02010_ ) );
INV_X1 _09597_ ( .A(_02010_ ), .ZN(\io_master_araddr [27] ) );
OR3_X1 _09598_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02011_ ) );
OAI211_X1 _09599_ ( .A(_01972_ ), .B(_02011_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01969_ ), .ZN(_02012_ ) );
INV_X1 _09600_ ( .A(\IF_ID_pc [30] ), .ZN(_02013_ ) );
OAI21_X1 _09601_ ( .A(_02012_ ), .B1(_02013_ ), .B2(_01981_ ), .ZN(\io_master_araddr [30] ) );
OR3_X1 _09602_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02014_ ) );
OAI211_X1 _09603_ ( .A(_01973_ ), .B(_02014_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01977_ ), .ZN(_02015_ ) );
OAI21_X1 _09604_ ( .A(_02015_ ), .B1(_01890_ ), .B2(_01981_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09605_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02016_ ) );
OAI211_X1 _09606_ ( .A(_01973_ ), .B(_02016_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01977_ ), .ZN(_02017_ ) );
INV_X1 _09607_ ( .A(\IF_ID_pc [18] ), .ZN(_02018_ ) );
OAI21_X1 _09608_ ( .A(_02017_ ), .B1(_02018_ ), .B2(_01981_ ), .ZN(\io_master_araddr [18] ) );
NOR4_X1 _09609_ ( .A1(\io_master_araddr [27] ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [20] ), .A4(\io_master_araddr [18] ), .ZN(_02019_ ) );
OR3_X1 _09610_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02020_ ) );
OAI211_X1 _09611_ ( .A(_01973_ ), .B(_02020_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01977_ ), .ZN(_02021_ ) );
OAI21_X1 _09612_ ( .A(_02021_ ), .B1(_01806_ ), .B2(_01981_ ), .ZN(\io_master_araddr [21] ) );
OR3_X1 _09613_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02022_ ) );
OAI211_X1 _09614_ ( .A(_01972_ ), .B(_02022_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01969_ ), .ZN(_02023_ ) );
OAI21_X1 _09615_ ( .A(_02023_ ), .B1(_01928_ ), .B2(_01981_ ), .ZN(\io_master_araddr [28] ) );
INV_X1 _09616_ ( .A(\EX_LS_dest_csreg_mem [24] ), .ZN(_02024_ ) );
BUF_X4 _09617_ ( .A(_01967_ ), .Z(_02025_ ) );
NAND4_X1 _09618_ ( .A1(_01999_ ), .A2(_02024_ ), .A3(_02001_ ), .A4(_02025_ ), .ZN(_02026_ ) );
OAI211_X1 _09619_ ( .A(_01973_ ), .B(_02026_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01977_ ), .ZN(_02027_ ) );
OAI21_X1 _09620_ ( .A(_02027_ ), .B1(_01903_ ), .B2(_01982_ ), .ZN(\io_master_araddr [24] ) );
OR3_X1 _09621_ ( .A1(_01974_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02028_ ) );
OAI211_X1 _09622_ ( .A(_01972_ ), .B(_02028_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01969_ ), .ZN(_02029_ ) );
OAI21_X1 _09623_ ( .A(_02029_ ), .B1(_01847_ ), .B2(_01981_ ), .ZN(\io_master_araddr [31] ) );
NOR4_X1 _09624_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [28] ), .A3(\io_master_araddr [24] ), .A4(\io_master_araddr [31] ), .ZN(_02030_ ) );
NAND2_X1 _09625_ ( .A1(_02019_ ), .A2(_02030_ ), .ZN(_02031_ ) );
CLKBUF_X2 _09626_ ( .A(_01966_ ), .Z(_02032_ ) );
CLKBUF_X2 _09627_ ( .A(_02032_ ), .Z(_02033_ ) );
CLKBUF_X2 _09628_ ( .A(_02033_ ), .Z(_02034_ ) );
CLKBUF_X2 _09629_ ( .A(_02034_ ), .Z(_02035_ ) );
NAND2_X1 _09630_ ( .A1(_02024_ ), .A2(_02000_ ), .ZN(_02036_ ) );
NOR3_X1 _09631_ ( .A1(_02036_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\EX_LS_dest_csreg_mem [26] ), .ZN(_02037_ ) );
INV_X1 _09632_ ( .A(_02037_ ), .ZN(_02038_ ) );
OR4_X1 _09633_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(_02038_ ), .A3(\EX_LS_dest_csreg_mem [30] ), .A4(\EX_LS_dest_csreg_mem [29] ), .ZN(_02039_ ) );
NOR2_X1 _09634_ ( .A1(_02039_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .ZN(_02040_ ) );
AND2_X2 _09635_ ( .A1(_02001_ ), .A2(_01967_ ), .ZN(_02041_ ) );
AND2_X1 _09636_ ( .A1(_02040_ ), .A2(_02041_ ), .ZN(_02042_ ) );
INV_X1 _09637_ ( .A(_02042_ ), .ZN(_02043_ ) );
NOR2_X1 _09638_ ( .A1(fanout_net_3 ), .A2(\EX_LS_dest_csreg_mem [1] ), .ZN(_02044_ ) );
INV_X1 _09639_ ( .A(_02044_ ), .ZN(_02045_ ) );
INV_X1 _09640_ ( .A(\EX_LS_typ [0] ), .ZN(_02046_ ) );
NOR2_X1 _09641_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .ZN(_02047_ ) );
NAND4_X1 _09642_ ( .A1(_02045_ ), .A2(\EX_LS_typ [2] ), .A3(_02046_ ), .A4(_02047_ ), .ZN(_02048_ ) );
NOR2_X1 _09643_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02049_ ) );
INV_X1 _09644_ ( .A(_02049_ ), .ZN(_02050_ ) );
AND2_X1 _09645_ ( .A1(fanout_net_3 ), .A2(\EX_LS_typ [1] ), .ZN(_02051_ ) );
INV_X1 _09646_ ( .A(_02051_ ), .ZN(_02052_ ) );
OAI21_X1 _09647_ ( .A(_02048_ ), .B1(_02050_ ), .B2(_02052_ ), .ZN(_02053_ ) );
INV_X1 _09648_ ( .A(\EX_LS_typ [4] ), .ZN(_02054_ ) );
AND2_X1 _09649_ ( .A1(_02041_ ), .A2(_02054_ ), .ZN(_02055_ ) );
NAND2_X1 _09650_ ( .A1(_02053_ ), .A2(_02055_ ), .ZN(_02056_ ) );
AND2_X1 _09651_ ( .A1(_02043_ ), .A2(_02056_ ), .ZN(_02057_ ) );
INV_X32 _09652_ ( .A(\EX_LS_flag [1] ), .ZN(_02058_ ) );
NOR2_X4 _09653_ ( .A1(_02058_ ), .A2(\EX_LS_flag [0] ), .ZN(_02059_ ) );
AND2_X1 _09654_ ( .A1(_02059_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02060_ ) );
AND2_X1 _09655_ ( .A1(_02040_ ), .A2(_02060_ ), .ZN(_02061_ ) );
NAND3_X1 _09656_ ( .A1(_02025_ ), .A2(_02054_ ), .A3(\EX_LS_typ [0] ), .ZN(_02062_ ) );
NOR3_X1 _09657_ ( .A1(_02062_ ), .A2(_02058_ ), .A3(\EX_LS_flag [0] ), .ZN(_02063_ ) );
INV_X1 _09658_ ( .A(_02063_ ), .ZN(_02064_ ) );
AND3_X1 _09659_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02065_ ) );
AOI22_X1 _09660_ ( .A1(_02045_ ), .A2(_02065_ ), .B1(_02051_ ), .B2(_02049_ ), .ZN(_02066_ ) );
NOR2_X1 _09661_ ( .A1(_02064_ ), .A2(_02066_ ), .ZN(_02067_ ) );
NOR2_X1 _09662_ ( .A1(_02061_ ), .A2(_02067_ ), .ZN(_02068_ ) );
AND2_X1 _09663_ ( .A1(_02057_ ), .A2(_02068_ ), .ZN(_02069_ ) );
AOI21_X1 _09664_ ( .A(_02035_ ), .B1(_01978_ ), .B2(_02069_ ), .ZN(_02070_ ) );
NOR2_X1 _09665_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02071_ ) );
AOI211_X1 _09666_ ( .A(_01965_ ), .B(_01964_ ), .C1(\myifu.state [0] ), .C2(_02071_ ), .ZN(_02072_ ) );
NOR4_X1 _09667_ ( .A1(_02006_ ), .A2(_02031_ ), .A3(_02070_ ), .A4(_02072_ ), .ZN(_02073_ ) );
OAI21_X1 _09668_ ( .A(_01602_ ), .B1(_02073_ ), .B2(\myclint.rvalid ), .ZN(_02074_ ) );
OR4_X4 _09669_ ( .A1(\io_master_araddr [29] ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [28] ), .A4(\io_master_araddr [31] ), .ZN(_02075_ ) );
INV_X1 _09670_ ( .A(_01997_ ), .ZN(\io_master_araddr [26] ) );
NAND2_X2 _09671_ ( .A1(_02010_ ), .A2(\io_master_araddr [25] ), .ZN(_02076_ ) );
NOR4_X4 _09672_ ( .A1(_02075_ ), .A2(\io_master_araddr [26] ), .A3(\io_master_araddr [24] ), .A4(_02076_ ), .ZN(_02077_ ) );
NOR4_X1 _09673_ ( .A1(\io_master_araddr [22] ), .A2(\io_master_araddr [19] ), .A3(\io_master_araddr [16] ), .A4(\io_master_araddr [21] ), .ZN(_02078_ ) );
NOR4_X1 _09674_ ( .A1(\io_master_araddr [17] ), .A2(\io_master_araddr [23] ), .A3(\io_master_araddr [20] ), .A4(\io_master_araddr [18] ), .ZN(_02079_ ) );
AND2_X4 _09675_ ( .A1(_02078_ ), .A2(_02079_ ), .ZN(_02080_ ) );
NAND3_X1 _09676_ ( .A1(_02077_ ), .A2(\myclint.rvalid ), .A3(_02080_ ), .ZN(_02081_ ) );
AOI211_X1 _09677_ ( .A(_01970_ ), .B(_02035_ ), .C1(_01978_ ), .C2(_02069_ ), .ZN(_02082_ ) );
AND3_X1 _09678_ ( .A1(_01961_ ), .A2(\myifu.state [0] ), .A3(_02071_ ), .ZN(_02083_ ) );
NOR4_X1 _09679_ ( .A1(_01964_ ), .A2(_01963_ ), .A3(_01965_ ), .A4(_02083_ ), .ZN(_02084_ ) );
NOR3_X1 _09680_ ( .A1(_02081_ ), .A2(_02082_ ), .A3(_02084_ ), .ZN(_02085_ ) );
NOR2_X1 _09681_ ( .A1(_02074_ ), .A2(_02085_ ), .ZN(_00064_ ) );
INV_X1 _09682_ ( .A(\LS_WB_wdata_csreg [5] ), .ZN(_02086_ ) );
NOR2_X1 _09683_ ( .A1(_02086_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00065_ ) );
INV_X1 _09684_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02087_ ) );
CLKBUF_X2 _09685_ ( .A(_02087_ ), .Z(_02088_ ) );
AND2_X1 _09686_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [4] ), .ZN(_00066_ ) );
AND2_X1 _09687_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00067_ ) );
AND2_X1 _09688_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00068_ ) );
AND2_X1 _09689_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00069_ ) );
INV_X1 _09690_ ( .A(\LS_WB_wdata_csreg [20] ), .ZN(_02089_ ) );
NOR2_X1 _09691_ ( .A1(_02089_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00070_ ) );
AND2_X1 _09692_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [19] ), .ZN(_00071_ ) );
INV_X1 _09693_ ( .A(\LS_WB_wdata_csreg [18] ), .ZN(_02090_ ) );
NOR2_X1 _09694_ ( .A1(_02090_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00072_ ) );
AND2_X1 _09695_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [17] ), .ZN(_00073_ ) );
AND2_X1 _09696_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00074_ ) );
AND2_X1 _09697_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00075_ ) );
AND2_X1 _09698_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00076_ ) );
AND2_X1 _09699_ ( .A1(_02088_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00077_ ) );
CLKBUF_X2 _09700_ ( .A(_02087_ ), .Z(_02091_ ) );
AND2_X1 _09701_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00078_ ) );
AND2_X1 _09702_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00079_ ) );
AND2_X1 _09703_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00080_ ) );
AND2_X1 _09704_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00081_ ) );
AND2_X1 _09705_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00082_ ) );
AND2_X1 _09706_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00083_ ) );
AND2_X1 _09707_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00084_ ) );
AND2_X1 _09708_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [6] ), .ZN(_00085_ ) );
AND2_X1 _09709_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00086_ ) );
AND2_X1 _09710_ ( .A1(_02091_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00087_ ) );
AND2_X1 _09711_ ( .A1(_02087_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00088_ ) );
AND2_X1 _09712_ ( .A1(_02087_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00089_ ) );
AND2_X1 _09713_ ( .A1(_02087_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00090_ ) );
AND2_X1 _09714_ ( .A1(_02087_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00091_ ) );
AND2_X1 _09715_ ( .A1(_02087_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00092_ ) );
CLKBUF_X2 _09716_ ( .A(_01559_ ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ) );
INV_X1 _09717_ ( .A(_02057_ ), .ZN(_02092_ ) );
INV_X1 _09718_ ( .A(_02068_ ), .ZN(_02093_ ) );
NOR2_X1 _09719_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02094_ ) );
NAND2_X1 _09720_ ( .A1(_02094_ ), .A2(_01559_ ), .ZN(_02095_ ) );
OR2_X1 _09721_ ( .A1(\myexu.pc_jump [26] ), .A2(\myexu.pc_jump [25] ), .ZN(_02096_ ) );
OR3_X1 _09722_ ( .A1(_02096_ ), .A2(\myexu.pc_jump [27] ), .A3(\myexu.pc_jump [24] ), .ZN(_02097_ ) );
OR4_X1 _09723_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02098_ ) );
NOR2_X1 _09724_ ( .A1(_02097_ ), .A2(_02098_ ), .ZN(_02099_ ) );
NOR2_X1 _09725_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02100_ ) );
INV_X1 _09726_ ( .A(_02100_ ), .ZN(_02101_ ) );
NOR3_X1 _09727_ ( .A1(_02099_ ), .A2(exception_quest_IDU ), .A3(_02101_ ), .ZN(_02102_ ) );
NOR4_X1 _09728_ ( .A1(_02092_ ), .A2(_02093_ ), .A3(_02095_ ), .A4(_02102_ ), .ZN(_00093_ ) );
AOI21_X1 _09729_ ( .A(_02095_ ), .B1(_02069_ ), .B2(exception_quest_IDU ), .ZN(_00094_ ) );
INV_X1 _09730_ ( .A(fanout_net_27 ), .ZN(_02103_ ) );
BUF_X4 _09731_ ( .A(_02103_ ), .Z(_02104_ ) );
BUF_X4 _09732_ ( .A(_02104_ ), .Z(_02105_ ) );
INV_X2 _09733_ ( .A(fanout_net_26 ), .ZN(_02106_ ) );
BUF_X4 _09734_ ( .A(_02106_ ), .Z(_02107_ ) );
BUF_X4 _09735_ ( .A(_02107_ ), .Z(_02108_ ) );
MUX2_X1 _09736_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02109_ ) );
AND2_X1 _09737_ ( .A1(_02109_ ), .A2(fanout_net_23 ), .ZN(_02110_ ) );
INV_X1 _09738_ ( .A(fanout_net_23 ), .ZN(_02111_ ) );
BUF_X4 _09739_ ( .A(_02111_ ), .Z(_02112_ ) );
BUF_X4 _09740_ ( .A(_02112_ ), .Z(_02113_ ) );
BUF_X4 _09741_ ( .A(_02113_ ), .Z(_02114_ ) );
BUF_X4 _09742_ ( .A(_02114_ ), .Z(_02115_ ) );
MUX2_X1 _09743_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02116_ ) );
AOI211_X1 _09744_ ( .A(_02108_ ), .B(_02110_ ), .C1(_02115_ ), .C2(_02116_ ), .ZN(_02117_ ) );
BUF_X4 _09745_ ( .A(_02108_ ), .Z(_02118_ ) );
MUX2_X1 _09746_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02119_ ) );
AND2_X1 _09747_ ( .A1(_02119_ ), .A2(fanout_net_23 ), .ZN(_02120_ ) );
MUX2_X1 _09748_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02121_ ) );
AOI21_X1 _09749_ ( .A(_02120_ ), .B1(_02115_ ), .B2(_02121_ ), .ZN(_02122_ ) );
AOI211_X1 _09750_ ( .A(_02105_ ), .B(_02117_ ), .C1(_02118_ ), .C2(_02122_ ), .ZN(_02123_ ) );
AND3_X1 _09751_ ( .A1(_02058_ ), .A2(\EX_LS_flag [0] ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02124_ ) );
AND2_X1 _09752_ ( .A1(_02058_ ), .A2(\EX_LS_flag [0] ), .ZN(_02125_ ) );
AOI211_X1 _09753_ ( .A(_02124_ ), .B(_02041_ ), .C1(\EX_LS_flag [2] ), .C2(_02125_ ), .ZN(_02126_ ) );
AND2_X4 _09754_ ( .A1(_02059_ ), .A2(\EX_LS_flag [2] ), .ZN(_02127_ ) );
BUF_X4 _09755_ ( .A(_02127_ ), .Z(_02128_ ) );
INV_X8 _09756_ ( .A(_02128_ ), .ZN(_02129_ ) );
NAND2_X2 _09757_ ( .A1(_02126_ ), .A2(_02129_ ), .ZN(_02130_ ) );
XNOR2_X1 _09758_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02131_ ) );
OR3_X1 _09759_ ( .A1(\EX_LS_dest_reg [2] ), .A2(\EX_LS_dest_reg [1] ), .A3(\EX_LS_dest_reg [0] ), .ZN(_02132_ ) );
OR2_X1 _09760_ ( .A1(\EX_LS_dest_reg [4] ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02133_ ) );
NOR2_X1 _09761_ ( .A1(_02132_ ), .A2(_02133_ ), .ZN(_02134_ ) );
INV_X1 _09762_ ( .A(_02134_ ), .ZN(_02135_ ) );
INV_X8 _09763_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02136_ ) );
NAND2_X1 _09764_ ( .A1(_02136_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02137_ ) );
NAND4_X4 _09765_ ( .A1(_02130_ ), .A2(_02131_ ), .A3(_02135_ ), .A4(_02137_ ), .ZN(_02138_ ) );
BUF_X4 _09766_ ( .A(_02138_ ), .Z(_02139_ ) );
CLKBUF_X2 _09767_ ( .A(_02139_ ), .Z(_02140_ ) );
XOR2_X1 _09768_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .Z(_02141_ ) );
XOR2_X1 _09769_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .Z(_02142_ ) );
INV_X1 _09770_ ( .A(\ID_EX_rs1 [3] ), .ZN(_02143_ ) );
OAI22_X1 _09771_ ( .A1(_02143_ ), .A2(\EX_LS_dest_reg [3] ), .B1(_02136_ ), .B2(\ID_EX_rs1 [1] ), .ZN(_02144_ ) );
INV_X1 _09772_ ( .A(\EX_LS_dest_reg [3] ), .ZN(_02145_ ) );
OAI21_X1 _09773_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02145_ ), .B2(\ID_EX_rs1 [3] ), .ZN(_02146_ ) );
OR4_X2 _09774_ ( .A1(_02141_ ), .A2(_02142_ ), .A3(_02144_ ), .A4(_02146_ ), .ZN(_02147_ ) );
BUF_X2 _09775_ ( .A(_02147_ ), .Z(_02148_ ) );
BUF_X2 _09776_ ( .A(_02148_ ), .Z(_02149_ ) );
BUF_X2 _09777_ ( .A(_02149_ ), .Z(_02150_ ) );
NOR2_X1 _09778_ ( .A1(_02140_ ), .A2(_02150_ ), .ZN(_02151_ ) );
OR2_X1 _09779_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02152_ ) );
BUF_X4 _09780_ ( .A(_02111_ ), .Z(_02153_ ) );
BUF_X4 _09781_ ( .A(_02153_ ), .Z(_02154_ ) );
BUF_X4 _09782_ ( .A(_02154_ ), .Z(_02155_ ) );
INV_X1 _09783_ ( .A(fanout_net_15 ), .ZN(_02156_ ) );
BUF_X4 _09784_ ( .A(_02156_ ), .Z(_02157_ ) );
BUF_X4 _09785_ ( .A(_02157_ ), .Z(_02158_ ) );
BUF_X4 _09786_ ( .A(_02158_ ), .Z(_02159_ ) );
BUF_X4 _09787_ ( .A(_02159_ ), .Z(_02160_ ) );
OAI211_X1 _09788_ ( .A(_02152_ ), .B(_02155_ ), .C1(_02160_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02161_ ) );
OR2_X1 _09789_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02162_ ) );
BUF_X4 _09790_ ( .A(_02157_ ), .Z(_02163_ ) );
BUF_X4 _09791_ ( .A(_02163_ ), .Z(_02164_ ) );
OAI211_X1 _09792_ ( .A(_02162_ ), .B(fanout_net_23 ), .C1(_02164_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02165_ ) );
AND3_X1 _09793_ ( .A1(_02161_ ), .A2(_02165_ ), .A3(fanout_net_26 ), .ZN(_02166_ ) );
OAI21_X1 _09794_ ( .A(fanout_net_23 ), .B1(fanout_net_15 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02167_ ) );
INV_X1 _09795_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02168_ ) );
AOI21_X1 _09796_ ( .A(_02167_ ), .B1(fanout_net_15 ), .B2(_02168_ ), .ZN(_02169_ ) );
MUX2_X1 _09797_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02170_ ) );
AOI21_X1 _09798_ ( .A(_02169_ ), .B1(_02115_ ), .B2(_02170_ ), .ZN(_02171_ ) );
AOI211_X1 _09799_ ( .A(fanout_net_27 ), .B(_02166_ ), .C1(_02118_ ), .C2(_02171_ ), .ZN(_02172_ ) );
OR3_X2 _09800_ ( .A1(_02123_ ), .A2(_02151_ ), .A3(_02172_ ), .ZN(_02173_ ) );
BUF_X2 _09801_ ( .A(_02138_ ), .Z(_02174_ ) );
BUF_X2 _09802_ ( .A(_02174_ ), .Z(_02175_ ) );
BUF_X2 _09803_ ( .A(_02175_ ), .Z(_02176_ ) );
OR3_X2 _09804_ ( .A1(_02176_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02150_ ), .ZN(_02177_ ) );
AND2_X2 _09805_ ( .A1(_02173_ ), .A2(_02177_ ), .ZN(_02178_ ) );
XOR2_X1 _09806_ ( .A(_02178_ ), .B(\ID_EX_imm [30] ), .Z(_02179_ ) );
BUF_X4 _09807_ ( .A(_02147_ ), .Z(_02180_ ) );
CLKBUF_X2 _09808_ ( .A(_02180_ ), .Z(_02181_ ) );
OR3_X1 _09809_ ( .A1(_02140_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02181_ ), .ZN(_02182_ ) );
OR2_X1 _09810_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02183_ ) );
BUF_X4 _09811_ ( .A(_02112_ ), .Z(_02184_ ) );
BUF_X4 _09812_ ( .A(_02184_ ), .Z(_02185_ ) );
BUF_X4 _09813_ ( .A(_02185_ ), .Z(_02186_ ) );
BUF_X4 _09814_ ( .A(_02163_ ), .Z(_02187_ ) );
BUF_X4 _09815_ ( .A(_02187_ ), .Z(_02188_ ) );
OAI211_X1 _09816_ ( .A(_02183_ ), .B(_02186_ ), .C1(_02188_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02189_ ) );
OR2_X1 _09817_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02190_ ) );
OAI211_X1 _09818_ ( .A(_02190_ ), .B(fanout_net_23 ), .C1(_02160_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02191_ ) );
BUF_X4 _09819_ ( .A(_02106_ ), .Z(_02192_ ) );
BUF_X4 _09820_ ( .A(_02192_ ), .Z(_02193_ ) );
NAND3_X1 _09821_ ( .A1(_02189_ ), .A2(_02191_ ), .A3(_02193_ ), .ZN(_02194_ ) );
MUX2_X1 _09822_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02195_ ) );
MUX2_X1 _09823_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02196_ ) );
MUX2_X1 _09824_ ( .A(_02195_ ), .B(_02196_ ), .S(_02155_ ), .Z(_02197_ ) );
OAI211_X1 _09825_ ( .A(_02105_ ), .B(_02194_ ), .C1(_02197_ ), .C2(_02118_ ), .ZN(_02198_ ) );
OR2_X1 _09826_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02199_ ) );
OAI211_X1 _09827_ ( .A(_02199_ ), .B(_02155_ ), .C1(_02160_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02200_ ) );
NOR2_X1 _09828_ ( .A1(_02188_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02201_ ) );
OAI21_X1 _09829_ ( .A(fanout_net_23 ), .B1(fanout_net_15 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02202_ ) );
OAI211_X1 _09830_ ( .A(_02200_ ), .B(fanout_net_26 ), .C1(_02201_ ), .C2(_02202_ ), .ZN(_02203_ ) );
MUX2_X1 _09831_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02204_ ) );
MUX2_X1 _09832_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02205_ ) );
MUX2_X1 _09833_ ( .A(_02204_ ), .B(_02205_ ), .S(fanout_net_23 ), .Z(_02206_ ) );
OAI211_X1 _09834_ ( .A(fanout_net_27 ), .B(_02203_ ), .C1(_02206_ ), .C2(fanout_net_26 ), .ZN(_02207_ ) );
OAI211_X1 _09835_ ( .A(_02198_ ), .B(_02207_ ), .C1(_02176_ ), .C2(_02181_ ), .ZN(_02208_ ) );
NAND2_X1 _09836_ ( .A1(_02182_ ), .A2(_02208_ ), .ZN(_02209_ ) );
XNOR2_X1 _09837_ ( .A(_02209_ ), .B(\ID_EX_imm [28] ), .ZN(_02210_ ) );
OR3_X1 _09838_ ( .A1(_02140_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02181_ ), .ZN(_02211_ ) );
INV_X1 _09839_ ( .A(\ID_EX_imm [27] ), .ZN(_02212_ ) );
OR2_X1 _09840_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02213_ ) );
BUF_X4 _09841_ ( .A(_02164_ ), .Z(_02214_ ) );
OAI211_X1 _09842_ ( .A(_02213_ ), .B(_02115_ ), .C1(_02214_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02215_ ) );
OR2_X1 _09843_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02216_ ) );
OAI211_X1 _09844_ ( .A(_02216_ ), .B(fanout_net_23 ), .C1(_02214_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02217_ ) );
NAND3_X1 _09845_ ( .A1(_02215_ ), .A2(_02217_ ), .A3(_02193_ ), .ZN(_02218_ ) );
MUX2_X1 _09846_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02219_ ) );
MUX2_X1 _09847_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02220_ ) );
MUX2_X1 _09848_ ( .A(_02219_ ), .B(_02220_ ), .S(_02186_ ), .Z(_02221_ ) );
OAI211_X1 _09849_ ( .A(_02105_ ), .B(_02218_ ), .C1(_02221_ ), .C2(_02118_ ), .ZN(_02222_ ) );
OR2_X1 _09850_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02223_ ) );
OAI211_X1 _09851_ ( .A(_02223_ ), .B(_02186_ ), .C1(_02188_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02224_ ) );
NOR2_X1 _09852_ ( .A1(_02214_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02225_ ) );
OAI21_X1 _09853_ ( .A(fanout_net_23 ), .B1(fanout_net_15 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02226_ ) );
OAI211_X1 _09854_ ( .A(_02224_ ), .B(fanout_net_26 ), .C1(_02225_ ), .C2(_02226_ ), .ZN(_02227_ ) );
MUX2_X1 _09855_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02228_ ) );
MUX2_X1 _09856_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02229_ ) );
MUX2_X1 _09857_ ( .A(_02228_ ), .B(_02229_ ), .S(fanout_net_23 ), .Z(_02230_ ) );
OAI211_X1 _09858_ ( .A(fanout_net_27 ), .B(_02227_ ), .C1(_02230_ ), .C2(fanout_net_26 ), .ZN(_02231_ ) );
OAI211_X1 _09859_ ( .A(_02222_ ), .B(_02231_ ), .C1(_02176_ ), .C2(_02150_ ), .ZN(_02232_ ) );
AND3_X1 _09860_ ( .A1(_02211_ ), .A2(_02212_ ), .A3(_02232_ ), .ZN(_02233_ ) );
AOI21_X1 _09861_ ( .A(_02212_ ), .B1(_02211_ ), .B2(_02232_ ), .ZN(_02234_ ) );
NOR2_X1 _09862_ ( .A1(_02233_ ), .A2(_02234_ ), .ZN(_02235_ ) );
OR3_X1 _09863_ ( .A1(_02140_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02181_ ), .ZN(_02236_ ) );
OR2_X1 _09864_ ( .A1(_02187_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02237_ ) );
OAI211_X1 _09865_ ( .A(_02237_ ), .B(_02115_ ), .C1(fanout_net_15 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02238_ ) );
OR2_X1 _09866_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02239_ ) );
OAI211_X1 _09867_ ( .A(_02239_ ), .B(fanout_net_23 ), .C1(_02188_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02240_ ) );
NAND3_X1 _09868_ ( .A1(_02238_ ), .A2(fanout_net_26 ), .A3(_02240_ ), .ZN(_02241_ ) );
MUX2_X1 _09869_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02242_ ) );
MUX2_X1 _09870_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_02243_ ) );
MUX2_X1 _09871_ ( .A(_02242_ ), .B(_02243_ ), .S(_02186_ ), .Z(_02244_ ) );
OAI211_X1 _09872_ ( .A(_02105_ ), .B(_02241_ ), .C1(_02244_ ), .C2(fanout_net_26 ), .ZN(_02245_ ) );
NOR2_X1 _09873_ ( .A1(_02160_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02246_ ) );
OAI21_X1 _09874_ ( .A(fanout_net_23 ), .B1(fanout_net_16 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02247_ ) );
NOR2_X1 _09875_ ( .A1(fanout_net_16 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02248_ ) );
OAI21_X1 _09876_ ( .A(_02186_ ), .B1(_02160_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02249_ ) );
OAI221_X1 _09877_ ( .A(_02193_ ), .B1(_02246_ ), .B2(_02247_ ), .C1(_02248_ ), .C2(_02249_ ), .ZN(_02250_ ) );
MUX2_X1 _09878_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02251_ ) );
MUX2_X1 _09879_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02252_ ) );
MUX2_X1 _09880_ ( .A(_02251_ ), .B(_02252_ ), .S(fanout_net_23 ), .Z(_02253_ ) );
OAI211_X1 _09881_ ( .A(fanout_net_27 ), .B(_02250_ ), .C1(_02253_ ), .C2(_02118_ ), .ZN(_02254_ ) );
OAI211_X1 _09882_ ( .A(_02245_ ), .B(_02254_ ), .C1(_02176_ ), .C2(_02150_ ), .ZN(_02255_ ) );
NAND2_X2 _09883_ ( .A1(_02236_ ), .A2(_02255_ ), .ZN(_02256_ ) );
INV_X1 _09884_ ( .A(\ID_EX_imm [26] ), .ZN(_02257_ ) );
XNOR2_X1 _09885_ ( .A(_02256_ ), .B(_02257_ ), .ZN(_02258_ ) );
BUF_X2 _09886_ ( .A(_02147_ ), .Z(_02259_ ) );
OR3_X1 _09887_ ( .A1(_02175_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02259_ ), .ZN(_02260_ ) );
OR2_X1 _09888_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02261_ ) );
OAI211_X1 _09889_ ( .A(_02261_ ), .B(_02114_ ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02262_ ) );
OR2_X1 _09890_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02263_ ) );
OAI211_X1 _09891_ ( .A(_02263_ ), .B(fanout_net_23 ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02264_ ) );
BUF_X4 _09892_ ( .A(_02106_ ), .Z(_02265_ ) );
BUF_X4 _09893_ ( .A(_02265_ ), .Z(_02266_ ) );
NAND3_X1 _09894_ ( .A1(_02262_ ), .A2(_02264_ ), .A3(_02266_ ), .ZN(_02267_ ) );
MUX2_X1 _09895_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02268_ ) );
MUX2_X1 _09896_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02269_ ) );
MUX2_X1 _09897_ ( .A(_02268_ ), .B(_02269_ ), .S(_02185_ ), .Z(_02270_ ) );
OAI211_X1 _09898_ ( .A(_02104_ ), .B(_02267_ ), .C1(_02270_ ), .C2(_02108_ ), .ZN(_02271_ ) );
OR2_X1 _09899_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02272_ ) );
OAI211_X1 _09900_ ( .A(_02272_ ), .B(fanout_net_23 ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02273_ ) );
OR2_X1 _09901_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02274_ ) );
OAI211_X1 _09902_ ( .A(_02274_ ), .B(_02185_ ), .C1(_02159_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02275_ ) );
NAND3_X1 _09903_ ( .A1(_02273_ ), .A2(_02275_ ), .A3(fanout_net_26 ), .ZN(_02276_ ) );
MUX2_X1 _09904_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02277_ ) );
MUX2_X1 _09905_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02278_ ) );
MUX2_X1 _09906_ ( .A(_02277_ ), .B(_02278_ ), .S(fanout_net_23 ), .Z(_02279_ ) );
OAI211_X1 _09907_ ( .A(fanout_net_27 ), .B(_02276_ ), .C1(_02279_ ), .C2(fanout_net_26 ), .ZN(_02280_ ) );
OAI211_X1 _09908_ ( .A(_02271_ ), .B(_02280_ ), .C1(_02140_ ), .C2(_02181_ ), .ZN(_02281_ ) );
NAND2_X2 _09909_ ( .A1(_02260_ ), .A2(_02281_ ), .ZN(_02282_ ) );
INV_X1 _09910_ ( .A(\ID_EX_imm [23] ), .ZN(_02283_ ) );
XNOR2_X1 _09911_ ( .A(_02282_ ), .B(_02283_ ), .ZN(_02284_ ) );
OR3_X1 _09912_ ( .A1(_02175_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02149_ ), .ZN(_02285_ ) );
OR2_X1 _09913_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02286_ ) );
OAI211_X1 _09914_ ( .A(_02286_ ), .B(_02114_ ), .C1(_02164_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02287_ ) );
OR2_X1 _09915_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02288_ ) );
OAI211_X1 _09916_ ( .A(_02288_ ), .B(fanout_net_23 ), .C1(_02164_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02289_ ) );
NAND3_X1 _09917_ ( .A1(_02287_ ), .A2(_02289_ ), .A3(_02108_ ), .ZN(_02290_ ) );
MUX2_X1 _09918_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02291_ ) );
MUX2_X1 _09919_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02292_ ) );
MUX2_X1 _09920_ ( .A(_02291_ ), .B(_02292_ ), .S(_02114_ ), .Z(_02293_ ) );
OAI211_X1 _09921_ ( .A(_02104_ ), .B(_02290_ ), .C1(_02293_ ), .C2(_02193_ ), .ZN(_02294_ ) );
OR2_X1 _09922_ ( .A1(_02163_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02295_ ) );
OAI211_X1 _09923_ ( .A(_02295_ ), .B(fanout_net_23 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02296_ ) );
OR2_X1 _09924_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02297_ ) );
OAI211_X1 _09925_ ( .A(_02297_ ), .B(_02114_ ), .C1(_02164_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02298_ ) );
NAND3_X1 _09926_ ( .A1(_02296_ ), .A2(fanout_net_26 ), .A3(_02298_ ), .ZN(_02299_ ) );
MUX2_X1 _09927_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02300_ ) );
MUX2_X1 _09928_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02301_ ) );
MUX2_X1 _09929_ ( .A(_02300_ ), .B(_02301_ ), .S(fanout_net_23 ), .Z(_02302_ ) );
OAI211_X1 _09930_ ( .A(fanout_net_27 ), .B(_02299_ ), .C1(_02302_ ), .C2(fanout_net_26 ), .ZN(_02303_ ) );
OAI211_X1 _09931_ ( .A(_02294_ ), .B(_02303_ ), .C1(_02140_ ), .C2(_02181_ ), .ZN(_02304_ ) );
NAND2_X2 _09932_ ( .A1(_02285_ ), .A2(_02304_ ), .ZN(_02305_ ) );
INV_X1 _09933_ ( .A(\ID_EX_imm [22] ), .ZN(_02306_ ) );
XNOR2_X1 _09934_ ( .A(_02305_ ), .B(_02306_ ), .ZN(_02307_ ) );
AND2_X1 _09935_ ( .A1(_02284_ ), .A2(_02307_ ), .ZN(_02308_ ) );
OR3_X1 _09936_ ( .A1(_02175_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02149_ ), .ZN(_02309_ ) );
OR2_X1 _09937_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02310_ ) );
OAI211_X1 _09938_ ( .A(_02310_ ), .B(_02155_ ), .C1(_02164_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02311_ ) );
OR2_X1 _09939_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02312_ ) );
OAI211_X1 _09940_ ( .A(_02312_ ), .B(fanout_net_23 ), .C1(_02164_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02313_ ) );
NAND3_X1 _09941_ ( .A1(_02311_ ), .A2(_02313_ ), .A3(fanout_net_26 ), .ZN(_02314_ ) );
MUX2_X1 _09942_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02315_ ) );
MUX2_X1 _09943_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02316_ ) );
MUX2_X1 _09944_ ( .A(_02315_ ), .B(_02316_ ), .S(_02114_ ), .Z(_02317_ ) );
OAI211_X1 _09945_ ( .A(_02105_ ), .B(_02314_ ), .C1(_02317_ ), .C2(fanout_net_26 ), .ZN(_02318_ ) );
NOR2_X1 _09946_ ( .A1(_02164_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02319_ ) );
OAI21_X1 _09947_ ( .A(fanout_net_23 ), .B1(fanout_net_16 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02320_ ) );
NOR2_X1 _09948_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02321_ ) );
OAI21_X1 _09949_ ( .A(_02114_ ), .B1(_02164_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02322_ ) );
OAI221_X1 _09950_ ( .A(_02108_ ), .B1(_02319_ ), .B2(_02320_ ), .C1(_02321_ ), .C2(_02322_ ), .ZN(_02323_ ) );
MUX2_X1 _09951_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02324_ ) );
MUX2_X1 _09952_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02325_ ) );
MUX2_X1 _09953_ ( .A(_02324_ ), .B(_02325_ ), .S(fanout_net_23 ), .Z(_02326_ ) );
OAI211_X1 _09954_ ( .A(fanout_net_27 ), .B(_02323_ ), .C1(_02326_ ), .C2(_02193_ ), .ZN(_02327_ ) );
OAI211_X1 _09955_ ( .A(_02318_ ), .B(_02327_ ), .C1(_02140_ ), .C2(_02181_ ), .ZN(_02328_ ) );
NAND2_X2 _09956_ ( .A1(_02309_ ), .A2(_02328_ ), .ZN(_02329_ ) );
INV_X1 _09957_ ( .A(\ID_EX_imm [20] ), .ZN(_02330_ ) );
XNOR2_X1 _09958_ ( .A(_02329_ ), .B(_02330_ ), .ZN(_02331_ ) );
OR3_X1 _09959_ ( .A1(_02175_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02259_ ), .ZN(_02332_ ) );
INV_X1 _09960_ ( .A(\ID_EX_imm [21] ), .ZN(_02333_ ) );
OR2_X1 _09961_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02334_ ) );
OAI211_X1 _09962_ ( .A(_02334_ ), .B(_02114_ ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02335_ ) );
OR2_X1 _09963_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02336_ ) );
OAI211_X1 _09964_ ( .A(_02336_ ), .B(fanout_net_23 ), .C1(_02159_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02337_ ) );
NAND3_X1 _09965_ ( .A1(_02335_ ), .A2(_02337_ ), .A3(_02266_ ), .ZN(_02338_ ) );
MUX2_X1 _09966_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02339_ ) );
MUX2_X1 _09967_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02340_ ) );
MUX2_X1 _09968_ ( .A(_02339_ ), .B(_02340_ ), .S(_02185_ ), .Z(_02341_ ) );
OAI211_X1 _09969_ ( .A(fanout_net_27 ), .B(_02338_ ), .C1(_02341_ ), .C2(_02108_ ), .ZN(_02342_ ) );
OR2_X1 _09970_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02343_ ) );
OAI211_X1 _09971_ ( .A(_02343_ ), .B(_02185_ ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02344_ ) );
OR2_X1 _09972_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02345_ ) );
OAI211_X1 _09973_ ( .A(_02345_ ), .B(fanout_net_23 ), .C1(_02159_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02346_ ) );
NAND3_X1 _09974_ ( .A1(_02344_ ), .A2(_02346_ ), .A3(_02266_ ), .ZN(_02347_ ) );
MUX2_X1 _09975_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02348_ ) );
MUX2_X1 _09976_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02349_ ) );
MUX2_X1 _09977_ ( .A(_02348_ ), .B(_02349_ ), .S(_02154_ ), .Z(_02350_ ) );
OAI211_X1 _09978_ ( .A(_02104_ ), .B(_02347_ ), .C1(_02350_ ), .C2(_02108_ ), .ZN(_02351_ ) );
OAI211_X1 _09979_ ( .A(_02342_ ), .B(_02351_ ), .C1(_02175_ ), .C2(_02149_ ), .ZN(_02352_ ) );
AND3_X1 _09980_ ( .A1(_02332_ ), .A2(_02333_ ), .A3(_02352_ ), .ZN(_02353_ ) );
AOI21_X1 _09981_ ( .A(_02333_ ), .B1(_02332_ ), .B2(_02352_ ), .ZN(_02354_ ) );
NOR2_X1 _09982_ ( .A1(_02353_ ), .A2(_02354_ ), .ZN(_02355_ ) );
AND2_X1 _09983_ ( .A1(_02331_ ), .A2(_02355_ ), .ZN(_02356_ ) );
AND2_X1 _09984_ ( .A1(_02308_ ), .A2(_02356_ ), .ZN(_02357_ ) );
INV_X1 _09985_ ( .A(_02357_ ), .ZN(_02358_ ) );
OR2_X1 _09986_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02359_ ) );
BUF_X4 _09987_ ( .A(_02158_ ), .Z(_02360_ ) );
OAI211_X1 _09988_ ( .A(_02359_ ), .B(_02154_ ), .C1(_02360_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02361_ ) );
OR2_X1 _09989_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02362_ ) );
OAI211_X1 _09990_ ( .A(_02362_ ), .B(fanout_net_23 ), .C1(_02360_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02363_ ) );
NAND3_X1 _09991_ ( .A1(_02361_ ), .A2(_02363_ ), .A3(_02192_ ), .ZN(_02364_ ) );
MUX2_X1 _09992_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02365_ ) );
MUX2_X1 _09993_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02366_ ) );
BUF_X4 _09994_ ( .A(_02112_ ), .Z(_02367_ ) );
MUX2_X1 _09995_ ( .A(_02365_ ), .B(_02366_ ), .S(_02367_ ), .Z(_02368_ ) );
OAI211_X1 _09996_ ( .A(fanout_net_27 ), .B(_02364_ ), .C1(_02368_ ), .C2(_02266_ ), .ZN(_02369_ ) );
MUX2_X1 _09997_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02370_ ) );
AND2_X1 _09998_ ( .A1(_02370_ ), .A2(fanout_net_23 ), .ZN(_02371_ ) );
MUX2_X1 _09999_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02372_ ) );
AOI211_X1 _10000_ ( .A(fanout_net_26 ), .B(_02371_ ), .C1(_02155_ ), .C2(_02372_ ), .ZN(_02373_ ) );
BUF_X4 _10001_ ( .A(_02103_ ), .Z(_02374_ ) );
MUX2_X1 _10002_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02375_ ) );
MUX2_X1 _10003_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02376_ ) );
MUX2_X1 _10004_ ( .A(_02375_ ), .B(_02376_ ), .S(_02184_ ), .Z(_02377_ ) );
OAI21_X1 _10005_ ( .A(_02374_ ), .B1(_02377_ ), .B2(_02192_ ), .ZN(_02378_ ) );
BUF_X2 _10006_ ( .A(_02138_ ), .Z(_02379_ ) );
OAI221_X1 _10007_ ( .A(_02369_ ), .B1(_02373_ ), .B2(_02378_ ), .C1(_02379_ ), .C2(_02259_ ), .ZN(_02380_ ) );
OR3_X1 _10008_ ( .A1(_02139_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02180_ ), .ZN(_02381_ ) );
NAND2_X1 _10009_ ( .A1(_02380_ ), .A2(_02381_ ), .ZN(_02382_ ) );
INV_X1 _10010_ ( .A(\ID_EX_imm [19] ), .ZN(_02383_ ) );
XNOR2_X1 _10011_ ( .A(_02382_ ), .B(_02383_ ), .ZN(_02384_ ) );
OR3_X1 _10012_ ( .A1(_02175_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02149_ ), .ZN(_02385_ ) );
OR2_X1 _10013_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02386_ ) );
OAI211_X1 _10014_ ( .A(_02386_ ), .B(_02114_ ), .C1(_02164_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02387_ ) );
OR2_X1 _10015_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02388_ ) );
OAI211_X1 _10016_ ( .A(_02388_ ), .B(fanout_net_23 ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02389_ ) );
NAND3_X1 _10017_ ( .A1(_02387_ ), .A2(_02389_ ), .A3(_02266_ ), .ZN(_02390_ ) );
MUX2_X1 _10018_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02391_ ) );
MUX2_X1 _10019_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02392_ ) );
MUX2_X1 _10020_ ( .A(_02391_ ), .B(_02392_ ), .S(_02185_ ), .Z(_02393_ ) );
OAI211_X1 _10021_ ( .A(_02104_ ), .B(_02390_ ), .C1(_02393_ ), .C2(_02108_ ), .ZN(_02394_ ) );
OR2_X1 _10022_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02395_ ) );
OAI211_X1 _10023_ ( .A(_02395_ ), .B(fanout_net_23 ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02396_ ) );
OR2_X1 _10024_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02397_ ) );
OAI211_X1 _10025_ ( .A(_02397_ ), .B(_02185_ ), .C1(_02187_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02398_ ) );
NAND3_X1 _10026_ ( .A1(_02396_ ), .A2(_02398_ ), .A3(fanout_net_26 ), .ZN(_02399_ ) );
MUX2_X1 _10027_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02400_ ) );
MUX2_X1 _10028_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02401_ ) );
MUX2_X1 _10029_ ( .A(_02400_ ), .B(_02401_ ), .S(fanout_net_23 ), .Z(_02402_ ) );
OAI211_X1 _10030_ ( .A(fanout_net_27 ), .B(_02399_ ), .C1(_02402_ ), .C2(fanout_net_26 ), .ZN(_02403_ ) );
OAI211_X1 _10031_ ( .A(_02394_ ), .B(_02403_ ), .C1(_02175_ ), .C2(_02149_ ), .ZN(_02404_ ) );
NAND2_X2 _10032_ ( .A1(_02385_ ), .A2(_02404_ ), .ZN(_02405_ ) );
INV_X1 _10033_ ( .A(\ID_EX_imm [18] ), .ZN(_02406_ ) );
XNOR2_X1 _10034_ ( .A(_02405_ ), .B(_02406_ ), .ZN(_02407_ ) );
AND2_X1 _10035_ ( .A1(_02384_ ), .A2(_02407_ ), .ZN(_02408_ ) );
OR3_X1 _10036_ ( .A1(_02174_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02148_ ), .ZN(_02409_ ) );
OR2_X1 _10037_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02410_ ) );
BUF_X4 _10038_ ( .A(_02157_ ), .Z(_02411_ ) );
OAI211_X1 _10039_ ( .A(_02410_ ), .B(_02184_ ), .C1(_02411_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02412_ ) );
OR2_X1 _10040_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02413_ ) );
OAI211_X1 _10041_ ( .A(_02413_ ), .B(fanout_net_24 ), .C1(_02158_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02414_ ) );
NAND3_X1 _10042_ ( .A1(_02412_ ), .A2(_02414_ ), .A3(_02106_ ), .ZN(_02415_ ) );
MUX2_X1 _10043_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02416_ ) );
MUX2_X1 _10044_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02417_ ) );
MUX2_X1 _10045_ ( .A(_02416_ ), .B(_02417_ ), .S(_02153_ ), .Z(_02418_ ) );
OAI211_X1 _10046_ ( .A(_02374_ ), .B(_02415_ ), .C1(_02418_ ), .C2(_02107_ ), .ZN(_02419_ ) );
OR2_X1 _10047_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02420_ ) );
OAI211_X1 _10048_ ( .A(_02420_ ), .B(fanout_net_24 ), .C1(_02158_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02421_ ) );
OR2_X1 _10049_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02422_ ) );
OAI211_X1 _10050_ ( .A(_02422_ ), .B(_02184_ ), .C1(_02158_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02423_ ) );
NAND3_X1 _10051_ ( .A1(_02421_ ), .A2(_02423_ ), .A3(fanout_net_26 ), .ZN(_02424_ ) );
MUX2_X1 _10052_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02425_ ) );
MUX2_X1 _10053_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02426_ ) );
MUX2_X1 _10054_ ( .A(_02425_ ), .B(_02426_ ), .S(fanout_net_24 ), .Z(_02427_ ) );
OAI211_X1 _10055_ ( .A(fanout_net_27 ), .B(_02424_ ), .C1(_02427_ ), .C2(fanout_net_26 ), .ZN(_02428_ ) );
OAI211_X1 _10056_ ( .A(_02419_ ), .B(_02428_ ), .C1(_02139_ ), .C2(_02180_ ), .ZN(_02429_ ) );
NAND2_X1 _10057_ ( .A1(_02409_ ), .A2(_02429_ ), .ZN(_02430_ ) );
INV_X1 _10058_ ( .A(\ID_EX_imm [17] ), .ZN(_02431_ ) );
XNOR2_X1 _10059_ ( .A(_02430_ ), .B(_02431_ ), .ZN(_02432_ ) );
OR3_X1 _10060_ ( .A1(_02140_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02181_ ), .ZN(_02433_ ) );
OR2_X1 _10061_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02434_ ) );
OAI211_X1 _10062_ ( .A(_02434_ ), .B(_02115_ ), .C1(_02214_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02435_ ) );
OR2_X1 _10063_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02436_ ) );
OAI211_X1 _10064_ ( .A(_02436_ ), .B(fanout_net_24 ), .C1(_02214_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02437_ ) );
NAND3_X1 _10065_ ( .A1(_02435_ ), .A2(_02437_ ), .A3(fanout_net_26 ), .ZN(_02438_ ) );
MUX2_X1 _10066_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02439_ ) );
MUX2_X1 _10067_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02440_ ) );
MUX2_X1 _10068_ ( .A(_02439_ ), .B(_02440_ ), .S(_02186_ ), .Z(_02441_ ) );
OAI211_X1 _10069_ ( .A(_02105_ ), .B(_02438_ ), .C1(_02441_ ), .C2(fanout_net_26 ), .ZN(_02442_ ) );
NOR2_X1 _10070_ ( .A1(_02188_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02443_ ) );
OAI21_X1 _10071_ ( .A(fanout_net_24 ), .B1(fanout_net_18 ), .B2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02444_ ) );
NOR2_X1 _10072_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02445_ ) );
OAI21_X1 _10073_ ( .A(_02186_ ), .B1(_02188_ ), .B2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02446_ ) );
OAI221_X1 _10074_ ( .A(_02193_ ), .B1(_02443_ ), .B2(_02444_ ), .C1(_02445_ ), .C2(_02446_ ), .ZN(_02447_ ) );
MUX2_X1 _10075_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02448_ ) );
MUX2_X1 _10076_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02449_ ) );
MUX2_X1 _10077_ ( .A(_02448_ ), .B(_02449_ ), .S(fanout_net_24 ), .Z(_02450_ ) );
OAI211_X1 _10078_ ( .A(fanout_net_27 ), .B(_02447_ ), .C1(_02450_ ), .C2(_02118_ ), .ZN(_02451_ ) );
OAI211_X1 _10079_ ( .A(_02442_ ), .B(_02451_ ), .C1(_02176_ ), .C2(_02150_ ), .ZN(_02452_ ) );
NAND2_X1 _10080_ ( .A1(_02433_ ), .A2(_02452_ ), .ZN(_02453_ ) );
BUF_X4 _10081_ ( .A(_02453_ ), .Z(_02454_ ) );
INV_X1 _10082_ ( .A(\ID_EX_imm [16] ), .ZN(_02455_ ) );
XNOR2_X1 _10083_ ( .A(_02454_ ), .B(_02455_ ), .ZN(_02456_ ) );
NAND3_X1 _10084_ ( .A1(_02408_ ), .A2(_02432_ ), .A3(_02456_ ), .ZN(_02457_ ) );
OR3_X1 _10085_ ( .A1(_02174_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02148_ ), .ZN(_02458_ ) );
OR2_X1 _10086_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02459_ ) );
OAI211_X1 _10087_ ( .A(_02459_ ), .B(_02113_ ), .C1(_02163_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02460_ ) );
OR2_X1 _10088_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02461_ ) );
OAI211_X1 _10089_ ( .A(_02461_ ), .B(fanout_net_24 ), .C1(_02411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02462_ ) );
NAND3_X1 _10090_ ( .A1(_02460_ ), .A2(_02462_ ), .A3(_02265_ ), .ZN(_02463_ ) );
MUX2_X1 _10091_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02464_ ) );
MUX2_X1 _10092_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02465_ ) );
MUX2_X1 _10093_ ( .A(_02464_ ), .B(_02465_ ), .S(_02184_ ), .Z(_02466_ ) );
OAI211_X1 _10094_ ( .A(_02374_ ), .B(_02463_ ), .C1(_02466_ ), .C2(_02192_ ), .ZN(_02467_ ) );
OR2_X1 _10095_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02468_ ) );
OAI211_X1 _10096_ ( .A(_02468_ ), .B(fanout_net_24 ), .C1(_02411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02469_ ) );
OR2_X1 _10097_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02470_ ) );
OAI211_X1 _10098_ ( .A(_02470_ ), .B(_02184_ ), .C1(_02411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02471_ ) );
NAND3_X1 _10099_ ( .A1(_02469_ ), .A2(_02471_ ), .A3(fanout_net_26 ), .ZN(_02472_ ) );
MUX2_X1 _10100_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02473_ ) );
MUX2_X1 _10101_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02474_ ) );
MUX2_X1 _10102_ ( .A(_02473_ ), .B(_02474_ ), .S(fanout_net_24 ), .Z(_02475_ ) );
OAI211_X1 _10103_ ( .A(fanout_net_27 ), .B(_02472_ ), .C1(_02475_ ), .C2(fanout_net_26 ), .ZN(_02476_ ) );
OAI211_X1 _10104_ ( .A(_02467_ ), .B(_02476_ ), .C1(_02139_ ), .C2(_02259_ ), .ZN(_02477_ ) );
NAND2_X2 _10105_ ( .A1(_02458_ ), .A2(_02477_ ), .ZN(_02478_ ) );
XNOR2_X1 _10106_ ( .A(_02478_ ), .B(\ID_EX_imm [1] ), .ZN(_02479_ ) );
INV_X1 _10107_ ( .A(\ID_EX_imm [0] ), .ZN(_02480_ ) );
OR3_X1 _10108_ ( .A1(_02138_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_02147_ ), .ZN(_02481_ ) );
OR2_X1 _10109_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(fanout_net_18 ), .ZN(_02482_ ) );
BUF_X4 _10110_ ( .A(_02156_ ), .Z(_02483_ ) );
OAI211_X1 _10111_ ( .A(_02482_ ), .B(_02153_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_02483_ ), .ZN(_02484_ ) );
OR2_X1 _10112_ ( .A1(fanout_net_18 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02485_ ) );
OAI211_X1 _10113_ ( .A(_02485_ ), .B(fanout_net_24 ), .C1(_02483_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02486_ ) );
NAND3_X1 _10114_ ( .A1(_02484_ ), .A2(_02486_ ), .A3(_02106_ ), .ZN(_02487_ ) );
MUX2_X1 _10115_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02488_ ) );
MUX2_X1 _10116_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02489_ ) );
MUX2_X1 _10117_ ( .A(_02488_ ), .B(_02489_ ), .S(_02112_ ), .Z(_02490_ ) );
OAI211_X1 _10118_ ( .A(_02103_ ), .B(_02487_ ), .C1(_02490_ ), .C2(_02265_ ), .ZN(_02491_ ) );
OR2_X1 _10119_ ( .A1(fanout_net_18 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02492_ ) );
OAI211_X1 _10120_ ( .A(_02492_ ), .B(fanout_net_24 ), .C1(_02483_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02493_ ) );
OR2_X1 _10121_ ( .A1(fanout_net_18 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02494_ ) );
OAI211_X1 _10122_ ( .A(_02494_ ), .B(_02153_ ), .C1(_02483_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02495_ ) );
NAND3_X1 _10123_ ( .A1(_02493_ ), .A2(_02495_ ), .A3(fanout_net_26 ), .ZN(_02496_ ) );
MUX2_X1 _10124_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02497_ ) );
MUX2_X1 _10125_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02498_ ) );
MUX2_X1 _10126_ ( .A(_02497_ ), .B(_02498_ ), .S(fanout_net_24 ), .Z(_02499_ ) );
OAI211_X1 _10127_ ( .A(fanout_net_27 ), .B(_02496_ ), .C1(_02499_ ), .C2(fanout_net_26 ), .ZN(_02500_ ) );
OAI211_X1 _10128_ ( .A(_02491_ ), .B(_02500_ ), .C1(_02174_ ), .C2(_02148_ ), .ZN(_02501_ ) );
NAND2_X1 _10129_ ( .A1(_02481_ ), .A2(_02501_ ), .ZN(_02502_ ) );
INV_X1 _10130_ ( .A(_02502_ ), .ZN(_02503_ ) );
NOR3_X1 _10131_ ( .A1(_02479_ ), .A2(_02480_ ), .A3(_02503_ ), .ZN(_02504_ ) );
AOI21_X1 _10132_ ( .A(_02504_ ), .B1(\ID_EX_imm [1] ), .B2(_02478_ ), .ZN(_02505_ ) );
OR3_X1 _10133_ ( .A1(_02379_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02259_ ), .ZN(_02506_ ) );
OR2_X1 _10134_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02507_ ) );
OAI211_X1 _10135_ ( .A(_02507_ ), .B(_02154_ ), .C1(_02159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02508_ ) );
OR2_X1 _10136_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02509_ ) );
OAI211_X1 _10137_ ( .A(_02509_ ), .B(fanout_net_24 ), .C1(_02360_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02510_ ) );
NAND3_X1 _10138_ ( .A1(_02508_ ), .A2(_02510_ ), .A3(fanout_net_26 ), .ZN(_02511_ ) );
MUX2_X1 _10139_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02512_ ) );
MUX2_X1 _10140_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02513_ ) );
MUX2_X1 _10141_ ( .A(_02512_ ), .B(_02513_ ), .S(_02154_ ), .Z(_02514_ ) );
OAI211_X1 _10142_ ( .A(_02104_ ), .B(_02511_ ), .C1(_02514_ ), .C2(fanout_net_26 ), .ZN(_02515_ ) );
NOR2_X1 _10143_ ( .A1(fanout_net_18 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02516_ ) );
OAI21_X1 _10144_ ( .A(_02113_ ), .B1(_02163_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02517_ ) );
INV_X1 _10145_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02518_ ) );
INV_X1 _10146_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02519_ ) );
MUX2_X1 _10147_ ( .A(_02518_ ), .B(_02519_ ), .S(fanout_net_18 ), .Z(_02520_ ) );
OAI221_X1 _10148_ ( .A(_02107_ ), .B1(_02516_ ), .B2(_02517_ ), .C1(_02520_ ), .C2(_02114_ ), .ZN(_02521_ ) );
MUX2_X1 _10149_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02522_ ) );
MUX2_X1 _10150_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02523_ ) );
MUX2_X1 _10151_ ( .A(_02522_ ), .B(_02523_ ), .S(fanout_net_24 ), .Z(_02524_ ) );
OAI211_X1 _10152_ ( .A(fanout_net_27 ), .B(_02521_ ), .C1(_02524_ ), .C2(_02108_ ), .ZN(_02525_ ) );
OAI211_X1 _10153_ ( .A(_02515_ ), .B(_02525_ ), .C1(_02175_ ), .C2(_02149_ ), .ZN(_02526_ ) );
NAND2_X1 _10154_ ( .A1(_02506_ ), .A2(_02526_ ), .ZN(_02527_ ) );
XNOR2_X1 _10155_ ( .A(_02527_ ), .B(\ID_EX_imm [3] ), .ZN(_02528_ ) );
OR3_X1 _10156_ ( .A1(_02379_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02259_ ), .ZN(_02529_ ) );
OR2_X1 _10157_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02530_ ) );
OAI211_X1 _10158_ ( .A(_02530_ ), .B(_02185_ ), .C1(_02159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02531_ ) );
OR2_X1 _10159_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02532_ ) );
OAI211_X1 _10160_ ( .A(_02532_ ), .B(fanout_net_24 ), .C1(_02159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02533_ ) );
NAND3_X1 _10161_ ( .A1(_02531_ ), .A2(_02533_ ), .A3(_02192_ ), .ZN(_02534_ ) );
MUX2_X1 _10162_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02535_ ) );
MUX2_X1 _10163_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02536_ ) );
MUX2_X1 _10164_ ( .A(_02535_ ), .B(_02536_ ), .S(_02154_ ), .Z(_02537_ ) );
OAI211_X1 _10165_ ( .A(_02104_ ), .B(_02534_ ), .C1(_02537_ ), .C2(_02108_ ), .ZN(_02538_ ) );
OR2_X1 _10166_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02539_ ) );
OAI211_X1 _10167_ ( .A(_02539_ ), .B(fanout_net_24 ), .C1(_02159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02540_ ) );
OR2_X1 _10168_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02541_ ) );
OAI211_X1 _10169_ ( .A(_02541_ ), .B(_02185_ ), .C1(_02159_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02542_ ) );
NAND3_X1 _10170_ ( .A1(_02540_ ), .A2(_02542_ ), .A3(fanout_net_26 ), .ZN(_02543_ ) );
MUX2_X1 _10171_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02544_ ) );
MUX2_X1 _10172_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02545_ ) );
MUX2_X1 _10173_ ( .A(_02544_ ), .B(_02545_ ), .S(fanout_net_24 ), .Z(_02546_ ) );
OAI211_X1 _10174_ ( .A(fanout_net_27 ), .B(_02543_ ), .C1(_02546_ ), .C2(fanout_net_26 ), .ZN(_02547_ ) );
OAI211_X1 _10175_ ( .A(_02538_ ), .B(_02547_ ), .C1(_02175_ ), .C2(_02149_ ), .ZN(_02548_ ) );
NAND2_X1 _10176_ ( .A1(_02529_ ), .A2(_02548_ ), .ZN(_02549_ ) );
XNOR2_X1 _10177_ ( .A(_02549_ ), .B(\ID_EX_imm [2] ), .ZN(_02550_ ) );
NOR3_X1 _10178_ ( .A1(_02505_ ), .A2(_02528_ ), .A3(_02550_ ), .ZN(_02551_ ) );
INV_X1 _10179_ ( .A(_02528_ ), .ZN(_02552_ ) );
AND2_X1 _10180_ ( .A1(_02549_ ), .A2(\ID_EX_imm [2] ), .ZN(_02553_ ) );
NAND2_X1 _10181_ ( .A1(_02552_ ), .A2(_02553_ ), .ZN(_02554_ ) );
INV_X1 _10182_ ( .A(_02527_ ), .ZN(_02555_ ) );
OAI21_X1 _10183_ ( .A(_02554_ ), .B1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B2(_02555_ ), .ZN(_02556_ ) );
NOR2_X1 _10184_ ( .A1(_02551_ ), .A2(_02556_ ), .ZN(_02557_ ) );
INV_X1 _10185_ ( .A(_02557_ ), .ZN(_02558_ ) );
OR3_X1 _10186_ ( .A1(_02174_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02148_ ), .ZN(_02559_ ) );
OR2_X1 _10187_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02560_ ) );
OAI211_X1 _10188_ ( .A(_02560_ ), .B(_02184_ ), .C1(_02411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02561_ ) );
OR2_X1 _10189_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02562_ ) );
OAI211_X1 _10190_ ( .A(_02562_ ), .B(fanout_net_24 ), .C1(_02411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02563_ ) );
NAND3_X1 _10191_ ( .A1(_02561_ ), .A2(_02563_ ), .A3(_02265_ ), .ZN(_02564_ ) );
MUX2_X1 _10192_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02565_ ) );
MUX2_X1 _10193_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02566_ ) );
MUX2_X1 _10194_ ( .A(_02565_ ), .B(_02566_ ), .S(_02184_ ), .Z(_02567_ ) );
OAI211_X1 _10195_ ( .A(fanout_net_27 ), .B(_02564_ ), .C1(_02567_ ), .C2(_02107_ ), .ZN(_02568_ ) );
OR2_X1 _10196_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02569_ ) );
OAI211_X1 _10197_ ( .A(_02569_ ), .B(_02184_ ), .C1(_02411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02570_ ) );
OR2_X1 _10198_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02571_ ) );
OAI211_X1 _10199_ ( .A(_02571_ ), .B(fanout_net_24 ), .C1(_02411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02572_ ) );
NAND3_X1 _10200_ ( .A1(_02570_ ), .A2(_02572_ ), .A3(_02265_ ), .ZN(_02573_ ) );
MUX2_X1 _10201_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02574_ ) );
MUX2_X1 _10202_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02575_ ) );
MUX2_X1 _10203_ ( .A(_02574_ ), .B(_02575_ ), .S(_02153_ ), .Z(_02576_ ) );
OAI211_X1 _10204_ ( .A(_02374_ ), .B(_02573_ ), .C1(_02576_ ), .C2(_02107_ ), .ZN(_02577_ ) );
OAI211_X4 _10205_ ( .A(_02568_ ), .B(_02577_ ), .C1(_02139_ ), .C2(_02180_ ), .ZN(_02578_ ) );
NAND2_X2 _10206_ ( .A1(_02559_ ), .A2(_02578_ ), .ZN(_02579_ ) );
XNOR2_X1 _10207_ ( .A(_02579_ ), .B(\ID_EX_imm [5] ), .ZN(_02580_ ) );
INV_X1 _10208_ ( .A(_02580_ ), .ZN(_02581_ ) );
OR3_X1 _10209_ ( .A1(_02139_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02180_ ), .ZN(_02582_ ) );
OR2_X1 _10210_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02583_ ) );
OAI211_X1 _10211_ ( .A(_02583_ ), .B(_02154_ ), .C1(_02360_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02584_ ) );
OR2_X1 _10212_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02585_ ) );
BUF_X4 _10213_ ( .A(_02483_ ), .Z(_02586_ ) );
OAI211_X1 _10214_ ( .A(_02585_ ), .B(fanout_net_24 ), .C1(_02586_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02587_ ) );
NAND3_X1 _10215_ ( .A1(_02584_ ), .A2(_02587_ ), .A3(_02107_ ), .ZN(_02588_ ) );
MUX2_X1 _10216_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02589_ ) );
MUX2_X1 _10217_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02590_ ) );
MUX2_X1 _10218_ ( .A(_02589_ ), .B(_02590_ ), .S(_02367_ ), .Z(_02591_ ) );
OAI211_X1 _10219_ ( .A(fanout_net_27 ), .B(_02588_ ), .C1(_02591_ ), .C2(_02266_ ), .ZN(_02592_ ) );
OR2_X1 _10220_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02593_ ) );
OAI211_X1 _10221_ ( .A(_02593_ ), .B(_02154_ ), .C1(_02360_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02594_ ) );
OR2_X1 _10222_ ( .A1(fanout_net_19 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02595_ ) );
OAI211_X1 _10223_ ( .A(_02595_ ), .B(fanout_net_24 ), .C1(_02586_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02596_ ) );
NAND3_X1 _10224_ ( .A1(_02594_ ), .A2(_02596_ ), .A3(_02107_ ), .ZN(_02597_ ) );
MUX2_X1 _10225_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02598_ ) );
MUX2_X1 _10226_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02599_ ) );
MUX2_X1 _10227_ ( .A(_02598_ ), .B(_02599_ ), .S(_02113_ ), .Z(_02600_ ) );
OAI211_X1 _10228_ ( .A(_02104_ ), .B(_02597_ ), .C1(_02600_ ), .C2(_02266_ ), .ZN(_02601_ ) );
OAI211_X1 _10229_ ( .A(_02592_ ), .B(_02601_ ), .C1(_02379_ ), .C2(_02149_ ), .ZN(_02602_ ) );
NAND2_X1 _10230_ ( .A1(_02582_ ), .A2(_02602_ ), .ZN(_02603_ ) );
INV_X1 _10231_ ( .A(\ID_EX_imm [4] ), .ZN(_02604_ ) );
XNOR2_X1 _10232_ ( .A(_02603_ ), .B(_02604_ ), .ZN(_02605_ ) );
OR3_X1 _10233_ ( .A1(_02379_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02180_ ), .ZN(_02606_ ) );
OR2_X1 _10234_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02607_ ) );
OAI211_X1 _10235_ ( .A(_02607_ ), .B(_02154_ ), .C1(_02360_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02608_ ) );
OR2_X1 _10236_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02609_ ) );
OAI211_X1 _10237_ ( .A(_02609_ ), .B(fanout_net_24 ), .C1(_02360_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02610_ ) );
NAND3_X1 _10238_ ( .A1(_02608_ ), .A2(_02610_ ), .A3(_02192_ ), .ZN(_02611_ ) );
MUX2_X1 _10239_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02612_ ) );
MUX2_X1 _10240_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02613_ ) );
MUX2_X1 _10241_ ( .A(_02612_ ), .B(_02613_ ), .S(_02367_ ), .Z(_02614_ ) );
OAI211_X1 _10242_ ( .A(_02104_ ), .B(_02611_ ), .C1(_02614_ ), .C2(_02266_ ), .ZN(_02615_ ) );
OR2_X1 _10243_ ( .A1(fanout_net_20 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02616_ ) );
OAI211_X1 _10244_ ( .A(_02616_ ), .B(fanout_net_24 ), .C1(_02360_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02617_ ) );
OR2_X1 _10245_ ( .A1(fanout_net_20 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02618_ ) );
OAI211_X1 _10246_ ( .A(_02618_ ), .B(_02154_ ), .C1(_02360_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02619_ ) );
NAND3_X1 _10247_ ( .A1(_02617_ ), .A2(_02619_ ), .A3(fanout_net_26 ), .ZN(_02620_ ) );
MUX2_X1 _10248_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02621_ ) );
MUX2_X1 _10249_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02622_ ) );
MUX2_X1 _10250_ ( .A(_02621_ ), .B(_02622_ ), .S(fanout_net_24 ), .Z(_02623_ ) );
OAI211_X1 _10251_ ( .A(fanout_net_27 ), .B(_02620_ ), .C1(_02623_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02624_ ) );
OAI211_X1 _10252_ ( .A(_02615_ ), .B(_02624_ ), .C1(_02379_ ), .C2(_02149_ ), .ZN(_02625_ ) );
NAND2_X2 _10253_ ( .A1(_02606_ ), .A2(_02625_ ), .ZN(_02626_ ) );
INV_X1 _10254_ ( .A(\ID_EX_imm [6] ), .ZN(_02627_ ) );
XNOR2_X1 _10255_ ( .A(_02626_ ), .B(_02627_ ), .ZN(_02628_ ) );
OR3_X1 _10256_ ( .A1(_02138_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02147_ ), .ZN(_02629_ ) );
INV_X1 _10257_ ( .A(\ID_EX_imm [7] ), .ZN(_02630_ ) );
OR2_X1 _10258_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02631_ ) );
OAI211_X1 _10259_ ( .A(_02631_ ), .B(_02153_ ), .C1(_02158_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02632_ ) );
OR2_X1 _10260_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02633_ ) );
OAI211_X1 _10261_ ( .A(_02633_ ), .B(fanout_net_24 ), .C1(_02158_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02634_ ) );
NAND3_X1 _10262_ ( .A1(_02632_ ), .A2(_02634_ ), .A3(_02106_ ), .ZN(_02635_ ) );
MUX2_X1 _10263_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02636_ ) );
MUX2_X1 _10264_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02637_ ) );
MUX2_X1 _10265_ ( .A(_02636_ ), .B(_02637_ ), .S(_02153_ ), .Z(_02638_ ) );
OAI211_X1 _10266_ ( .A(_02374_ ), .B(_02635_ ), .C1(_02638_ ), .C2(_02107_ ), .ZN(_02639_ ) );
OR2_X1 _10267_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02640_ ) );
OAI211_X1 _10268_ ( .A(_02640_ ), .B(fanout_net_24 ), .C1(_02158_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02641_ ) );
OR2_X1 _10269_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02642_ ) );
OAI211_X1 _10270_ ( .A(_02642_ ), .B(_02153_ ), .C1(_02158_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02643_ ) );
NAND3_X1 _10271_ ( .A1(_02641_ ), .A2(_02643_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02644_ ) );
MUX2_X1 _10272_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02645_ ) );
MUX2_X1 _10273_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02646_ ) );
MUX2_X1 _10274_ ( .A(_02645_ ), .B(_02646_ ), .S(fanout_net_24 ), .Z(_02647_ ) );
OAI211_X1 _10275_ ( .A(fanout_net_27 ), .B(_02644_ ), .C1(_02647_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02648_ ) );
OAI211_X1 _10276_ ( .A(_02639_ ), .B(_02648_ ), .C1(_02174_ ), .C2(_02148_ ), .ZN(_02649_ ) );
NAND3_X1 _10277_ ( .A1(_02629_ ), .A2(_02630_ ), .A3(_02649_ ), .ZN(_02650_ ) );
NAND2_X1 _10278_ ( .A1(_02629_ ), .A2(_02649_ ), .ZN(_02651_ ) );
NAND2_X1 _10279_ ( .A1(_02651_ ), .A2(\ID_EX_imm [7] ), .ZN(_02652_ ) );
AND3_X1 _10280_ ( .A1(_02628_ ), .A2(_02650_ ), .A3(_02652_ ), .ZN(_02653_ ) );
NAND4_X1 _10281_ ( .A1(_02558_ ), .A2(_02581_ ), .A3(_02605_ ), .A4(_02653_ ), .ZN(_02654_ ) );
AND4_X1 _10282_ ( .A1(\ID_EX_imm [6] ), .A2(_02652_ ), .A3(_02626_ ), .A4(_02650_ ), .ZN(_02655_ ) );
INV_X4 _10283_ ( .A(_02603_ ), .ZN(_02656_ ) );
NOR3_X1 _10284_ ( .A1(_02580_ ), .A2(_02604_ ), .A3(_02656_ ), .ZN(_02657_ ) );
AOI21_X1 _10285_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02559_ ), .B2(_02578_ ), .ZN(_02658_ ) );
NOR2_X1 _10286_ ( .A1(_02657_ ), .A2(_02658_ ), .ZN(_02659_ ) );
INV_X1 _10287_ ( .A(_02659_ ), .ZN(_02660_ ) );
AOI221_X4 _10288_ ( .A(_02655_ ), .B1(\ID_EX_imm [7] ), .B2(_02651_ ), .C1(_02660_ ), .C2(_02653_ ), .ZN(_02661_ ) );
NAND2_X1 _10289_ ( .A1(_02654_ ), .A2(_02661_ ), .ZN(_02662_ ) );
OR3_X1 _10290_ ( .A1(_02139_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02180_ ), .ZN(_02663_ ) );
OR2_X1 _10291_ ( .A1(_02483_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02664_ ) );
OAI211_X1 _10292_ ( .A(_02664_ ), .B(fanout_net_24 ), .C1(fanout_net_20 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02665_ ) );
OR2_X1 _10293_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02666_ ) );
OAI211_X1 _10294_ ( .A(_02666_ ), .B(_02367_ ), .C1(_02586_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02667_ ) );
NAND3_X1 _10295_ ( .A1(_02665_ ), .A2(_02192_ ), .A3(_02667_ ), .ZN(_02668_ ) );
MUX2_X1 _10296_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02669_ ) );
MUX2_X1 _10297_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02670_ ) );
MUX2_X1 _10298_ ( .A(_02669_ ), .B(_02670_ ), .S(_02367_ ), .Z(_02671_ ) );
OAI211_X1 _10299_ ( .A(_02104_ ), .B(_02668_ ), .C1(_02671_ ), .C2(_02266_ ), .ZN(_02672_ ) );
OR2_X1 _10300_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02673_ ) );
OAI211_X1 _10301_ ( .A(_02673_ ), .B(fanout_net_24 ), .C1(_02360_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02674_ ) );
OR2_X1 _10302_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02675_ ) );
OAI211_X1 _10303_ ( .A(_02675_ ), .B(_02367_ ), .C1(_02586_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02676_ ) );
NAND3_X1 _10304_ ( .A1(_02674_ ), .A2(_02676_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02677_ ) );
MUX2_X1 _10305_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02678_ ) );
MUX2_X1 _10306_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02679_ ) );
MUX2_X1 _10307_ ( .A(_02678_ ), .B(_02679_ ), .S(fanout_net_24 ), .Z(_02680_ ) );
OAI211_X1 _10308_ ( .A(fanout_net_27 ), .B(_02677_ ), .C1(_02680_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02681_ ) );
OAI211_X1 _10309_ ( .A(_02672_ ), .B(_02681_ ), .C1(_02379_ ), .C2(_02259_ ), .ZN(_02682_ ) );
NAND2_X2 _10310_ ( .A1(_02663_ ), .A2(_02682_ ), .ZN(_02683_ ) );
INV_X1 _10311_ ( .A(\ID_EX_imm [15] ), .ZN(_02684_ ) );
XNOR2_X1 _10312_ ( .A(_02683_ ), .B(_02684_ ), .ZN(_02685_ ) );
OR3_X1 _10313_ ( .A1(_02139_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02180_ ), .ZN(_02686_ ) );
OR2_X1 _10314_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02687_ ) );
OAI211_X1 _10315_ ( .A(_02687_ ), .B(_02367_ ), .C1(_02586_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02688_ ) );
OR2_X1 _10316_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02689_ ) );
OAI211_X1 _10317_ ( .A(_02689_ ), .B(fanout_net_25 ), .C1(_02586_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02690_ ) );
NAND3_X1 _10318_ ( .A1(_02688_ ), .A2(_02690_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02691_ ) );
MUX2_X1 _10319_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02692_ ) );
MUX2_X1 _10320_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02693_ ) );
MUX2_X1 _10321_ ( .A(_02692_ ), .B(_02693_ ), .S(_02113_ ), .Z(_02694_ ) );
OAI211_X1 _10322_ ( .A(_02374_ ), .B(_02691_ ), .C1(_02694_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02695_ ) );
NOR2_X1 _10323_ ( .A1(_02411_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02696_ ) );
OAI21_X1 _10324_ ( .A(fanout_net_25 ), .B1(fanout_net_20 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02697_ ) );
NOR2_X1 _10325_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02698_ ) );
OAI21_X1 _10326_ ( .A(_02113_ ), .B1(_02163_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02699_ ) );
OAI221_X1 _10327_ ( .A(_02265_ ), .B1(_02696_ ), .B2(_02697_ ), .C1(_02698_ ), .C2(_02699_ ), .ZN(_02700_ ) );
MUX2_X1 _10328_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02701_ ) );
MUX2_X1 _10329_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02702_ ) );
MUX2_X1 _10330_ ( .A(_02701_ ), .B(_02702_ ), .S(fanout_net_25 ), .Z(_02703_ ) );
OAI211_X1 _10331_ ( .A(fanout_net_27 ), .B(_02700_ ), .C1(_02703_ ), .C2(_02192_ ), .ZN(_02704_ ) );
OAI211_X1 _10332_ ( .A(_02695_ ), .B(_02704_ ), .C1(_02379_ ), .C2(_02259_ ), .ZN(_02705_ ) );
NAND2_X2 _10333_ ( .A1(_02686_ ), .A2(_02705_ ), .ZN(_02706_ ) );
BUF_X4 _10334_ ( .A(_02706_ ), .Z(_02707_ ) );
INV_X1 _10335_ ( .A(\ID_EX_imm [14] ), .ZN(_02708_ ) );
XNOR2_X1 _10336_ ( .A(_02707_ ), .B(_02708_ ), .ZN(_02709_ ) );
AND2_X1 _10337_ ( .A1(_02685_ ), .A2(_02709_ ), .ZN(_02710_ ) );
OR3_X1 _10338_ ( .A1(_02174_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02148_ ), .ZN(_02711_ ) );
OR2_X1 _10339_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02712_ ) );
OAI211_X1 _10340_ ( .A(_02712_ ), .B(_02367_ ), .C1(_02586_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02713_ ) );
OR2_X1 _10341_ ( .A1(fanout_net_20 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02714_ ) );
OAI211_X1 _10342_ ( .A(_02714_ ), .B(fanout_net_25 ), .C1(_02163_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02715_ ) );
NAND3_X1 _10343_ ( .A1(_02713_ ), .A2(_02715_ ), .A3(_02107_ ), .ZN(_02716_ ) );
MUX2_X1 _10344_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02717_ ) );
MUX2_X1 _10345_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02718_ ) );
MUX2_X1 _10346_ ( .A(_02717_ ), .B(_02718_ ), .S(_02113_ ), .Z(_02719_ ) );
OAI211_X1 _10347_ ( .A(_02374_ ), .B(_02716_ ), .C1(_02719_ ), .C2(_02192_ ), .ZN(_02720_ ) );
OR2_X1 _10348_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02721_ ) );
OAI211_X1 _10349_ ( .A(_02721_ ), .B(fanout_net_25 ), .C1(_02163_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02722_ ) );
OR2_X1 _10350_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02723_ ) );
OAI211_X1 _10351_ ( .A(_02723_ ), .B(_02113_ ), .C1(_02163_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02724_ ) );
NAND3_X1 _10352_ ( .A1(_02722_ ), .A2(_02724_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02725_ ) );
MUX2_X1 _10353_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02726_ ) );
MUX2_X1 _10354_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02727_ ) );
MUX2_X1 _10355_ ( .A(_02726_ ), .B(_02727_ ), .S(fanout_net_25 ), .Z(_02728_ ) );
OAI211_X1 _10356_ ( .A(fanout_net_27 ), .B(_02725_ ), .C1(_02728_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02729_ ) );
OAI211_X1 _10357_ ( .A(_02720_ ), .B(_02729_ ), .C1(_02379_ ), .C2(_02259_ ), .ZN(_02730_ ) );
NAND2_X2 _10358_ ( .A1(_02711_ ), .A2(_02730_ ), .ZN(_02731_ ) );
INV_X1 _10359_ ( .A(\ID_EX_imm [12] ), .ZN(_02732_ ) );
XNOR2_X1 _10360_ ( .A(_02731_ ), .B(_02732_ ), .ZN(_02733_ ) );
OR3_X1 _10361_ ( .A1(_02138_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02147_ ), .ZN(_02734_ ) );
INV_X1 _10362_ ( .A(\ID_EX_imm [13] ), .ZN(_02735_ ) );
OR2_X1 _10363_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02736_ ) );
OAI211_X1 _10364_ ( .A(_02736_ ), .B(_02112_ ), .C1(_02157_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02737_ ) );
OR2_X1 _10365_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02738_ ) );
OAI211_X1 _10366_ ( .A(_02738_ ), .B(fanout_net_25 ), .C1(_02157_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02739_ ) );
NAND3_X1 _10367_ ( .A1(_02737_ ), .A2(_02739_ ), .A3(_02106_ ), .ZN(_02740_ ) );
MUX2_X1 _10368_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02741_ ) );
MUX2_X1 _10369_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02742_ ) );
MUX2_X1 _10370_ ( .A(_02741_ ), .B(_02742_ ), .S(_02111_ ), .Z(_02743_ ) );
OAI211_X1 _10371_ ( .A(_02103_ ), .B(_02740_ ), .C1(_02743_ ), .C2(_02106_ ), .ZN(_02744_ ) );
OR2_X1 _10372_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02745_ ) );
OAI211_X1 _10373_ ( .A(_02745_ ), .B(fanout_net_25 ), .C1(_02157_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02746_ ) );
OR2_X1 _10374_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02747_ ) );
OAI211_X1 _10375_ ( .A(_02747_ ), .B(_02111_ ), .C1(_02157_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02748_ ) );
NAND3_X1 _10376_ ( .A1(_02746_ ), .A2(_02748_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02749_ ) );
MUX2_X1 _10377_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02750_ ) );
MUX2_X1 _10378_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02751_ ) );
MUX2_X1 _10379_ ( .A(_02750_ ), .B(_02751_ ), .S(fanout_net_25 ), .Z(_02752_ ) );
OAI211_X1 _10380_ ( .A(fanout_net_27 ), .B(_02749_ ), .C1(_02752_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02753_ ) );
OAI211_X1 _10381_ ( .A(_02744_ ), .B(_02753_ ), .C1(_02138_ ), .C2(_02147_ ), .ZN(_02754_ ) );
AND3_X1 _10382_ ( .A1(_02734_ ), .A2(_02735_ ), .A3(_02754_ ), .ZN(_02755_ ) );
AOI21_X1 _10383_ ( .A(_02735_ ), .B1(_02734_ ), .B2(_02754_ ), .ZN(_02756_ ) );
NOR2_X1 _10384_ ( .A1(_02755_ ), .A2(_02756_ ), .ZN(_02757_ ) );
AND2_X1 _10385_ ( .A1(_02733_ ), .A2(_02757_ ), .ZN(_02758_ ) );
AND2_X1 _10386_ ( .A1(_02710_ ), .A2(_02758_ ), .ZN(_02759_ ) );
OR3_X1 _10387_ ( .A1(_02139_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02180_ ), .ZN(_02760_ ) );
OR2_X1 _10388_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02761_ ) );
OAI211_X1 _10389_ ( .A(_02761_ ), .B(_02367_ ), .C1(_02586_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02762_ ) );
OR2_X1 _10390_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02763_ ) );
OAI211_X1 _10391_ ( .A(_02763_ ), .B(fanout_net_25 ), .C1(_02586_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02764_ ) );
NAND3_X1 _10392_ ( .A1(_02762_ ), .A2(_02764_ ), .A3(_02107_ ), .ZN(_02765_ ) );
MUX2_X1 _10393_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02766_ ) );
MUX2_X1 _10394_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02767_ ) );
MUX2_X1 _10395_ ( .A(_02766_ ), .B(_02767_ ), .S(_02113_ ), .Z(_02768_ ) );
OAI211_X1 _10396_ ( .A(_02374_ ), .B(_02765_ ), .C1(_02768_ ), .C2(_02266_ ), .ZN(_02769_ ) );
OR2_X1 _10397_ ( .A1(_02483_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02770_ ) );
OAI211_X1 _10398_ ( .A(_02770_ ), .B(fanout_net_25 ), .C1(fanout_net_21 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02771_ ) );
OR2_X1 _10399_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02772_ ) );
OAI211_X1 _10400_ ( .A(_02772_ ), .B(_02367_ ), .C1(_02586_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02773_ ) );
NAND3_X1 _10401_ ( .A1(_02771_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02773_ ), .ZN(_02774_ ) );
MUX2_X1 _10402_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02775_ ) );
MUX2_X1 _10403_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02776_ ) );
MUX2_X1 _10404_ ( .A(_02775_ ), .B(_02776_ ), .S(fanout_net_25 ), .Z(_02777_ ) );
OAI211_X1 _10405_ ( .A(fanout_net_27 ), .B(_02774_ ), .C1(_02777_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02778_ ) );
OAI211_X1 _10406_ ( .A(_02769_ ), .B(_02778_ ), .C1(_02379_ ), .C2(_02259_ ), .ZN(_02779_ ) );
NAND2_X1 _10407_ ( .A1(_02760_ ), .A2(_02779_ ), .ZN(_02780_ ) );
INV_X1 _10408_ ( .A(\ID_EX_imm [8] ), .ZN(_02781_ ) );
XNOR2_X1 _10409_ ( .A(_02780_ ), .B(_02781_ ), .ZN(_02782_ ) );
OR2_X1 _10410_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02783_ ) );
OAI211_X1 _10411_ ( .A(_02783_ ), .B(_02113_ ), .C1(_02163_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02784_ ) );
OR2_X1 _10412_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02785_ ) );
OAI211_X1 _10413_ ( .A(_02785_ ), .B(fanout_net_25 ), .C1(_02411_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02786_ ) );
NAND3_X1 _10414_ ( .A1(_02784_ ), .A2(_02786_ ), .A3(_02265_ ), .ZN(_02787_ ) );
MUX2_X1 _10415_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02788_ ) );
MUX2_X1 _10416_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02789_ ) );
MUX2_X1 _10417_ ( .A(_02788_ ), .B(_02789_ ), .S(_02184_ ), .Z(_02790_ ) );
OAI211_X1 _10418_ ( .A(fanout_net_27 ), .B(_02787_ ), .C1(_02790_ ), .C2(_02192_ ), .ZN(_02791_ ) );
MUX2_X1 _10419_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02792_ ) );
AND2_X1 _10420_ ( .A1(_02792_ ), .A2(fanout_net_25 ), .ZN(_02793_ ) );
MUX2_X1 _10421_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02794_ ) );
AOI211_X1 _10422_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_02793_ ), .C1(_02185_ ), .C2(_02794_ ), .ZN(_02795_ ) );
MUX2_X1 _10423_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02796_ ) );
MUX2_X1 _10424_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02797_ ) );
MUX2_X1 _10425_ ( .A(_02796_ ), .B(_02797_ ), .S(_02112_ ), .Z(_02798_ ) );
OAI21_X1 _10426_ ( .A(_02374_ ), .B1(_02798_ ), .B2(_02265_ ), .ZN(_02799_ ) );
OAI221_X1 _10427_ ( .A(_02791_ ), .B1(_02795_ ), .B2(_02799_ ), .C1(_02139_ ), .C2(_02180_ ), .ZN(_02800_ ) );
OR3_X1 _10428_ ( .A1(_02174_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02148_ ), .ZN(_02801_ ) );
NAND2_X2 _10429_ ( .A1(_02800_ ), .A2(_02801_ ), .ZN(_02802_ ) );
AND2_X1 _10430_ ( .A1(_02802_ ), .A2(\ID_EX_imm [9] ), .ZN(_02803_ ) );
INV_X1 _10431_ ( .A(_02803_ ), .ZN(_02804_ ) );
INV_X1 _10432_ ( .A(\ID_EX_imm [9] ), .ZN(_02805_ ) );
NAND3_X1 _10433_ ( .A1(_02800_ ), .A2(_02801_ ), .A3(_02805_ ), .ZN(_02806_ ) );
AND3_X1 _10434_ ( .A1(_02782_ ), .A2(_02804_ ), .A3(_02806_ ), .ZN(_02807_ ) );
OR3_X1 _10435_ ( .A1(_02138_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02147_ ), .ZN(_02808_ ) );
OR2_X1 _10436_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02809_ ) );
OAI211_X1 _10437_ ( .A(_02809_ ), .B(_02153_ ), .C1(_02158_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02810_ ) );
OR2_X1 _10438_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02811_ ) );
OAI211_X1 _10439_ ( .A(_02811_ ), .B(fanout_net_25 ), .C1(_02483_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02812_ ) );
NAND3_X1 _10440_ ( .A1(_02810_ ), .A2(_02812_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02813_ ) );
MUX2_X1 _10441_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02814_ ) );
MUX2_X1 _10442_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02815_ ) );
MUX2_X1 _10443_ ( .A(_02814_ ), .B(_02815_ ), .S(_02112_ ), .Z(_02816_ ) );
OAI211_X1 _10444_ ( .A(_02374_ ), .B(_02813_ ), .C1(_02816_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02817_ ) );
NOR2_X1 _10445_ ( .A1(_02157_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02818_ ) );
OAI21_X1 _10446_ ( .A(fanout_net_25 ), .B1(fanout_net_22 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02819_ ) );
NOR2_X1 _10447_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02820_ ) );
OAI21_X1 _10448_ ( .A(_02112_ ), .B1(_02483_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02821_ ) );
OAI221_X1 _10449_ ( .A(_02106_ ), .B1(_02818_ ), .B2(_02819_ ), .C1(_02820_ ), .C2(_02821_ ), .ZN(_02822_ ) );
MUX2_X1 _10450_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02823_ ) );
MUX2_X1 _10451_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02824_ ) );
MUX2_X1 _10452_ ( .A(_02823_ ), .B(_02824_ ), .S(fanout_net_25 ), .Z(_02825_ ) );
OAI211_X1 _10453_ ( .A(fanout_net_27 ), .B(_02822_ ), .C1(_02825_ ), .C2(_02265_ ), .ZN(_02826_ ) );
OAI211_X1 _10454_ ( .A(_02817_ ), .B(_02826_ ), .C1(_02174_ ), .C2(_02148_ ), .ZN(_02827_ ) );
NAND2_X1 _10455_ ( .A1(_02808_ ), .A2(_02827_ ), .ZN(_02828_ ) );
INV_X1 _10456_ ( .A(\ID_EX_imm [10] ), .ZN(_02829_ ) );
XNOR2_X1 _10457_ ( .A(_02828_ ), .B(_02829_ ), .ZN(_02830_ ) );
OR3_X1 _10458_ ( .A1(_02138_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_02147_ ), .ZN(_02831_ ) );
OR2_X1 _10459_ ( .A1(_02156_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02832_ ) );
OAI211_X1 _10460_ ( .A(_02832_ ), .B(_02153_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02833_ ) );
OR2_X1 _10461_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02834_ ) );
OAI211_X1 _10462_ ( .A(_02834_ ), .B(fanout_net_25 ), .C1(_02483_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02835_ ) );
NAND3_X1 _10463_ ( .A1(_02833_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02835_ ), .ZN(_02836_ ) );
MUX2_X1 _10464_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02837_ ) );
MUX2_X1 _10465_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02838_ ) );
MUX2_X1 _10466_ ( .A(_02837_ ), .B(_02838_ ), .S(_02112_ ), .Z(_02839_ ) );
OAI211_X1 _10467_ ( .A(_02103_ ), .B(_02836_ ), .C1(_02839_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02840_ ) );
NOR2_X1 _10468_ ( .A1(_02157_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02841_ ) );
OAI21_X1 _10469_ ( .A(fanout_net_25 ), .B1(fanout_net_22 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02842_ ) );
NOR2_X1 _10470_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02843_ ) );
OAI21_X1 _10471_ ( .A(_02112_ ), .B1(_02157_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02844_ ) );
OAI221_X1 _10472_ ( .A(_02106_ ), .B1(_02841_ ), .B2(_02842_ ), .C1(_02843_ ), .C2(_02844_ ), .ZN(_02845_ ) );
MUX2_X1 _10473_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02846_ ) );
MUX2_X1 _10474_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02847_ ) );
MUX2_X1 _10475_ ( .A(_02846_ ), .B(_02847_ ), .S(fanout_net_25 ), .Z(_02848_ ) );
OAI211_X1 _10476_ ( .A(fanout_net_27 ), .B(_02845_ ), .C1(_02848_ ), .C2(_02265_ ), .ZN(_02849_ ) );
OAI211_X1 _10477_ ( .A(_02840_ ), .B(_02849_ ), .C1(_02174_ ), .C2(_02148_ ), .ZN(_02850_ ) );
NAND2_X2 _10478_ ( .A1(_02831_ ), .A2(_02850_ ), .ZN(_02851_ ) );
INV_X1 _10479_ ( .A(\ID_EX_imm [11] ), .ZN(_02852_ ) );
XNOR2_X1 _10480_ ( .A(_02851_ ), .B(_02852_ ), .ZN(_02853_ ) );
AND2_X1 _10481_ ( .A1(_02830_ ), .A2(_02853_ ), .ZN(_02854_ ) );
AND2_X1 _10482_ ( .A1(_02807_ ), .A2(_02854_ ), .ZN(_02855_ ) );
AND3_X1 _10483_ ( .A1(_02662_ ), .A2(_02759_ ), .A3(_02855_ ), .ZN(_02856_ ) );
INV_X1 _10484_ ( .A(_02856_ ), .ZN(_02857_ ) );
XNOR2_X1 _10485_ ( .A(_02802_ ), .B(\ID_EX_imm [9] ), .ZN(_02858_ ) );
NAND2_X1 _10486_ ( .A1(_02780_ ), .A2(\ID_EX_imm [8] ), .ZN(_02859_ ) );
OAI21_X1 _10487_ ( .A(_02804_ ), .B1(_02858_ ), .B2(_02859_ ), .ZN(_02860_ ) );
AND2_X1 _10488_ ( .A1(_02854_ ), .A2(_02860_ ), .ZN(_02861_ ) );
AOI21_X1 _10489_ ( .A(_02852_ ), .B1(_02831_ ), .B2(_02850_ ), .ZN(_02862_ ) );
AND2_X1 _10490_ ( .A1(_02828_ ), .A2(\ID_EX_imm [10] ), .ZN(_02863_ ) );
AND2_X1 _10491_ ( .A1(_02853_ ), .A2(_02863_ ), .ZN(_02864_ ) );
NOR3_X1 _10492_ ( .A1(_02861_ ), .A2(_02862_ ), .A3(_02864_ ), .ZN(_02865_ ) );
INV_X1 _10493_ ( .A(_02865_ ), .ZN(_02866_ ) );
NAND2_X1 _10494_ ( .A1(_02866_ ), .A2(_02759_ ), .ZN(_02867_ ) );
OAI211_X1 _10495_ ( .A(\ID_EX_imm [14] ), .B(_02707_ ), .C1(_02683_ ), .C2(\ID_EX_imm [15] ), .ZN(_02868_ ) );
NAND2_X1 _10496_ ( .A1(_02731_ ), .A2(\ID_EX_imm [12] ), .ZN(_02869_ ) );
NOR3_X1 _10497_ ( .A1(_02869_ ), .A2(_02755_ ), .A3(_02756_ ), .ZN(_02870_ ) );
OR2_X1 _10498_ ( .A1(_02870_ ), .A2(_02756_ ), .ZN(_02871_ ) );
AOI22_X1 _10499_ ( .A1(_02871_ ), .A2(_02710_ ), .B1(\ID_EX_imm [15] ), .B2(_02683_ ), .ZN(_02872_ ) );
AND3_X1 _10500_ ( .A1(_02867_ ), .A2(_02868_ ), .A3(_02872_ ), .ZN(_02873_ ) );
AOI211_X1 _10501_ ( .A(_02358_ ), .B(_02457_ ), .C1(_02857_ ), .C2(_02873_ ), .ZN(_02874_ ) );
INV_X1 _10502_ ( .A(_02874_ ), .ZN(_02875_ ) );
AND2_X1 _10503_ ( .A1(_02454_ ), .A2(\ID_EX_imm [16] ), .ZN(_02876_ ) );
AND2_X1 _10504_ ( .A1(_02432_ ), .A2(_02876_ ), .ZN(_02877_ ) );
AOI21_X1 _10505_ ( .A(_02877_ ), .B1(\ID_EX_imm [17] ), .B2(_02430_ ), .ZN(_02878_ ) );
INV_X1 _10506_ ( .A(_02878_ ), .ZN(_02879_ ) );
AND2_X1 _10507_ ( .A1(_02879_ ), .A2(_02408_ ), .ZN(_02880_ ) );
AOI21_X1 _10508_ ( .A(_02383_ ), .B1(_02380_ ), .B2(_02381_ ), .ZN(_02881_ ) );
AND2_X1 _10509_ ( .A1(_02405_ ), .A2(\ID_EX_imm [18] ), .ZN(_02882_ ) );
AND2_X1 _10510_ ( .A1(_02384_ ), .A2(_02882_ ), .ZN(_02883_ ) );
NOR3_X1 _10511_ ( .A1(_02880_ ), .A2(_02881_ ), .A3(_02883_ ), .ZN(_02884_ ) );
NOR2_X1 _10512_ ( .A1(_02884_ ), .A2(_02358_ ), .ZN(_02885_ ) );
AND2_X1 _10513_ ( .A1(_02282_ ), .A2(\ID_EX_imm [23] ), .ZN(_02886_ ) );
NAND2_X1 _10514_ ( .A1(_02329_ ), .A2(\ID_EX_imm [20] ), .ZN(_02887_ ) );
NOR3_X1 _10515_ ( .A1(_02887_ ), .A2(_02353_ ), .A3(_02354_ ), .ZN(_02888_ ) );
OR2_X1 _10516_ ( .A1(_02888_ ), .A2(_02354_ ), .ZN(_02889_ ) );
AND2_X1 _10517_ ( .A1(_02889_ ), .A2(_02308_ ), .ZN(_02890_ ) );
AND2_X1 _10518_ ( .A1(_02305_ ), .A2(\ID_EX_imm [22] ), .ZN(_02891_ ) );
AND2_X1 _10519_ ( .A1(_02284_ ), .A2(_02891_ ), .ZN(_02892_ ) );
NOR4_X1 _10520_ ( .A1(_02885_ ), .A2(_02886_ ), .A3(_02890_ ), .A4(_02892_ ), .ZN(_02893_ ) );
NAND2_X1 _10521_ ( .A1(_02875_ ), .A2(_02893_ ), .ZN(_02894_ ) );
OR3_X1 _10522_ ( .A1(_02176_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02150_ ), .ZN(_02895_ ) );
OR2_X1 _10523_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02896_ ) );
OAI211_X1 _10524_ ( .A(_02896_ ), .B(_02115_ ), .C1(_02214_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02897_ ) );
OR2_X1 _10525_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02898_ ) );
OAI211_X1 _10526_ ( .A(_02898_ ), .B(fanout_net_25 ), .C1(_02214_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02899_ ) );
NAND3_X1 _10527_ ( .A1(_02897_ ), .A2(_02899_ ), .A3(_02118_ ), .ZN(_02900_ ) );
MUX2_X1 _10528_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02901_ ) );
MUX2_X1 _10529_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02902_ ) );
MUX2_X1 _10530_ ( .A(_02901_ ), .B(_02902_ ), .S(_02115_ ), .Z(_02903_ ) );
OAI211_X1 _10531_ ( .A(_02105_ ), .B(_02900_ ), .C1(_02903_ ), .C2(_02118_ ), .ZN(_02904_ ) );
OR2_X1 _10532_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02905_ ) );
OAI211_X1 _10533_ ( .A(_02905_ ), .B(_02115_ ), .C1(_02214_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02906_ ) );
NOR2_X1 _10534_ ( .A1(_02214_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02907_ ) );
OAI21_X1 _10535_ ( .A(fanout_net_25 ), .B1(fanout_net_22 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02908_ ) );
OAI211_X1 _10536_ ( .A(_02906_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_02907_ ), .C2(_02908_ ), .ZN(_02909_ ) );
MUX2_X1 _10537_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02910_ ) );
MUX2_X1 _10538_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02911_ ) );
MUX2_X1 _10539_ ( .A(_02910_ ), .B(_02911_ ), .S(fanout_net_25 ), .Z(_02912_ ) );
OAI211_X1 _10540_ ( .A(fanout_net_27 ), .B(_02909_ ), .C1(_02912_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02913_ ) );
OAI211_X1 _10541_ ( .A(_02904_ ), .B(_02913_ ), .C1(_02176_ ), .C2(_02150_ ), .ZN(_02914_ ) );
NAND2_X2 _10542_ ( .A1(_02895_ ), .A2(_02914_ ), .ZN(_02915_ ) );
INV_X1 _10543_ ( .A(\ID_EX_imm [24] ), .ZN(_02916_ ) );
XNOR2_X1 _10544_ ( .A(_02915_ ), .B(_02916_ ), .ZN(_02917_ ) );
OR3_X1 _10545_ ( .A1(_02140_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02181_ ), .ZN(_02918_ ) );
OR2_X1 _10546_ ( .A1(_02159_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02919_ ) );
OAI211_X1 _10547_ ( .A(_02919_ ), .B(fanout_net_25 ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02920_ ) );
OR2_X1 _10548_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02921_ ) );
OAI211_X1 _10549_ ( .A(_02921_ ), .B(_02186_ ), .C1(_02160_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02922_ ) );
NAND3_X1 _10550_ ( .A1(_02920_ ), .A2(_02193_ ), .A3(_02922_ ), .ZN(_02923_ ) );
MUX2_X1 _10551_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02924_ ) );
MUX2_X1 _10552_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02925_ ) );
MUX2_X1 _10553_ ( .A(_02924_ ), .B(_02925_ ), .S(_02155_ ), .Z(_02926_ ) );
OAI211_X1 _10554_ ( .A(_02105_ ), .B(_02923_ ), .C1(_02926_ ), .C2(_02118_ ), .ZN(_02927_ ) );
OR2_X1 _10555_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02928_ ) );
OAI211_X1 _10556_ ( .A(_02928_ ), .B(_02155_ ), .C1(_02160_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02929_ ) );
NOR2_X1 _10557_ ( .A1(_02188_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02930_ ) );
OAI21_X1 _10558_ ( .A(fanout_net_25 ), .B1(fanout_net_22 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02931_ ) );
OAI211_X1 _10559_ ( .A(_02929_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_02930_ ), .C2(_02931_ ), .ZN(_02932_ ) );
MUX2_X1 _10560_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02933_ ) );
MUX2_X1 _10561_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02934_ ) );
MUX2_X1 _10562_ ( .A(_02933_ ), .B(_02934_ ), .S(fanout_net_25 ), .Z(_02935_ ) );
OAI211_X1 _10563_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02932_ ), .C1(_02935_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02936_ ) );
OAI211_X1 _10564_ ( .A(_02927_ ), .B(_02936_ ), .C1(_02176_ ), .C2(_02150_ ), .ZN(_02937_ ) );
NAND2_X1 _10565_ ( .A1(_02918_ ), .A2(_02937_ ), .ZN(_02938_ ) );
INV_X1 _10566_ ( .A(\ID_EX_imm [25] ), .ZN(_02939_ ) );
XNOR2_X1 _10567_ ( .A(_02938_ ), .B(_02939_ ), .ZN(_02940_ ) );
AND3_X1 _10568_ ( .A1(_02894_ ), .A2(_02917_ ), .A3(_02940_ ), .ZN(_02941_ ) );
AND2_X1 _10569_ ( .A1(_02938_ ), .A2(\ID_EX_imm [25] ), .ZN(_02942_ ) );
AND3_X1 _10570_ ( .A1(_02918_ ), .A2(_02939_ ), .A3(_02937_ ), .ZN(_02943_ ) );
NAND2_X1 _10571_ ( .A1(_02915_ ), .A2(\ID_EX_imm [24] ), .ZN(_02944_ ) );
OR3_X1 _10572_ ( .A1(_02942_ ), .A2(_02943_ ), .A3(_02944_ ), .ZN(_02945_ ) );
INV_X1 _10573_ ( .A(_02938_ ), .ZN(_02946_ ) );
OAI21_X1 _10574_ ( .A(_02945_ ), .B1(_02939_ ), .B2(_02946_ ), .ZN(_02947_ ) );
OAI211_X1 _10575_ ( .A(_02235_ ), .B(_02258_ ), .C1(_02941_ ), .C2(_02947_ ), .ZN(_02948_ ) );
NAND2_X1 _10576_ ( .A1(_02256_ ), .A2(\ID_EX_imm [26] ), .ZN(_02949_ ) );
NOR3_X1 _10577_ ( .A1(_02949_ ), .A2(_02233_ ), .A3(_02234_ ), .ZN(_02950_ ) );
NOR2_X1 _10578_ ( .A1(_02950_ ), .A2(_02234_ ), .ZN(_02951_ ) );
AOI21_X1 _10579_ ( .A(_02210_ ), .B1(_02948_ ), .B2(_02951_ ), .ZN(_02952_ ) );
OR3_X1 _10580_ ( .A1(_02140_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02181_ ), .ZN(_02953_ ) );
OR2_X1 _10581_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02954_ ) );
OAI211_X1 _10582_ ( .A(_02954_ ), .B(_02115_ ), .C1(_02214_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02955_ ) );
OR2_X1 _10583_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02956_ ) );
OAI211_X1 _10584_ ( .A(_02956_ ), .B(fanout_net_25 ), .C1(_02188_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02957_ ) );
NAND3_X1 _10585_ ( .A1(_02955_ ), .A2(_02957_ ), .A3(_02193_ ), .ZN(_02958_ ) );
MUX2_X1 _10586_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02959_ ) );
MUX2_X1 _10587_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02960_ ) );
MUX2_X1 _10588_ ( .A(_02959_ ), .B(_02960_ ), .S(_02186_ ), .Z(_02961_ ) );
OAI211_X1 _10589_ ( .A(_02105_ ), .B(_02958_ ), .C1(_02961_ ), .C2(_02118_ ), .ZN(_02962_ ) );
OR2_X1 _10590_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02963_ ) );
OAI211_X1 _10591_ ( .A(_02963_ ), .B(fanout_net_25 ), .C1(_02188_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02964_ ) );
OR2_X1 _10592_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02965_ ) );
OAI211_X1 _10593_ ( .A(_02965_ ), .B(_02186_ ), .C1(_02188_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02966_ ) );
NAND3_X1 _10594_ ( .A1(_02964_ ), .A2(_02966_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02967_ ) );
MUX2_X1 _10595_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02968_ ) );
MUX2_X1 _10596_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02969_ ) );
MUX2_X1 _10597_ ( .A(_02968_ ), .B(_02969_ ), .S(fanout_net_25 ), .Z(_02970_ ) );
OAI211_X1 _10598_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02967_ ), .C1(_02970_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02971_ ) );
OAI211_X1 _10599_ ( .A(_02962_ ), .B(_02971_ ), .C1(_02176_ ), .C2(_02150_ ), .ZN(_02972_ ) );
NAND2_X2 _10600_ ( .A1(_02953_ ), .A2(_02972_ ), .ZN(_02973_ ) );
INV_X1 _10601_ ( .A(\ID_EX_imm [29] ), .ZN(_02974_ ) );
XNOR2_X1 _10602_ ( .A(_02973_ ), .B(_02974_ ), .ZN(_02975_ ) );
NAND2_X1 _10603_ ( .A1(_02952_ ), .A2(_02975_ ), .ZN(_02976_ ) );
AOI21_X1 _10604_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02182_ ), .B2(_02208_ ), .ZN(_02977_ ) );
INV_X1 _10605_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02978_ ) );
AOI22_X1 _10606_ ( .A1(_02975_ ), .A2(_02977_ ), .B1(_02978_ ), .B2(_02973_ ), .ZN(_02979_ ) );
AOI21_X1 _10607_ ( .A(_02179_ ), .B1(_02976_ ), .B2(_02979_ ), .ZN(_02980_ ) );
AOI21_X1 _10608_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02173_ ), .B2(_02177_ ), .ZN(_02981_ ) );
NOR2_X1 _10609_ ( .A1(_02980_ ), .A2(_02981_ ), .ZN(_02982_ ) );
NAND2_X1 _10610_ ( .A1(_02151_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_02983_ ) );
OR2_X1 _10611_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02984_ ) );
OAI211_X1 _10612_ ( .A(_02984_ ), .B(_02155_ ), .C1(_02160_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02985_ ) );
OR2_X1 _10613_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02986_ ) );
OAI211_X1 _10614_ ( .A(_02986_ ), .B(fanout_net_25 ), .C1(_02160_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02987_ ) );
NAND3_X1 _10615_ ( .A1(_02985_ ), .A2(_02987_ ), .A3(_02193_ ), .ZN(_02988_ ) );
MUX2_X1 _10616_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02989_ ) );
MUX2_X1 _10617_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02990_ ) );
MUX2_X1 _10618_ ( .A(_02989_ ), .B(_02990_ ), .S(_02155_ ), .Z(_02991_ ) );
OAI211_X1 _10619_ ( .A(_02105_ ), .B(_02988_ ), .C1(_02991_ ), .C2(_02193_ ), .ZN(_02992_ ) );
OR2_X1 _10620_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02993_ ) );
OAI211_X1 _10621_ ( .A(_02993_ ), .B(_02155_ ), .C1(_02160_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02994_ ) );
INV_X1 _10622_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02995_ ) );
NAND2_X1 _10623_ ( .A1(_02995_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .ZN(_02996_ ) );
OAI211_X1 _10624_ ( .A(_02996_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02997_ ) );
NAND3_X1 _10625_ ( .A1(_02994_ ), .A2(_02997_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02998_ ) );
MUX2_X1 _10626_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02999_ ) );
MUX2_X1 _10627_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03000_ ) );
MUX2_X1 _10628_ ( .A(_02999_ ), .B(_03000_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03001_ ) );
OAI211_X1 _10629_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02998_ ), .C1(_03001_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03002_ ) );
NAND2_X1 _10630_ ( .A1(_02992_ ), .A2(_03002_ ), .ZN(_03003_ ) );
OAI21_X1 _10631_ ( .A(_03003_ ), .B1(_02176_ ), .B2(_02150_ ), .ZN(_03004_ ) );
AND2_X1 _10632_ ( .A1(_02983_ ), .A2(_03004_ ), .ZN(_03005_ ) );
BUF_X4 _10633_ ( .A(_03005_ ), .Z(_03006_ ) );
XNOR2_X1 _10634_ ( .A(_03006_ ), .B(\ID_EX_imm [31] ), .ZN(_03007_ ) );
XNOR2_X1 _10635_ ( .A(_02982_ ), .B(_03007_ ), .ZN(_03008_ ) );
AND2_X2 _10636_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_03009_ ) );
BUF_X4 _10637_ ( .A(_03009_ ), .Z(_03010_ ) );
NOR2_X1 _10638_ ( .A1(_03008_ ), .A2(_03010_ ), .ZN(_00096_ ) );
NAND2_X1 _10639_ ( .A1(_02976_ ), .A2(_02979_ ), .ZN(_03011_ ) );
XNOR2_X1 _10640_ ( .A(_03011_ ), .B(_02179_ ), .ZN(_03012_ ) );
INV_X1 _10641_ ( .A(_03009_ ), .ZN(_03013_ ) );
CLKBUF_X2 _10642_ ( .A(_03013_ ), .Z(_03014_ ) );
AND2_X1 _10643_ ( .A1(_03012_ ), .A2(_03014_ ), .ZN(_00097_ ) );
AOI21_X1 _10644_ ( .A(_02457_ ), .B1(_02857_ ), .B2(_02873_ ), .ZN(_03015_ ) );
INV_X1 _10645_ ( .A(_02884_ ), .ZN(_03016_ ) );
OAI21_X1 _10646_ ( .A(_02331_ ), .B1(_03015_ ), .B2(_03016_ ), .ZN(_03017_ ) );
NAND2_X1 _10647_ ( .A1(_03017_ ), .A2(_02887_ ), .ZN(_03018_ ) );
XNOR2_X1 _10648_ ( .A(_03018_ ), .B(_02355_ ), .ZN(_03019_ ) );
NOR2_X1 _10649_ ( .A1(_03019_ ), .A2(_03010_ ), .ZN(_00098_ ) );
OR3_X1 _10650_ ( .A1(_03015_ ), .A2(_02331_ ), .A3(_03016_ ), .ZN(_03020_ ) );
AND3_X1 _10651_ ( .A1(_03020_ ), .A2(_03014_ ), .A3(_03017_ ), .ZN(_00099_ ) );
INV_X1 _10652_ ( .A(_02456_ ), .ZN(_03021_ ) );
AOI21_X1 _10653_ ( .A(_03021_ ), .B1(_02857_ ), .B2(_02873_ ), .ZN(_03022_ ) );
AND2_X1 _10654_ ( .A1(_03022_ ), .A2(_02432_ ), .ZN(_03023_ ) );
OAI21_X1 _10655_ ( .A(_02407_ ), .B1(_03023_ ), .B2(_02879_ ), .ZN(_03024_ ) );
INV_X1 _10656_ ( .A(_02882_ ), .ZN(_03025_ ) );
NAND2_X1 _10657_ ( .A1(_03024_ ), .A2(_03025_ ), .ZN(_03026_ ) );
XNOR2_X1 _10658_ ( .A(_03026_ ), .B(_02384_ ), .ZN(_03027_ ) );
NOR2_X1 _10659_ ( .A1(_03027_ ), .A2(_03010_ ), .ZN(_00100_ ) );
NOR2_X1 _10660_ ( .A1(_03023_ ), .A2(_02879_ ), .ZN(_03028_ ) );
XNOR2_X1 _10661_ ( .A(_03028_ ), .B(_02407_ ), .ZN(_03029_ ) );
AND2_X1 _10662_ ( .A1(_03029_ ), .A2(_03014_ ), .ZN(_00101_ ) );
OR2_X1 _10663_ ( .A1(_03022_ ), .A2(_02876_ ), .ZN(_03030_ ) );
XNOR2_X1 _10664_ ( .A(_03030_ ), .B(_02432_ ), .ZN(_03031_ ) );
NOR2_X1 _10665_ ( .A1(_03031_ ), .A2(_03010_ ), .ZN(_00102_ ) );
AND3_X1 _10666_ ( .A1(_02857_ ), .A2(_02873_ ), .A3(_03021_ ), .ZN(_03032_ ) );
NOR3_X1 _10667_ ( .A1(_03032_ ), .A2(_03022_ ), .A3(_03009_ ), .ZN(_00103_ ) );
INV_X1 _10668_ ( .A(_02758_ ), .ZN(_03033_ ) );
INV_X1 _10669_ ( .A(_02855_ ), .ZN(_03034_ ) );
AOI21_X1 _10670_ ( .A(_03034_ ), .B1(_02654_ ), .B2(_02661_ ), .ZN(_03035_ ) );
INV_X1 _10671_ ( .A(_03035_ ), .ZN(_03036_ ) );
AOI21_X1 _10672_ ( .A(_03033_ ), .B1(_03036_ ), .B2(_02865_ ), .ZN(_03037_ ) );
OR2_X1 _10673_ ( .A1(_03037_ ), .A2(_02871_ ), .ZN(_03038_ ) );
AND2_X1 _10674_ ( .A1(_03038_ ), .A2(_02709_ ), .ZN(_03039_ ) );
AND2_X1 _10675_ ( .A1(_02707_ ), .A2(\ID_EX_imm [14] ), .ZN(_03040_ ) );
OR2_X1 _10676_ ( .A1(_03039_ ), .A2(_03040_ ), .ZN(_03041_ ) );
XNOR2_X1 _10677_ ( .A(_03041_ ), .B(_02685_ ), .ZN(_03042_ ) );
NOR2_X1 _10678_ ( .A1(_03042_ ), .A2(_03010_ ), .ZN(_00104_ ) );
XOR2_X1 _10679_ ( .A(_03038_ ), .B(_02709_ ), .Z(_03043_ ) );
AND2_X1 _10680_ ( .A1(_03043_ ), .A2(_03014_ ), .ZN(_00105_ ) );
OAI21_X1 _10681_ ( .A(_02733_ ), .B1(_03035_ ), .B2(_02866_ ), .ZN(_03044_ ) );
NAND2_X1 _10682_ ( .A1(_03044_ ), .A2(_02869_ ), .ZN(_03045_ ) );
XNOR2_X1 _10683_ ( .A(_03045_ ), .B(_02757_ ), .ZN(_03046_ ) );
NOR2_X1 _10684_ ( .A1(_03046_ ), .A2(_03010_ ), .ZN(_00106_ ) );
OR3_X1 _10685_ ( .A1(_03035_ ), .A2(_02733_ ), .A3(_02866_ ), .ZN(_03047_ ) );
AND3_X1 _10686_ ( .A1(_03047_ ), .A2(_03014_ ), .A3(_03044_ ), .ZN(_00107_ ) );
OR2_X1 _10687_ ( .A1(_02952_ ), .A2(_02977_ ), .ZN(_03048_ ) );
XNOR2_X1 _10688_ ( .A(_03048_ ), .B(_02975_ ), .ZN(_03049_ ) );
NOR2_X1 _10689_ ( .A1(_03049_ ), .A2(_03010_ ), .ZN(_00108_ ) );
AND3_X1 _10690_ ( .A1(_02948_ ), .A2(_02951_ ), .A3(_02210_ ), .ZN(_03050_ ) );
NOR3_X1 _10691_ ( .A1(_03050_ ), .A2(_02952_ ), .A3(_03009_ ), .ZN(_00109_ ) );
OAI21_X1 _10692_ ( .A(_02258_ ), .B1(_02941_ ), .B2(_02947_ ), .ZN(_03051_ ) );
NAND2_X1 _10693_ ( .A1(_03051_ ), .A2(_02949_ ), .ZN(_03052_ ) );
XNOR2_X1 _10694_ ( .A(_03052_ ), .B(_02235_ ), .ZN(_03053_ ) );
NOR2_X1 _10695_ ( .A1(_03053_ ), .A2(_03010_ ), .ZN(_00110_ ) );
OR3_X1 _10696_ ( .A1(_02941_ ), .A2(_02258_ ), .A3(_02947_ ), .ZN(_03054_ ) );
AND3_X1 _10697_ ( .A1(_03054_ ), .A2(_03014_ ), .A3(_03051_ ), .ZN(_00111_ ) );
NAND2_X1 _10698_ ( .A1(_02894_ ), .A2(_02917_ ), .ZN(_03055_ ) );
NAND2_X1 _10699_ ( .A1(_03055_ ), .A2(_02944_ ), .ZN(_03056_ ) );
XNOR2_X1 _10700_ ( .A(_03056_ ), .B(_02940_ ), .ZN(_03057_ ) );
NOR2_X1 _10701_ ( .A1(_03057_ ), .A2(_03010_ ), .ZN(_00112_ ) );
XOR2_X1 _10702_ ( .A(_02894_ ), .B(_02917_ ), .Z(_03058_ ) );
AND2_X1 _10703_ ( .A1(_03058_ ), .A2(_03014_ ), .ZN(_00113_ ) );
OAI21_X1 _10704_ ( .A(_02356_ ), .B1(_03015_ ), .B2(_03016_ ), .ZN(_03059_ ) );
INV_X1 _10705_ ( .A(_03059_ ), .ZN(_03060_ ) );
OR2_X1 _10706_ ( .A1(_03060_ ), .A2(_02889_ ), .ZN(_03061_ ) );
AND2_X1 _10707_ ( .A1(_03061_ ), .A2(_02307_ ), .ZN(_03062_ ) );
OR2_X1 _10708_ ( .A1(_03062_ ), .A2(_02891_ ), .ZN(_03063_ ) );
XNOR2_X1 _10709_ ( .A(_03063_ ), .B(_02284_ ), .ZN(_03064_ ) );
NOR2_X1 _10710_ ( .A1(_03064_ ), .A2(_03010_ ), .ZN(_00114_ ) );
XOR2_X1 _10711_ ( .A(_03061_ ), .B(_02307_ ), .Z(_03065_ ) );
AND2_X1 _10712_ ( .A1(_03065_ ), .A2(_03014_ ), .ZN(_00115_ ) );
INV_X1 _10713_ ( .A(\IF_ID_inst [31] ), .ZN(_03066_ ) );
NOR2_X1 _10714_ ( .A1(fanout_net_2 ), .A2(excp_written ), .ZN(_03067_ ) );
AND2_X1 _10715_ ( .A1(_02094_ ), .A2(_03067_ ), .ZN(_03068_ ) );
INV_X2 _10716_ ( .A(_03068_ ), .ZN(_03069_ ) );
BUF_X4 _10717_ ( .A(_03069_ ), .Z(_03070_ ) );
AND2_X1 _10718_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_03071_ ) );
NOR2_X1 _10719_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_03072_ ) );
AND2_X1 _10720_ ( .A1(_03071_ ), .A2(_03072_ ), .ZN(_03073_ ) );
CLKBUF_X2 _10721_ ( .A(_03073_ ), .Z(_03074_ ) );
BUF_X2 _10722_ ( .A(_03074_ ), .Z(_03075_ ) );
AND4_X1 _10723_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03076_ ) );
AND2_X1 _10724_ ( .A1(_03075_ ), .A2(_03076_ ), .ZN(_03077_ ) );
INV_X1 _10725_ ( .A(_03077_ ), .ZN(_03078_ ) );
INV_X1 _10726_ ( .A(\IF_ID_inst [6] ), .ZN(_03079_ ) );
NOR2_X1 _10727_ ( .A1(_03079_ ), .A2(\IF_ID_inst [12] ), .ZN(_03080_ ) );
AND2_X1 _10728_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03081_ ) );
AND3_X1 _10729_ ( .A1(_03080_ ), .A2(\IF_ID_inst [13] ), .A3(_03081_ ), .ZN(_03082_ ) );
NAND2_X2 _10730_ ( .A1(_03082_ ), .A2(_03075_ ), .ZN(_03083_ ) );
AOI211_X1 _10731_ ( .A(_03066_ ), .B(_03070_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00194_ ) );
INV_X1 _10732_ ( .A(\IF_ID_inst [30] ), .ZN(_03084_ ) );
AOI211_X1 _10733_ ( .A(_03084_ ), .B(_03070_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00195_ ) );
INV_X1 _10734_ ( .A(\IF_ID_inst [21] ), .ZN(_03085_ ) );
AOI211_X1 _10735_ ( .A(_03085_ ), .B(_03070_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00196_ ) );
BUF_X4 _10736_ ( .A(_03069_ ), .Z(_03086_ ) );
AND2_X2 _10737_ ( .A1(_03078_ ), .A2(_03083_ ), .ZN(_03087_ ) );
INV_X1 _10738_ ( .A(_03087_ ), .ZN(_03088_ ) );
INV_X1 _10739_ ( .A(\IF_ID_inst [20] ), .ZN(_03089_ ) );
AOI21_X1 _10740_ ( .A(_03086_ ), .B1(_03088_ ), .B2(_03089_ ), .ZN(_00197_ ) );
INV_X1 _10741_ ( .A(\IF_ID_inst [29] ), .ZN(_03090_ ) );
AOI21_X1 _10742_ ( .A(_03086_ ), .B1(_03088_ ), .B2(_03090_ ), .ZN(_00198_ ) );
INV_X1 _10743_ ( .A(\IF_ID_inst [28] ), .ZN(_03091_ ) );
AOI21_X1 _10744_ ( .A(_03086_ ), .B1(_03088_ ), .B2(_03091_ ), .ZN(_00199_ ) );
INV_X1 _10745_ ( .A(\IF_ID_inst [27] ), .ZN(_03092_ ) );
AOI211_X1 _10746_ ( .A(_03092_ ), .B(_03070_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00200_ ) );
INV_X1 _10747_ ( .A(\IF_ID_inst [26] ), .ZN(_03093_ ) );
AOI21_X1 _10748_ ( .A(_03086_ ), .B1(_03088_ ), .B2(_03093_ ), .ZN(_00201_ ) );
INV_X1 _10749_ ( .A(\IF_ID_inst [25] ), .ZN(_03094_ ) );
BUF_X4 _10750_ ( .A(_03069_ ), .Z(_03095_ ) );
AOI211_X1 _10751_ ( .A(_03094_ ), .B(_03095_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00202_ ) );
INV_X1 _10752_ ( .A(\IF_ID_inst [24] ), .ZN(_03096_ ) );
AOI211_X1 _10753_ ( .A(_03096_ ), .B(_03095_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00203_ ) );
INV_X1 _10754_ ( .A(\IF_ID_inst [23] ), .ZN(_03097_ ) );
AOI211_X1 _10755_ ( .A(_03097_ ), .B(_03095_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00204_ ) );
INV_X1 _10756_ ( .A(\IF_ID_inst [22] ), .ZN(_03098_ ) );
AOI211_X1 _10757_ ( .A(_03098_ ), .B(_03095_ ), .C1(_03078_ ), .C2(_03083_ ), .ZN(_00205_ ) );
CLKBUF_X2 _10758_ ( .A(_03067_ ), .Z(_03099_ ) );
CLKBUF_X2 _10759_ ( .A(_03099_ ), .Z(_03100_ ) );
AND3_X1 _10760_ ( .A1(_02094_ ), .A2(_03100_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00206_ ) );
AND3_X1 _10761_ ( .A1(_02094_ ), .A2(_03067_ ), .A3(\myidu.state [2] ), .ZN(_00207_ ) );
INV_X1 _10762_ ( .A(\IF_ID_inst [5] ), .ZN(_03101_ ) );
NOR2_X1 _10763_ ( .A1(_03101_ ), .A2(\IF_ID_inst [4] ), .ZN(_03102_ ) );
AND2_X1 _10764_ ( .A1(_03080_ ), .A2(_03102_ ), .ZN(_03103_ ) );
AND2_X1 _10765_ ( .A1(_03103_ ), .A2(_03074_ ), .ZN(_03104_ ) );
NAND2_X1 _10766_ ( .A1(_03104_ ), .A2(\IF_ID_inst [14] ), .ZN(_03105_ ) );
INV_X1 _10767_ ( .A(\IF_ID_inst [12] ), .ZN(_03106_ ) );
NOR2_X1 _10768_ ( .A1(_03106_ ), .A2(\IF_ID_inst [6] ), .ZN(_03107_ ) );
NOR2_X1 _10769_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03108_ ) );
NOR2_X1 _10770_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03109_ ) );
AND3_X1 _10771_ ( .A1(_03107_ ), .A2(_03108_ ), .A3(_03109_ ), .ZN(_03110_ ) );
AND3_X1 _10772_ ( .A1(_03071_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_03111_ ) );
AND2_X1 _10773_ ( .A1(_03110_ ), .A2(_03111_ ), .ZN(_03112_ ) );
INV_X1 _10774_ ( .A(\IF_ID_inst [11] ), .ZN(_03113_ ) );
INV_X1 _10775_ ( .A(\IF_ID_inst [10] ), .ZN(_03114_ ) );
NOR2_X1 _10776_ ( .A1(\IF_ID_inst [9] ), .A2(\IF_ID_inst [8] ), .ZN(_03115_ ) );
AND4_X1 _10777_ ( .A1(_03113_ ), .A2(_03075_ ), .A3(_03114_ ), .A4(_03115_ ), .ZN(_03116_ ) );
INV_X1 _10778_ ( .A(\IF_ID_inst [7] ), .ZN(_03117_ ) );
INV_X1 _10779_ ( .A(\IF_ID_inst [14] ), .ZN(_03118_ ) );
INV_X1 _10780_ ( .A(\IF_ID_inst [13] ), .ZN(_03119_ ) );
AND4_X1 _10781_ ( .A1(_03118_ ), .A2(_03119_ ), .A3(\IF_ID_inst [4] ), .A4(\IF_ID_inst [5] ), .ZN(_03120_ ) );
INV_X1 _10782_ ( .A(\IF_ID_inst [15] ), .ZN(_03121_ ) );
AND4_X1 _10783_ ( .A1(_03117_ ), .A2(_03120_ ), .A3(_03121_ ), .A4(_03080_ ), .ZN(_03122_ ) );
AND2_X1 _10784_ ( .A1(_03116_ ), .A2(_03122_ ), .ZN(_03123_ ) );
NAND4_X1 _10785_ ( .A1(_03089_ ), .A2(_03097_ ), .A3(_03098_ ), .A4(\IF_ID_inst [29] ), .ZN(_03124_ ) );
NAND4_X1 _10786_ ( .A1(_03084_ ), .A2(_03066_ ), .A3(\IF_ID_inst [21] ), .A4(\IF_ID_inst [28] ), .ZN(_03125_ ) );
NOR2_X1 _10787_ ( .A1(_03124_ ), .A2(_03125_ ), .ZN(_03126_ ) );
NAND3_X1 _10788_ ( .A1(_03093_ ), .A2(_03094_ ), .A3(_03096_ ), .ZN(_03127_ ) );
NOR2_X1 _10789_ ( .A1(_03127_ ), .A2(\IF_ID_inst [27] ), .ZN(_03128_ ) );
NOR2_X1 _10790_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [18] ), .ZN(_03129_ ) );
NOR2_X1 _10791_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_03130_ ) );
AND2_X1 _10792_ ( .A1(_03129_ ), .A2(_03130_ ), .ZN(_03131_ ) );
AND3_X1 _10793_ ( .A1(_03126_ ), .A2(_03128_ ), .A3(_03131_ ), .ZN(_03132_ ) );
AOI221_X4 _10794_ ( .A(_03112_ ), .B1(_03108_ ), .B2(_03104_ ), .C1(_03123_ ), .C2(_03132_ ), .ZN(_03133_ ) );
AND3_X1 _10795_ ( .A1(_03074_ ), .A2(\IF_ID_inst [12] ), .A3(\IF_ID_inst [6] ), .ZN(_03134_ ) );
NAND3_X1 _10796_ ( .A1(_03134_ ), .A2(_03119_ ), .A3(_03102_ ), .ZN(_03135_ ) );
NOR4_X1 _10797_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .A4(\IF_ID_inst [31] ), .ZN(_03136_ ) );
AND2_X1 _10798_ ( .A1(_03128_ ), .A2(_03136_ ), .ZN(_03137_ ) );
AND3_X1 _10799_ ( .A1(_03116_ ), .A2(_03122_ ), .A3(_03137_ ), .ZN(_03138_ ) );
AND3_X1 _10800_ ( .A1(_03131_ ), .A2(_03097_ ), .A3(_03098_ ), .ZN(_03139_ ) );
AND3_X1 _10801_ ( .A1(_03139_ ), .A2(_03085_ ), .A3(\IF_ID_inst [20] ), .ZN(_03140_ ) );
AND2_X1 _10802_ ( .A1(_03134_ ), .A2(_03102_ ), .ZN(_03141_ ) );
AND2_X2 _10803_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03142_ ) );
AOI22_X1 _10804_ ( .A1(_03138_ ), .A2(_03140_ ), .B1(_03141_ ), .B2(_03142_ ), .ZN(_03143_ ) );
AND4_X1 _10805_ ( .A1(_03105_ ), .A2(_03133_ ), .A3(_03135_ ), .A4(_03143_ ), .ZN(_03144_ ) );
CLKBUF_X2 _10806_ ( .A(_03068_ ), .Z(_03145_ ) );
NOR2_X1 _10807_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03146_ ) );
AND3_X1 _10808_ ( .A1(_03074_ ), .A2(_03102_ ), .A3(_03146_ ), .ZN(_03147_ ) );
NOR2_X1 _10809_ ( .A1(_03119_ ), .A2(\IF_ID_inst [14] ), .ZN(_03148_ ) );
AND2_X1 _10810_ ( .A1(_03147_ ), .A2(_03148_ ), .ZN(_03149_ ) );
INV_X1 _10811_ ( .A(_03149_ ), .ZN(_03150_ ) );
AND3_X1 _10812_ ( .A1(_03074_ ), .A2(_03102_ ), .A3(_03107_ ), .ZN(_03151_ ) );
OAI21_X1 _10813_ ( .A(_03108_ ), .B1(_03147_ ), .B2(_03151_ ), .ZN(_03152_ ) );
AND2_X2 _10814_ ( .A1(_03150_ ), .A2(_03152_ ), .ZN(_03153_ ) );
AND4_X1 _10815_ ( .A1(\IF_ID_inst [11] ), .A2(_03144_ ), .A3(_03145_ ), .A4(_03153_ ), .ZN(_00208_ ) );
AND4_X1 _10816_ ( .A1(\IF_ID_inst [10] ), .A2(_03144_ ), .A3(_03145_ ), .A4(_03153_ ), .ZN(_00209_ ) );
AND4_X1 _10817_ ( .A1(\IF_ID_inst [9] ), .A2(_03144_ ), .A3(_03145_ ), .A4(_03153_ ), .ZN(_00210_ ) );
AND4_X1 _10818_ ( .A1(\IF_ID_inst [8] ), .A2(_03144_ ), .A3(_03145_ ), .A4(_03153_ ), .ZN(_00211_ ) );
AND4_X1 _10819_ ( .A1(\IF_ID_inst [7] ), .A2(_03144_ ), .A3(_03145_ ), .A4(_03153_ ), .ZN(_00212_ ) );
NOR4_X1 _10820_ ( .A1(_03124_ ), .A2(_03125_ ), .A3(_03127_ ), .A4(\IF_ID_inst [27] ), .ZN(_03154_ ) );
AND3_X1 _10821_ ( .A1(_03116_ ), .A2(_03122_ ), .A3(_03154_ ), .ZN(_03155_ ) );
AND2_X1 _10822_ ( .A1(_03155_ ), .A2(_03131_ ), .ZN(_03156_ ) );
INV_X1 _10823_ ( .A(_03156_ ), .ZN(_03157_ ) );
INV_X1 _10824_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03158_ ) );
AND2_X1 _10825_ ( .A1(_03102_ ), .A2(_03158_ ), .ZN(_03159_ ) );
AND2_X2 _10826_ ( .A1(_03159_ ), .A2(_03111_ ), .ZN(_03160_ ) );
BUF_X2 _10827_ ( .A(_03160_ ), .Z(_03161_ ) );
BUF_X2 _10828_ ( .A(_03161_ ), .Z(_03162_ ) );
NAND3_X1 _10829_ ( .A1(\IF_ID_inst [2] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [1] ), .ZN(_03163_ ) );
NOR2_X1 _10830_ ( .A1(_03163_ ), .A2(\IF_ID_inst [3] ), .ZN(_03164_ ) );
INV_X1 _10831_ ( .A(\IF_ID_inst [4] ), .ZN(_03165_ ) );
NOR2_X1 _10832_ ( .A1(_03165_ ), .A2(\IF_ID_inst [6] ), .ZN(_03166_ ) );
AND2_X1 _10833_ ( .A1(_03164_ ), .A2(_03166_ ), .ZN(_03167_ ) );
NOR2_X2 _10834_ ( .A1(_03162_ ), .A2(_03167_ ), .ZN(_03168_ ) );
NAND2_X1 _10835_ ( .A1(_03157_ ), .A2(_03168_ ), .ZN(_03169_ ) );
INV_X1 _10836_ ( .A(\IF_ID_inst [19] ), .ZN(_03170_ ) );
AND3_X1 _10837_ ( .A1(_03109_ ), .A2(\IF_ID_inst [12] ), .A3(_03079_ ), .ZN(_03171_ ) );
AND2_X1 _10838_ ( .A1(_03111_ ), .A2(_03171_ ), .ZN(_03172_ ) );
NAND2_X1 _10839_ ( .A1(_03172_ ), .A2(_03108_ ), .ZN(_03173_ ) );
CLKBUF_X2 _10840_ ( .A(_03081_ ), .Z(_03174_ ) );
AND4_X1 _10841_ ( .A1(\IF_ID_inst [6] ), .A2(_03075_ ), .A3(_03117_ ), .A4(_03174_ ), .ZN(_03175_ ) );
AND3_X1 _10842_ ( .A1(_03115_ ), .A2(_03113_ ), .A3(_03114_ ), .ZN(_03176_ ) );
NOR4_X1 _10843_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_03177_ ) );
NAND3_X1 _10844_ ( .A1(_03175_ ), .A2(_03176_ ), .A3(_03177_ ), .ZN(_03178_ ) );
NAND4_X1 _10845_ ( .A1(_03137_ ), .A2(_03139_ ), .A3(_03085_ ), .A4(\IF_ID_inst [20] ), .ZN(_03179_ ) );
OAI21_X1 _10846_ ( .A(_03173_ ), .B1(_03178_ ), .B2(_03179_ ), .ZN(_03180_ ) );
NOR4_X1 _10847_ ( .A1(_03169_ ), .A2(_03170_ ), .A3(_03095_ ), .A4(_03180_ ), .ZN(_00213_ ) );
INV_X1 _10848_ ( .A(\IF_ID_inst [18] ), .ZN(_03181_ ) );
NOR4_X1 _10849_ ( .A1(_03169_ ), .A2(_03181_ ), .A3(_03095_ ), .A4(_03180_ ), .ZN(_00214_ ) );
INV_X1 _10850_ ( .A(\IF_ID_inst [17] ), .ZN(_03182_ ) );
NOR4_X1 _10851_ ( .A1(_03169_ ), .A2(_03182_ ), .A3(_03095_ ), .A4(_03180_ ), .ZN(_00215_ ) );
XNOR2_X1 _10852_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_03183_ ) );
XNOR2_X1 _10853_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_03184_ ) );
XNOR2_X1 _10854_ ( .A(fanout_net_7 ), .B(\myexu.pc_jump [3] ), .ZN(_03185_ ) );
XNOR2_X1 _10855_ ( .A(\myexu.pc_jump [2] ), .B(\IF_ID_pc [2] ), .ZN(_03186_ ) );
AND4_X1 _10856_ ( .A1(_03183_ ), .A2(_03184_ ), .A3(_03185_ ), .A4(_03186_ ), .ZN(_03187_ ) );
XNOR2_X1 _10857_ ( .A(fanout_net_11 ), .B(\myexu.pc_jump [4] ), .ZN(_03188_ ) );
XNOR2_X1 _10858_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_03189_ ) );
XNOR2_X1 _10859_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_03190_ ) );
XNOR2_X1 _10860_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_03191_ ) );
AND4_X1 _10861_ ( .A1(_03188_ ), .A2(_03189_ ), .A3(_03190_ ), .A4(_03191_ ), .ZN(_03192_ ) );
XNOR2_X1 _10862_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_03193_ ) );
XNOR2_X1 _10863_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_03194_ ) );
XNOR2_X1 _10864_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_03195_ ) );
XNOR2_X1 _10865_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_03196_ ) );
AND4_X1 _10866_ ( .A1(_03193_ ), .A2(_03194_ ), .A3(_03195_ ), .A4(_03196_ ), .ZN(_03197_ ) );
XNOR2_X1 _10867_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_03198_ ) );
XNOR2_X1 _10868_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_03199_ ) );
XNOR2_X1 _10869_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_03200_ ) );
XNOR2_X1 _10870_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_03201_ ) );
AND4_X1 _10871_ ( .A1(_03198_ ), .A2(_03199_ ), .A3(_03200_ ), .A4(_03201_ ), .ZN(_03202_ ) );
AND4_X1 _10872_ ( .A1(_03187_ ), .A2(_03192_ ), .A3(_03197_ ), .A4(_03202_ ), .ZN(_03203_ ) );
XNOR2_X1 _10873_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_03204_ ) );
XNOR2_X1 _10874_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_03205_ ) );
XNOR2_X1 _10875_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_03206_ ) );
XNOR2_X1 _10876_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_03207_ ) );
AND4_X1 _10877_ ( .A1(_03204_ ), .A2(_03205_ ), .A3(_03206_ ), .A4(_03207_ ), .ZN(_03208_ ) );
XNOR2_X1 _10878_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_03209_ ) );
XNOR2_X1 _10879_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_03210_ ) );
XNOR2_X1 _10880_ ( .A(\IF_ID_pc [25] ), .B(\myexu.pc_jump [25] ), .ZN(_03211_ ) );
XNOR2_X1 _10881_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_03212_ ) );
AND4_X1 _10882_ ( .A1(_03209_ ), .A2(_03210_ ), .A3(_03211_ ), .A4(_03212_ ), .ZN(_03213_ ) );
XNOR2_X1 _10883_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_03214_ ) );
XNOR2_X1 _10884_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_03215_ ) );
XNOR2_X1 _10885_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_03216_ ) );
XNOR2_X1 _10886_ ( .A(\IF_ID_pc [21] ), .B(\myexu.pc_jump [21] ), .ZN(_03217_ ) );
AND4_X1 _10887_ ( .A1(_03214_ ), .A2(_03215_ ), .A3(_03216_ ), .A4(_03217_ ), .ZN(_03218_ ) );
XNOR2_X1 _10888_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_03219_ ) );
XNOR2_X1 _10889_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_03220_ ) );
XNOR2_X1 _10890_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_03221_ ) );
XNOR2_X1 _10891_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_03222_ ) );
AND4_X1 _10892_ ( .A1(_03219_ ), .A2(_03220_ ), .A3(_03221_ ), .A4(_03222_ ), .ZN(_03223_ ) );
AND4_X1 _10893_ ( .A1(_03208_ ), .A2(_03213_ ), .A3(_03218_ ), .A4(_03223_ ), .ZN(_03224_ ) );
AND2_X1 _10894_ ( .A1(_03203_ ), .A2(_03224_ ), .ZN(_03225_ ) );
INV_X1 _10895_ ( .A(check_quest ), .ZN(_03226_ ) );
NOR2_X2 _10896_ ( .A1(_03225_ ), .A2(_03226_ ), .ZN(_03227_ ) );
INV_X1 _10897_ ( .A(\myifu.state [1] ), .ZN(_03228_ ) );
NOR2_X1 _10898_ ( .A1(_03228_ ), .A2(\myifu.to_reset ), .ZN(_03229_ ) );
INV_X1 _10899_ ( .A(_03229_ ), .ZN(_03230_ ) );
NOR2_X1 _10900_ ( .A1(_03227_ ), .A2(_03230_ ), .ZN(_03231_ ) );
AND2_X1 _10901_ ( .A1(_03231_ ), .A2(IDU_ready_IFU ), .ZN(_03232_ ) );
INV_X1 _10902_ ( .A(_03232_ ), .ZN(_03233_ ) );
BUF_X4 _10903_ ( .A(_03233_ ), .Z(_03234_ ) );
AND2_X2 _10904_ ( .A1(_03075_ ), .A2(_03107_ ), .ZN(_03235_ ) );
NOR2_X1 _10905_ ( .A1(_03165_ ), .A2(\IF_ID_inst [5] ), .ZN(_03236_ ) );
AND2_X1 _10906_ ( .A1(_03235_ ), .A2(_03236_ ), .ZN(_03237_ ) );
NOR3_X1 _10907_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_03238_ ) );
AND3_X1 _10908_ ( .A1(_03238_ ), .A2(_03092_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03239_ ) );
NOR2_X1 _10909_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_03240_ ) );
AND2_X1 _10910_ ( .A1(_03108_ ), .A2(_03240_ ), .ZN(_03241_ ) );
AND2_X1 _10911_ ( .A1(_03239_ ), .A2(_03241_ ), .ZN(_03242_ ) );
NOR2_X1 _10912_ ( .A1(_03084_ ), .A2(\IF_ID_inst [29] ), .ZN(_03243_ ) );
NOR2_X1 _10913_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_03244_ ) );
AND3_X1 _10914_ ( .A1(_03243_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_03244_ ), .ZN(_03245_ ) );
NOR2_X1 _10915_ ( .A1(_03118_ ), .A2(\IF_ID_inst [13] ), .ZN(_03246_ ) );
AND2_X1 _10916_ ( .A1(_03246_ ), .A2(_03240_ ), .ZN(_03247_ ) );
AND2_X1 _10917_ ( .A1(_03245_ ), .A2(_03247_ ), .ZN(_03248_ ) );
NOR2_X1 _10918_ ( .A1(_03242_ ), .A2(_03248_ ), .ZN(_03249_ ) );
INV_X1 _10919_ ( .A(_03249_ ), .ZN(_03250_ ) );
AND2_X1 _10920_ ( .A1(_03239_ ), .A2(_03247_ ), .ZN(_03251_ ) );
OAI21_X1 _10921_ ( .A(_03237_ ), .B1(_03250_ ), .B2(_03251_ ), .ZN(_03252_ ) );
AND2_X2 _10922_ ( .A1(_03238_ ), .A2(_03092_ ), .ZN(_03253_ ) );
INV_X1 _10923_ ( .A(_03253_ ), .ZN(_03254_ ) );
NAND4_X1 _10924_ ( .A1(_03240_ ), .A2(_03118_ ), .A3(\IF_ID_inst [13] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03255_ ) );
NOR2_X1 _10925_ ( .A1(_03254_ ), .A2(_03255_ ), .ZN(_03256_ ) );
AND2_X2 _10926_ ( .A1(_03074_ ), .A2(_03146_ ), .ZN(_03257_ ) );
NAND3_X1 _10927_ ( .A1(_03256_ ), .A2(_03174_ ), .A3(_03257_ ), .ZN(_03258_ ) );
NAND4_X1 _10928_ ( .A1(_03257_ ), .A2(_03081_ ), .A3(_03241_ ), .A4(_03245_ ), .ZN(_03259_ ) );
AND2_X1 _10929_ ( .A1(_03258_ ), .A2(_03259_ ), .ZN(_03260_ ) );
NAND2_X1 _10930_ ( .A1(_03252_ ), .A2(_03260_ ), .ZN(_03261_ ) );
OR2_X1 _10931_ ( .A1(_03141_ ), .A2(_03104_ ), .ZN(_03262_ ) );
INV_X1 _10932_ ( .A(_03148_ ), .ZN(_03263_ ) );
AND2_X2 _10933_ ( .A1(_03262_ ), .A2(_03263_ ), .ZN(_03264_ ) );
INV_X1 _10934_ ( .A(_03153_ ), .ZN(_03265_ ) );
NOR3_X1 _10935_ ( .A1(_03261_ ), .A2(_03264_ ), .A3(_03265_ ), .ZN(_03266_ ) );
AND3_X1 _10936_ ( .A1(_03081_ ), .A2(_03071_ ), .A3(_03072_ ), .ZN(_03267_ ) );
NAND4_X1 _10937_ ( .A1(_03238_ ), .A2(_03092_ ), .A3(_03142_ ), .A4(_03240_ ), .ZN(_03268_ ) );
INV_X1 _10938_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03269_ ) );
NOR2_X1 _10939_ ( .A1(_03268_ ), .A2(_03269_ ), .ZN(_03270_ ) );
OAI211_X1 _10940_ ( .A(_03079_ ), .B(_03267_ ), .C1(_03270_ ), .C2(_03106_ ), .ZN(_03271_ ) );
INV_X1 _10941_ ( .A(_03270_ ), .ZN(_03272_ ) );
OAI211_X1 _10942_ ( .A(_03253_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .C1(_03247_ ), .C2(_03241_ ), .ZN(_03273_ ) );
AOI21_X1 _10943_ ( .A(_03271_ ), .B1(_03272_ ), .B2(_03273_ ), .ZN(_03274_ ) );
AND2_X1 _10944_ ( .A1(_03267_ ), .A2(_03107_ ), .ZN(_03275_ ) );
AND4_X1 _10945_ ( .A1(\IF_ID_inst [14] ), .A2(_03240_ ), .A3(_03119_ ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03276_ ) );
AND2_X1 _10946_ ( .A1(_03253_ ), .A2(_03276_ ), .ZN(_03277_ ) );
OAI21_X1 _10947_ ( .A(_03275_ ), .B1(_03256_ ), .B2(_03277_ ), .ZN(_03278_ ) );
INV_X1 _10948_ ( .A(_03278_ ), .ZN(_03279_ ) );
AND3_X1 _10949_ ( .A1(_03253_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_03241_ ), .ZN(_03280_ ) );
OAI21_X1 _10950_ ( .A(_03275_ ), .B1(_03280_ ), .B2(_03248_ ), .ZN(_03281_ ) );
INV_X1 _10951_ ( .A(_03281_ ), .ZN(_03282_ ) );
NOR3_X1 _10952_ ( .A1(_03274_ ), .A2(_03279_ ), .A3(_03282_ ), .ZN(_03283_ ) );
AND2_X1 _10953_ ( .A1(_03266_ ), .A2(_03283_ ), .ZN(_03284_ ) );
AND2_X1 _10954_ ( .A1(_03257_ ), .A2(_03236_ ), .ZN(_03285_ ) );
AND2_X1 _10955_ ( .A1(_03285_ ), .A2(_03148_ ), .ZN(_03286_ ) );
NAND3_X1 _10956_ ( .A1(_03235_ ), .A2(\IF_ID_inst [13] ), .A3(_03236_ ), .ZN(_03287_ ) );
NOR2_X1 _10957_ ( .A1(_03287_ ), .A2(\IF_ID_inst [14] ), .ZN(_03288_ ) );
NOR2_X1 _10958_ ( .A1(_03286_ ), .A2(_03288_ ), .ZN(_03289_ ) );
AND2_X1 _10959_ ( .A1(_03171_ ), .A2(_03075_ ), .ZN(_03290_ ) );
NAND2_X1 _10960_ ( .A1(_03290_ ), .A2(_03119_ ), .ZN(_03291_ ) );
AND3_X1 _10961_ ( .A1(_03103_ ), .A2(_03108_ ), .A3(_03164_ ), .ZN(_03292_ ) );
INV_X1 _10962_ ( .A(_03292_ ), .ZN(_03293_ ) );
INV_X1 _10963_ ( .A(_03142_ ), .ZN(_03294_ ) );
NAND3_X1 _10964_ ( .A1(_03257_ ), .A2(_03294_ ), .A3(_03109_ ), .ZN(_03295_ ) );
NAND4_X1 _10965_ ( .A1(_03289_ ), .A2(_03291_ ), .A3(_03293_ ), .A4(_03295_ ), .ZN(_03296_ ) );
NAND2_X1 _10966_ ( .A1(_03285_ ), .A2(_03263_ ), .ZN(_03297_ ) );
NAND4_X1 _10967_ ( .A1(_03071_ ), .A2(_03072_ ), .A3(\IF_ID_inst [4] ), .A4(_03101_ ), .ZN(_03298_ ) );
INV_X1 _10968_ ( .A(_03107_ ), .ZN(_03299_ ) );
OR3_X1 _10969_ ( .A1(_03298_ ), .A2(_03299_ ), .A3(_03294_ ), .ZN(_03300_ ) );
NAND2_X1 _10970_ ( .A1(_03297_ ), .A2(_03300_ ), .ZN(_03301_ ) );
NOR2_X2 _10971_ ( .A1(_03296_ ), .A2(_03301_ ), .ZN(_03302_ ) );
AND3_X1 _10972_ ( .A1(_03284_ ), .A2(_03087_ ), .A3(_03302_ ), .ZN(_03303_ ) );
NOR2_X1 _10973_ ( .A1(_03169_ ), .A2(_03180_ ), .ZN(_03304_ ) );
AND2_X1 _10974_ ( .A1(_03303_ ), .A2(_03304_ ), .ZN(_03305_ ) );
AOI211_X1 _10975_ ( .A(_03234_ ), .B(_03305_ ), .C1(\IF_ID_inst [18] ), .C2(_03304_ ), .ZN(_03306_ ) );
BUF_X4 _10976_ ( .A(_03305_ ), .Z(_03307_ ) );
NOR2_X1 _10977_ ( .A1(_03307_ ), .A2(_03234_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _10978_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_03308_ ) );
AOI211_X1 _10979_ ( .A(_03069_ ), .B(_03306_ ), .C1(_02143_ ), .C2(_03308_ ), .ZN(_00216_ ) );
INV_X1 _10980_ ( .A(\IF_ID_inst [16] ), .ZN(_03309_ ) );
NOR4_X1 _10981_ ( .A1(_03169_ ), .A2(_03309_ ), .A3(_03095_ ), .A4(_03180_ ), .ZN(_00217_ ) );
INV_X1 _10982_ ( .A(_03304_ ), .ZN(_03310_ ) );
OR4_X1 _10983_ ( .A1(_03182_ ), .A2(_03303_ ), .A3(_03310_ ), .A4(_03233_ ), .ZN(_03311_ ) );
OAI21_X1 _10984_ ( .A(\ID_EX_rs1 [2] ), .B1(_03307_ ), .B2(_03234_ ), .ZN(_03312_ ) );
AOI21_X1 _10985_ ( .A(_03086_ ), .B1(_03311_ ), .B2(_03312_ ), .ZN(_00218_ ) );
NOR4_X1 _10986_ ( .A1(_03169_ ), .A2(_03121_ ), .A3(_03095_ ), .A4(_03180_ ), .ZN(_00219_ ) );
OR4_X1 _10987_ ( .A1(_03309_ ), .A2(_03303_ ), .A3(_03310_ ), .A4(_03233_ ), .ZN(_03313_ ) );
OAI21_X1 _10988_ ( .A(\ID_EX_rs1 [1] ), .B1(_03307_ ), .B2(_03234_ ), .ZN(_03314_ ) );
AOI21_X1 _10989_ ( .A(_03086_ ), .B1(_03313_ ), .B2(_03314_ ), .ZN(_00220_ ) );
NAND2_X1 _10990_ ( .A1(_03138_ ), .A2(_03140_ ), .ZN(_03315_ ) );
NAND2_X1 _10991_ ( .A1(_03315_ ), .A2(_03087_ ), .ZN(_03316_ ) );
NOR2_X1 _10992_ ( .A1(_03298_ ), .A2(_03299_ ), .ZN(_03317_ ) );
AOI22_X1 _10993_ ( .A1(_03285_ ), .A2(\IF_ID_inst [14] ), .B1(\IF_ID_inst [13] ), .B2(_03317_ ), .ZN(_03318_ ) );
NAND3_X1 _10994_ ( .A1(_03257_ ), .A2(_03119_ ), .A3(_03109_ ), .ZN(_03319_ ) );
AND2_X1 _10995_ ( .A1(_03319_ ), .A2(_03291_ ), .ZN(_03320_ ) );
NAND2_X1 _10996_ ( .A1(_03318_ ), .A2(_03320_ ), .ZN(_03321_ ) );
AND2_X1 _10997_ ( .A1(_03285_ ), .A2(_03108_ ), .ZN(_03322_ ) );
AND2_X1 _10998_ ( .A1(_03257_ ), .A2(_03109_ ), .ZN(_03323_ ) );
NAND2_X1 _10999_ ( .A1(_03323_ ), .A2(_03148_ ), .ZN(_03324_ ) );
NOR2_X1 _11000_ ( .A1(_03292_ ), .A2(_03162_ ), .ZN(_03325_ ) );
NAND2_X1 _11001_ ( .A1(_03324_ ), .A2(_03325_ ), .ZN(_03326_ ) );
NOR4_X1 _11002_ ( .A1(_03316_ ), .A2(_03321_ ), .A3(_03322_ ), .A4(_03326_ ), .ZN(_03327_ ) );
NOR2_X1 _11003_ ( .A1(_03286_ ), .A2(_03167_ ), .ZN(_03328_ ) );
NAND2_X1 _11004_ ( .A1(_03280_ ), .A2(_03317_ ), .ZN(_03329_ ) );
NAND3_X1 _11005_ ( .A1(_03317_ ), .A2(_03245_ ), .A3(_03247_ ), .ZN(_03330_ ) );
NAND3_X1 _11006_ ( .A1(_03317_ ), .A2(_03253_ ), .A3(_03276_ ), .ZN(_03331_ ) );
AND3_X1 _11007_ ( .A1(_03329_ ), .A2(_03330_ ), .A3(_03331_ ), .ZN(_03332_ ) );
AOI21_X1 _11008_ ( .A(_03112_ ), .B1(_03155_ ), .B2(_03131_ ), .ZN(_03333_ ) );
AND3_X1 _11009_ ( .A1(_03328_ ), .A2(_03332_ ), .A3(_03333_ ), .ZN(_03334_ ) );
AND4_X1 _11010_ ( .A1(\IF_ID_inst [24] ), .A2(_03327_ ), .A3(_03145_ ), .A4(_03334_ ), .ZN(_00221_ ) );
OR4_X1 _11011_ ( .A1(_03121_ ), .A2(_03303_ ), .A3(_03310_ ), .A4(_03233_ ), .ZN(_03335_ ) );
OAI21_X1 _11012_ ( .A(\ID_EX_rs1 [0] ), .B1(_03307_ ), .B2(_03234_ ), .ZN(_03336_ ) );
AOI21_X1 _11013_ ( .A(_03086_ ), .B1(_03335_ ), .B2(_03336_ ), .ZN(_00222_ ) );
AND4_X1 _11014_ ( .A1(\IF_ID_inst [23] ), .A2(_03327_ ), .A3(_03145_ ), .A4(_03334_ ), .ZN(_00223_ ) );
AND4_X1 _11015_ ( .A1(\IF_ID_inst [22] ), .A2(_03327_ ), .A3(_03068_ ), .A4(_03334_ ), .ZN(_00224_ ) );
AND2_X1 _11016_ ( .A1(_03327_ ), .A2(_03334_ ), .ZN(_03337_ ) );
AOI221_X4 _11017_ ( .A(_03233_ ), .B1(\IF_ID_inst [23] ), .B2(_03337_ ), .C1(_03303_ ), .C2(_03304_ ), .ZN(_03338_ ) );
INV_X1 _11018_ ( .A(\ID_EX_rs2 [3] ), .ZN(_03339_ ) );
AOI211_X1 _11019_ ( .A(_03069_ ), .B(_03338_ ), .C1(_03308_ ), .C2(_03339_ ), .ZN(_00225_ ) );
AND4_X1 _11020_ ( .A1(\IF_ID_inst [21] ), .A2(_03327_ ), .A3(_03068_ ), .A4(_03334_ ), .ZN(_00226_ ) );
INV_X1 _11021_ ( .A(_03307_ ), .ZN(_03340_ ) );
NAND4_X1 _11022_ ( .A1(_03340_ ), .A2(\IF_ID_inst [22] ), .A3(_03232_ ), .A4(_03337_ ), .ZN(_03341_ ) );
OAI21_X1 _11023_ ( .A(\ID_EX_rs2 [2] ), .B1(_03307_ ), .B2(_03234_ ), .ZN(_03342_ ) );
AOI21_X1 _11024_ ( .A(_03086_ ), .B1(_03341_ ), .B2(_03342_ ), .ZN(_00227_ ) );
AND4_X1 _11025_ ( .A1(\IF_ID_inst [20] ), .A2(_03327_ ), .A3(_03068_ ), .A4(_03334_ ), .ZN(_00228_ ) );
AOI221_X4 _11026_ ( .A(_03233_ ), .B1(\IF_ID_inst [21] ), .B2(_03337_ ), .C1(_03303_ ), .C2(_03304_ ), .ZN(_03343_ ) );
INV_X1 _11027_ ( .A(\ID_EX_rs2 [1] ), .ZN(_03344_ ) );
AOI211_X1 _11028_ ( .A(_03069_ ), .B(_03343_ ), .C1(_03308_ ), .C2(_03344_ ), .ZN(_00229_ ) );
INV_X1 _11029_ ( .A(IDU_valid_EXU ), .ZN(_03345_ ) );
AND4_X1 _11030_ ( .A1(_03345_ ), .A2(_03110_ ), .A3(_03068_ ), .A4(_03111_ ), .ZN(_00230_ ) );
NAND4_X1 _11031_ ( .A1(_03340_ ), .A2(\IF_ID_inst [20] ), .A3(_03232_ ), .A4(_03337_ ), .ZN(_03346_ ) );
OAI21_X1 _11032_ ( .A(\ID_EX_rs2 [0] ), .B1(_03307_ ), .B2(_03234_ ), .ZN(_03347_ ) );
AOI21_X1 _11033_ ( .A(_03086_ ), .B1(_03346_ ), .B2(_03347_ ), .ZN(_00231_ ) );
INV_X1 _11034_ ( .A(\ID_EX_typ [7] ), .ZN(_03348_ ) );
INV_X1 _11035_ ( .A(\ID_EX_rd [3] ), .ZN(_03349_ ) );
NOR2_X1 _11036_ ( .A1(_03349_ ), .A2(\IF_ID_inst [18] ), .ZN(_03350_ ) );
OAI22_X1 _11037_ ( .A1(\ID_EX_rd [3] ), .A2(_03181_ ), .B1(_03309_ ), .B2(\ID_EX_rd [1] ), .ZN(_03351_ ) );
AOI211_X1 _11038_ ( .A(_03350_ ), .B(_03351_ ), .C1(\ID_EX_rd [1] ), .C2(_03309_ ), .ZN(_03352_ ) );
AND2_X1 _11039_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03353_ ) );
XNOR2_X1 _11040_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_03354_ ) );
AND4_X1 _11041_ ( .A1(_03348_ ), .A2(_03352_ ), .A3(_03353_ ), .A4(_03354_ ), .ZN(_03355_ ) );
XNOR2_X1 _11042_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_03356_ ) );
XNOR2_X1 _11043_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_03357_ ) );
NAND3_X1 _11044_ ( .A1(_03355_ ), .A2(_03356_ ), .A3(_03357_ ), .ZN(_03358_ ) );
INV_X1 _11045_ ( .A(_03302_ ), .ZN(_03359_ ) );
OAI21_X1 _11046_ ( .A(_03358_ ), .B1(_03359_ ), .B2(_03088_ ), .ZN(_03360_ ) );
XNOR2_X1 _11047_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_03361_ ) );
CLKBUF_X2 _11048_ ( .A(_03353_ ), .Z(_03362_ ) );
AND3_X1 _11049_ ( .A1(_03361_ ), .A2(_03348_ ), .A3(_03362_ ), .ZN(_03363_ ) );
XNOR2_X1 _11050_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_03364_ ) );
XNOR2_X1 _11051_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_03365_ ) );
AND2_X1 _11052_ ( .A1(_03364_ ), .A2(_03365_ ), .ZN(_03366_ ) );
XNOR2_X1 _11053_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_03367_ ) );
XNOR2_X1 _11054_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_03368_ ) );
NAND4_X1 _11055_ ( .A1(_03363_ ), .A2(_03366_ ), .A3(_03367_ ), .A4(_03368_ ), .ZN(_03369_ ) );
NAND2_X1 _11056_ ( .A1(_03358_ ), .A2(_03369_ ), .ZN(_03370_ ) );
AND3_X1 _11057_ ( .A1(_03140_ ), .A2(_03122_ ), .A3(_03116_ ), .ZN(_03371_ ) );
AOI21_X1 _11058_ ( .A(_03112_ ), .B1(_03371_ ), .B2(_03137_ ), .ZN(_03372_ ) );
NAND4_X1 _11059_ ( .A1(_03370_ ), .A2(_03372_ ), .A3(_03157_ ), .A4(_03168_ ), .ZN(_03373_ ) );
NAND3_X1 _11060_ ( .A1(_03302_ ), .A2(_03373_ ), .A3(_03087_ ), .ZN(_03374_ ) );
AND3_X1 _11061_ ( .A1(_02094_ ), .A2(_03067_ ), .A3(IDU_ready_IFU ), .ZN(_03375_ ) );
AND3_X1 _11062_ ( .A1(_03360_ ), .A2(_03374_ ), .A3(_03375_ ), .ZN(_00232_ ) );
AND2_X1 _11063_ ( .A1(_03123_ ), .A2(_03132_ ), .ZN(_03376_ ) );
OR2_X1 _11064_ ( .A1(_03376_ ), .A2(_03112_ ), .ZN(_03377_ ) );
NOR4_X1 _11065_ ( .A1(_03377_ ), .A2(_03264_ ), .A3(_03162_ ), .A4(_03292_ ), .ZN(_03378_ ) );
NAND4_X1 _11066_ ( .A1(_03122_ ), .A2(_03089_ ), .A3(_03075_ ), .A4(_03176_ ), .ZN(_03379_ ) );
NAND3_X1 _11067_ ( .A1(_03137_ ), .A2(_03085_ ), .A3(_03139_ ), .ZN(_03380_ ) );
NOR2_X1 _11068_ ( .A1(_03379_ ), .A2(_03380_ ), .ZN(_03381_ ) );
NOR2_X1 _11069_ ( .A1(_03381_ ), .A2(_03088_ ), .ZN(_03382_ ) );
AOI21_X1 _11070_ ( .A(_03086_ ), .B1(_03378_ ), .B2(_03382_ ), .ZN(_00233_ ) );
AND2_X1 _11071_ ( .A1(_03290_ ), .A2(_03246_ ), .ZN(_03383_ ) );
INV_X1 _11072_ ( .A(_03383_ ), .ZN(_03384_ ) );
NAND3_X1 _11073_ ( .A1(_03171_ ), .A2(_03075_ ), .A3(_03108_ ), .ZN(_03385_ ) );
AND4_X1 _11074_ ( .A1(_03153_ ), .A2(_03384_ ), .A3(_03295_ ), .A4(_03385_ ), .ZN(_03386_ ) );
AOI21_X1 _11075_ ( .A(_03070_ ), .B1(_03386_ ), .B2(_03382_ ), .ZN(_00234_ ) );
AND3_X1 _11076_ ( .A1(_03250_ ), .A2(_03174_ ), .A3(_03235_ ), .ZN(_03387_ ) );
NAND3_X1 _11077_ ( .A1(_03256_ ), .A2(_03174_ ), .A3(_03235_ ), .ZN(_03388_ ) );
NAND3_X1 _11078_ ( .A1(_03251_ ), .A2(_03174_ ), .A3(_03235_ ), .ZN(_03389_ ) );
NAND2_X1 _11079_ ( .A1(_03388_ ), .A2(_03389_ ), .ZN(_03390_ ) );
NOR2_X1 _11080_ ( .A1(_03387_ ), .A2(_03390_ ), .ZN(_03391_ ) );
NOR3_X1 _11081_ ( .A1(_03269_ ), .A2(\IF_ID_inst [26] ), .A3(\IF_ID_inst [25] ), .ZN(_03392_ ) );
AND3_X1 _11082_ ( .A1(_03253_ ), .A2(_03142_ ), .A3(_03392_ ), .ZN(_03393_ ) );
NOR2_X1 _11083_ ( .A1(_03251_ ), .A2(_03393_ ), .ZN(_03394_ ) );
INV_X1 _11084_ ( .A(_03394_ ), .ZN(_03395_ ) );
AND3_X1 _11085_ ( .A1(_03393_ ), .A2(_03174_ ), .A3(_03235_ ), .ZN(_03396_ ) );
AND2_X1 _11086_ ( .A1(_03257_ ), .A2(_03174_ ), .ZN(_03397_ ) );
OAI22_X1 _11087_ ( .A1(_03395_ ), .A2(_03242_ ), .B1(_03396_ ), .B2(_03397_ ), .ZN(_03398_ ) );
NAND2_X1 _11088_ ( .A1(_03391_ ), .A2(_03398_ ), .ZN(_03399_ ) );
NAND3_X1 _11089_ ( .A1(_03320_ ), .A2(_03258_ ), .A3(_03259_ ), .ZN(_03400_ ) );
AND3_X1 _11090_ ( .A1(_03139_ ), .A2(_03085_ ), .A3(_03089_ ), .ZN(_03401_ ) );
AND2_X1 _11091_ ( .A1(_03138_ ), .A2(_03401_ ), .ZN(_03402_ ) );
NOR4_X1 _11092_ ( .A1(_03399_ ), .A2(_03400_ ), .A3(_03326_ ), .A4(_03402_ ), .ZN(_03403_ ) );
AND2_X1 _11093_ ( .A1(_03297_ ), .A2(_03287_ ), .ZN(_03404_ ) );
AND3_X1 _11094_ ( .A1(_03328_ ), .A2(_03332_ ), .A3(_03404_ ), .ZN(_03405_ ) );
AOI21_X1 _11095_ ( .A(_03070_ ), .B1(_03403_ ), .B2(_03405_ ), .ZN(_00235_ ) );
INV_X1 _11096_ ( .A(_03112_ ), .ZN(_03406_ ) );
AOI21_X1 _11097_ ( .A(_03070_ ), .B1(_03405_ ), .B2(_03406_ ), .ZN(_00236_ ) );
AND3_X1 _11098_ ( .A1(_03256_ ), .A2(_03174_ ), .A3(_03257_ ), .ZN(_03407_ ) );
AND4_X1 _11099_ ( .A1(_03174_ ), .A2(_03257_ ), .A3(_03241_ ), .A4(_03245_ ), .ZN(_03408_ ) );
NOR4_X1 _11100_ ( .A1(_03376_ ), .A2(_03149_ ), .A3(_03407_ ), .A4(_03408_ ), .ZN(_03409_ ) );
AOI21_X1 _11101_ ( .A(_03070_ ), .B1(_03409_ ), .B2(_03328_ ), .ZN(_00237_ ) );
NAND2_X1 _11102_ ( .A1(_03317_ ), .A2(_03148_ ), .ZN(_03410_ ) );
AND4_X1 _11103_ ( .A1(_03324_ ), .A2(_03278_ ), .A3(_03281_ ), .A4(_03410_ ), .ZN(_03411_ ) );
AOI21_X1 _11104_ ( .A(_03167_ ), .B1(_03147_ ), .B2(_03148_ ), .ZN(_03412_ ) );
AND3_X1 _11105_ ( .A1(_03075_ ), .A2(\IF_ID_inst [13] ), .A3(_03076_ ), .ZN(_03413_ ) );
AOI21_X1 _11106_ ( .A(_03413_ ), .B1(_03141_ ), .B2(\IF_ID_inst [14] ), .ZN(_03414_ ) );
NAND4_X1 _11107_ ( .A1(_03411_ ), .A2(_03332_ ), .A3(_03412_ ), .A4(_03414_ ), .ZN(_03415_ ) );
AND2_X1 _11108_ ( .A1(_03415_ ), .A2(_03145_ ), .ZN(_00238_ ) );
AND2_X1 _11109_ ( .A1(_03395_ ), .A2(_03397_ ), .ZN(_03416_ ) );
NAND3_X1 _11110_ ( .A1(_03248_ ), .A2(_03235_ ), .A3(_03236_ ), .ZN(_03417_ ) );
NAND4_X1 _11111_ ( .A1(_03235_ ), .A2(_03236_ ), .A3(_03239_ ), .A4(_03247_ ), .ZN(_03418_ ) );
NAND2_X1 _11112_ ( .A1(_03417_ ), .A2(_03418_ ), .ZN(_03419_ ) );
AND2_X1 _11113_ ( .A1(_03285_ ), .A2(\IF_ID_inst [14] ), .ZN(_03420_ ) );
NAND4_X1 _11114_ ( .A1(_03235_ ), .A2(_03174_ ), .A3(_03245_ ), .A4(_03247_ ), .ZN(_03421_ ) );
NAND3_X1 _11115_ ( .A1(_03421_ ), .A2(_03105_ ), .A3(_03083_ ), .ZN(_03422_ ) );
NOR4_X1 _11116_ ( .A1(_03416_ ), .A2(_03419_ ), .A3(_03420_ ), .A4(_03422_ ), .ZN(_03423_ ) );
AND3_X1 _11117_ ( .A1(_03079_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_03424_ ) );
NAND2_X1 _11118_ ( .A1(_03164_ ), .A2(_03424_ ), .ZN(_03425_ ) );
NOR2_X1 _11119_ ( .A1(_03149_ ), .A2(_03383_ ), .ZN(_03426_ ) );
NAND3_X1 _11120_ ( .A1(_03235_ ), .A2(_03108_ ), .A3(_03102_ ), .ZN(_03427_ ) );
AND2_X1 _11121_ ( .A1(_03427_ ), .A2(_03385_ ), .ZN(_03428_ ) );
AND4_X1 _11122_ ( .A1(_03425_ ), .A2(_03426_ ), .A3(_03389_ ), .A4(_03428_ ), .ZN(_03429_ ) );
AOI21_X1 _11123_ ( .A(_03070_ ), .B1(_03423_ ), .B2(_03429_ ), .ZN(_00239_ ) );
AOI221_X4 _11124_ ( .A(_03292_ ), .B1(_03142_ ), .B2(_03141_ ), .C1(_03371_ ), .C2(_03137_ ), .ZN(_03430_ ) );
NAND3_X1 _11125_ ( .A1(_03075_ ), .A2(_03076_ ), .A3(_03246_ ), .ZN(_03431_ ) );
NAND2_X1 _11126_ ( .A1(_03141_ ), .A2(_03108_ ), .ZN(_03432_ ) );
NAND4_X1 _11127_ ( .A1(_03267_ ), .A2(\IF_ID_inst [14] ), .A3(\IF_ID_inst [13] ), .A4(_03080_ ), .ZN(_03433_ ) );
AND4_X1 _11128_ ( .A1(_03431_ ), .A2(_03432_ ), .A3(_03150_ ), .A4(_03433_ ), .ZN(_03434_ ) );
NAND2_X1 _11129_ ( .A1(_03323_ ), .A2(_03246_ ), .ZN(_03435_ ) );
AND4_X1 _11130_ ( .A1(_03152_ ), .A2(_03435_ ), .A3(_03384_ ), .A4(_03330_ ), .ZN(_03436_ ) );
AND2_X1 _11131_ ( .A1(_03267_ ), .A2(_03146_ ), .ZN(_03437_ ) );
NAND4_X1 _11132_ ( .A1(_03437_ ), .A2(_03148_ ), .A3(_03253_ ), .A4(_03392_ ), .ZN(_03438_ ) );
AND3_X1 _11133_ ( .A1(_03281_ ), .A2(_03329_ ), .A3(_03438_ ), .ZN(_03439_ ) );
AND4_X1 _11134_ ( .A1(_03430_ ), .A2(_03434_ ), .A3(_03436_ ), .A4(_03439_ ), .ZN(_03440_ ) );
NAND3_X1 _11135_ ( .A1(_03285_ ), .A2(\IF_ID_inst [14] ), .A3(_03119_ ), .ZN(_03441_ ) );
OAI21_X1 _11136_ ( .A(_03142_ ), .B1(_03104_ ), .B2(_03077_ ), .ZN(_03442_ ) );
AOI22_X1 _11137_ ( .A1(_03437_ ), .A2(_03277_ ), .B1(_03275_ ), .B2(_03270_ ), .ZN(_03443_ ) );
AND4_X1 _11138_ ( .A1(_03300_ ), .A2(_03441_ ), .A3(_03442_ ), .A4(_03443_ ), .ZN(_03444_ ) );
AOI21_X1 _11139_ ( .A(_03070_ ), .B1(_03440_ ), .B2(_03444_ ), .ZN(_00240_ ) );
INV_X1 _11140_ ( .A(_03225_ ), .ZN(_03445_ ) );
INV_X1 _11141_ ( .A(\myifu.to_reset ), .ZN(_03446_ ) );
BUF_X4 _11142_ ( .A(_03446_ ), .Z(_03447_ ) );
NAND4_X1 _11143_ ( .A1(_03445_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_03447_ ), .ZN(_03448_ ) );
NAND2_X1 _11144_ ( .A1(\mtvec [0] ), .A2(\myifu.to_reset ), .ZN(_03449_ ) );
AOI21_X1 _11145_ ( .A(fanout_net_2 ), .B1(_03448_ ), .B2(_03449_ ), .ZN(_00244_ ) );
INV_X1 _11146_ ( .A(_03227_ ), .ZN(_03450_ ) );
BUF_X4 _11147_ ( .A(_03450_ ), .Z(_03451_ ) );
AND4_X1 _11148_ ( .A1(\IF_ID_inst [31] ), .A2(_03165_ ), .A3(_03158_ ), .A4(\IF_ID_inst [5] ), .ZN(_03452_ ) );
AND2_X2 _11149_ ( .A1(_03073_ ), .A2(_03452_ ), .ZN(_03453_ ) );
AOI21_X1 _11150_ ( .A(_03453_ ), .B1(_03162_ ), .B2(\IF_ID_inst [31] ), .ZN(_03454_ ) );
AND2_X1 _11151_ ( .A1(_03453_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03455_ ) );
NOR2_X1 _11152_ ( .A1(_03454_ ), .A2(_03455_ ), .ZN(_03456_ ) );
BUF_X4 _11153_ ( .A(_03456_ ), .Z(_03457_ ) );
BUF_X4 _11154_ ( .A(_03457_ ), .Z(_03458_ ) );
XNOR2_X1 _11155_ ( .A(_03458_ ), .B(_01801_ ), .ZN(_03459_ ) );
INV_X1 _11156_ ( .A(_03459_ ), .ZN(_03460_ ) );
AND2_X1 _11157_ ( .A1(_03162_ ), .A2(\IF_ID_inst [19] ), .ZN(_03461_ ) );
INV_X1 _11158_ ( .A(_03453_ ), .ZN(_03462_ ) );
MUX2_X1 _11159_ ( .A(_03269_ ), .B(_03461_ ), .S(_03462_ ), .Z(_03463_ ) );
XNOR2_X1 _11160_ ( .A(_03463_ ), .B(_01939_ ), .ZN(_03464_ ) );
XNOR2_X1 _11161_ ( .A(_03456_ ), .B(_01890_ ), .ZN(_03465_ ) );
AND2_X1 _11162_ ( .A1(_03464_ ), .A2(_03465_ ), .ZN(_03466_ ) );
AND2_X1 _11163_ ( .A1(_03161_ ), .A2(\IF_ID_inst [18] ), .ZN(_03467_ ) );
NAND4_X1 _11164_ ( .A1(_03102_ ), .A2(_03158_ ), .A3(_03071_ ), .A4(_03072_ ), .ZN(_03468_ ) );
NOR2_X1 _11165_ ( .A1(_03468_ ), .A2(_03066_ ), .ZN(_03469_ ) );
INV_X1 _11166_ ( .A(_03469_ ), .ZN(_03470_ ) );
MUX2_X1 _11167_ ( .A(_03269_ ), .B(_03467_ ), .S(_03470_ ), .Z(_03471_ ) );
XNOR2_X1 _11168_ ( .A(_03471_ ), .B(_02018_ ), .ZN(_03472_ ) );
AND2_X1 _11169_ ( .A1(_03162_ ), .A2(\IF_ID_inst [17] ), .ZN(_03473_ ) );
MUX2_X1 _11170_ ( .A(_03269_ ), .B(_03473_ ), .S(_03462_ ), .Z(_03474_ ) );
XNOR2_X1 _11171_ ( .A(_03474_ ), .B(_01824_ ), .ZN(_03475_ ) );
AND2_X1 _11172_ ( .A1(_03472_ ), .A2(_03475_ ), .ZN(_03476_ ) );
AND2_X1 _11173_ ( .A1(_03160_ ), .A2(\IF_ID_inst [15] ), .ZN(_03477_ ) );
MUX2_X1 _11174_ ( .A(_03269_ ), .B(_03477_ ), .S(_03462_ ), .Z(_03478_ ) );
INV_X1 _11175_ ( .A(\IF_ID_pc [15] ), .ZN(_03479_ ) );
XNOR2_X1 _11176_ ( .A(_03478_ ), .B(_03479_ ), .ZN(_03480_ ) );
AND2_X1 _11177_ ( .A1(_03469_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03481_ ) );
INV_X1 _11178_ ( .A(_03481_ ), .ZN(_03482_ ) );
AND2_X1 _11179_ ( .A1(_03161_ ), .A2(\IF_ID_inst [16] ), .ZN(_03483_ ) );
OAI21_X1 _11180_ ( .A(_03482_ ), .B1(_03483_ ), .B2(_03469_ ), .ZN(_03484_ ) );
NAND2_X1 _11181_ ( .A1(_03484_ ), .A2(_01859_ ), .ZN(_03485_ ) );
OR2_X1 _11182_ ( .A1(_03484_ ), .A2(_01859_ ), .ZN(_03486_ ) );
NAND3_X1 _11183_ ( .A1(_03480_ ), .A2(_03485_ ), .A3(_03486_ ), .ZN(_03487_ ) );
AND2_X1 _11184_ ( .A1(_03160_ ), .A2(\IF_ID_inst [13] ), .ZN(_03488_ ) );
MUX2_X1 _11185_ ( .A(_03269_ ), .B(_03488_ ), .S(_03462_ ), .Z(_03489_ ) );
XNOR2_X1 _11186_ ( .A(_03489_ ), .B(_01949_ ), .ZN(_03490_ ) );
INV_X1 _11187_ ( .A(_03490_ ), .ZN(_03491_ ) );
AND2_X1 _11188_ ( .A1(_03160_ ), .A2(\IF_ID_inst [14] ), .ZN(_03492_ ) );
MUX2_X1 _11189_ ( .A(_03269_ ), .B(_03492_ ), .S(_03462_ ), .Z(_03493_ ) );
XNOR2_X1 _11190_ ( .A(_03493_ ), .B(\IF_ID_pc [14] ), .ZN(_03494_ ) );
OR3_X1 _11191_ ( .A1(_03487_ ), .A2(_03491_ ), .A3(_03494_ ), .ZN(_03495_ ) );
NAND2_X1 _11192_ ( .A1(_03161_ ), .A2(\IF_ID_inst [20] ), .ZN(_03496_ ) );
OAI21_X1 _11193_ ( .A(_03496_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03462_ ), .ZN(_03497_ ) );
XNOR2_X1 _11194_ ( .A(_03497_ ), .B(_01923_ ), .ZN(_03498_ ) );
AOI21_X1 _11195_ ( .A(_03453_ ), .B1(_03161_ ), .B2(\IF_ID_inst [12] ), .ZN(_03499_ ) );
NOR3_X1 _11196_ ( .A1(_03499_ ), .A2(_03481_ ), .A3(_01832_ ), .ZN(_03500_ ) );
INV_X1 _11197_ ( .A(_03500_ ), .ZN(_03501_ ) );
OAI21_X1 _11198_ ( .A(_01832_ ), .B1(_03499_ ), .B2(_03455_ ), .ZN(_03502_ ) );
AND3_X1 _11199_ ( .A1(_03498_ ), .A2(_03501_ ), .A3(_03502_ ), .ZN(_03503_ ) );
INV_X1 _11200_ ( .A(_03503_ ), .ZN(_03504_ ) );
AND2_X1 _11201_ ( .A1(_03160_ ), .A2(\IF_ID_inst [29] ), .ZN(_03505_ ) );
INV_X1 _11202_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03506_ ) );
AOI21_X1 _11203_ ( .A(_03505_ ), .B1(_03506_ ), .B2(_03453_ ), .ZN(_03507_ ) );
XNOR2_X1 _11204_ ( .A(_03507_ ), .B(\IF_ID_pc [9] ), .ZN(_03508_ ) );
INV_X1 _11205_ ( .A(_03508_ ), .ZN(_03509_ ) );
INV_X1 _11206_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03510_ ) );
AND3_X1 _11207_ ( .A1(_03074_ ), .A2(_03452_ ), .A3(_03510_ ), .ZN(_03511_ ) );
AOI21_X1 _11208_ ( .A(_03511_ ), .B1(\IF_ID_inst [30] ), .B2(_03161_ ), .ZN(_03512_ ) );
XNOR2_X1 _11209_ ( .A(_03512_ ), .B(_01863_ ), .ZN(_03513_ ) );
OR3_X1 _11210_ ( .A1(_03504_ ), .A2(_03509_ ), .A3(_03513_ ), .ZN(_03514_ ) );
AND2_X1 _11211_ ( .A1(_03162_ ), .A2(\IF_ID_inst [28] ), .ZN(_03515_ ) );
INV_X1 _11212_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03516_ ) );
AOI21_X1 _11213_ ( .A(_03515_ ), .B1(_03516_ ), .B2(_03453_ ), .ZN(_03517_ ) );
XNOR2_X1 _11214_ ( .A(_03517_ ), .B(\IF_ID_pc [8] ), .ZN(_03518_ ) );
AND2_X1 _11215_ ( .A1(_03162_ ), .A2(\IF_ID_inst [27] ), .ZN(_03519_ ) );
INV_X1 _11216_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03520_ ) );
AOI21_X1 _11217_ ( .A(_03519_ ), .B1(_03520_ ), .B2(_03453_ ), .ZN(_03521_ ) );
XNOR2_X1 _11218_ ( .A(_03521_ ), .B(\IF_ID_pc [7] ), .ZN(_03522_ ) );
AND2_X1 _11219_ ( .A1(_03161_ ), .A2(\IF_ID_inst [25] ), .ZN(_03523_ ) );
INV_X1 _11220_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03524_ ) );
AND3_X1 _11221_ ( .A1(_03074_ ), .A2(_03452_ ), .A3(_03524_ ), .ZN(_03525_ ) );
NOR2_X1 _11222_ ( .A1(_03523_ ), .A2(_03525_ ), .ZN(_03526_ ) );
INV_X1 _11223_ ( .A(\IF_ID_pc [5] ), .ZN(_03527_ ) );
XNOR2_X1 _11224_ ( .A(_03526_ ), .B(_03527_ ), .ZN(_03528_ ) );
INV_X1 _11225_ ( .A(_03528_ ), .ZN(_03529_ ) );
INV_X1 _11226_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03530_ ) );
AND3_X1 _11227_ ( .A1(_03074_ ), .A2(_03452_ ), .A3(_03530_ ), .ZN(_03531_ ) );
AOI21_X1 _11228_ ( .A(_03531_ ), .B1(\IF_ID_inst [26] ), .B2(_03161_ ), .ZN(_03532_ ) );
XNOR2_X1 _11229_ ( .A(_03532_ ), .B(\IF_ID_pc [6] ), .ZN(_03533_ ) );
NAND2_X1 _11230_ ( .A1(_03529_ ), .A2(_03533_ ), .ZN(_03534_ ) );
INV_X1 _11231_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03535_ ) );
NOR3_X1 _11232_ ( .A1(_03468_ ), .A2(_03066_ ), .A3(_03535_ ), .ZN(_03536_ ) );
AOI21_X1 _11233_ ( .A(_03536_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .B2(_03160_ ), .ZN(_03537_ ) );
XOR2_X1 _11234_ ( .A(_03537_ ), .B(\IF_ID_pc [2] ), .Z(_03538_ ) );
INV_X1 _11235_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03539_ ) );
AND3_X1 _11236_ ( .A1(_03073_ ), .A2(_03452_ ), .A3(_03539_ ), .ZN(_03540_ ) );
AOI21_X1 _11237_ ( .A(_03540_ ), .B1(\IF_ID_inst [21] ), .B2(_03160_ ), .ZN(_03541_ ) );
INV_X1 _11238_ ( .A(\IF_ID_pc [1] ), .ZN(_03542_ ) );
NOR2_X1 _11239_ ( .A1(_03541_ ), .A2(_03542_ ), .ZN(_03543_ ) );
AND2_X1 _11240_ ( .A1(_03538_ ), .A2(_03543_ ), .ZN(_03544_ ) );
AND2_X1 _11241_ ( .A1(_03537_ ), .A2(\IF_ID_pc [2] ), .ZN(_03545_ ) );
NOR2_X1 _11242_ ( .A1(_03544_ ), .A2(_03545_ ), .ZN(_03546_ ) );
AOI21_X1 _11243_ ( .A(_03469_ ), .B1(_03161_ ), .B2(\IF_ID_inst [23] ), .ZN(_03547_ ) );
INV_X1 _11244_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03548_ ) );
NOR3_X1 _11245_ ( .A1(_03468_ ), .A2(_03066_ ), .A3(_03548_ ), .ZN(_03549_ ) );
NOR2_X1 _11246_ ( .A1(_03547_ ), .A2(_03549_ ), .ZN(_03550_ ) );
XNOR2_X1 _11247_ ( .A(_03550_ ), .B(fanout_net_7 ), .ZN(_03551_ ) );
OR2_X1 _11248_ ( .A1(_03546_ ), .A2(_03551_ ), .ZN(_03552_ ) );
OR3_X1 _11249_ ( .A1(_03547_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(_03549_ ), .ZN(_03553_ ) );
NAND2_X1 _11250_ ( .A1(_03552_ ), .A2(_03553_ ), .ZN(_03554_ ) );
INV_X1 _11251_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_03555_ ) );
NAND3_X1 _11252_ ( .A1(_03074_ ), .A2(_03452_ ), .A3(_03555_ ), .ZN(_03556_ ) );
INV_X1 _11253_ ( .A(_03161_ ), .ZN(_03557_ ) );
OAI21_X1 _11254_ ( .A(_03556_ ), .B1(_03557_ ), .B2(_03096_ ), .ZN(_03558_ ) );
OAI21_X1 _11255_ ( .A(_03554_ ), .B1(fanout_net_11 ), .B2(_03558_ ), .ZN(_03559_ ) );
NAND2_X1 _11256_ ( .A1(_03558_ ), .A2(fanout_net_11 ), .ZN(_03560_ ) );
AOI21_X1 _11257_ ( .A(_03534_ ), .B1(_03559_ ), .B2(_03560_ ), .ZN(_03561_ ) );
NOR2_X1 _11258_ ( .A1(_03532_ ), .A2(_01908_ ), .ZN(_03562_ ) );
NOR2_X1 _11259_ ( .A1(_03526_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03563_ ) );
AND2_X1 _11260_ ( .A1(_03532_ ), .A2(_01908_ ), .ZN(_03564_ ) );
INV_X1 _11261_ ( .A(_03564_ ), .ZN(_03565_ ) );
AOI21_X1 _11262_ ( .A(_03562_ ), .B1(_03563_ ), .B2(_03565_ ), .ZN(_03566_ ) );
INV_X1 _11263_ ( .A(_03566_ ), .ZN(_03567_ ) );
OAI211_X1 _11264_ ( .A(_03518_ ), .B(_03522_ ), .C1(_03561_ ), .C2(_03567_ ), .ZN(_03568_ ) );
NOR2_X1 _11265_ ( .A1(_03517_ ), .A2(_01810_ ), .ZN(_03569_ ) );
NOR2_X1 _11266_ ( .A1(_03521_ ), .A2(_01789_ ), .ZN(_03570_ ) );
AOI21_X1 _11267_ ( .A(_03569_ ), .B1(_03518_ ), .B2(_03570_ ), .ZN(_03571_ ) );
AOI211_X1 _11268_ ( .A(_03495_ ), .B(_03514_ ), .C1(_03568_ ), .C2(_03571_ ), .ZN(_03572_ ) );
NOR2_X1 _11269_ ( .A1(_03484_ ), .A2(_01859_ ), .ZN(_03573_ ) );
OR2_X1 _11270_ ( .A1(_03512_ ), .A2(_01863_ ), .ZN(_03574_ ) );
MUX2_X1 _11271_ ( .A(_03506_ ), .B(_03505_ ), .S(_03470_ ), .Z(_03575_ ) );
AND2_X1 _11272_ ( .A1(_03575_ ), .A2(\IF_ID_pc [9] ), .ZN(_03576_ ) );
INV_X1 _11273_ ( .A(_03576_ ), .ZN(_03577_ ) );
OAI21_X1 _11274_ ( .A(_03574_ ), .B1(_03577_ ), .B2(_03513_ ), .ZN(_03578_ ) );
NAND2_X1 _11275_ ( .A1(_03578_ ), .A2(_03503_ ), .ZN(_03579_ ) );
NAND4_X1 _11276_ ( .A1(_03501_ ), .A2(\IF_ID_pc [11] ), .A3(_03502_ ), .A4(_03497_ ), .ZN(_03580_ ) );
AND3_X1 _11277_ ( .A1(_03579_ ), .A2(_03501_ ), .A3(_03580_ ), .ZN(_03581_ ) );
NOR2_X1 _11278_ ( .A1(_03581_ ), .A2(_03495_ ), .ZN(_03582_ ) );
OAI21_X1 _11279_ ( .A(_03482_ ), .B1(_03488_ ), .B2(_03469_ ), .ZN(_03583_ ) );
OR3_X1 _11280_ ( .A1(_03494_ ), .A2(_01949_ ), .A3(_03583_ ), .ZN(_03584_ ) );
NAND2_X1 _11281_ ( .A1(_03493_ ), .A2(\IF_ID_pc [14] ), .ZN(_03585_ ) );
AOI21_X1 _11282_ ( .A(_03487_ ), .B1(_03584_ ), .B2(_03585_ ), .ZN(_03586_ ) );
AND4_X1 _11283_ ( .A1(\IF_ID_pc [15] ), .A2(_03486_ ), .A3(_03485_ ), .A4(_03478_ ), .ZN(_03587_ ) );
OR4_X1 _11284_ ( .A1(_03573_ ), .A2(_03582_ ), .A3(_03586_ ), .A4(_03587_ ), .ZN(_03588_ ) );
OAI211_X1 _11285_ ( .A(_03466_ ), .B(_03476_ ), .C1(_03572_ ), .C2(_03588_ ), .ZN(_03589_ ) );
OAI211_X1 _11286_ ( .A(_03463_ ), .B(\IF_ID_pc [19] ), .C1(\IF_ID_pc [20] ), .C2(_03456_ ), .ZN(_03590_ ) );
INV_X1 _11287_ ( .A(_03456_ ), .ZN(_03591_ ) );
OAI21_X1 _11288_ ( .A(_03590_ ), .B1(_01890_ ), .B2(_03591_ ), .ZN(_03592_ ) );
AND2_X1 _11289_ ( .A1(_03474_ ), .A2(\IF_ID_pc [17] ), .ZN(_03593_ ) );
AND2_X1 _11290_ ( .A1(_03472_ ), .A2(_03593_ ), .ZN(_03594_ ) );
AOI21_X1 _11291_ ( .A(_03594_ ), .B1(\IF_ID_pc [18] ), .B2(_03471_ ), .ZN(_03595_ ) );
INV_X1 _11292_ ( .A(_03595_ ), .ZN(_03596_ ) );
AOI21_X1 _11293_ ( .A(_03592_ ), .B1(_03596_ ), .B2(_03466_ ), .ZN(_03597_ ) );
AND2_X1 _11294_ ( .A1(_03589_ ), .A2(_03597_ ), .ZN(_03598_ ) );
XNOR2_X1 _11295_ ( .A(_03456_ ), .B(_01903_ ), .ZN(_03599_ ) );
XNOR2_X1 _11296_ ( .A(_03456_ ), .B(_01785_ ), .ZN(_03600_ ) );
AND2_X1 _11297_ ( .A1(_03599_ ), .A2(_03600_ ), .ZN(_03601_ ) );
INV_X1 _11298_ ( .A(_03601_ ), .ZN(_03602_ ) );
XNOR2_X1 _11299_ ( .A(_03457_ ), .B(\IF_ID_pc [22] ), .ZN(_03603_ ) );
XNOR2_X1 _11300_ ( .A(_03457_ ), .B(_01806_ ), .ZN(_03604_ ) );
INV_X1 _11301_ ( .A(_03604_ ), .ZN(_03605_ ) );
NOR4_X1 _11302_ ( .A1(_03598_ ), .A2(_03602_ ), .A3(_03603_ ), .A4(_03605_ ), .ZN(_03606_ ) );
AND2_X1 _11303_ ( .A1(_03457_ ), .A2(\IF_ID_pc [22] ), .ZN(_03607_ ) );
AND2_X1 _11304_ ( .A1(_03457_ ), .A2(\IF_ID_pc [21] ), .ZN(_03608_ ) );
OAI21_X1 _11305_ ( .A(_03601_ ), .B1(_03607_ ), .B2(_03608_ ), .ZN(_03609_ ) );
NAND2_X1 _11306_ ( .A1(_03457_ ), .A2(\IF_ID_pc [24] ), .ZN(_03610_ ) );
NAND2_X1 _11307_ ( .A1(_03457_ ), .A2(\IF_ID_pc [23] ), .ZN(_03611_ ) );
NAND3_X1 _11308_ ( .A1(_03609_ ), .A2(_03610_ ), .A3(_03611_ ), .ZN(_03612_ ) );
NOR2_X1 _11309_ ( .A1(_03606_ ), .A2(_03612_ ), .ZN(_03613_ ) );
INV_X1 _11310_ ( .A(_03613_ ), .ZN(_03614_ ) );
XNOR2_X1 _11311_ ( .A(_03457_ ), .B(_02004_ ), .ZN(_03615_ ) );
AND2_X1 _11312_ ( .A1(_03614_ ), .A2(_03615_ ), .ZN(_03616_ ) );
XNOR2_X1 _11313_ ( .A(_03458_ ), .B(_01928_ ), .ZN(_03617_ ) );
XOR2_X1 _11314_ ( .A(_03457_ ), .B(\IF_ID_pc [27] ), .Z(_03618_ ) );
XOR2_X1 _11315_ ( .A(_03457_ ), .B(\IF_ID_pc [26] ), .Z(_03619_ ) );
NAND4_X1 _11316_ ( .A1(_03616_ ), .A2(_03617_ ), .A3(_03618_ ), .A4(_03619_ ), .ZN(_03620_ ) );
OAI21_X1 _11317_ ( .A(_03458_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_03621_ ) );
INV_X1 _11318_ ( .A(_03621_ ), .ZN(_03622_ ) );
NAND3_X1 _11319_ ( .A1(_03618_ ), .A2(_03617_ ), .A3(_03622_ ), .ZN(_03623_ ) );
NAND2_X1 _11320_ ( .A1(_03458_ ), .A2(\IF_ID_pc [28] ), .ZN(_03624_ ) );
AND2_X1 _11321_ ( .A1(_03458_ ), .A2(\IF_ID_pc [27] ), .ZN(_03625_ ) );
INV_X1 _11322_ ( .A(_03625_ ), .ZN(_03626_ ) );
AND3_X1 _11323_ ( .A1(_03623_ ), .A2(_03624_ ), .A3(_03626_ ), .ZN(_03627_ ) );
AOI21_X1 _11324_ ( .A(_03460_ ), .B1(_03620_ ), .B2(_03627_ ), .ZN(_03628_ ) );
NOR3_X1 _11325_ ( .A1(_03454_ ), .A2(_03481_ ), .A3(_01801_ ), .ZN(_03629_ ) );
OR2_X1 _11326_ ( .A1(_03628_ ), .A2(_03629_ ), .ZN(_03630_ ) );
XNOR2_X1 _11327_ ( .A(_03458_ ), .B(_02013_ ), .ZN(_03631_ ) );
OAI21_X1 _11328_ ( .A(_03451_ ), .B1(_03630_ ), .B2(_03631_ ), .ZN(_03632_ ) );
AOI21_X1 _11329_ ( .A(_03632_ ), .B1(_03630_ ), .B2(_03631_ ), .ZN(_03633_ ) );
BUF_X4 _11330_ ( .A(_03227_ ), .Z(_03634_ ) );
AOI211_X1 _11331_ ( .A(\myifu.to_reset ), .B(_03633_ ), .C1(\myexu.pc_jump [30] ), .C2(_03634_ ), .ZN(_03635_ ) );
BUF_X4 _11332_ ( .A(_03447_ ), .Z(_03636_ ) );
NOR2_X1 _11333_ ( .A1(_03636_ ), .A2(\mtvec [30] ), .ZN(_03637_ ) );
NOR3_X1 _11334_ ( .A1(_03635_ ), .A2(fanout_net_2 ), .A3(_03637_ ), .ZN(_00245_ ) );
BUF_X4 _11335_ ( .A(_03451_ ), .Z(_03638_ ) );
BUF_X4 _11336_ ( .A(_03638_ ), .Z(_03639_ ) );
AND3_X1 _11337_ ( .A1(_03589_ ), .A2(_03605_ ), .A3(_03597_ ), .ZN(_03640_ ) );
AOI21_X1 _11338_ ( .A(_03605_ ), .B1(_03589_ ), .B2(_03597_ ), .ZN(_03641_ ) );
OAI21_X1 _11339_ ( .A(_03639_ ), .B1(_03640_ ), .B2(_03641_ ), .ZN(_03642_ ) );
BUF_X4 _11340_ ( .A(_03638_ ), .Z(_03643_ ) );
OAI211_X1 _11341_ ( .A(_03642_ ), .B(_03636_ ), .C1(\myexu.pc_jump [21] ), .C2(_03643_ ), .ZN(_03644_ ) );
NAND2_X1 _11342_ ( .A1(\mtvec [21] ), .A2(\myifu.to_reset ), .ZN(_03645_ ) );
AOI21_X1 _11343_ ( .A(fanout_net_2 ), .B1(_03644_ ), .B2(_03645_ ), .ZN(_00246_ ) );
AND2_X1 _11344_ ( .A1(_03463_ ), .A2(\IF_ID_pc [19] ), .ZN(_03646_ ) );
NOR2_X1 _11345_ ( .A1(_03572_ ), .A2(_03588_ ), .ZN(_03647_ ) );
INV_X1 _11346_ ( .A(_03647_ ), .ZN(_03648_ ) );
AND2_X1 _11347_ ( .A1(_03648_ ), .A2(_03476_ ), .ZN(_03649_ ) );
NOR2_X1 _11348_ ( .A1(_03649_ ), .A2(_03596_ ), .ZN(_03650_ ) );
INV_X1 _11349_ ( .A(_03650_ ), .ZN(_03651_ ) );
AOI21_X1 _11350_ ( .A(_03646_ ), .B1(_03651_ ), .B2(_03464_ ), .ZN(_03652_ ) );
XNOR2_X1 _11351_ ( .A(_03652_ ), .B(_03465_ ), .ZN(_03653_ ) );
MUX2_X1 _11352_ ( .A(\myexu.pc_jump [20] ), .B(_03653_ ), .S(_03451_ ), .Z(_03654_ ) );
MUX2_X1 _11353_ ( .A(\mtvec [20] ), .B(_03654_ ), .S(_03447_ ), .Z(_03655_ ) );
AND2_X1 _11354_ ( .A1(_03655_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(_00247_ ) );
XNOR2_X1 _11355_ ( .A(_03650_ ), .B(_03464_ ), .ZN(_03656_ ) );
MUX2_X1 _11356_ ( .A(\myexu.pc_jump [19] ), .B(_03656_ ), .S(_03451_ ), .Z(_03657_ ) );
MUX2_X1 _11357_ ( .A(\mtvec [19] ), .B(_03657_ ), .S(_03447_ ), .Z(_03658_ ) );
AND2_X1 _11358_ ( .A1(_03658_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(_00248_ ) );
OAI21_X1 _11359_ ( .A(_03475_ ), .B1(_03572_ ), .B2(_03588_ ), .ZN(_03659_ ) );
INV_X1 _11360_ ( .A(_03593_ ), .ZN(_03660_ ) );
AND2_X1 _11361_ ( .A1(_03659_ ), .A2(_03660_ ), .ZN(_03661_ ) );
XNOR2_X1 _11362_ ( .A(_03661_ ), .B(_03472_ ), .ZN(_03662_ ) );
MUX2_X1 _11363_ ( .A(\myexu.pc_jump [18] ), .B(_03662_ ), .S(_03451_ ), .Z(_03663_ ) );
MUX2_X1 _11364_ ( .A(\mtvec [18] ), .B(_03663_ ), .S(_03447_ ), .Z(_03664_ ) );
AND2_X1 _11365_ ( .A1(_03664_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(_00249_ ) );
XOR2_X1 _11366_ ( .A(_03647_ ), .B(_03475_ ), .Z(_03665_ ) );
NAND2_X1 _11367_ ( .A1(_03665_ ), .A2(_03639_ ), .ZN(_03666_ ) );
BUF_X4 _11368_ ( .A(_03447_ ), .Z(_03667_ ) );
OAI211_X1 _11369_ ( .A(_03666_ ), .B(_03667_ ), .C1(\myexu.pc_jump [17] ), .C2(_03643_ ), .ZN(_03668_ ) );
NAND2_X1 _11370_ ( .A1(\mtvec [17] ), .A2(\myifu.to_reset ), .ZN(_03669_ ) );
AOI21_X1 _11371_ ( .A(fanout_net_2 ), .B1(_03668_ ), .B2(_03669_ ), .ZN(_00250_ ) );
AND2_X1 _11372_ ( .A1(_03568_ ), .A2(_03571_ ), .ZN(_03670_ ) );
OR2_X1 _11373_ ( .A1(_03670_ ), .A2(_03514_ ), .ZN(_03671_ ) );
AOI211_X1 _11374_ ( .A(_03491_ ), .B(_03494_ ), .C1(_03671_ ), .C2(_03581_ ), .ZN(_03672_ ) );
NAND2_X1 _11375_ ( .A1(_03584_ ), .A2(_03585_ ), .ZN(_03673_ ) );
OAI21_X1 _11376_ ( .A(_03480_ ), .B1(_03672_ ), .B2(_03673_ ), .ZN(_03674_ ) );
AND2_X1 _11377_ ( .A1(_03478_ ), .A2(\IF_ID_pc [15] ), .ZN(_03675_ ) );
INV_X1 _11378_ ( .A(_03675_ ), .ZN(_03676_ ) );
AND4_X1 _11379_ ( .A1(_03485_ ), .A2(_03674_ ), .A3(_03486_ ), .A4(_03676_ ), .ZN(_03677_ ) );
AOI22_X1 _11380_ ( .A1(_03674_ ), .A2(_03676_ ), .B1(_03485_ ), .B2(_03486_ ), .ZN(_03678_ ) );
OR3_X1 _11381_ ( .A1(_03677_ ), .A2(_03227_ ), .A3(_03678_ ), .ZN(_03679_ ) );
OAI211_X1 _11382_ ( .A(_03679_ ), .B(_03667_ ), .C1(\myexu.pc_jump [16] ), .C2(_03643_ ), .ZN(_03680_ ) );
NAND2_X1 _11383_ ( .A1(\mtvec [16] ), .A2(\myifu.to_reset ), .ZN(_03681_ ) );
AOI21_X1 _11384_ ( .A(fanout_net_2 ), .B1(_03680_ ), .B2(_03681_ ), .ZN(_00251_ ) );
OR2_X1 _11385_ ( .A1(_03672_ ), .A2(_03673_ ), .ZN(_03682_ ) );
XNOR2_X1 _11386_ ( .A(_03682_ ), .B(_03480_ ), .ZN(_03683_ ) );
NAND2_X1 _11387_ ( .A1(_03683_ ), .A2(_03639_ ), .ZN(_03684_ ) );
OAI211_X1 _11388_ ( .A(_03684_ ), .B(_03667_ ), .C1(\myexu.pc_jump [15] ), .C2(_03643_ ), .ZN(_03685_ ) );
NAND2_X1 _11389_ ( .A1(\mtvec [15] ), .A2(\myifu.to_reset ), .ZN(_03686_ ) );
AOI21_X1 _11390_ ( .A(fanout_net_2 ), .B1(_03685_ ), .B2(_03686_ ), .ZN(_00252_ ) );
AND2_X1 _11391_ ( .A1(_03671_ ), .A2(_03581_ ), .ZN(_03687_ ) );
NOR2_X1 _11392_ ( .A1(_03687_ ), .A2(_03491_ ), .ZN(_03688_ ) );
AND2_X1 _11393_ ( .A1(_03489_ ), .A2(\IF_ID_pc [13] ), .ZN(_03689_ ) );
OAI21_X1 _11394_ ( .A(_03494_ ), .B1(_03688_ ), .B2(_03689_ ), .ZN(_03690_ ) );
OR3_X1 _11395_ ( .A1(_03688_ ), .A2(_03689_ ), .A3(_03494_ ), .ZN(_03691_ ) );
AOI21_X1 _11396_ ( .A(_03227_ ), .B1(_03690_ ), .B2(_03691_ ), .ZN(_03692_ ) );
AOI211_X1 _11397_ ( .A(\myifu.to_reset ), .B(_03692_ ), .C1(\myexu.pc_jump [14] ), .C2(_03634_ ), .ZN(_03693_ ) );
NOR2_X1 _11398_ ( .A1(_03636_ ), .A2(\mtvec [14] ), .ZN(_03694_ ) );
NOR3_X1 _11399_ ( .A1(_03693_ ), .A2(fanout_net_2 ), .A3(_03694_ ), .ZN(_00253_ ) );
OAI21_X1 _11400_ ( .A(_03451_ ), .B1(_03687_ ), .B2(_03491_ ), .ZN(_03695_ ) );
AOI21_X1 _11401_ ( .A(_03695_ ), .B1(_03491_ ), .B2(_03687_ ), .ZN(_03696_ ) );
AOI211_X1 _11402_ ( .A(\myifu.to_reset ), .B(_03696_ ), .C1(\myexu.pc_jump [13] ), .C2(_03634_ ), .ZN(_03697_ ) );
NOR2_X1 _11403_ ( .A1(_03636_ ), .A2(\mtvec [13] ), .ZN(_03698_ ) );
NOR3_X1 _11404_ ( .A1(_03697_ ), .A2(fanout_net_2 ), .A3(_03698_ ), .ZN(_00254_ ) );
AOI211_X1 _11405_ ( .A(_03509_ ), .B(_03513_ ), .C1(_03568_ ), .C2(_03571_ ), .ZN(_03699_ ) );
OAI21_X1 _11406_ ( .A(_03498_ ), .B1(_03699_ ), .B2(_03578_ ), .ZN(_03700_ ) );
NAND2_X1 _11407_ ( .A1(_03497_ ), .A2(\IF_ID_pc [11] ), .ZN(_03701_ ) );
AND2_X1 _11408_ ( .A1(_03700_ ), .A2(_03701_ ), .ZN(_03702_ ) );
AND2_X1 _11409_ ( .A1(_03501_ ), .A2(_03502_ ), .ZN(_03703_ ) );
XNOR2_X1 _11410_ ( .A(_03702_ ), .B(_03703_ ), .ZN(_03704_ ) );
MUX2_X1 _11411_ ( .A(\myexu.pc_jump [12] ), .B(_03704_ ), .S(_03451_ ), .Z(_03705_ ) );
MUX2_X1 _11412_ ( .A(\mtvec [12] ), .B(_03705_ ), .S(_03447_ ), .Z(_03706_ ) );
AND2_X1 _11413_ ( .A1(_03706_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(_00255_ ) );
AND3_X1 _11414_ ( .A1(_03620_ ), .A2(_03627_ ), .A3(_03460_ ), .ZN(_03707_ ) );
OAI21_X1 _11415_ ( .A(_03638_ ), .B1(_03707_ ), .B2(_03628_ ), .ZN(_03708_ ) );
OAI211_X1 _11416_ ( .A(_03708_ ), .B(_03667_ ), .C1(\myexu.pc_jump [29] ), .C2(_03643_ ), .ZN(_03709_ ) );
NAND2_X1 _11417_ ( .A1(\mtvec [29] ), .A2(\myifu.to_reset ), .ZN(_03710_ ) );
AOI21_X1 _11418_ ( .A(fanout_net_2 ), .B1(_03709_ ), .B2(_03710_ ), .ZN(_00256_ ) );
OR3_X1 _11419_ ( .A1(_03699_ ), .A2(_03498_ ), .A3(_03578_ ), .ZN(_03711_ ) );
AND3_X1 _11420_ ( .A1(_03711_ ), .A2(_03638_ ), .A3(_03700_ ), .ZN(_03712_ ) );
AOI211_X1 _11421_ ( .A(\myifu.to_reset ), .B(_03712_ ), .C1(\myexu.pc_jump [11] ), .C2(_03634_ ), .ZN(_03713_ ) );
NOR2_X1 _11422_ ( .A1(_03636_ ), .A2(\mtvec [11] ), .ZN(_03714_ ) );
NOR3_X1 _11423_ ( .A1(_03713_ ), .A2(fanout_net_2 ), .A3(_03714_ ), .ZN(_00257_ ) );
NOR2_X1 _11424_ ( .A1(_03670_ ), .A2(_03509_ ), .ZN(_03715_ ) );
NOR2_X1 _11425_ ( .A1(_03715_ ), .A2(_03576_ ), .ZN(_03716_ ) );
AOI21_X1 _11426_ ( .A(_03227_ ), .B1(_03716_ ), .B2(_03513_ ), .ZN(_03717_ ) );
OR2_X1 _11427_ ( .A1(_03716_ ), .A2(_03513_ ), .ZN(_03718_ ) );
AOI221_X4 _11428_ ( .A(\myifu.to_reset ), .B1(\myexu.pc_jump [10] ), .B2(_03227_ ), .C1(_03717_ ), .C2(_03718_ ), .ZN(_03719_ ) );
NOR2_X1 _11429_ ( .A1(_03636_ ), .A2(\mtvec [10] ), .ZN(_03720_ ) );
NOR3_X1 _11430_ ( .A1(_03719_ ), .A2(fanout_net_2 ), .A3(_03720_ ), .ZN(_00258_ ) );
XNOR2_X1 _11431_ ( .A(_03670_ ), .B(_03508_ ), .ZN(_03721_ ) );
MUX2_X1 _11432_ ( .A(\myexu.pc_jump [9] ), .B(_03721_ ), .S(_03451_ ), .Z(_03722_ ) );
MUX2_X1 _11433_ ( .A(\mtvec [9] ), .B(_03722_ ), .S(_03446_ ), .Z(_03723_ ) );
AND2_X1 _11434_ ( .A1(_03723_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(_00259_ ) );
OAI21_X1 _11435_ ( .A(_03522_ ), .B1(_03561_ ), .B2(_03567_ ), .ZN(_03724_ ) );
INV_X1 _11436_ ( .A(_03570_ ), .ZN(_03725_ ) );
NAND2_X1 _11437_ ( .A1(_03724_ ), .A2(_03725_ ), .ZN(_03726_ ) );
XNOR2_X1 _11438_ ( .A(_03726_ ), .B(_03518_ ), .ZN(_03727_ ) );
NOR2_X1 _11439_ ( .A1(_03727_ ), .A2(_03227_ ), .ZN(_03728_ ) );
AOI211_X1 _11440_ ( .A(\myifu.to_reset ), .B(_03728_ ), .C1(\myexu.pc_jump [8] ), .C2(_03634_ ), .ZN(_03729_ ) );
NOR2_X1 _11441_ ( .A1(_03636_ ), .A2(\mtvec [8] ), .ZN(_03730_ ) );
NOR3_X1 _11442_ ( .A1(_03729_ ), .A2(fanout_net_2 ), .A3(_03730_ ), .ZN(_00260_ ) );
NOR2_X1 _11443_ ( .A1(_03561_ ), .A2(_03567_ ), .ZN(_03731_ ) );
XOR2_X1 _11444_ ( .A(_03731_ ), .B(_03522_ ), .Z(_03732_ ) );
NAND2_X1 _11445_ ( .A1(_03732_ ), .A2(_03639_ ), .ZN(_03733_ ) );
OAI211_X1 _11446_ ( .A(_03733_ ), .B(_03667_ ), .C1(\myexu.pc_jump [7] ), .C2(_03643_ ), .ZN(_03734_ ) );
NAND2_X1 _11447_ ( .A1(\mtvec [7] ), .A2(\myifu.to_reset ), .ZN(_03735_ ) );
AOI21_X1 _11448_ ( .A(fanout_net_2 ), .B1(_03734_ ), .B2(_03735_ ), .ZN(_00261_ ) );
AOI21_X1 _11449_ ( .A(_03528_ ), .B1(_03559_ ), .B2(_03560_ ), .ZN(_03736_ ) );
NOR2_X1 _11450_ ( .A1(_03736_ ), .A2(_03563_ ), .ZN(_03737_ ) );
XNOR2_X1 _11451_ ( .A(_03737_ ), .B(_03533_ ), .ZN(_03738_ ) );
MUX2_X1 _11452_ ( .A(\myexu.pc_jump [6] ), .B(_03738_ ), .S(_03451_ ), .Z(_03739_ ) );
MUX2_X1 _11453_ ( .A(\mtvec [6] ), .B(_03739_ ), .S(_03446_ ), .Z(_03740_ ) );
AND2_X1 _11454_ ( .A1(_03740_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(_00262_ ) );
AND3_X1 _11455_ ( .A1(_03559_ ), .A2(_03560_ ), .A3(_03528_ ), .ZN(_03741_ ) );
OAI21_X1 _11456_ ( .A(_03638_ ), .B1(_03736_ ), .B2(_03741_ ), .ZN(_03742_ ) );
OAI211_X1 _11457_ ( .A(_03742_ ), .B(_03667_ ), .C1(\myexu.pc_jump [5] ), .C2(_03643_ ), .ZN(_03743_ ) );
NAND2_X1 _11458_ ( .A1(\mtvec [5] ), .A2(\myifu.to_reset ), .ZN(_03744_ ) );
AOI21_X1 _11459_ ( .A(fanout_net_2 ), .B1(_03743_ ), .B2(_03744_ ), .ZN(_00263_ ) );
AND2_X1 _11460_ ( .A1(\mtvec [4] ), .A2(\myifu.to_reset ), .ZN(_03745_ ) );
XNOR2_X1 _11461_ ( .A(_03558_ ), .B(fanout_net_11 ), .ZN(_03746_ ) );
XNOR2_X1 _11462_ ( .A(_03554_ ), .B(_03746_ ), .ZN(_03747_ ) );
MUX2_X1 _11463_ ( .A(\myexu.pc_jump [4] ), .B(_03747_ ), .S(_03451_ ), .Z(_03748_ ) );
AOI21_X1 _11464_ ( .A(_03745_ ), .B1(_03748_ ), .B2(_03447_ ), .ZN(_03749_ ) );
NOR2_X1 _11465_ ( .A1(_03749_ ), .A2(fanout_net_2 ), .ZN(_00264_ ) );
XOR2_X1 _11466_ ( .A(_03546_ ), .B(_03551_ ), .Z(_03750_ ) );
MUX2_X1 _11467_ ( .A(\myexu.pc_jump [3] ), .B(_03750_ ), .S(_03450_ ), .Z(_03751_ ) );
AND2_X1 _11468_ ( .A1(_03751_ ), .A2(_03446_ ), .ZN(_03752_ ) );
AOI21_X1 _11469_ ( .A(_03752_ ), .B1(\mtvec [3] ), .B2(\myifu.to_reset ), .ZN(_03753_ ) );
NOR2_X1 _11470_ ( .A1(_03753_ ), .A2(fanout_net_2 ), .ZN(_00265_ ) );
AND2_X1 _11471_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
OAI21_X1 _11472_ ( .A(_01559_ ), .B1(\myifu.pc_$_SDFFE_PP1P__Q_E ), .B2(fanout_net_11 ), .ZN(_03754_ ) );
AOI21_X1 _11473_ ( .A(_03754_ ), .B1(_03749_ ), .B2(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_00266_ ) );
NOR2_X1 _11474_ ( .A1(_03538_ ), .A2(_03543_ ), .ZN(_03755_ ) );
OAI21_X1 _11475_ ( .A(_03638_ ), .B1(_03544_ ), .B2(_03755_ ), .ZN(_03756_ ) );
OAI211_X1 _11476_ ( .A(_03756_ ), .B(_03667_ ), .C1(\myexu.pc_jump [2] ), .C2(_03639_ ), .ZN(_03757_ ) );
NAND2_X1 _11477_ ( .A1(\mtvec [2] ), .A2(\myifu.to_reset ), .ZN(_03758_ ) );
AOI21_X1 _11478_ ( .A(fanout_net_2 ), .B1(_03757_ ), .B2(_03758_ ), .ZN(_00267_ ) );
OAI21_X1 _11479_ ( .A(_01559_ ), .B1(\myifu.pc_$_SDFFE_PP1P__Q_E ), .B2(fanout_net_7 ), .ZN(_03759_ ) );
AOI21_X1 _11480_ ( .A(_03759_ ), .B1(_03753_ ), .B2(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_00268_ ) );
AND3_X1 _11481_ ( .A1(_03614_ ), .A2(_03619_ ), .A3(_03615_ ), .ZN(_03760_ ) );
OAI21_X1 _11482_ ( .A(_03618_ ), .B1(_03760_ ), .B2(_03622_ ), .ZN(_03761_ ) );
AND2_X1 _11483_ ( .A1(_03761_ ), .A2(_03626_ ), .ZN(_03762_ ) );
XNOR2_X1 _11484_ ( .A(_03762_ ), .B(_03617_ ), .ZN(_03763_ ) );
MUX2_X1 _11485_ ( .A(\myexu.pc_jump [28] ), .B(_03763_ ), .S(_03450_ ), .Z(_03764_ ) );
MUX2_X1 _11486_ ( .A(\mtvec [28] ), .B(_03764_ ), .S(_03446_ ), .Z(_03765_ ) );
AND2_X1 _11487_ ( .A1(_03765_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(_00269_ ) );
XNOR2_X1 _11488_ ( .A(_03541_ ), .B(_03542_ ), .ZN(_03766_ ) );
AOI21_X1 _11489_ ( .A(_03766_ ), .B1(check_quest ), .B2(_03445_ ), .ZN(_03767_ ) );
AOI211_X1 _11490_ ( .A(\myifu.to_reset ), .B(_03767_ ), .C1(\myexu.pc_jump [1] ), .C2(_03634_ ), .ZN(_03768_ ) );
NOR2_X1 _11491_ ( .A1(_03636_ ), .A2(\mtvec [1] ), .ZN(_03769_ ) );
NOR3_X1 _11492_ ( .A1(_03768_ ), .A2(fanout_net_2 ), .A3(_03769_ ), .ZN(_00270_ ) );
OAI211_X1 _11493_ ( .A(_03619_ ), .B(_03615_ ), .C1(_03606_ ), .C2(_03612_ ), .ZN(_03770_ ) );
AND2_X1 _11494_ ( .A1(_03770_ ), .A2(_03621_ ), .ZN(_03771_ ) );
XNOR2_X1 _11495_ ( .A(_03771_ ), .B(_03618_ ), .ZN(_03772_ ) );
OR2_X1 _11496_ ( .A1(_03772_ ), .A2(_03227_ ), .ZN(_03773_ ) );
OAI211_X1 _11497_ ( .A(_03773_ ), .B(_03667_ ), .C1(\myexu.pc_jump [27] ), .C2(_03639_ ), .ZN(_03774_ ) );
NAND2_X1 _11498_ ( .A1(\mtvec [27] ), .A2(\myifu.to_reset ), .ZN(_03775_ ) );
AOI21_X1 _11499_ ( .A(fanout_net_2 ), .B1(_03774_ ), .B2(_03775_ ), .ZN(_00271_ ) );
AND2_X1 _11500_ ( .A1(_03458_ ), .A2(\IF_ID_pc [25] ), .ZN(_03776_ ) );
OR3_X1 _11501_ ( .A1(_03616_ ), .A2(_03776_ ), .A3(_03619_ ), .ZN(_03777_ ) );
OAI21_X1 _11502_ ( .A(_03619_ ), .B1(_03616_ ), .B2(_03776_ ), .ZN(_03778_ ) );
AND3_X1 _11503_ ( .A1(_03777_ ), .A2(_03638_ ), .A3(_03778_ ), .ZN(_03779_ ) );
AOI211_X1 _11504_ ( .A(\myifu.to_reset ), .B(_03779_ ), .C1(\myexu.pc_jump [26] ), .C2(_03634_ ), .ZN(_03780_ ) );
NOR2_X1 _11505_ ( .A1(_03636_ ), .A2(\mtvec [26] ), .ZN(_03781_ ) );
NOR3_X1 _11506_ ( .A1(_03780_ ), .A2(reset ), .A3(_03781_ ), .ZN(_00272_ ) );
NOR3_X1 _11507_ ( .A1(_03606_ ), .A2(_03612_ ), .A3(_03615_ ), .ZN(_03782_ ) );
OAI21_X1 _11508_ ( .A(_03638_ ), .B1(_03616_ ), .B2(_03782_ ), .ZN(_03783_ ) );
OAI211_X1 _11509_ ( .A(_03783_ ), .B(_03667_ ), .C1(\myexu.pc_jump [25] ), .C2(_03639_ ), .ZN(_03784_ ) );
NAND2_X1 _11510_ ( .A1(\mtvec [25] ), .A2(\myifu.to_reset ), .ZN(_03785_ ) );
AOI21_X1 _11511_ ( .A(reset ), .B1(_03784_ ), .B2(_03785_ ), .ZN(_00273_ ) );
NOR2_X1 _11512_ ( .A1(_03641_ ), .A2(_03608_ ), .ZN(_03786_ ) );
AOI21_X1 _11513_ ( .A(_03786_ ), .B1(_01980_ ), .B2(_03591_ ), .ZN(_03787_ ) );
OAI21_X1 _11514_ ( .A(_03600_ ), .B1(_03787_ ), .B2(_03607_ ), .ZN(_03788_ ) );
AND3_X1 _11515_ ( .A1(_03788_ ), .A2(_03611_ ), .A3(_03599_ ), .ZN(_03789_ ) );
AOI21_X1 _11516_ ( .A(_03599_ ), .B1(_03788_ ), .B2(_03611_ ), .ZN(_03790_ ) );
OR3_X1 _11517_ ( .A1(_03789_ ), .A2(_03790_ ), .A3(_03227_ ), .ZN(_03791_ ) );
OAI211_X1 _11518_ ( .A(_03791_ ), .B(_03667_ ), .C1(\myexu.pc_jump [24] ), .C2(_03639_ ), .ZN(_03792_ ) );
NAND2_X1 _11519_ ( .A1(\mtvec [24] ), .A2(\myifu.to_reset ), .ZN(_03793_ ) );
AOI21_X1 _11520_ ( .A(reset ), .B1(_03792_ ), .B2(_03793_ ), .ZN(_00274_ ) );
OR3_X1 _11521_ ( .A1(_03787_ ), .A2(_03600_ ), .A3(_03607_ ), .ZN(_03794_ ) );
AND3_X1 _11522_ ( .A1(_03794_ ), .A2(_03638_ ), .A3(_03788_ ), .ZN(_03795_ ) );
AOI211_X1 _11523_ ( .A(\myifu.to_reset ), .B(_03795_ ), .C1(\myexu.pc_jump [23] ), .C2(_03634_ ), .ZN(_03796_ ) );
NOR2_X1 _11524_ ( .A1(_03636_ ), .A2(\mtvec [23] ), .ZN(_03797_ ) );
NOR3_X1 _11525_ ( .A1(_03796_ ), .A2(reset ), .A3(_03797_ ), .ZN(_00275_ ) );
XNOR2_X1 _11526_ ( .A(_03786_ ), .B(_03603_ ), .ZN(_03798_ ) );
NAND2_X1 _11527_ ( .A1(_03798_ ), .A2(_03639_ ), .ZN(_03799_ ) );
OAI211_X1 _11528_ ( .A(_03799_ ), .B(_03447_ ), .C1(\myexu.pc_jump [22] ), .C2(_03639_ ), .ZN(_03800_ ) );
NAND2_X1 _11529_ ( .A1(\mtvec [22] ), .A2(\myifu.to_reset ), .ZN(_03801_ ) );
AOI21_X1 _11530_ ( .A(reset ), .B1(_03800_ ), .B2(_03801_ ), .ZN(_00276_ ) );
NAND2_X1 _11531_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_03802_ ) );
OAI22_X1 _11532_ ( .A1(_03628_ ), .A2(_03629_ ), .B1(\IF_ID_pc [30] ), .B2(_03458_ ), .ZN(_03803_ ) );
NAND2_X1 _11533_ ( .A1(_03458_ ), .A2(\IF_ID_pc [30] ), .ZN(_03804_ ) );
NAND2_X1 _11534_ ( .A1(_03803_ ), .A2(_03804_ ), .ZN(_03805_ ) );
XNOR2_X1 _11535_ ( .A(_03458_ ), .B(\IF_ID_pc [31] ), .ZN(_03806_ ) );
OAI21_X1 _11536_ ( .A(_03638_ ), .B1(_03805_ ), .B2(_03806_ ), .ZN(_03807_ ) );
AOI21_X1 _11537_ ( .A(_03807_ ), .B1(_03805_ ), .B2(_03806_ ), .ZN(_03808_ ) );
OAI21_X1 _11538_ ( .A(_03447_ ), .B1(_03643_ ), .B2(\myexu.pc_jump [31] ), .ZN(_03809_ ) );
OAI211_X1 _11539_ ( .A(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .B(_03802_ ), .C1(_03808_ ), .C2(_03809_ ), .ZN(_00277_ ) );
NOR2_X1 _11540_ ( .A1(_02006_ ), .A2(_02031_ ), .ZN(_03810_ ) );
INV_X1 _11541_ ( .A(_03810_ ), .ZN(_03811_ ) );
NOR2_X1 _11542_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_03812_ ) );
NOR2_X1 _11543_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_03813_ ) );
INV_X1 _11544_ ( .A(\io_master_rid [1] ), .ZN(_03814_ ) );
NAND4_X1 _11545_ ( .A1(_03812_ ), .A2(_03813_ ), .A3(_03814_ ), .A4(\io_master_rid [0] ), .ZN(_03815_ ) );
AOI21_X1 _11546_ ( .A(_01982_ ), .B1(_03811_ ), .B2(_03815_ ), .ZN(_03816_ ) );
AND2_X4 _11547_ ( .A1(_02077_ ), .A2(_02080_ ), .ZN(_03817_ ) );
BUF_X4 _11548_ ( .A(_03817_ ), .Z(_03818_ ) );
BUF_X2 _11549_ ( .A(_03818_ ), .Z(_03819_ ) );
BUF_X2 _11550_ ( .A(_03819_ ), .Z(_03820_ ) );
NOR2_X1 _11551_ ( .A1(_03820_ ), .A2(io_master_rlast ), .ZN(_03821_ ) );
INV_X1 _11552_ ( .A(_03821_ ), .ZN(_03822_ ) );
AND3_X1 _11553_ ( .A1(_02077_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .A3(_02080_ ), .ZN(_03823_ ) );
AOI21_X1 _11554_ ( .A(io_master_rvalid ), .B1(_02077_ ), .B2(_02080_ ), .ZN(_03824_ ) );
NOR2_X1 _11555_ ( .A1(_03823_ ), .A2(_03824_ ), .ZN(_03825_ ) );
NAND3_X1 _11556_ ( .A1(_03816_ ), .A2(_03822_ ), .A3(_03825_ ), .ZN(_03826_ ) );
INV_X1 _11557_ ( .A(\myifu.tmp_offset [2] ), .ZN(_03827_ ) );
AND3_X1 _11558_ ( .A1(_03826_ ), .A2(_01602_ ), .A3(_03827_ ), .ZN(_00278_ ) );
NOR3_X1 _11559_ ( .A1(reset ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00279_ ) );
AND3_X1 _11560_ ( .A1(_02094_ ), .A2(_03228_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_03828_ ) );
INV_X1 _11561_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_03829_ ) );
MUX2_X1 _11562_ ( .A(_02094_ ), .B(_03829_ ), .S(\myifu.to_reset ), .Z(_03830_ ) );
AOI211_X1 _11563_ ( .A(reset ), .B(_03828_ ), .C1(_03830_ ), .C2(\myifu.state [1] ), .ZN(_00280_ ) );
INV_X1 _11564_ ( .A(_02060_ ), .ZN(_03831_ ) );
NOR2_X1 _11565_ ( .A1(_02068_ ), .A2(_03831_ ), .ZN(_03832_ ) );
INV_X1 _11566_ ( .A(_03832_ ), .ZN(_03833_ ) );
BUF_X2 _11567_ ( .A(_03833_ ), .Z(_03834_ ) );
BUF_X4 _11568_ ( .A(_02128_ ), .Z(_03835_ ) );
MUX2_X1 _11569_ ( .A(\LS_WB_waddr_csreg [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_03835_ ), .Z(_03836_ ) );
BUF_X4 _11570_ ( .A(_02059_ ), .Z(_03837_ ) );
NOR2_X1 _11571_ ( .A1(\EX_LS_flag [2] ), .A2(\EX_LS_flag [1] ), .ZN(_03838_ ) );
NOR2_X1 _11572_ ( .A1(_03837_ ), .A2(_03838_ ), .ZN(_03839_ ) );
NOR2_X1 _11573_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_03840_ ) );
AND2_X2 _11574_ ( .A1(_03840_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_03841_ ) );
NOR2_X1 _11575_ ( .A1(_03839_ ), .A2(_03841_ ), .ZN(_03842_ ) );
BUF_X4 _11576_ ( .A(_03842_ ), .Z(_03843_ ) );
BUF_X2 _11577_ ( .A(_03843_ ), .Z(_03844_ ) );
AND3_X1 _11578_ ( .A1(_03834_ ), .A2(_03836_ ), .A3(_03844_ ), .ZN(_00283_ ) );
NOR2_X1 _11579_ ( .A1(_02041_ ), .A2(_03841_ ), .ZN(_03845_ ) );
AND2_X1 _11580_ ( .A1(_03833_ ), .A2(_03845_ ), .ZN(_03846_ ) );
INV_X1 _11581_ ( .A(_03846_ ), .ZN(_03847_ ) );
NAND3_X1 _11582_ ( .A1(_03837_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_03848_ ) );
BUF_X4 _11583_ ( .A(_02025_ ), .Z(_03849_ ) );
NAND2_X1 _11584_ ( .A1(_03849_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03850_ ) );
AOI21_X1 _11585_ ( .A(_03847_ ), .B1(_03848_ ), .B2(_03850_ ), .ZN(_00284_ ) );
NAND3_X1 _11586_ ( .A1(_03837_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_03851_ ) );
NAND2_X1 _11587_ ( .A1(_03849_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_03852_ ) );
AOI21_X1 _11588_ ( .A(_03847_ ), .B1(_03851_ ), .B2(_03852_ ), .ZN(_00285_ ) );
NAND3_X1 _11589_ ( .A1(_03837_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_03853_ ) );
NAND2_X1 _11590_ ( .A1(_03849_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_03854_ ) );
AOI21_X1 _11591_ ( .A(_03847_ ), .B1(_03853_ ), .B2(_03854_ ), .ZN(_00286_ ) );
NAND3_X1 _11592_ ( .A1(_03837_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_03855_ ) );
NAND2_X1 _11593_ ( .A1(_03849_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03856_ ) );
AOI21_X1 _11594_ ( .A(_03847_ ), .B1(_03855_ ), .B2(_03856_ ), .ZN(_00287_ ) );
NAND3_X1 _11595_ ( .A1(_03837_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_03857_ ) );
NAND2_X1 _11596_ ( .A1(_03849_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_03858_ ) );
AOI21_X1 _11597_ ( .A(_03847_ ), .B1(_03857_ ), .B2(_03858_ ), .ZN(_00288_ ) );
NAND3_X1 _11598_ ( .A1(_03837_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_03859_ ) );
NAND2_X1 _11599_ ( .A1(_03849_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_03860_ ) );
AOI21_X1 _11600_ ( .A(_03847_ ), .B1(_03859_ ), .B2(_03860_ ), .ZN(_00289_ ) );
NAND3_X1 _11601_ ( .A1(_03837_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_flag [2] ), .ZN(_03861_ ) );
NAND2_X1 _11602_ ( .A1(_03849_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_03862_ ) );
AOI21_X1 _11603_ ( .A(_03847_ ), .B1(_03861_ ), .B2(_03862_ ), .ZN(_00290_ ) );
NOR4_X1 _11604_ ( .A1(_03849_ ), .A2(_02058_ ), .A3(\EX_LS_dest_csreg_mem [9] ), .A4(\EX_LS_flag [0] ), .ZN(_03863_ ) );
NOR2_X1 _11605_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_03864_ ) );
OAI221_X1 _11606_ ( .A(_03845_ ), .B1(_03863_ ), .B2(_03864_ ), .C1(_02068_ ), .C2(_03831_ ), .ZN(_00291_ ) );
NOR4_X1 _11607_ ( .A1(_03849_ ), .A2(_02058_ ), .A3(\EX_LS_dest_csreg_mem [8] ), .A4(\EX_LS_flag [0] ), .ZN(_03865_ ) );
NOR2_X1 _11608_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_03866_ ) );
OAI221_X1 _11609_ ( .A(_03845_ ), .B1(_03865_ ), .B2(_03866_ ), .C1(_02068_ ), .C2(_03831_ ), .ZN(_00292_ ) );
NOR4_X1 _11610_ ( .A1(_03849_ ), .A2(_02058_ ), .A3(\EX_LS_dest_csreg_mem [6] ), .A4(\EX_LS_flag [0] ), .ZN(_03867_ ) );
NOR2_X1 _11611_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_03868_ ) );
OAI221_X1 _11612_ ( .A(_03845_ ), .B1(_03867_ ), .B2(_03868_ ), .C1(_02068_ ), .C2(_03831_ ), .ZN(_00293_ ) );
NOR4_X1 _11613_ ( .A1(_02025_ ), .A2(_02058_ ), .A3(fanout_net_3 ), .A4(\EX_LS_flag [0] ), .ZN(_03869_ ) );
NOR2_X1 _11614_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_03870_ ) );
OAI221_X1 _11615_ ( .A(_03845_ ), .B1(_03869_ ), .B2(_03870_ ), .C1(_02068_ ), .C2(_03831_ ), .ZN(_00294_ ) );
INV_X1 _11616_ ( .A(\mysc.state [2] ), .ZN(_03871_ ) );
NOR2_X1 _11617_ ( .A1(_03871_ ), .A2(reset ), .ZN(_00302_ ) );
INV_X1 _11618_ ( .A(\ID_EX_typ [6] ), .ZN(_03872_ ) );
NAND2_X1 _11619_ ( .A1(_03872_ ), .A2(\ID_EX_typ [7] ), .ZN(_03873_ ) );
OR3_X1 _11620_ ( .A1(_03873_ ), .A2(\ID_EX_typ [5] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03874_ ) );
INV_X1 _11621_ ( .A(\ID_EX_typ [5] ), .ZN(_03875_ ) );
NOR2_X1 _11622_ ( .A1(_03873_ ), .A2(_03875_ ), .ZN(_03876_ ) );
BUF_X4 _11623_ ( .A(_03876_ ), .Z(_03877_ ) );
INV_X2 _11624_ ( .A(_03877_ ), .ZN(_03878_ ) );
BUF_X4 _11625_ ( .A(_03878_ ), .Z(_03879_ ) );
OAI21_X1 _11626_ ( .A(_03874_ ), .B1(_03879_ ), .B2(fanout_net_4 ), .ZN(_03880_ ) );
NOR2_X1 _11627_ ( .A1(_03345_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
NAND2_X1 _11628_ ( .A1(_03880_ ), .A2(\myexu.state_$_ANDNOT__B_Y ), .ZN(_03881_ ) );
INV_X1 _11629_ ( .A(\myec.state [1] ), .ZN(_03882_ ) );
NAND2_X1 _11630_ ( .A1(_03882_ ), .A2(\myec.state [0] ), .ZN(_03883_ ) );
AND2_X2 _11631_ ( .A1(_03883_ ), .A2(_03067_ ), .ZN(_03884_ ) );
BUF_X4 _11632_ ( .A(_03884_ ), .Z(_03885_ ) );
INV_X1 _11633_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_03886_ ) );
OAI22_X1 _11634_ ( .A1(_03886_ ), .A2(_03873_ ), .B1(_03226_ ), .B2(check_assert ), .ZN(_03887_ ) );
AND3_X1 _11635_ ( .A1(_03881_ ), .A2(_03885_ ), .A3(_03887_ ), .ZN(_00095_ ) );
CLKBUF_X2 _11636_ ( .A(_03883_ ), .Z(_03888_ ) );
CLKBUF_X2 _11637_ ( .A(_03888_ ), .Z(_03889_ ) );
AND3_X1 _11638_ ( .A1(_03889_ ), .A2(\ID_EX_rd [4] ), .A3(_03100_ ), .ZN(_00116_ ) );
AND3_X1 _11639_ ( .A1(_03889_ ), .A2(\ID_EX_rd [3] ), .A3(_03100_ ), .ZN(_00117_ ) );
AND3_X1 _11640_ ( .A1(_03889_ ), .A2(\ID_EX_rd [2] ), .A3(_03100_ ), .ZN(_00118_ ) );
AND3_X1 _11641_ ( .A1(_03889_ ), .A2(\ID_EX_rd [1] ), .A3(_03100_ ), .ZN(_00119_ ) );
AND3_X1 _11642_ ( .A1(_03889_ ), .A2(\ID_EX_rd [0] ), .A3(_03100_ ), .ZN(_00120_ ) );
INV_X2 _11643_ ( .A(_03885_ ), .ZN(_03890_ ) );
BUF_X4 _11644_ ( .A(_03890_ ), .Z(_03891_ ) );
XNOR2_X1 _11645_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_03892_ ) );
XNOR2_X1 _11646_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_03893_ ) );
XNOR2_X1 _11647_ ( .A(\EX_LS_dest_csreg_mem [1] ), .B(\ID_EX_csr [1] ), .ZN(_03894_ ) );
XNOR2_X1 _11648_ ( .A(fanout_net_3 ), .B(\ID_EX_csr [0] ), .ZN(_03895_ ) );
AND4_X1 _11649_ ( .A1(_03892_ ), .A2(_03893_ ), .A3(_03894_ ), .A4(_03895_ ), .ZN(_03896_ ) );
XOR2_X1 _11650_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .Z(_03897_ ) );
INV_X1 _11651_ ( .A(_02059_ ), .ZN(_03898_ ) );
NOR3_X1 _11652_ ( .A1(_03897_ ), .A2(_02025_ ), .A3(_03898_ ), .ZN(_03899_ ) );
XNOR2_X1 _11653_ ( .A(\EX_LS_dest_csreg_mem [8] ), .B(\ID_EX_csr [8] ), .ZN(_03900_ ) );
XNOR2_X1 _11654_ ( .A(\EX_LS_dest_csreg_mem [9] ), .B(\ID_EX_csr [9] ), .ZN(_03901_ ) );
NAND4_X1 _11655_ ( .A1(_03896_ ), .A2(_03899_ ), .A3(_03900_ ), .A4(_03901_ ), .ZN(_03902_ ) );
XNOR2_X1 _11656_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_03903_ ) );
XNOR2_X1 _11657_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_03904_ ) );
XNOR2_X1 _11658_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_03905_ ) );
AND3_X1 _11659_ ( .A1(_03903_ ), .A2(_03904_ ), .A3(_03905_ ), .ZN(_03906_ ) );
INV_X1 _11660_ ( .A(\EX_LS_dest_csreg_mem [3] ), .ZN(_03907_ ) );
NAND2_X1 _11661_ ( .A1(_03907_ ), .A2(\ID_EX_csr [3] ), .ZN(_03908_ ) );
INV_X1 _11662_ ( .A(\ID_EX_csr [3] ), .ZN(_03909_ ) );
NAND2_X1 _11663_ ( .A1(_03909_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .ZN(_03910_ ) );
XNOR2_X1 _11664_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_03911_ ) );
NAND4_X1 _11665_ ( .A1(_03906_ ), .A2(_03908_ ), .A3(_03910_ ), .A4(_03911_ ), .ZN(_03912_ ) );
NOR2_X1 _11666_ ( .A1(_03902_ ), .A2(_03912_ ), .ZN(_03913_ ) );
INV_X1 _11667_ ( .A(_03913_ ), .ZN(_03914_ ) );
INV_X1 _11668_ ( .A(\ID_EX_csr [1] ), .ZN(_03915_ ) );
NOR2_X1 _11669_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_03916_ ) );
NOR2_X1 _11670_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_03917_ ) );
AND2_X1 _11671_ ( .A1(_03916_ ), .A2(_03917_ ), .ZN(_03918_ ) );
BUF_X4 _11672_ ( .A(_03918_ ), .Z(_03919_ ) );
AND4_X2 _11673_ ( .A1(_03915_ ), .A2(_03919_ ), .A3(\ID_EX_csr [0] ), .A4(_03909_ ), .ZN(_03920_ ) );
INV_X1 _11674_ ( .A(\ID_EX_csr [11] ), .ZN(_03921_ ) );
NAND3_X1 _11675_ ( .A1(_03921_ ), .A2(\ID_EX_csr [9] ), .A3(\ID_EX_csr [8] ), .ZN(_03922_ ) );
NOR2_X1 _11676_ ( .A1(_03922_ ), .A2(\ID_EX_csr [10] ), .ZN(_03923_ ) );
BUF_X4 _11677_ ( .A(_03923_ ), .Z(_03924_ ) );
NAND4_X1 _11678_ ( .A1(_03920_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [30] ), .A4(_03924_ ), .ZN(_03925_ ) );
INV_X1 _11679_ ( .A(\ID_EX_csr [7] ), .ZN(_03926_ ) );
NAND3_X1 _11680_ ( .A1(_03917_ ), .A2(_03926_ ), .A3(\ID_EX_csr [6] ), .ZN(_03927_ ) );
NOR3_X2 _11681_ ( .A1(_03927_ ), .A2(\ID_EX_csr [10] ), .A3(_03922_ ), .ZN(_03928_ ) );
BUF_X4 _11682_ ( .A(_03928_ ), .Z(_03929_ ) );
NAND3_X1 _11683_ ( .A1(_03915_ ), .A2(_03909_ ), .A3(\ID_EX_csr [0] ), .ZN(_03930_ ) );
NOR2_X2 _11684_ ( .A1(_03930_ ), .A2(\ID_EX_csr [2] ), .ZN(_03931_ ) );
BUF_X4 _11685_ ( .A(_03931_ ), .Z(_03932_ ) );
NAND3_X1 _11686_ ( .A1(_03929_ ), .A2(\mepc [30] ), .A3(_03932_ ), .ZN(_03933_ ) );
NOR2_X1 _11687_ ( .A1(\ID_EX_csr [3] ), .A2(\ID_EX_csr [2] ), .ZN(_03934_ ) );
INV_X1 _11688_ ( .A(\ID_EX_csr [0] ), .ZN(_03935_ ) );
AND3_X2 _11689_ ( .A1(_03934_ ), .A2(_03915_ ), .A3(_03935_ ), .ZN(_03936_ ) );
AND2_X2 _11690_ ( .A1(_03936_ ), .A2(_03919_ ), .ZN(_03937_ ) );
BUF_X2 _11691_ ( .A(_03923_ ), .Z(_03938_ ) );
NAND3_X1 _11692_ ( .A1(_03937_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_03938_ ), .ZN(_03939_ ) );
AND3_X1 _11693_ ( .A1(_03925_ ), .A2(_03933_ ), .A3(_03939_ ), .ZN(_03940_ ) );
INV_X1 _11694_ ( .A(\ID_EX_csr [2] ), .ZN(_03941_ ) );
NAND3_X1 _11695_ ( .A1(_03909_ ), .A2(_03941_ ), .A3(\ID_EX_csr [1] ), .ZN(_03942_ ) );
NOR2_X2 _11696_ ( .A1(_03942_ ), .A2(\ID_EX_csr [0] ), .ZN(_03943_ ) );
AND2_X1 _11697_ ( .A1(_03928_ ), .A2(_03943_ ), .ZN(_03944_ ) );
BUF_X4 _11698_ ( .A(_03931_ ), .Z(_03945_ ) );
AND2_X1 _11699_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_03946_ ) );
AND3_X1 _11700_ ( .A1(_03946_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_03947_ ) );
INV_X1 _11701_ ( .A(\ID_EX_csr [5] ), .ZN(_03948_ ) );
AND3_X1 _11702_ ( .A1(_03916_ ), .A2(_03948_ ), .A3(\ID_EX_csr [4] ), .ZN(_03949_ ) );
AND2_X1 _11703_ ( .A1(_03947_ ), .A2(_03949_ ), .ZN(_03950_ ) );
AOI22_X1 _11704_ ( .A1(_03944_ ), .A2(\mycsreg.CSReg[3][30] ), .B1(_03945_ ), .B2(_03950_ ), .ZN(_03951_ ) );
NAND3_X1 _11705_ ( .A1(_03914_ ), .A2(_03940_ ), .A3(_03951_ ), .ZN(_03952_ ) );
OR3_X1 _11706_ ( .A1(_03902_ ), .A2(_03912_ ), .A3(\EX_LS_result_csreg_mem [30] ), .ZN(_03953_ ) );
AND2_X1 _11707_ ( .A1(_03952_ ), .A2(_03953_ ), .ZN(_03954_ ) );
AND2_X1 _11708_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_03955_ ) );
AND2_X1 _11709_ ( .A1(_03955_ ), .A2(\ID_EX_pc [4] ), .ZN(_03956_ ) );
AND2_X1 _11710_ ( .A1(_03956_ ), .A2(\ID_EX_pc [5] ), .ZN(_03957_ ) );
AND2_X1 _11711_ ( .A1(_03957_ ), .A2(\ID_EX_pc [6] ), .ZN(_03958_ ) );
AND2_X1 _11712_ ( .A1(_03958_ ), .A2(\ID_EX_pc [7] ), .ZN(_03959_ ) );
AND2_X1 _11713_ ( .A1(_03959_ ), .A2(\ID_EX_pc [8] ), .ZN(_03960_ ) );
AND2_X2 _11714_ ( .A1(_03960_ ), .A2(\ID_EX_pc [9] ), .ZN(_03961_ ) );
AND2_X1 _11715_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_03962_ ) );
AND2_X1 _11716_ ( .A1(_03961_ ), .A2(_03962_ ), .ZN(_03963_ ) );
AND3_X1 _11717_ ( .A1(_03963_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_03964_ ) );
AND3_X1 _11718_ ( .A1(_03964_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_03965_ ) );
AND3_X1 _11719_ ( .A1(_03965_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_03966_ ) );
AND3_X1 _11720_ ( .A1(_03966_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_03967_ ) );
AND3_X1 _11721_ ( .A1(_03967_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_03968_ ) );
AND3_X1 _11722_ ( .A1(_03968_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_03969_ ) );
AND3_X1 _11723_ ( .A1(_03969_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_03970_ ) );
AND3_X1 _11724_ ( .A1(_03970_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_03971_ ) );
NAND3_X1 _11725_ ( .A1(_03971_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_03972_ ) );
XNOR2_X1 _11726_ ( .A(_03972_ ), .B(\ID_EX_pc [30] ), .ZN(_03973_ ) );
NOR2_X1 _11727_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_03974_ ) );
XOR2_X1 _11728_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_03975_ ) );
XOR2_X1 _11729_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_03976_ ) );
AND2_X1 _11730_ ( .A1(_03975_ ), .A2(_03976_ ), .ZN(_03977_ ) );
XOR2_X1 _11731_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_03978_ ) );
AND2_X1 _11732_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_03979_ ) );
NOR2_X1 _11733_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_03980_ ) );
NOR2_X1 _11734_ ( .A1(_03979_ ), .A2(_03980_ ), .ZN(_03981_ ) );
AND2_X1 _11735_ ( .A1(_03978_ ), .A2(_03981_ ), .ZN(_03982_ ) );
AND2_X1 _11736_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03983_ ) );
NOR2_X1 _11737_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03984_ ) );
XOR2_X1 _11738_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_03985_ ) );
XOR2_X1 _11739_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_03986_ ) );
AND2_X1 _11740_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_03987_ ) );
AND2_X1 _11741_ ( .A1(_03986_ ), .A2(_03987_ ), .ZN(_03988_ ) );
AND2_X1 _11742_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_03989_ ) );
OAI21_X1 _11743_ ( .A(_03985_ ), .B1(_03988_ ), .B2(_03989_ ), .ZN(_03990_ ) );
NAND2_X1 _11744_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_03991_ ) );
AOI21_X1 _11745_ ( .A(_03984_ ), .B1(_03990_ ), .B2(_03991_ ), .ZN(_03992_ ) );
AND2_X1 _11746_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03993_ ) );
OR2_X1 _11747_ ( .A1(_03992_ ), .A2(_03993_ ), .ZN(_03994_ ) );
XOR2_X1 _11748_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_03995_ ) );
AOI221_X4 _11749_ ( .A(_03983_ ), .B1(\ID_EX_pc [5] ), .B2(\ID_EX_imm [5] ), .C1(_03994_ ), .C2(_03995_ ), .ZN(_03996_ ) );
NOR2_X1 _11750_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03997_ ) );
NOR2_X1 _11751_ ( .A1(_03996_ ), .A2(_03997_ ), .ZN(_03998_ ) );
XOR2_X1 _11752_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_03999_ ) );
NAND2_X1 _11753_ ( .A1(_03998_ ), .A2(_03999_ ), .ZN(_04000_ ) );
NAND2_X1 _11754_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_04001_ ) );
NAND2_X1 _11755_ ( .A1(_04000_ ), .A2(_04001_ ), .ZN(_04002_ ) );
OAI21_X1 _11756_ ( .A(_04002_ ), .B1(\ID_EX_pc [7] ), .B2(\ID_EX_imm [7] ), .ZN(_04003_ ) );
AND2_X1 _11757_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04004_ ) );
INV_X1 _11758_ ( .A(_04004_ ), .ZN(_04005_ ) );
NAND2_X1 _11759_ ( .A1(_04003_ ), .A2(_04005_ ), .ZN(_04006_ ) );
XOR2_X1 _11760_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_04007_ ) );
XOR2_X1 _11761_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_04008_ ) );
NAND2_X1 _11762_ ( .A1(_04007_ ), .A2(_04008_ ), .ZN(_04009_ ) );
XOR2_X1 _11763_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_04010_ ) );
INV_X1 _11764_ ( .A(_04010_ ), .ZN(_04011_ ) );
XNOR2_X1 _11765_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .ZN(_04012_ ) );
NOR3_X1 _11766_ ( .A1(_04009_ ), .A2(_04011_ ), .A3(_04012_ ), .ZN(_04013_ ) );
XOR2_X1 _11767_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_04014_ ) );
XOR2_X1 _11768_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_04015_ ) );
AND2_X1 _11769_ ( .A1(_04014_ ), .A2(_04015_ ), .ZN(_04016_ ) );
XOR2_X1 _11770_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_04017_ ) );
XOR2_X1 _11771_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_04018_ ) );
AND2_X1 _11772_ ( .A1(_04017_ ), .A2(_04018_ ), .ZN(_04019_ ) );
AND2_X1 _11773_ ( .A1(_04016_ ), .A2(_04019_ ), .ZN(_04020_ ) );
NAND3_X1 _11774_ ( .A1(_04006_ ), .A2(_04013_ ), .A3(_04020_ ), .ZN(_04021_ ) );
AND2_X1 _11775_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_04022_ ) );
AND2_X1 _11776_ ( .A1(_04014_ ), .A2(_04022_ ), .ZN(_04023_ ) );
AOI21_X1 _11777_ ( .A(_04023_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_04024_ ) );
AND2_X1 _11778_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_04025_ ) );
AND2_X1 _11779_ ( .A1(_04018_ ), .A2(_04025_ ), .ZN(_04026_ ) );
AOI21_X1 _11780_ ( .A(_04026_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_04027_ ) );
INV_X1 _11781_ ( .A(_04016_ ), .ZN(_04028_ ) );
OAI21_X1 _11782_ ( .A(_04024_ ), .B1(_04027_ ), .B2(_04028_ ), .ZN(_04029_ ) );
AND2_X1 _11783_ ( .A1(_04029_ ), .A2(_04013_ ), .ZN(_04030_ ) );
AND2_X1 _11784_ ( .A1(\ID_EX_pc [15] ), .A2(\ID_EX_imm [15] ), .ZN(_04031_ ) );
NAND2_X1 _11785_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_04032_ ) );
NOR2_X1 _11786_ ( .A1(_04012_ ), .A2(_04032_ ), .ZN(_04033_ ) );
AOI21_X1 _11787_ ( .A(_04033_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_04034_ ) );
NOR2_X1 _11788_ ( .A1(_04034_ ), .A2(_04009_ ), .ZN(_04035_ ) );
AND2_X1 _11789_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04036_ ) );
AND2_X1 _11790_ ( .A1(_04007_ ), .A2(_04036_ ), .ZN(_04037_ ) );
NOR4_X1 _11791_ ( .A1(_04030_ ), .A2(_04031_ ), .A3(_04035_ ), .A4(_04037_ ), .ZN(_04038_ ) );
AND2_X1 _11792_ ( .A1(_04021_ ), .A2(_04038_ ), .ZN(_04039_ ) );
XOR2_X1 _11793_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_04040_ ) );
XOR2_X1 _11794_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_04041_ ) );
NAND2_X1 _11795_ ( .A1(_04040_ ), .A2(_04041_ ), .ZN(_04042_ ) );
XOR2_X1 _11796_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_04043_ ) );
INV_X1 _11797_ ( .A(_04043_ ), .ZN(_04044_ ) );
XNOR2_X1 _11798_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .ZN(_04045_ ) );
NOR2_X1 _11799_ ( .A1(_04044_ ), .A2(_04045_ ), .ZN(_04046_ ) );
INV_X1 _11800_ ( .A(_04046_ ), .ZN(_04047_ ) );
XOR2_X1 _11801_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_04048_ ) );
XOR2_X1 _11802_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_04049_ ) );
AND2_X1 _11803_ ( .A1(_04048_ ), .A2(_04049_ ), .ZN(_04050_ ) );
XOR2_X1 _11804_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_04051_ ) );
XOR2_X1 _11805_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_04052_ ) );
NAND3_X1 _11806_ ( .A1(_04050_ ), .A2(_04051_ ), .A3(_04052_ ), .ZN(_04053_ ) );
NOR4_X1 _11807_ ( .A1(_04039_ ), .A2(_04042_ ), .A3(_04047_ ), .A4(_04053_ ), .ZN(_04054_ ) );
AND2_X1 _11808_ ( .A1(\ID_EX_pc [23] ), .A2(\ID_EX_imm [23] ), .ZN(_04055_ ) );
AND2_X1 _11809_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_04056_ ) );
AND2_X1 _11810_ ( .A1(_04051_ ), .A2(_04056_ ), .ZN(_04057_ ) );
AOI21_X1 _11811_ ( .A(_04057_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_04058_ ) );
INV_X1 _11812_ ( .A(_04058_ ), .ZN(_04059_ ) );
AND2_X1 _11813_ ( .A1(_04059_ ), .A2(_04050_ ), .ZN(_04060_ ) );
AND2_X1 _11814_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_imm [19] ), .ZN(_04061_ ) );
AND2_X1 _11815_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_04062_ ) );
AND2_X1 _11816_ ( .A1(_04048_ ), .A2(_04062_ ), .ZN(_04063_ ) );
NOR3_X1 _11817_ ( .A1(_04060_ ), .A2(_04061_ ), .A3(_04063_ ), .ZN(_04064_ ) );
NOR3_X1 _11818_ ( .A1(_04064_ ), .A2(_04042_ ), .A3(_04047_ ), .ZN(_04065_ ) );
NAND2_X1 _11819_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_04066_ ) );
NOR2_X1 _11820_ ( .A1(_04045_ ), .A2(_04066_ ), .ZN(_04067_ ) );
AOI21_X1 _11821_ ( .A(_04067_ ), .B1(\ID_EX_pc [21] ), .B2(\ID_EX_imm [21] ), .ZN(_04068_ ) );
NOR2_X1 _11822_ ( .A1(_04068_ ), .A2(_04042_ ), .ZN(_04069_ ) );
AND2_X1 _11823_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_04070_ ) );
AND2_X1 _11824_ ( .A1(_04040_ ), .A2(_04070_ ), .ZN(_04071_ ) );
OR4_X1 _11825_ ( .A1(_04055_ ), .A2(_04065_ ), .A3(_04069_ ), .A4(_04071_ ), .ZN(_04072_ ) );
OAI211_X1 _11826_ ( .A(_03977_ ), .B(_03982_ ), .C1(_04054_ ), .C2(_04072_ ), .ZN(_04073_ ) );
AND3_X1 _11827_ ( .A1(_03975_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_04074_ ) );
NAND2_X1 _11828_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_04075_ ) );
OR3_X1 _11829_ ( .A1(_03979_ ), .A2(_03980_ ), .A3(_04075_ ), .ZN(_04076_ ) );
INV_X1 _11830_ ( .A(\ID_EX_pc [25] ), .ZN(_04077_ ) );
OAI21_X1 _11831_ ( .A(_04076_ ), .B1(_04077_ ), .B2(_02939_ ), .ZN(_04078_ ) );
AOI221_X4 _11832_ ( .A(_04074_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .C1(_03977_ ), .C2(_04078_ ), .ZN(_04079_ ) );
NAND2_X1 _11833_ ( .A1(_04073_ ), .A2(_04079_ ), .ZN(_04080_ ) );
XOR2_X1 _11834_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_04081_ ) );
NAND2_X1 _11835_ ( .A1(_04080_ ), .A2(_04081_ ), .ZN(_04082_ ) );
NAND2_X1 _11836_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_04083_ ) );
AOI21_X1 _11837_ ( .A(_03974_ ), .B1(_04082_ ), .B2(_04083_ ), .ZN(_04084_ ) );
AND2_X1 _11838_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_04085_ ) );
OR2_X1 _11839_ ( .A1(_04084_ ), .A2(_04085_ ), .ZN(_04086_ ) );
XOR2_X1 _11840_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_04087_ ) );
XOR2_X1 _11841_ ( .A(_04086_ ), .B(_04087_ ), .Z(_04088_ ) );
NOR2_X1 _11842_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_4 ), .ZN(_04089_ ) );
AND2_X1 _11843_ ( .A1(_04089_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04090_ ) );
INV_X1 _11844_ ( .A(_04090_ ), .ZN(_04091_ ) );
XOR2_X2 _11845_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .Z(_04092_ ) );
INV_X2 _11846_ ( .A(_04092_ ), .ZN(_04093_ ) );
XNOR2_X1 _11847_ ( .A(\EX_LS_dest_reg [3] ), .B(\ID_EX_rs2 [3] ), .ZN(_04094_ ) );
XNOR2_X1 _11848_ ( .A(\EX_LS_dest_reg [1] ), .B(\ID_EX_rs2 [1] ), .ZN(_04095_ ) );
XNOR2_X1 _11849_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_04096_ ) );
XNOR2_X1 _11850_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_04097_ ) );
AND4_X1 _11851_ ( .A1(_04094_ ), .A2(_04095_ ), .A3(_04096_ ), .A4(_04097_ ), .ZN(_04098_ ) );
NAND4_X4 _11852_ ( .A1(_02130_ ), .A2(_02135_ ), .A3(_04093_ ), .A4(_04098_ ), .ZN(_04099_ ) );
BUF_X8 _11853_ ( .A(_04099_ ), .Z(_04100_ ) );
INV_X1 _11854_ ( .A(\EX_LS_result_reg [9] ), .ZN(_04101_ ) );
INV_X1 _11855_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .ZN(_04102_ ) );
BUF_X2 _11856_ ( .A(_04102_ ), .Z(_04103_ ) );
OR3_X1 _11857_ ( .A1(_04100_ ), .A2(_04101_ ), .A3(_04103_ ), .ZN(_04104_ ) );
INV_X1 _11858_ ( .A(fanout_net_40 ), .ZN(_04105_ ) );
BUF_X4 _11859_ ( .A(_04105_ ), .Z(_04106_ ) );
INV_X1 _11860_ ( .A(fanout_net_28 ), .ZN(_04107_ ) );
CLKBUF_X2 _11861_ ( .A(_04107_ ), .Z(_04108_ ) );
OR2_X1 _11862_ ( .A1(_04108_ ), .A2(\myreg.Reg[1][9] ), .ZN(_04109_ ) );
INV_X1 _11863_ ( .A(fanout_net_36 ), .ZN(_04110_ ) );
BUF_X4 _11864_ ( .A(_04110_ ), .Z(_04111_ ) );
BUF_X4 _11865_ ( .A(_04111_ ), .Z(_04112_ ) );
OAI211_X1 _11866_ ( .A(_04109_ ), .B(_04112_ ), .C1(fanout_net_28 ), .C2(\myreg.Reg[0][9] ), .ZN(_04113_ ) );
INV_X1 _11867_ ( .A(fanout_net_39 ), .ZN(_04114_ ) );
BUF_X4 _11868_ ( .A(_04114_ ), .Z(_04115_ ) );
OR2_X1 _11869_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[2][9] ), .ZN(_04116_ ) );
BUF_X2 _11870_ ( .A(_04107_ ), .Z(_04117_ ) );
BUF_X2 _11871_ ( .A(_04117_ ), .Z(_04118_ ) );
OAI211_X1 _11872_ ( .A(_04116_ ), .B(fanout_net_36 ), .C1(_04118_ ), .C2(\myreg.Reg[3][9] ), .ZN(_04119_ ) );
NAND3_X1 _11873_ ( .A1(_04113_ ), .A2(_04115_ ), .A3(_04119_ ), .ZN(_04120_ ) );
MUX2_X1 _11874_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_28 ), .Z(_04121_ ) );
MUX2_X1 _11875_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_28 ), .Z(_04122_ ) );
BUF_X4 _11876_ ( .A(_04111_ ), .Z(_04123_ ) );
MUX2_X1 _11877_ ( .A(_04121_ ), .B(_04122_ ), .S(_04123_ ), .Z(_04124_ ) );
BUF_X4 _11878_ ( .A(_04114_ ), .Z(_04125_ ) );
BUF_X4 _11879_ ( .A(_04125_ ), .Z(_04126_ ) );
OAI211_X1 _11880_ ( .A(_04106_ ), .B(_04120_ ), .C1(_04124_ ), .C2(_04126_ ), .ZN(_04127_ ) );
OR2_X1 _11881_ ( .A1(_04108_ ), .A2(\myreg.Reg[15][9] ), .ZN(_04128_ ) );
OAI211_X1 _11882_ ( .A(_04128_ ), .B(fanout_net_36 ), .C1(fanout_net_28 ), .C2(\myreg.Reg[14][9] ), .ZN(_04129_ ) );
OR2_X1 _11883_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[12][9] ), .ZN(_04130_ ) );
OAI211_X1 _11884_ ( .A(_04130_ ), .B(_04123_ ), .C1(_04118_ ), .C2(\myreg.Reg[13][9] ), .ZN(_04131_ ) );
NAND3_X1 _11885_ ( .A1(_04129_ ), .A2(fanout_net_39 ), .A3(_04131_ ), .ZN(_04132_ ) );
MUX2_X1 _11886_ ( .A(\myreg.Reg[8][9] ), .B(\myreg.Reg[9][9] ), .S(fanout_net_28 ), .Z(_04133_ ) );
MUX2_X1 _11887_ ( .A(\myreg.Reg[10][9] ), .B(\myreg.Reg[11][9] ), .S(fanout_net_28 ), .Z(_04134_ ) );
MUX2_X1 _11888_ ( .A(_04133_ ), .B(_04134_ ), .S(fanout_net_36 ), .Z(_04135_ ) );
OAI211_X1 _11889_ ( .A(fanout_net_40 ), .B(_04132_ ), .C1(_04135_ ), .C2(fanout_net_39 ), .ZN(_04136_ ) );
NAND2_X1 _11890_ ( .A1(_04127_ ), .A2(_04136_ ), .ZN(_04137_ ) );
BUF_X2 _11891_ ( .A(_04102_ ), .Z(_04138_ ) );
OAI21_X1 _11892_ ( .A(_04137_ ), .B1(_04100_ ), .B2(_04138_ ), .ZN(_04139_ ) );
AND2_X1 _11893_ ( .A1(_04104_ ), .A2(_04139_ ), .ZN(_04140_ ) );
AND2_X1 _11894_ ( .A1(_04140_ ), .A2(_02802_ ), .ZN(_04141_ ) );
NOR2_X1 _11895_ ( .A1(_04140_ ), .A2(_02802_ ), .ZN(_04142_ ) );
NOR2_X1 _11896_ ( .A1(_04141_ ), .A2(_04142_ ), .ZN(_04143_ ) );
INV_X1 _11897_ ( .A(_02780_ ), .ZN(_04144_ ) );
BUF_X2 _11898_ ( .A(_04100_ ), .Z(_04145_ ) );
INV_X1 _11899_ ( .A(\EX_LS_result_reg [8] ), .ZN(_04146_ ) );
OR3_X4 _11900_ ( .A1(_04145_ ), .A2(_04146_ ), .A3(_04138_ ), .ZN(_04147_ ) );
BUF_X4 _11901_ ( .A(_04106_ ), .Z(_04148_ ) );
OR2_X1 _11902_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[0][8] ), .ZN(_04149_ ) );
BUF_X4 _11903_ ( .A(_04112_ ), .Z(_04150_ ) );
BUF_X2 _11904_ ( .A(_04117_ ), .Z(_04151_ ) );
BUF_X4 _11905_ ( .A(_04151_ ), .Z(_04152_ ) );
BUF_X2 _11906_ ( .A(_04152_ ), .Z(_04153_ ) );
OAI211_X1 _11907_ ( .A(_04149_ ), .B(_04150_ ), .C1(_04153_ ), .C2(\myreg.Reg[1][8] ), .ZN(_04154_ ) );
OR2_X1 _11908_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[2][8] ), .ZN(_04155_ ) );
OAI211_X1 _11909_ ( .A(_04155_ ), .B(fanout_net_36 ), .C1(_04153_ ), .C2(\myreg.Reg[3][8] ), .ZN(_04156_ ) );
BUF_X4 _11910_ ( .A(_04115_ ), .Z(_04157_ ) );
NAND3_X1 _11911_ ( .A1(_04154_ ), .A2(_04156_ ), .A3(_04157_ ), .ZN(_04158_ ) );
MUX2_X1 _11912_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_28 ), .Z(_04159_ ) );
MUX2_X1 _11913_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_28 ), .Z(_04160_ ) );
MUX2_X1 _11914_ ( .A(_04159_ ), .B(_04160_ ), .S(_04150_ ), .Z(_04161_ ) );
OAI211_X1 _11915_ ( .A(_04148_ ), .B(_04158_ ), .C1(_04161_ ), .C2(_04157_ ), .ZN(_04162_ ) );
OR2_X1 _11916_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[14][8] ), .ZN(_04163_ ) );
OAI211_X1 _11917_ ( .A(_04163_ ), .B(fanout_net_36 ), .C1(_04153_ ), .C2(\myreg.Reg[15][8] ), .ZN(_04164_ ) );
OR2_X1 _11918_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[12][8] ), .ZN(_04165_ ) );
OAI211_X1 _11919_ ( .A(_04165_ ), .B(_04150_ ), .C1(_04153_ ), .C2(\myreg.Reg[13][8] ), .ZN(_04166_ ) );
NAND3_X1 _11920_ ( .A1(_04164_ ), .A2(_04166_ ), .A3(fanout_net_39 ), .ZN(_04167_ ) );
MUX2_X1 _11921_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_28 ), .Z(_04168_ ) );
MUX2_X1 _11922_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_28 ), .Z(_04169_ ) );
MUX2_X1 _11923_ ( .A(_04168_ ), .B(_04169_ ), .S(fanout_net_36 ), .Z(_04170_ ) );
OAI211_X1 _11924_ ( .A(fanout_net_40 ), .B(_04167_ ), .C1(_04170_ ), .C2(fanout_net_39 ), .ZN(_04171_ ) );
NAND2_X1 _11925_ ( .A1(_04162_ ), .A2(_04171_ ), .ZN(_04172_ ) );
BUF_X4 _11926_ ( .A(_04103_ ), .Z(_04173_ ) );
OAI21_X1 _11927_ ( .A(_04172_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04174_ ) );
AND2_X1 _11928_ ( .A1(_04147_ ), .A2(_04174_ ), .ZN(_04175_ ) );
XNOR2_X2 _11929_ ( .A(_04144_ ), .B(_04175_ ), .ZN(_04176_ ) );
AND2_X1 _11930_ ( .A1(_04143_ ), .A2(_04176_ ), .ZN(_04177_ ) );
NOR2_X1 _11931_ ( .A1(_04108_ ), .A2(\myreg.Reg[11][11] ), .ZN(_04178_ ) );
OAI21_X1 _11932_ ( .A(fanout_net_36 ), .B1(fanout_net_28 ), .B2(\myreg.Reg[10][11] ), .ZN(_04179_ ) );
NOR2_X1 _11933_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[8][11] ), .ZN(_04180_ ) );
OAI21_X1 _11934_ ( .A(_04111_ ), .B1(_04108_ ), .B2(\myreg.Reg[9][11] ), .ZN(_04181_ ) );
OAI221_X1 _11935_ ( .A(_04114_ ), .B1(_04178_ ), .B2(_04179_ ), .C1(_04180_ ), .C2(_04181_ ), .ZN(_04182_ ) );
MUX2_X1 _11936_ ( .A(\myreg.Reg[12][11] ), .B(\myreg.Reg[13][11] ), .S(fanout_net_28 ), .Z(_04183_ ) );
MUX2_X1 _11937_ ( .A(\myreg.Reg[14][11] ), .B(\myreg.Reg[15][11] ), .S(fanout_net_28 ), .Z(_04184_ ) );
MUX2_X1 _11938_ ( .A(_04183_ ), .B(_04184_ ), .S(fanout_net_36 ), .Z(_04185_ ) );
OAI211_X1 _11939_ ( .A(fanout_net_40 ), .B(_04182_ ), .C1(_04185_ ), .C2(_04125_ ), .ZN(_04186_ ) );
OR2_X1 _11940_ ( .A1(_04117_ ), .A2(\myreg.Reg[5][11] ), .ZN(_04187_ ) );
OAI211_X1 _11941_ ( .A(_04187_ ), .B(_04111_ ), .C1(fanout_net_28 ), .C2(\myreg.Reg[4][11] ), .ZN(_04188_ ) );
OR2_X1 _11942_ ( .A1(_04117_ ), .A2(\myreg.Reg[7][11] ), .ZN(_04189_ ) );
OAI211_X1 _11943_ ( .A(_04189_ ), .B(fanout_net_36 ), .C1(fanout_net_28 ), .C2(\myreg.Reg[6][11] ), .ZN(_04190_ ) );
NAND3_X1 _11944_ ( .A1(_04188_ ), .A2(_04190_ ), .A3(fanout_net_39 ), .ZN(_04191_ ) );
MUX2_X1 _11945_ ( .A(\myreg.Reg[2][11] ), .B(\myreg.Reg[3][11] ), .S(fanout_net_28 ), .Z(_04192_ ) );
MUX2_X1 _11946_ ( .A(\myreg.Reg[0][11] ), .B(\myreg.Reg[1][11] ), .S(fanout_net_28 ), .Z(_04193_ ) );
MUX2_X1 _11947_ ( .A(_04192_ ), .B(_04193_ ), .S(_04111_ ), .Z(_04194_ ) );
OAI211_X1 _11948_ ( .A(_04105_ ), .B(_04191_ ), .C1(_04194_ ), .C2(fanout_net_39 ), .ZN(_04195_ ) );
NAND2_X1 _11949_ ( .A1(_04186_ ), .A2(_04195_ ), .ZN(_04196_ ) );
OAI21_X1 _11950_ ( .A(_04196_ ), .B1(_04099_ ), .B2(_04102_ ), .ZN(_04197_ ) );
BUF_X4 _11951_ ( .A(_02130_ ), .Z(_04198_ ) );
OAI21_X1 _11952_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02136_ ), .B2(\ID_EX_rs2 [1] ), .ZN(_04199_ ) );
AOI211_X4 _11953_ ( .A(_04199_ ), .B(_02134_ ), .C1(_02136_ ), .C2(\ID_EX_rs2 [1] ), .ZN(_04200_ ) );
AND4_X2 _11954_ ( .A1(_04094_ ), .A2(_04093_ ), .A3(_04096_ ), .A4(_04097_ ), .ZN(_04201_ ) );
NAND4_X1 _11955_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [11] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04202_ ) );
AND2_X1 _11956_ ( .A1(_04197_ ), .A2(_04202_ ), .ZN(_04203_ ) );
XOR2_X1 _11957_ ( .A(_02851_ ), .B(_04203_ ), .Z(_04204_ ) );
INV_X1 _11958_ ( .A(_02828_ ), .ZN(_04205_ ) );
OR2_X1 _11959_ ( .A1(_04117_ ), .A2(\myreg.Reg[9][10] ), .ZN(_04206_ ) );
BUF_X4 _11960_ ( .A(_04110_ ), .Z(_04207_ ) );
OAI211_X1 _11961_ ( .A(_04206_ ), .B(_04207_ ), .C1(fanout_net_28 ), .C2(\myreg.Reg[8][10] ), .ZN(_04208_ ) );
OR2_X1 _11962_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[10][10] ), .ZN(_04209_ ) );
OAI211_X1 _11963_ ( .A(_04209_ ), .B(fanout_net_36 ), .C1(_04151_ ), .C2(\myreg.Reg[11][10] ), .ZN(_04210_ ) );
NAND3_X1 _11964_ ( .A1(_04208_ ), .A2(_04114_ ), .A3(_04210_ ), .ZN(_04211_ ) );
MUX2_X1 _11965_ ( .A(\myreg.Reg[14][10] ), .B(\myreg.Reg[15][10] ), .S(fanout_net_28 ), .Z(_04212_ ) );
MUX2_X1 _11966_ ( .A(\myreg.Reg[12][10] ), .B(\myreg.Reg[13][10] ), .S(fanout_net_28 ), .Z(_04213_ ) );
MUX2_X1 _11967_ ( .A(_04212_ ), .B(_04213_ ), .S(_04111_ ), .Z(_04214_ ) );
OAI211_X1 _11968_ ( .A(fanout_net_40 ), .B(_04211_ ), .C1(_04214_ ), .C2(_04125_ ), .ZN(_04215_ ) );
MUX2_X1 _11969_ ( .A(\myreg.Reg[2][10] ), .B(\myreg.Reg[3][10] ), .S(fanout_net_28 ), .Z(_04216_ ) );
AND2_X1 _11970_ ( .A1(_04216_ ), .A2(fanout_net_36 ), .ZN(_04217_ ) );
BUF_X4 _11971_ ( .A(_04207_ ), .Z(_04218_ ) );
MUX2_X1 _11972_ ( .A(\myreg.Reg[0][10] ), .B(\myreg.Reg[1][10] ), .S(fanout_net_29 ), .Z(_04219_ ) );
AOI211_X1 _11973_ ( .A(fanout_net_39 ), .B(_04217_ ), .C1(_04218_ ), .C2(_04219_ ), .ZN(_04220_ ) );
MUX2_X1 _11974_ ( .A(\myreg.Reg[6][10] ), .B(\myreg.Reg[7][10] ), .S(fanout_net_29 ), .Z(_04221_ ) );
MUX2_X1 _11975_ ( .A(\myreg.Reg[4][10] ), .B(\myreg.Reg[5][10] ), .S(fanout_net_29 ), .Z(_04222_ ) );
MUX2_X1 _11976_ ( .A(_04221_ ), .B(_04222_ ), .S(_04111_ ), .Z(_04223_ ) );
OAI21_X1 _11977_ ( .A(_04105_ ), .B1(_04223_ ), .B2(_04125_ ), .ZN(_04224_ ) );
OAI21_X1 _11978_ ( .A(_04215_ ), .B1(_04220_ ), .B2(_04224_ ), .ZN(_04225_ ) );
OAI21_X1 _11979_ ( .A(_04225_ ), .B1(_04103_ ), .B2(_04100_ ), .ZN(_04226_ ) );
NAND4_X1 _11980_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [10] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04227_ ) );
AND2_X1 _11981_ ( .A1(_04226_ ), .A2(_04227_ ), .ZN(_04228_ ) );
XNOR2_X1 _11982_ ( .A(_04205_ ), .B(_04228_ ), .ZN(_04229_ ) );
AND3_X1 _11983_ ( .A1(_04177_ ), .A2(_04204_ ), .A3(_04229_ ), .ZN(_04230_ ) );
INV_X1 _11984_ ( .A(_02683_ ), .ZN(_04231_ ) );
INV_X1 _11985_ ( .A(\EX_LS_result_reg [15] ), .ZN(_04232_ ) );
OR3_X1 _11986_ ( .A1(_04100_ ), .A2(_04232_ ), .A3(_04103_ ), .ZN(_04233_ ) );
OR2_X1 _11987_ ( .A1(_04108_ ), .A2(\myreg.Reg[3][15] ), .ZN(_04234_ ) );
OAI211_X1 _11988_ ( .A(_04234_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[2][15] ), .ZN(_04235_ ) );
OR2_X1 _11989_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][15] ), .ZN(_04236_ ) );
OAI211_X1 _11990_ ( .A(_04236_ ), .B(_04112_ ), .C1(_04152_ ), .C2(\myreg.Reg[1][15] ), .ZN(_04237_ ) );
NAND3_X1 _11991_ ( .A1(_04235_ ), .A2(_04115_ ), .A3(_04237_ ), .ZN(_04238_ ) );
MUX2_X1 _11992_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_29 ), .Z(_04239_ ) );
MUX2_X1 _11993_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_29 ), .Z(_04240_ ) );
MUX2_X1 _11994_ ( .A(_04239_ ), .B(_04240_ ), .S(_04123_ ), .Z(_04241_ ) );
OAI211_X1 _11995_ ( .A(_04106_ ), .B(_04238_ ), .C1(_04241_ ), .C2(_04126_ ), .ZN(_04242_ ) );
OR2_X1 _11996_ ( .A1(_04108_ ), .A2(\myreg.Reg[15][15] ), .ZN(_04243_ ) );
OAI211_X1 _11997_ ( .A(_04243_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[14][15] ), .ZN(_04244_ ) );
OR2_X1 _11998_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[12][15] ), .ZN(_04245_ ) );
OAI211_X1 _11999_ ( .A(_04245_ ), .B(_04123_ ), .C1(_04118_ ), .C2(\myreg.Reg[13][15] ), .ZN(_04246_ ) );
NAND3_X1 _12000_ ( .A1(_04244_ ), .A2(fanout_net_39 ), .A3(_04246_ ), .ZN(_04247_ ) );
MUX2_X1 _12001_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_29 ), .Z(_04248_ ) );
MUX2_X1 _12002_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_29 ), .Z(_04249_ ) );
MUX2_X1 _12003_ ( .A(_04248_ ), .B(_04249_ ), .S(fanout_net_36 ), .Z(_04250_ ) );
OAI211_X1 _12004_ ( .A(fanout_net_40 ), .B(_04247_ ), .C1(_04250_ ), .C2(fanout_net_39 ), .ZN(_04251_ ) );
NAND2_X1 _12005_ ( .A1(_04242_ ), .A2(_04251_ ), .ZN(_04252_ ) );
BUF_X2 _12006_ ( .A(_04099_ ), .Z(_04253_ ) );
OAI21_X1 _12007_ ( .A(_04252_ ), .B1(_04253_ ), .B2(_04138_ ), .ZN(_04254_ ) );
AND2_X1 _12008_ ( .A1(_04233_ ), .A2(_04254_ ), .ZN(_04255_ ) );
XNOR2_X1 _12009_ ( .A(_04231_ ), .B(_04255_ ), .ZN(_04256_ ) );
NOR2_X1 _12010_ ( .A1(_04152_ ), .A2(\myreg.Reg[11][14] ), .ZN(_04257_ ) );
OAI21_X1 _12011_ ( .A(fanout_net_36 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[10][14] ), .ZN(_04258_ ) );
NOR2_X1 _12012_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][14] ), .ZN(_04259_ ) );
OAI21_X1 _12013_ ( .A(_04112_ ), .B1(_04152_ ), .B2(\myreg.Reg[9][14] ), .ZN(_04260_ ) );
OAI221_X1 _12014_ ( .A(_04115_ ), .B1(_04257_ ), .B2(_04258_ ), .C1(_04259_ ), .C2(_04260_ ), .ZN(_04261_ ) );
MUX2_X1 _12015_ ( .A(\myreg.Reg[12][14] ), .B(\myreg.Reg[13][14] ), .S(fanout_net_29 ), .Z(_04262_ ) );
MUX2_X1 _12016_ ( .A(\myreg.Reg[14][14] ), .B(\myreg.Reg[15][14] ), .S(fanout_net_29 ), .Z(_04263_ ) );
MUX2_X1 _12017_ ( .A(_04262_ ), .B(_04263_ ), .S(fanout_net_36 ), .Z(_04264_ ) );
BUF_X4 _12018_ ( .A(_04125_ ), .Z(_04265_ ) );
OAI211_X1 _12019_ ( .A(fanout_net_40 ), .B(_04261_ ), .C1(_04264_ ), .C2(_04265_ ), .ZN(_04266_ ) );
OR2_X1 _12020_ ( .A1(_04151_ ), .A2(\myreg.Reg[5][14] ), .ZN(_04267_ ) );
BUF_X4 _12021_ ( .A(_04207_ ), .Z(_04268_ ) );
OAI211_X1 _12022_ ( .A(_04267_ ), .B(_04268_ ), .C1(fanout_net_29 ), .C2(\myreg.Reg[4][14] ), .ZN(_04269_ ) );
OR2_X1 _12023_ ( .A1(_04151_ ), .A2(\myreg.Reg[7][14] ), .ZN(_04270_ ) );
OAI211_X1 _12024_ ( .A(_04270_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[6][14] ), .ZN(_04271_ ) );
NAND3_X1 _12025_ ( .A1(_04269_ ), .A2(_04271_ ), .A3(fanout_net_39 ), .ZN(_04272_ ) );
MUX2_X1 _12026_ ( .A(\myreg.Reg[2][14] ), .B(\myreg.Reg[3][14] ), .S(fanout_net_29 ), .Z(_04273_ ) );
MUX2_X1 _12027_ ( .A(\myreg.Reg[0][14] ), .B(\myreg.Reg[1][14] ), .S(fanout_net_29 ), .Z(_04274_ ) );
MUX2_X1 _12028_ ( .A(_04273_ ), .B(_04274_ ), .S(_04112_ ), .Z(_04275_ ) );
OAI211_X1 _12029_ ( .A(_04106_ ), .B(_04272_ ), .C1(_04275_ ), .C2(fanout_net_39 ), .ZN(_04276_ ) );
NAND2_X1 _12030_ ( .A1(_04266_ ), .A2(_04276_ ), .ZN(_04277_ ) );
OAI21_X1 _12031_ ( .A(_04277_ ), .B1(_04253_ ), .B2(_04138_ ), .ZN(_04278_ ) );
NAND4_X1 _12032_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [14] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04279_ ) );
AND2_X1 _12033_ ( .A1(_04278_ ), .A2(_04279_ ), .ZN(_04280_ ) );
XOR2_X2 _12034_ ( .A(_02707_ ), .B(_04280_ ), .Z(_04281_ ) );
AND2_X1 _12035_ ( .A1(_04256_ ), .A2(_04281_ ), .ZN(_04282_ ) );
NAND2_X1 _12036_ ( .A1(_02734_ ), .A2(_02754_ ), .ZN(_04283_ ) );
INV_X1 _12037_ ( .A(_04283_ ), .ZN(_04284_ ) );
INV_X1 _12038_ ( .A(\EX_LS_result_reg [13] ), .ZN(_04285_ ) );
OR3_X1 _12039_ ( .A1(_04099_ ), .A2(_04285_ ), .A3(_04102_ ), .ZN(_04286_ ) );
OR2_X1 _12040_ ( .A1(_04107_ ), .A2(\myreg.Reg[3][13] ), .ZN(_04287_ ) );
OAI211_X1 _12041_ ( .A(_04287_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[2][13] ), .ZN(_04288_ ) );
OR2_X1 _12042_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][13] ), .ZN(_04289_ ) );
OAI211_X1 _12043_ ( .A(_04289_ ), .B(_04111_ ), .C1(_04117_ ), .C2(\myreg.Reg[1][13] ), .ZN(_04290_ ) );
NAND3_X1 _12044_ ( .A1(_04288_ ), .A2(_04114_ ), .A3(_04290_ ), .ZN(_04291_ ) );
MUX2_X1 _12045_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_29 ), .Z(_04292_ ) );
MUX2_X1 _12046_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_29 ), .Z(_04293_ ) );
MUX2_X1 _12047_ ( .A(_04292_ ), .B(_04293_ ), .S(_04111_ ), .Z(_04294_ ) );
OAI211_X1 _12048_ ( .A(_04105_ ), .B(_04291_ ), .C1(_04294_ ), .C2(_04125_ ), .ZN(_04295_ ) );
OR2_X1 _12049_ ( .A1(_04107_ ), .A2(\myreg.Reg[15][13] ), .ZN(_04296_ ) );
OAI211_X1 _12050_ ( .A(_04296_ ), .B(fanout_net_36 ), .C1(fanout_net_29 ), .C2(\myreg.Reg[14][13] ), .ZN(_04297_ ) );
OR2_X1 _12051_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[12][13] ), .ZN(_04298_ ) );
OAI211_X1 _12052_ ( .A(_04298_ ), .B(_04111_ ), .C1(_04117_ ), .C2(\myreg.Reg[13][13] ), .ZN(_04299_ ) );
NAND3_X1 _12053_ ( .A1(_04297_ ), .A2(fanout_net_39 ), .A3(_04299_ ), .ZN(_04300_ ) );
MUX2_X1 _12054_ ( .A(\myreg.Reg[8][13] ), .B(\myreg.Reg[9][13] ), .S(fanout_net_29 ), .Z(_04301_ ) );
MUX2_X1 _12055_ ( .A(\myreg.Reg[10][13] ), .B(\myreg.Reg[11][13] ), .S(fanout_net_29 ), .Z(_04302_ ) );
MUX2_X1 _12056_ ( .A(_04301_ ), .B(_04302_ ), .S(fanout_net_36 ), .Z(_04303_ ) );
OAI211_X1 _12057_ ( .A(fanout_net_40 ), .B(_04300_ ), .C1(_04303_ ), .C2(fanout_net_39 ), .ZN(_04304_ ) );
NAND2_X1 _12058_ ( .A1(_04295_ ), .A2(_04304_ ), .ZN(_04305_ ) );
OAI21_X1 _12059_ ( .A(_04305_ ), .B1(_04099_ ), .B2(_04102_ ), .ZN(_04306_ ) );
AND2_X1 _12060_ ( .A1(_04286_ ), .A2(_04306_ ), .ZN(_04307_ ) );
XNOR2_X1 _12061_ ( .A(_04284_ ), .B(_04307_ ), .ZN(_04308_ ) );
BUF_X2 _12062_ ( .A(_04117_ ), .Z(_04309_ ) );
BUF_X4 _12063_ ( .A(_04309_ ), .Z(_04310_ ) );
NOR2_X1 _12064_ ( .A1(_04310_ ), .A2(\myreg.Reg[11][12] ), .ZN(_04311_ ) );
OAI21_X1 _12065_ ( .A(fanout_net_36 ), .B1(fanout_net_29 ), .B2(\myreg.Reg[10][12] ), .ZN(_04312_ ) );
NOR2_X1 _12066_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[8][12] ), .ZN(_04313_ ) );
BUF_X4 _12067_ ( .A(_04207_ ), .Z(_04314_ ) );
OAI21_X1 _12068_ ( .A(_04314_ ), .B1(_04310_ ), .B2(\myreg.Reg[9][12] ), .ZN(_04315_ ) );
OAI221_X1 _12069_ ( .A(_04126_ ), .B1(_04311_ ), .B2(_04312_ ), .C1(_04313_ ), .C2(_04315_ ), .ZN(_04316_ ) );
MUX2_X1 _12070_ ( .A(\myreg.Reg[12][12] ), .B(\myreg.Reg[13][12] ), .S(fanout_net_29 ), .Z(_04317_ ) );
MUX2_X1 _12071_ ( .A(\myreg.Reg[14][12] ), .B(\myreg.Reg[15][12] ), .S(fanout_net_30 ), .Z(_04318_ ) );
MUX2_X1 _12072_ ( .A(_04317_ ), .B(_04318_ ), .S(fanout_net_36 ), .Z(_04319_ ) );
OAI211_X1 _12073_ ( .A(fanout_net_40 ), .B(_04316_ ), .C1(_04319_ ), .C2(_04157_ ), .ZN(_04320_ ) );
OR2_X1 _12074_ ( .A1(_04118_ ), .A2(\myreg.Reg[5][12] ), .ZN(_04321_ ) );
OAI211_X1 _12075_ ( .A(_04321_ ), .B(_04314_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[4][12] ), .ZN(_04322_ ) );
OR2_X1 _12076_ ( .A1(_04118_ ), .A2(\myreg.Reg[7][12] ), .ZN(_04323_ ) );
OAI211_X1 _12077_ ( .A(_04323_ ), .B(fanout_net_36 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[6][12] ), .ZN(_04324_ ) );
NAND3_X1 _12078_ ( .A1(_04322_ ), .A2(_04324_ ), .A3(fanout_net_39 ), .ZN(_04325_ ) );
MUX2_X1 _12079_ ( .A(\myreg.Reg[2][12] ), .B(\myreg.Reg[3][12] ), .S(fanout_net_30 ), .Z(_04326_ ) );
MUX2_X1 _12080_ ( .A(\myreg.Reg[0][12] ), .B(\myreg.Reg[1][12] ), .S(fanout_net_30 ), .Z(_04327_ ) );
MUX2_X1 _12081_ ( .A(_04326_ ), .B(_04327_ ), .S(_04218_ ), .Z(_04328_ ) );
OAI211_X1 _12082_ ( .A(_04148_ ), .B(_04325_ ), .C1(_04328_ ), .C2(fanout_net_39 ), .ZN(_04329_ ) );
NAND2_X1 _12083_ ( .A1(_04320_ ), .A2(_04329_ ), .ZN(_04330_ ) );
OAI21_X1 _12084_ ( .A(_04330_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04331_ ) );
NAND4_X1 _12085_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [12] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04332_ ) );
AND2_X1 _12086_ ( .A1(_04331_ ), .A2(_04332_ ), .ZN(_04333_ ) );
XOR2_X1 _12087_ ( .A(_02731_ ), .B(_04333_ ), .Z(_04334_ ) );
AND2_X1 _12088_ ( .A1(_04308_ ), .A2(_04334_ ), .ZN(_04335_ ) );
AND2_X1 _12089_ ( .A1(_04282_ ), .A2(_04335_ ), .ZN(_04336_ ) );
AND2_X1 _12090_ ( .A1(_04230_ ), .A2(_04336_ ), .ZN(_04337_ ) );
INV_X1 _12091_ ( .A(_04337_ ), .ZN(_04338_ ) );
INV_X1 _12092_ ( .A(_02478_ ), .ZN(_04339_ ) );
INV_X1 _12093_ ( .A(\EX_LS_result_reg [1] ), .ZN(_04340_ ) );
OR3_X1 _12094_ ( .A1(_04100_ ), .A2(_04340_ ), .A3(_04103_ ), .ZN(_04341_ ) );
OR2_X1 _12095_ ( .A1(_04151_ ), .A2(\myreg.Reg[1][1] ), .ZN(_04342_ ) );
OAI211_X1 _12096_ ( .A(_04342_ ), .B(_04268_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[0][1] ), .ZN(_04343_ ) );
OR2_X1 _12097_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[2][1] ), .ZN(_04344_ ) );
OAI211_X1 _12098_ ( .A(_04344_ ), .B(fanout_net_36 ), .C1(_04152_ ), .C2(\myreg.Reg[3][1] ), .ZN(_04345_ ) );
NAND3_X1 _12099_ ( .A1(_04343_ ), .A2(_04115_ ), .A3(_04345_ ), .ZN(_04346_ ) );
MUX2_X1 _12100_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(fanout_net_30 ), .Z(_04347_ ) );
MUX2_X1 _12101_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(fanout_net_30 ), .Z(_04348_ ) );
MUX2_X1 _12102_ ( .A(_04347_ ), .B(_04348_ ), .S(_04112_ ), .Z(_04349_ ) );
OAI211_X1 _12103_ ( .A(_04106_ ), .B(_04346_ ), .C1(_04349_ ), .C2(_04126_ ), .ZN(_04350_ ) );
OR2_X1 _12104_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[14][1] ), .ZN(_04351_ ) );
BUF_X2 _12105_ ( .A(_04151_ ), .Z(_04352_ ) );
OAI211_X1 _12106_ ( .A(_04351_ ), .B(fanout_net_36 ), .C1(_04352_ ), .C2(\myreg.Reg[15][1] ), .ZN(_04353_ ) );
OR2_X1 _12107_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[12][1] ), .ZN(_04354_ ) );
OAI211_X1 _12108_ ( .A(_04354_ ), .B(_04112_ ), .C1(_04152_ ), .C2(\myreg.Reg[13][1] ), .ZN(_04355_ ) );
NAND3_X1 _12109_ ( .A1(_04353_ ), .A2(_04355_ ), .A3(fanout_net_39 ), .ZN(_04356_ ) );
MUX2_X1 _12110_ ( .A(\myreg.Reg[8][1] ), .B(\myreg.Reg[9][1] ), .S(fanout_net_30 ), .Z(_04357_ ) );
MUX2_X1 _12111_ ( .A(\myreg.Reg[10][1] ), .B(\myreg.Reg[11][1] ), .S(fanout_net_30 ), .Z(_04358_ ) );
MUX2_X1 _12112_ ( .A(_04357_ ), .B(_04358_ ), .S(fanout_net_36 ), .Z(_04359_ ) );
OAI211_X1 _12113_ ( .A(fanout_net_40 ), .B(_04356_ ), .C1(_04359_ ), .C2(fanout_net_39 ), .ZN(_04360_ ) );
NAND2_X1 _12114_ ( .A1(_04350_ ), .A2(_04360_ ), .ZN(_04361_ ) );
OAI21_X1 _12115_ ( .A(_04361_ ), .B1(_04253_ ), .B2(_04138_ ), .ZN(_04362_ ) );
AND2_X1 _12116_ ( .A1(_04341_ ), .A2(_04362_ ), .ZN(_04363_ ) );
XNOR2_X1 _12117_ ( .A(_04339_ ), .B(_04363_ ), .ZN(_04364_ ) );
NOR2_X1 _12118_ ( .A1(_04151_ ), .A2(\myreg.Reg[3][0] ), .ZN(_04365_ ) );
OAI21_X1 _12119_ ( .A(fanout_net_36 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[2][0] ), .ZN(_04366_ ) );
NOR2_X1 _12120_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[0][0] ), .ZN(_04367_ ) );
OAI21_X1 _12121_ ( .A(_04207_ ), .B1(_04151_ ), .B2(\myreg.Reg[1][0] ), .ZN(_04368_ ) );
OAI221_X1 _12122_ ( .A(_04114_ ), .B1(_04365_ ), .B2(_04366_ ), .C1(_04367_ ), .C2(_04368_ ), .ZN(_04369_ ) );
MUX2_X1 _12123_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_30 ), .Z(_04370_ ) );
MUX2_X1 _12124_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_30 ), .Z(_04371_ ) );
MUX2_X1 _12125_ ( .A(_04370_ ), .B(_04371_ ), .S(_04207_ ), .Z(_04372_ ) );
OAI211_X1 _12126_ ( .A(_04105_ ), .B(_04369_ ), .C1(_04372_ ), .C2(_04125_ ), .ZN(_04373_ ) );
OR2_X1 _12127_ ( .A1(_04117_ ), .A2(\myreg.Reg[9][0] ), .ZN(_04374_ ) );
OAI211_X1 _12128_ ( .A(_04374_ ), .B(_04207_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[8][0] ), .ZN(_04375_ ) );
OR2_X1 _12129_ ( .A1(_04117_ ), .A2(\myreg.Reg[11][0] ), .ZN(_04376_ ) );
OAI211_X1 _12130_ ( .A(_04376_ ), .B(fanout_net_36 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[10][0] ), .ZN(_04377_ ) );
NAND3_X1 _12131_ ( .A1(_04375_ ), .A2(_04377_ ), .A3(_04114_ ), .ZN(_04378_ ) );
MUX2_X1 _12132_ ( .A(\myreg.Reg[14][0] ), .B(\myreg.Reg[15][0] ), .S(fanout_net_30 ), .Z(_04379_ ) );
MUX2_X1 _12133_ ( .A(\myreg.Reg[12][0] ), .B(\myreg.Reg[13][0] ), .S(fanout_net_30 ), .Z(_04380_ ) );
MUX2_X1 _12134_ ( .A(_04379_ ), .B(_04380_ ), .S(_04207_ ), .Z(_04381_ ) );
OAI211_X1 _12135_ ( .A(fanout_net_40 ), .B(_04378_ ), .C1(_04381_ ), .C2(_04125_ ), .ZN(_04382_ ) );
NAND2_X1 _12136_ ( .A1(_04373_ ), .A2(_04382_ ), .ZN(_04383_ ) );
OAI21_X1 _12137_ ( .A(_04383_ ), .B1(_04100_ ), .B2(_04103_ ), .ZN(_04384_ ) );
NAND4_X1 _12138_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [0] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04385_ ) );
AND2_X1 _12139_ ( .A1(_04384_ ), .A2(_04385_ ), .ZN(_04386_ ) );
NOR2_X1 _12140_ ( .A1(_02502_ ), .A2(_04386_ ), .ZN(_04387_ ) );
INV_X1 _12141_ ( .A(_04387_ ), .ZN(_04388_ ) );
NAND2_X1 _12142_ ( .A1(_04364_ ), .A2(_04388_ ), .ZN(_04389_ ) );
INV_X1 _12143_ ( .A(_02549_ ), .ZN(_04390_ ) );
AOI22_X1 _12144_ ( .A1(_02145_ ), .A2(\ID_EX_rs2 [3] ), .B1(_03344_ ), .B2(\EX_LS_dest_reg [1] ), .ZN(_04391_ ) );
NAND3_X1 _12145_ ( .A1(_04093_ ), .A2(_04097_ ), .A3(_04391_ ), .ZN(_04392_ ) );
AOI211_X2 _12146_ ( .A(_04102_ ), .B(_04392_ ), .C1(\EX_LS_dest_reg [3] ), .C2(_03339_ ), .ZN(_04393_ ) );
NAND2_X2 _12147_ ( .A1(_04393_ ), .A2(_04198_ ), .ZN(_04394_ ) );
OAI221_X1 _12148_ ( .A(_04096_ ), .B1(\EX_LS_dest_reg [1] ), .B2(_03344_ ), .C1(_02132_ ), .C2(_02133_ ), .ZN(_04395_ ) );
OR3_X1 _12149_ ( .A1(_04394_ ), .A2(\EX_LS_result_reg [2] ), .A3(_04395_ ), .ZN(_04396_ ) );
OR2_X1 _12150_ ( .A1(_04118_ ), .A2(\myreg.Reg[7][2] ), .ZN(_04397_ ) );
OAI211_X1 _12151_ ( .A(_04397_ ), .B(fanout_net_36 ), .C1(fanout_net_30 ), .C2(\myreg.Reg[6][2] ), .ZN(_04398_ ) );
OR2_X1 _12152_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[4][2] ), .ZN(_04399_ ) );
BUF_X2 _12153_ ( .A(_04309_ ), .Z(_04400_ ) );
OAI211_X1 _12154_ ( .A(_04399_ ), .B(_04314_ ), .C1(_04400_ ), .C2(\myreg.Reg[5][2] ), .ZN(_04401_ ) );
NAND3_X1 _12155_ ( .A1(_04398_ ), .A2(fanout_net_39 ), .A3(_04401_ ), .ZN(_04402_ ) );
MUX2_X1 _12156_ ( .A(\myreg.Reg[2][2] ), .B(\myreg.Reg[3][2] ), .S(fanout_net_30 ), .Z(_04403_ ) );
MUX2_X1 _12157_ ( .A(\myreg.Reg[0][2] ), .B(\myreg.Reg[1][2] ), .S(fanout_net_30 ), .Z(_04404_ ) );
MUX2_X1 _12158_ ( .A(_04403_ ), .B(_04404_ ), .S(_04218_ ), .Z(_04405_ ) );
OAI211_X1 _12159_ ( .A(_04148_ ), .B(_04402_ ), .C1(_04405_ ), .C2(fanout_net_39 ), .ZN(_04406_ ) );
NOR2_X1 _12160_ ( .A1(_04310_ ), .A2(\myreg.Reg[11][2] ), .ZN(_04407_ ) );
OAI21_X1 _12161_ ( .A(fanout_net_37 ), .B1(fanout_net_30 ), .B2(\myreg.Reg[10][2] ), .ZN(_04408_ ) );
NOR2_X1 _12162_ ( .A1(fanout_net_30 ), .A2(\myreg.Reg[8][2] ), .ZN(_04409_ ) );
OAI21_X1 _12163_ ( .A(_04218_ ), .B1(_04310_ ), .B2(\myreg.Reg[9][2] ), .ZN(_04410_ ) );
OAI221_X1 _12164_ ( .A(_04126_ ), .B1(_04407_ ), .B2(_04408_ ), .C1(_04409_ ), .C2(_04410_ ), .ZN(_04411_ ) );
MUX2_X1 _12165_ ( .A(\myreg.Reg[12][2] ), .B(\myreg.Reg[13][2] ), .S(fanout_net_30 ), .Z(_04412_ ) );
MUX2_X1 _12166_ ( .A(\myreg.Reg[14][2] ), .B(\myreg.Reg[15][2] ), .S(fanout_net_30 ), .Z(_04413_ ) );
MUX2_X1 _12167_ ( .A(_04412_ ), .B(_04413_ ), .S(fanout_net_37 ), .Z(_04414_ ) );
OAI211_X1 _12168_ ( .A(fanout_net_40 ), .B(_04411_ ), .C1(_04414_ ), .C2(_04157_ ), .ZN(_04415_ ) );
CLKBUF_X2 _12169_ ( .A(_04394_ ), .Z(_04416_ ) );
CLKBUF_X2 _12170_ ( .A(_04395_ ), .Z(_04417_ ) );
OAI211_X1 _12171_ ( .A(_04406_ ), .B(_04415_ ), .C1(_04416_ ), .C2(_04417_ ), .ZN(_04418_ ) );
NAND2_X1 _12172_ ( .A1(_04396_ ), .A2(_04418_ ), .ZN(_04419_ ) );
XNOR2_X1 _12173_ ( .A(_04390_ ), .B(_04419_ ), .ZN(_04420_ ) );
INV_X1 _12174_ ( .A(_04420_ ), .ZN(_04421_ ) );
OR3_X1 _12175_ ( .A1(_04416_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04417_ ), .ZN(_04422_ ) );
BUF_X4 _12176_ ( .A(_04148_ ), .Z(_04423_ ) );
OR2_X1 _12177_ ( .A1(_04352_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04424_ ) );
OAI211_X1 _12178_ ( .A(_04424_ ), .B(_04150_ ), .C1(fanout_net_30 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04425_ ) );
OR2_X1 _12179_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04426_ ) );
OAI211_X1 _12180_ ( .A(_04426_ ), .B(fanout_net_37 ), .C1(_04153_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04427_ ) );
NAND3_X1 _12181_ ( .A1(_04425_ ), .A2(fanout_net_39 ), .A3(_04427_ ), .ZN(_04428_ ) );
MUX2_X1 _12182_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04429_ ) );
MUX2_X1 _12183_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04430_ ) );
MUX2_X1 _12184_ ( .A(_04429_ ), .B(_04430_ ), .S(_04150_ ), .Z(_04431_ ) );
OAI211_X1 _12185_ ( .A(_04423_ ), .B(_04428_ ), .C1(_04431_ ), .C2(fanout_net_39 ), .ZN(_04432_ ) );
NOR2_X1 _12186_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04433_ ) );
OAI21_X1 _12187_ ( .A(_04314_ ), .B1(_04400_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04434_ ) );
MUX2_X1 _12188_ ( .A(_02518_ ), .B(_02519_ ), .S(fanout_net_31 ), .Z(_04435_ ) );
BUF_X4 _12189_ ( .A(_04314_ ), .Z(_04436_ ) );
OAI221_X1 _12190_ ( .A(_04265_ ), .B1(_04433_ ), .B2(_04434_ ), .C1(_04435_ ), .C2(_04436_ ), .ZN(_04437_ ) );
MUX2_X1 _12191_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04438_ ) );
MUX2_X1 _12192_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04439_ ) );
MUX2_X1 _12193_ ( .A(_04438_ ), .B(_04439_ ), .S(fanout_net_37 ), .Z(_04440_ ) );
OAI211_X1 _12194_ ( .A(fanout_net_40 ), .B(_04437_ ), .C1(_04440_ ), .C2(_04157_ ), .ZN(_04441_ ) );
OAI211_X1 _12195_ ( .A(_04432_ ), .B(_04441_ ), .C1(_04416_ ), .C2(_04417_ ), .ZN(_04442_ ) );
NAND2_X1 _12196_ ( .A1(_04422_ ), .A2(_04442_ ), .ZN(_04443_ ) );
XNOR2_X1 _12197_ ( .A(_04443_ ), .B(_02527_ ), .ZN(_04444_ ) );
INV_X1 _12198_ ( .A(_04444_ ), .ZN(_04445_ ) );
NOR4_X1 _12199_ ( .A1(_04338_ ), .A2(_04389_ ), .A3(_04421_ ), .A4(_04445_ ), .ZN(_04446_ ) );
NOR2_X1 _12200_ ( .A1(_04099_ ), .A2(_04102_ ), .ZN(_04447_ ) );
NAND2_X1 _12201_ ( .A1(_04447_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_04448_ ) );
BUF_X2 _12202_ ( .A(_04310_ ), .Z(_04449_ ) );
OR2_X1 _12203_ ( .A1(_04449_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04450_ ) );
BUF_X4 _12204_ ( .A(_04436_ ), .Z(_04451_ ) );
OAI211_X1 _12205_ ( .A(_04450_ ), .B(_04451_ ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04452_ ) );
BUF_X4 _12206_ ( .A(_04157_ ), .Z(_04453_ ) );
NAND2_X1 _12207_ ( .A1(_02168_ ), .A2(fanout_net_31 ), .ZN(_04454_ ) );
OAI211_X1 _12208_ ( .A(_04454_ ), .B(fanout_net_37 ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04455_ ) );
NAND3_X1 _12209_ ( .A1(_04452_ ), .A2(_04453_ ), .A3(_04455_ ), .ZN(_04456_ ) );
MUX2_X1 _12210_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04457_ ) );
MUX2_X1 _12211_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04458_ ) );
BUF_X4 _12212_ ( .A(_04150_ ), .Z(_04459_ ) );
MUX2_X1 _12213_ ( .A(_04457_ ), .B(_04458_ ), .S(_04459_ ), .Z(_04460_ ) );
BUF_X4 _12214_ ( .A(_04453_ ), .Z(_04461_ ) );
OAI211_X1 _12215_ ( .A(_04423_ ), .B(_04456_ ), .C1(_04460_ ), .C2(_04461_ ), .ZN(_04462_ ) );
OR2_X1 _12216_ ( .A1(fanout_net_31 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04463_ ) );
BUF_X2 _12217_ ( .A(_04153_ ), .Z(_04464_ ) );
OAI211_X1 _12218_ ( .A(_04463_ ), .B(fanout_net_37 ), .C1(_04464_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04465_ ) );
OR2_X1 _12219_ ( .A1(fanout_net_31 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04466_ ) );
OAI211_X1 _12220_ ( .A(_04466_ ), .B(_04459_ ), .C1(_04464_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04467_ ) );
NAND3_X1 _12221_ ( .A1(_04465_ ), .A2(_04467_ ), .A3(fanout_net_39 ), .ZN(_04468_ ) );
MUX2_X1 _12222_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04469_ ) );
MUX2_X1 _12223_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04470_ ) );
MUX2_X1 _12224_ ( .A(_04469_ ), .B(_04470_ ), .S(fanout_net_37 ), .Z(_04471_ ) );
OAI211_X1 _12225_ ( .A(fanout_net_40 ), .B(_04468_ ), .C1(_04471_ ), .C2(fanout_net_39 ), .ZN(_04472_ ) );
NAND2_X1 _12226_ ( .A1(_04462_ ), .A2(_04472_ ), .ZN(_04473_ ) );
OAI21_X1 _12227_ ( .A(_04473_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04474_ ) );
AND2_X1 _12228_ ( .A1(_04448_ ), .A2(_04474_ ), .ZN(_04475_ ) );
INV_X1 _12229_ ( .A(_04475_ ), .ZN(_04476_ ) );
XNOR2_X1 _12230_ ( .A(_02178_ ), .B(_04476_ ), .ZN(_04477_ ) );
BUF_X2 _12231_ ( .A(_04153_ ), .Z(_04478_ ) );
OR2_X1 _12232_ ( .A1(_04478_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04479_ ) );
OAI211_X1 _12233_ ( .A(_04479_ ), .B(fanout_net_37 ), .C1(fanout_net_31 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04480_ ) );
OR2_X1 _12234_ ( .A1(fanout_net_31 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04481_ ) );
OAI211_X1 _12235_ ( .A(_04481_ ), .B(_04451_ ), .C1(_04464_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04482_ ) );
NAND3_X1 _12236_ ( .A1(_04480_ ), .A2(_04461_ ), .A3(_04482_ ), .ZN(_04483_ ) );
MUX2_X1 _12237_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04484_ ) );
MUX2_X1 _12238_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04485_ ) );
MUX2_X1 _12239_ ( .A(_04484_ ), .B(_04485_ ), .S(_04451_ ), .Z(_04486_ ) );
OAI211_X1 _12240_ ( .A(_04423_ ), .B(_04483_ ), .C1(_04486_ ), .C2(_04461_ ), .ZN(_04487_ ) );
OR2_X1 _12241_ ( .A1(_04478_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04488_ ) );
OAI211_X1 _12242_ ( .A(_04488_ ), .B(_04451_ ), .C1(fanout_net_31 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04489_ ) );
NAND2_X1 _12243_ ( .A1(_02995_ ), .A2(fanout_net_31 ), .ZN(_04490_ ) );
OAI211_X1 _12244_ ( .A(_04490_ ), .B(fanout_net_37 ), .C1(fanout_net_31 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04491_ ) );
NAND3_X1 _12245_ ( .A1(_04489_ ), .A2(fanout_net_39 ), .A3(_04491_ ), .ZN(_04492_ ) );
MUX2_X1 _12246_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04493_ ) );
MUX2_X1 _12247_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04494_ ) );
MUX2_X1 _12248_ ( .A(_04493_ ), .B(_04494_ ), .S(fanout_net_37 ), .Z(_04495_ ) );
OAI211_X1 _12249_ ( .A(fanout_net_40 ), .B(_04492_ ), .C1(_04495_ ), .C2(fanout_net_39 ), .ZN(_04496_ ) );
AOI21_X1 _12250_ ( .A(_04447_ ), .B1(_04487_ ), .B2(_04496_ ), .ZN(_04497_ ) );
AND2_X1 _12251_ ( .A1(_04447_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04498_ ) );
NOR2_X1 _12252_ ( .A1(_04497_ ), .A2(_04498_ ), .ZN(_04499_ ) );
XNOR2_X1 _12253_ ( .A(_04499_ ), .B(_03006_ ), .ZN(_04500_ ) );
OR3_X1 _12254_ ( .A1(_04416_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_04417_ ), .ZN(_04501_ ) );
OR2_X1 _12255_ ( .A1(_04449_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04502_ ) );
OAI211_X1 _12256_ ( .A(_04502_ ), .B(_04459_ ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04503_ ) );
OR2_X1 _12257_ ( .A1(_04449_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04504_ ) );
OAI211_X1 _12258_ ( .A(_04504_ ), .B(fanout_net_37 ), .C1(fanout_net_31 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04505_ ) );
NAND3_X1 _12259_ ( .A1(_04503_ ), .A2(_04505_ ), .A3(fanout_net_39 ), .ZN(_04506_ ) );
MUX2_X1 _12260_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04507_ ) );
MUX2_X1 _12261_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_31 ), .Z(_04508_ ) );
MUX2_X1 _12262_ ( .A(_04507_ ), .B(_04508_ ), .S(_04459_ ), .Z(_04509_ ) );
OAI211_X1 _12263_ ( .A(_04423_ ), .B(_04506_ ), .C1(_04509_ ), .C2(fanout_net_39 ), .ZN(_04510_ ) );
NOR2_X1 _12264_ ( .A1(_04478_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04511_ ) );
OAI21_X1 _12265_ ( .A(fanout_net_37 ), .B1(fanout_net_31 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04512_ ) );
NOR2_X1 _12266_ ( .A1(fanout_net_32 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04513_ ) );
OAI21_X1 _12267_ ( .A(_04459_ ), .B1(_04478_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04514_ ) );
OAI221_X1 _12268_ ( .A(_04453_ ), .B1(_04511_ ), .B2(_04512_ ), .C1(_04513_ ), .C2(_04514_ ), .ZN(_04515_ ) );
MUX2_X1 _12269_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04516_ ) );
MUX2_X1 _12270_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04517_ ) );
MUX2_X1 _12271_ ( .A(_04516_ ), .B(_04517_ ), .S(fanout_net_37 ), .Z(_04518_ ) );
OAI211_X1 _12272_ ( .A(fanout_net_40 ), .B(_04515_ ), .C1(_04518_ ), .C2(_04461_ ), .ZN(_04519_ ) );
OAI211_X1 _12273_ ( .A(_04510_ ), .B(_04519_ ), .C1(_04416_ ), .C2(_04417_ ), .ZN(_04520_ ) );
NAND2_X1 _12274_ ( .A1(_04501_ ), .A2(_04520_ ), .ZN(_04521_ ) );
XNOR2_X1 _12275_ ( .A(_04521_ ), .B(_02209_ ), .ZN(_04522_ ) );
NAND2_X1 _12276_ ( .A1(_04447_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04523_ ) );
OR2_X1 _12277_ ( .A1(_04400_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04524_ ) );
OAI211_X1 _12278_ ( .A(_04524_ ), .B(_04436_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04525_ ) );
OR2_X1 _12279_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04526_ ) );
OAI211_X1 _12280_ ( .A(_04526_ ), .B(fanout_net_37 ), .C1(_04449_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04527_ ) );
NAND3_X1 _12281_ ( .A1(_04525_ ), .A2(_04453_ ), .A3(_04527_ ), .ZN(_04528_ ) );
MUX2_X1 _12282_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04529_ ) );
MUX2_X1 _12283_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04530_ ) );
MUX2_X1 _12284_ ( .A(_04529_ ), .B(_04530_ ), .S(_04436_ ), .Z(_04531_ ) );
OAI211_X1 _12285_ ( .A(_04423_ ), .B(_04528_ ), .C1(_04531_ ), .C2(_04453_ ), .ZN(_04532_ ) );
OR2_X1 _12286_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04533_ ) );
OAI211_X1 _12287_ ( .A(_04533_ ), .B(fanout_net_37 ), .C1(_04449_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04534_ ) );
OR2_X1 _12288_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04535_ ) );
OAI211_X1 _12289_ ( .A(_04535_ ), .B(_04436_ ), .C1(_04449_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04536_ ) );
NAND3_X1 _12290_ ( .A1(_04534_ ), .A2(_04536_ ), .A3(fanout_net_39 ), .ZN(_04537_ ) );
MUX2_X1 _12291_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04538_ ) );
MUX2_X1 _12292_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04539_ ) );
MUX2_X1 _12293_ ( .A(_04538_ ), .B(_04539_ ), .S(fanout_net_37 ), .Z(_04540_ ) );
OAI211_X1 _12294_ ( .A(fanout_net_40 ), .B(_04537_ ), .C1(_04540_ ), .C2(fanout_net_39 ), .ZN(_04541_ ) );
NAND2_X1 _12295_ ( .A1(_04532_ ), .A2(_04541_ ), .ZN(_04542_ ) );
OAI21_X1 _12296_ ( .A(_04542_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04543_ ) );
AND2_X1 _12297_ ( .A1(_04523_ ), .A2(_04543_ ), .ZN(_04544_ ) );
XNOR2_X1 _12298_ ( .A(_04544_ ), .B(_02973_ ), .ZN(_04545_ ) );
AND2_X1 _12299_ ( .A1(_04522_ ), .A2(_04545_ ), .ZN(_04546_ ) );
AND3_X1 _12300_ ( .A1(_04477_ ), .A2(_04500_ ), .A3(_04546_ ), .ZN(_04547_ ) );
NOR2_X1 _12301_ ( .A1(_04416_ ), .A2(_04417_ ), .ZN(_04548_ ) );
INV_X1 _12302_ ( .A(_04548_ ), .ZN(_04549_ ) );
OR2_X1 _12303_ ( .A1(_04449_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04550_ ) );
OAI211_X1 _12304_ ( .A(_04550_ ), .B(_04459_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04551_ ) );
OR2_X1 _12305_ ( .A1(_04153_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04552_ ) );
OAI211_X1 _12306_ ( .A(_04552_ ), .B(fanout_net_37 ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04553_ ) );
NAND3_X1 _12307_ ( .A1(_04551_ ), .A2(_04553_ ), .A3(_04453_ ), .ZN(_04554_ ) );
MUX2_X1 _12308_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04555_ ) );
MUX2_X1 _12309_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04556_ ) );
MUX2_X1 _12310_ ( .A(_04555_ ), .B(_04556_ ), .S(_04459_ ), .Z(_04557_ ) );
OAI211_X1 _12311_ ( .A(fanout_net_40 ), .B(_04554_ ), .C1(_04557_ ), .C2(_04461_ ), .ZN(_04558_ ) );
OR2_X1 _12312_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04559_ ) );
OAI211_X1 _12313_ ( .A(_04559_ ), .B(_04459_ ), .C1(_04478_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04560_ ) );
NOR2_X1 _12314_ ( .A1(_04464_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04561_ ) );
OAI21_X1 _12315_ ( .A(fanout_net_37 ), .B1(fanout_net_32 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04562_ ) );
OAI211_X1 _12316_ ( .A(_04560_ ), .B(_04453_ ), .C1(_04561_ ), .C2(_04562_ ), .ZN(_04563_ ) );
MUX2_X1 _12317_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04564_ ) );
MUX2_X1 _12318_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04565_ ) );
MUX2_X1 _12319_ ( .A(_04564_ ), .B(_04565_ ), .S(_04459_ ), .Z(_04566_ ) );
OAI211_X1 _12320_ ( .A(_04423_ ), .B(_04563_ ), .C1(_04566_ ), .C2(_04461_ ), .ZN(_04567_ ) );
NAND3_X1 _12321_ ( .A1(_04549_ ), .A2(_04558_ ), .A3(_04567_ ), .ZN(_04568_ ) );
INV_X1 _12322_ ( .A(\EX_LS_result_reg [26] ), .ZN(_04569_ ) );
OR3_X1 _12323_ ( .A1(_04416_ ), .A2(_04569_ ), .A3(_04417_ ), .ZN(_04570_ ) );
NAND2_X1 _12324_ ( .A1(_04568_ ), .A2(_04570_ ), .ZN(_04571_ ) );
XNOR2_X1 _12325_ ( .A(_04571_ ), .B(_02256_ ), .ZN(_04572_ ) );
INV_X1 _12326_ ( .A(_04572_ ), .ZN(_04573_ ) );
OR2_X1 _12327_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04574_ ) );
OAI211_X1 _12328_ ( .A(_04574_ ), .B(_04459_ ), .C1(_04478_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04575_ ) );
OR2_X1 _12329_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04576_ ) );
OAI211_X1 _12330_ ( .A(_04576_ ), .B(fanout_net_37 ), .C1(_04478_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04577_ ) );
NAND3_X1 _12331_ ( .A1(_04575_ ), .A2(_04577_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04578_ ) );
MUX2_X1 _12332_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04579_ ) );
MUX2_X1 _12333_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04580_ ) );
MUX2_X1 _12334_ ( .A(_04579_ ), .B(_04580_ ), .S(_04436_ ), .Z(_04581_ ) );
OAI211_X1 _12335_ ( .A(_04423_ ), .B(_04578_ ), .C1(_04581_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04582_ ) );
NOR2_X1 _12336_ ( .A1(_04449_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04583_ ) );
OAI21_X1 _12337_ ( .A(fanout_net_37 ), .B1(fanout_net_32 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04584_ ) );
NOR2_X1 _12338_ ( .A1(fanout_net_32 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04585_ ) );
OAI21_X1 _12339_ ( .A(_04436_ ), .B1(_04478_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04586_ ) );
OAI221_X1 _12340_ ( .A(_04453_ ), .B1(_04583_ ), .B2(_04584_ ), .C1(_04585_ ), .C2(_04586_ ), .ZN(_04587_ ) );
MUX2_X1 _12341_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04588_ ) );
MUX2_X1 _12342_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04589_ ) );
MUX2_X1 _12343_ ( .A(_04588_ ), .B(_04589_ ), .S(fanout_net_37 ), .Z(_04590_ ) );
OAI211_X1 _12344_ ( .A(fanout_net_40 ), .B(_04587_ ), .C1(_04590_ ), .C2(_04453_ ), .ZN(_04591_ ) );
NAND3_X1 _12345_ ( .A1(_04549_ ), .A2(_04582_ ), .A3(_04591_ ), .ZN(_04592_ ) );
INV_X1 _12346_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04593_ ) );
OR3_X1 _12347_ ( .A1(_04416_ ), .A2(_04593_ ), .A3(_04417_ ), .ZN(_04594_ ) );
NAND2_X1 _12348_ ( .A1(_04592_ ), .A2(_04594_ ), .ZN(_04595_ ) );
NAND2_X1 _12349_ ( .A1(_02211_ ), .A2(_02232_ ), .ZN(_04596_ ) );
INV_X1 _12350_ ( .A(_04596_ ), .ZN(_04597_ ) );
XNOR2_X1 _12351_ ( .A(_04595_ ), .B(_04597_ ), .ZN(_04598_ ) );
NOR2_X1 _12352_ ( .A1(_04573_ ), .A2(_04598_ ), .ZN(_04599_ ) );
OR2_X1 _12353_ ( .A1(_04464_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04600_ ) );
OAI211_X1 _12354_ ( .A(_04600_ ), .B(_04451_ ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04601_ ) );
OR2_X1 _12355_ ( .A1(_04478_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04602_ ) );
OAI211_X1 _12356_ ( .A(_04602_ ), .B(fanout_net_37 ), .C1(fanout_net_32 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04603_ ) );
NAND3_X1 _12357_ ( .A1(_04601_ ), .A2(_04603_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04604_ ) );
MUX2_X1 _12358_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_32 ), .Z(_04605_ ) );
MUX2_X1 _12359_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04606_ ) );
MUX2_X1 _12360_ ( .A(_04605_ ), .B(_04606_ ), .S(_04451_ ), .Z(_04607_ ) );
OAI211_X1 _12361_ ( .A(_04423_ ), .B(_04604_ ), .C1(_04607_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04608_ ) );
NOR2_X1 _12362_ ( .A1(_04464_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04609_ ) );
OAI21_X1 _12363_ ( .A(fanout_net_37 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04610_ ) );
NOR2_X1 _12364_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04611_ ) );
OAI21_X1 _12365_ ( .A(_04451_ ), .B1(_04464_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04612_ ) );
OAI221_X1 _12366_ ( .A(_04461_ ), .B1(_04609_ ), .B2(_04610_ ), .C1(_04611_ ), .C2(_04612_ ), .ZN(_04613_ ) );
MUX2_X1 _12367_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04614_ ) );
MUX2_X1 _12368_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04615_ ) );
MUX2_X1 _12369_ ( .A(_04614_ ), .B(_04615_ ), .S(fanout_net_37 ), .Z(_04616_ ) );
OAI211_X1 _12370_ ( .A(fanout_net_40 ), .B(_04613_ ), .C1(_04616_ ), .C2(_04461_ ), .ZN(_04617_ ) );
NAND3_X1 _12371_ ( .A1(_04549_ ), .A2(_04608_ ), .A3(_04617_ ), .ZN(_04618_ ) );
INV_X1 _12372_ ( .A(\EX_LS_result_reg [24] ), .ZN(_04619_ ) );
OR3_X1 _12373_ ( .A1(_04416_ ), .A2(_04619_ ), .A3(_04417_ ), .ZN(_04620_ ) );
AND2_X1 _12374_ ( .A1(_04618_ ), .A2(_04620_ ), .ZN(_04621_ ) );
INV_X1 _12375_ ( .A(_02915_ ), .ZN(_04622_ ) );
XNOR2_X1 _12376_ ( .A(_04621_ ), .B(_04622_ ), .ZN(_04623_ ) );
OR2_X1 _12377_ ( .A1(_04464_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04624_ ) );
OAI211_X1 _12378_ ( .A(_04624_ ), .B(_04451_ ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04625_ ) );
OR2_X1 _12379_ ( .A1(_04478_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04626_ ) );
OAI211_X1 _12380_ ( .A(_04626_ ), .B(fanout_net_37 ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04627_ ) );
NAND3_X1 _12381_ ( .A1(_04625_ ), .A2(_04627_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04628_ ) );
MUX2_X1 _12382_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04629_ ) );
MUX2_X1 _12383_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04630_ ) );
MUX2_X1 _12384_ ( .A(_04629_ ), .B(_04630_ ), .S(_04451_ ), .Z(_04631_ ) );
OAI211_X1 _12385_ ( .A(_04423_ ), .B(_04628_ ), .C1(_04631_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04632_ ) );
NOR2_X1 _12386_ ( .A1(_04464_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04633_ ) );
OAI21_X1 _12387_ ( .A(fanout_net_37 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04634_ ) );
NOR2_X1 _12388_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04635_ ) );
OAI21_X1 _12389_ ( .A(_04451_ ), .B1(_04464_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04636_ ) );
OAI221_X1 _12390_ ( .A(_04461_ ), .B1(_04633_ ), .B2(_04634_ ), .C1(_04635_ ), .C2(_04636_ ), .ZN(_04637_ ) );
MUX2_X1 _12391_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04638_ ) );
MUX2_X1 _12392_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04639_ ) );
MUX2_X1 _12393_ ( .A(_04638_ ), .B(_04639_ ), .S(fanout_net_37 ), .Z(_04640_ ) );
OAI211_X1 _12394_ ( .A(fanout_net_40 ), .B(_04637_ ), .C1(_04640_ ), .C2(_04461_ ), .ZN(_04641_ ) );
NAND3_X1 _12395_ ( .A1(_04549_ ), .A2(_04632_ ), .A3(_04641_ ), .ZN(_04642_ ) );
INV_X1 _12396_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04643_ ) );
OR3_X1 _12397_ ( .A1(_04416_ ), .A2(_04643_ ), .A3(_04417_ ), .ZN(_04644_ ) );
NAND2_X1 _12398_ ( .A1(_04642_ ), .A2(_04644_ ), .ZN(_04645_ ) );
NAND2_X1 _12399_ ( .A1(_04645_ ), .A2(_02946_ ), .ZN(_04646_ ) );
NAND3_X1 _12400_ ( .A1(_04642_ ), .A2(_02938_ ), .A3(_04644_ ), .ZN(_04647_ ) );
AND2_X1 _12401_ ( .A1(_04646_ ), .A2(_04647_ ), .ZN(_04648_ ) );
AND2_X1 _12402_ ( .A1(_04623_ ), .A2(_04648_ ), .ZN(_04649_ ) );
AND3_X1 _12403_ ( .A1(_04547_ ), .A2(_04599_ ), .A3(_04649_ ), .ZN(_04650_ ) );
INV_X1 _12404_ ( .A(_02382_ ), .ZN(_04651_ ) );
INV_X1 _12405_ ( .A(\EX_LS_result_reg [19] ), .ZN(_04652_ ) );
OR3_X1 _12406_ ( .A1(_04100_ ), .A2(_04652_ ), .A3(_04103_ ), .ZN(_04653_ ) );
OR2_X1 _12407_ ( .A1(_04108_ ), .A2(\myreg.Reg[1][19] ), .ZN(_04654_ ) );
OAI211_X1 _12408_ ( .A(_04654_ ), .B(_04112_ ), .C1(fanout_net_33 ), .C2(\myreg.Reg[0][19] ), .ZN(_04655_ ) );
OR2_X1 _12409_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[2][19] ), .ZN(_04656_ ) );
OAI211_X1 _12410_ ( .A(_04656_ ), .B(fanout_net_37 ), .C1(_04152_ ), .C2(\myreg.Reg[3][19] ), .ZN(_04657_ ) );
NAND3_X1 _12411_ ( .A1(_04655_ ), .A2(_04115_ ), .A3(_04657_ ), .ZN(_04658_ ) );
MUX2_X1 _12412_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_33 ), .Z(_04659_ ) );
MUX2_X1 _12413_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_33 ), .Z(_04660_ ) );
MUX2_X1 _12414_ ( .A(_04659_ ), .B(_04660_ ), .S(_04123_ ), .Z(_04661_ ) );
OAI211_X1 _12415_ ( .A(_04106_ ), .B(_04658_ ), .C1(_04661_ ), .C2(_04126_ ), .ZN(_04662_ ) );
OR2_X1 _12416_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[14][19] ), .ZN(_04663_ ) );
OAI211_X1 _12417_ ( .A(_04663_ ), .B(fanout_net_37 ), .C1(_04152_ ), .C2(\myreg.Reg[15][19] ), .ZN(_04664_ ) );
OR2_X1 _12418_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[12][19] ), .ZN(_04665_ ) );
OAI211_X1 _12419_ ( .A(_04665_ ), .B(_04123_ ), .C1(_04152_ ), .C2(\myreg.Reg[13][19] ), .ZN(_04666_ ) );
NAND3_X1 _12420_ ( .A1(_04664_ ), .A2(_04666_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04667_ ) );
MUX2_X1 _12421_ ( .A(\myreg.Reg[8][19] ), .B(\myreg.Reg[9][19] ), .S(fanout_net_33 ), .Z(_04668_ ) );
MUX2_X1 _12422_ ( .A(\myreg.Reg[10][19] ), .B(\myreg.Reg[11][19] ), .S(fanout_net_33 ), .Z(_04669_ ) );
MUX2_X1 _12423_ ( .A(_04668_ ), .B(_04669_ ), .S(fanout_net_37 ), .Z(_04670_ ) );
OAI211_X1 _12424_ ( .A(fanout_net_40 ), .B(_04667_ ), .C1(_04670_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04671_ ) );
NAND2_X1 _12425_ ( .A1(_04662_ ), .A2(_04671_ ), .ZN(_04672_ ) );
OAI21_X1 _12426_ ( .A(_04672_ ), .B1(_04253_ ), .B2(_04138_ ), .ZN(_04673_ ) );
AND2_X1 _12427_ ( .A1(_04653_ ), .A2(_04673_ ), .ZN(_04674_ ) );
XNOR2_X1 _12428_ ( .A(_04651_ ), .B(_04674_ ), .ZN(_04675_ ) );
NOR2_X1 _12429_ ( .A1(_04310_ ), .A2(\myreg.Reg[11][18] ), .ZN(_04676_ ) );
OAI21_X1 _12430_ ( .A(fanout_net_38 ), .B1(fanout_net_33 ), .B2(\myreg.Reg[10][18] ), .ZN(_04677_ ) );
NOR2_X1 _12431_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[8][18] ), .ZN(_04678_ ) );
OAI21_X1 _12432_ ( .A(_04314_ ), .B1(_04310_ ), .B2(\myreg.Reg[9][18] ), .ZN(_04679_ ) );
OAI221_X1 _12433_ ( .A(_04265_ ), .B1(_04676_ ), .B2(_04677_ ), .C1(_04678_ ), .C2(_04679_ ), .ZN(_04680_ ) );
MUX2_X1 _12434_ ( .A(\myreg.Reg[12][18] ), .B(\myreg.Reg[13][18] ), .S(fanout_net_33 ), .Z(_04681_ ) );
MUX2_X1 _12435_ ( .A(\myreg.Reg[14][18] ), .B(\myreg.Reg[15][18] ), .S(fanout_net_33 ), .Z(_04682_ ) );
MUX2_X1 _12436_ ( .A(_04681_ ), .B(_04682_ ), .S(fanout_net_38 ), .Z(_04683_ ) );
OAI211_X1 _12437_ ( .A(fanout_net_40 ), .B(_04680_ ), .C1(_04683_ ), .C2(_04157_ ), .ZN(_04684_ ) );
OR2_X1 _12438_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[4][18] ), .ZN(_04685_ ) );
OAI211_X1 _12439_ ( .A(_04685_ ), .B(_04314_ ), .C1(_04400_ ), .C2(\myreg.Reg[5][18] ), .ZN(_04686_ ) );
OR2_X1 _12440_ ( .A1(fanout_net_33 ), .A2(\myreg.Reg[6][18] ), .ZN(_04687_ ) );
OAI211_X1 _12441_ ( .A(_04687_ ), .B(fanout_net_38 ), .C1(_04400_ ), .C2(\myreg.Reg[7][18] ), .ZN(_04688_ ) );
NAND3_X1 _12442_ ( .A1(_04686_ ), .A2(_04688_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04689_ ) );
MUX2_X1 _12443_ ( .A(\myreg.Reg[2][18] ), .B(\myreg.Reg[3][18] ), .S(fanout_net_33 ), .Z(_04690_ ) );
MUX2_X1 _12444_ ( .A(\myreg.Reg[0][18] ), .B(\myreg.Reg[1][18] ), .S(fanout_net_33 ), .Z(_04691_ ) );
MUX2_X1 _12445_ ( .A(_04690_ ), .B(_04691_ ), .S(_04314_ ), .Z(_04692_ ) );
OAI211_X1 _12446_ ( .A(_04148_ ), .B(_04689_ ), .C1(_04692_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04693_ ) );
NAND2_X1 _12447_ ( .A1(_04684_ ), .A2(_04693_ ), .ZN(_04694_ ) );
OAI21_X1 _12448_ ( .A(_04694_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04695_ ) );
NAND4_X1 _12449_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [18] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04696_ ) );
AND2_X1 _12450_ ( .A1(_04695_ ), .A2(_04696_ ), .ZN(_04697_ ) );
XOR2_X1 _12451_ ( .A(_02405_ ), .B(_04697_ ), .Z(_04698_ ) );
AND2_X1 _12452_ ( .A1(_04675_ ), .A2(_04698_ ), .ZN(_04699_ ) );
NOR2_X1 _12453_ ( .A1(_04449_ ), .A2(\myreg.Reg[11][16] ), .ZN(_04700_ ) );
OAI21_X1 _12454_ ( .A(fanout_net_38 ), .B1(fanout_net_33 ), .B2(\myreg.Reg[10][16] ), .ZN(_04701_ ) );
NOR2_X1 _12455_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[8][16] ), .ZN(_04702_ ) );
OAI21_X1 _12456_ ( .A(_04436_ ), .B1(_04449_ ), .B2(\myreg.Reg[9][16] ), .ZN(_04703_ ) );
OAI221_X1 _12457_ ( .A(_04157_ ), .B1(_04700_ ), .B2(_04701_ ), .C1(_04702_ ), .C2(_04703_ ), .ZN(_04704_ ) );
MUX2_X1 _12458_ ( .A(\myreg.Reg[12][16] ), .B(\myreg.Reg[13][16] ), .S(fanout_net_34 ), .Z(_04705_ ) );
MUX2_X1 _12459_ ( .A(\myreg.Reg[14][16] ), .B(\myreg.Reg[15][16] ), .S(fanout_net_34 ), .Z(_04706_ ) );
MUX2_X1 _12460_ ( .A(_04705_ ), .B(_04706_ ), .S(fanout_net_38 ), .Z(_04707_ ) );
OAI211_X1 _12461_ ( .A(fanout_net_40 ), .B(_04704_ ), .C1(_04707_ ), .C2(_04453_ ), .ZN(_04708_ ) );
OR2_X1 _12462_ ( .A1(_04153_ ), .A2(\myreg.Reg[5][16] ), .ZN(_04709_ ) );
OAI211_X1 _12463_ ( .A(_04709_ ), .B(_04436_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[4][16] ), .ZN(_04710_ ) );
OR2_X1 _12464_ ( .A1(_04400_ ), .A2(\myreg.Reg[7][16] ), .ZN(_04711_ ) );
OAI211_X1 _12465_ ( .A(_04711_ ), .B(fanout_net_38 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[6][16] ), .ZN(_04712_ ) );
NAND3_X1 _12466_ ( .A1(_04710_ ), .A2(_04712_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04713_ ) );
MUX2_X1 _12467_ ( .A(\myreg.Reg[2][16] ), .B(\myreg.Reg[3][16] ), .S(fanout_net_34 ), .Z(_04714_ ) );
MUX2_X1 _12468_ ( .A(\myreg.Reg[0][16] ), .B(\myreg.Reg[1][16] ), .S(fanout_net_34 ), .Z(_04715_ ) );
MUX2_X1 _12469_ ( .A(_04714_ ), .B(_04715_ ), .S(_04436_ ), .Z(_04716_ ) );
OAI211_X1 _12470_ ( .A(_04423_ ), .B(_04713_ ), .C1(_04716_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04717_ ) );
NAND2_X1 _12471_ ( .A1(_04708_ ), .A2(_04717_ ), .ZN(_04718_ ) );
OAI21_X1 _12472_ ( .A(_04718_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04719_ ) );
NAND4_X1 _12473_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [16] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04720_ ) );
AND2_X1 _12474_ ( .A1(_04719_ ), .A2(_04720_ ), .ZN(_04721_ ) );
XOR2_X1 _12475_ ( .A(_02454_ ), .B(_04721_ ), .Z(_04722_ ) );
INV_X1 _12476_ ( .A(_02430_ ), .ZN(_04723_ ) );
INV_X1 _12477_ ( .A(\EX_LS_result_reg [17] ), .ZN(_04724_ ) );
OR3_X1 _12478_ ( .A1(_04100_ ), .A2(_04724_ ), .A3(_04103_ ), .ZN(_04725_ ) );
OR2_X1 _12479_ ( .A1(_04309_ ), .A2(\myreg.Reg[3][17] ), .ZN(_04726_ ) );
OAI211_X1 _12480_ ( .A(_04726_ ), .B(fanout_net_38 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[2][17] ), .ZN(_04727_ ) );
OR2_X1 _12481_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[0][17] ), .ZN(_04728_ ) );
OAI211_X1 _12482_ ( .A(_04728_ ), .B(_04268_ ), .C1(_04352_ ), .C2(\myreg.Reg[1][17] ), .ZN(_04729_ ) );
NAND3_X1 _12483_ ( .A1(_04727_ ), .A2(_04115_ ), .A3(_04729_ ), .ZN(_04730_ ) );
MUX2_X1 _12484_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_34 ), .Z(_04731_ ) );
MUX2_X1 _12485_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_34 ), .Z(_04732_ ) );
MUX2_X1 _12486_ ( .A(_04731_ ), .B(_04732_ ), .S(_04268_ ), .Z(_04733_ ) );
OAI211_X1 _12487_ ( .A(_04106_ ), .B(_04730_ ), .C1(_04733_ ), .C2(_04265_ ), .ZN(_04734_ ) );
OR2_X1 _12488_ ( .A1(_04309_ ), .A2(\myreg.Reg[15][17] ), .ZN(_04735_ ) );
OAI211_X1 _12489_ ( .A(_04735_ ), .B(fanout_net_38 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[14][17] ), .ZN(_04736_ ) );
OR2_X1 _12490_ ( .A1(_04151_ ), .A2(\myreg.Reg[13][17] ), .ZN(_04737_ ) );
OAI211_X1 _12491_ ( .A(_04737_ ), .B(_04268_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[12][17] ), .ZN(_04738_ ) );
NAND3_X1 _12492_ ( .A1(_04736_ ), .A2(_04738_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04739_ ) );
MUX2_X1 _12493_ ( .A(\myreg.Reg[8][17] ), .B(\myreg.Reg[9][17] ), .S(fanout_net_34 ), .Z(_04740_ ) );
MUX2_X1 _12494_ ( .A(\myreg.Reg[10][17] ), .B(\myreg.Reg[11][17] ), .S(fanout_net_34 ), .Z(_04741_ ) );
MUX2_X1 _12495_ ( .A(_04740_ ), .B(_04741_ ), .S(fanout_net_38 ), .Z(_04742_ ) );
OAI211_X1 _12496_ ( .A(fanout_net_40 ), .B(_04739_ ), .C1(_04742_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04743_ ) );
NAND2_X1 _12497_ ( .A1(_04734_ ), .A2(_04743_ ), .ZN(_04744_ ) );
OAI21_X1 _12498_ ( .A(_04744_ ), .B1(_04253_ ), .B2(_04138_ ), .ZN(_04745_ ) );
AND2_X1 _12499_ ( .A1(_04725_ ), .A2(_04745_ ), .ZN(_04746_ ) );
XNOR2_X1 _12500_ ( .A(_04723_ ), .B(_04746_ ), .ZN(_04747_ ) );
AND3_X1 _12501_ ( .A1(_04699_ ), .A2(_04722_ ), .A3(_04747_ ), .ZN(_04748_ ) );
INV_X1 _12502_ ( .A(_02305_ ), .ZN(_04749_ ) );
INV_X1 _12503_ ( .A(\EX_LS_result_reg [22] ), .ZN(_04750_ ) );
OR3_X1 _12504_ ( .A1(_04253_ ), .A2(_04750_ ), .A3(_04138_ ), .ZN(_04751_ ) );
OR2_X1 _12505_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[0][22] ), .ZN(_04752_ ) );
OAI211_X1 _12506_ ( .A(_04752_ ), .B(_04314_ ), .C1(_04400_ ), .C2(\myreg.Reg[1][22] ), .ZN(_04753_ ) );
OR2_X1 _12507_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[2][22] ), .ZN(_04754_ ) );
OAI211_X1 _12508_ ( .A(_04754_ ), .B(fanout_net_38 ), .C1(_04400_ ), .C2(\myreg.Reg[3][22] ), .ZN(_04755_ ) );
NAND3_X1 _12509_ ( .A1(_04753_ ), .A2(_04755_ ), .A3(_04265_ ), .ZN(_04756_ ) );
MUX2_X1 _12510_ ( .A(\myreg.Reg[6][22] ), .B(\myreg.Reg[7][22] ), .S(fanout_net_34 ), .Z(_04757_ ) );
MUX2_X1 _12511_ ( .A(\myreg.Reg[4][22] ), .B(\myreg.Reg[5][22] ), .S(fanout_net_34 ), .Z(_04758_ ) );
MUX2_X1 _12512_ ( .A(_04757_ ), .B(_04758_ ), .S(_04218_ ), .Z(_04759_ ) );
OAI211_X1 _12513_ ( .A(_04148_ ), .B(_04756_ ), .C1(_04759_ ), .C2(_04157_ ), .ZN(_04760_ ) );
OR2_X1 _12514_ ( .A1(_04118_ ), .A2(\myreg.Reg[15][22] ), .ZN(_04761_ ) );
OAI211_X1 _12515_ ( .A(_04761_ ), .B(fanout_net_38 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[14][22] ), .ZN(_04762_ ) );
OR2_X1 _12516_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[12][22] ), .ZN(_04763_ ) );
OAI211_X1 _12517_ ( .A(_04763_ ), .B(_04314_ ), .C1(_04310_ ), .C2(\myreg.Reg[13][22] ), .ZN(_04764_ ) );
NAND3_X1 _12518_ ( .A1(_04762_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04764_ ), .ZN(_04765_ ) );
MUX2_X1 _12519_ ( .A(\myreg.Reg[8][22] ), .B(\myreg.Reg[9][22] ), .S(fanout_net_34 ), .Z(_04766_ ) );
MUX2_X1 _12520_ ( .A(\myreg.Reg[10][22] ), .B(\myreg.Reg[11][22] ), .S(fanout_net_34 ), .Z(_04767_ ) );
MUX2_X1 _12521_ ( .A(_04766_ ), .B(_04767_ ), .S(fanout_net_38 ), .Z(_04768_ ) );
OAI211_X1 _12522_ ( .A(fanout_net_40 ), .B(_04765_ ), .C1(_04768_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04769_ ) );
NAND2_X1 _12523_ ( .A1(_04760_ ), .A2(_04769_ ), .ZN(_04770_ ) );
OAI21_X1 _12524_ ( .A(_04770_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04771_ ) );
AND2_X1 _12525_ ( .A1(_04751_ ), .A2(_04771_ ), .ZN(_04772_ ) );
XNOR2_X1 _12526_ ( .A(_04749_ ), .B(_04772_ ), .ZN(_04773_ ) );
OR2_X1 _12527_ ( .A1(_04309_ ), .A2(\myreg.Reg[1][23] ), .ZN(_04774_ ) );
OAI211_X1 _12528_ ( .A(_04774_ ), .B(_04218_ ), .C1(fanout_net_34 ), .C2(\myreg.Reg[0][23] ), .ZN(_04775_ ) );
OR2_X1 _12529_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[2][23] ), .ZN(_04776_ ) );
OAI211_X1 _12530_ ( .A(_04776_ ), .B(fanout_net_38 ), .C1(_04310_ ), .C2(\myreg.Reg[3][23] ), .ZN(_04777_ ) );
NAND3_X1 _12531_ ( .A1(_04775_ ), .A2(_04126_ ), .A3(_04777_ ), .ZN(_04778_ ) );
MUX2_X1 _12532_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_34 ), .Z(_04779_ ) );
MUX2_X1 _12533_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_34 ), .Z(_04780_ ) );
MUX2_X1 _12534_ ( .A(_04779_ ), .B(_04780_ ), .S(_04268_ ), .Z(_04781_ ) );
OAI211_X1 _12535_ ( .A(_04148_ ), .B(_04778_ ), .C1(_04781_ ), .C2(_04265_ ), .ZN(_04782_ ) );
OR2_X1 _12536_ ( .A1(_04309_ ), .A2(\myreg.Reg[15][23] ), .ZN(_04783_ ) );
OAI211_X1 _12537_ ( .A(_04783_ ), .B(fanout_net_38 ), .C1(fanout_net_34 ), .C2(\myreg.Reg[14][23] ), .ZN(_04784_ ) );
OR2_X1 _12538_ ( .A1(fanout_net_34 ), .A2(\myreg.Reg[12][23] ), .ZN(_04785_ ) );
OAI211_X1 _12539_ ( .A(_04785_ ), .B(_04218_ ), .C1(_04352_ ), .C2(\myreg.Reg[13][23] ), .ZN(_04786_ ) );
NAND3_X1 _12540_ ( .A1(_04784_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04786_ ), .ZN(_04787_ ) );
MUX2_X1 _12541_ ( .A(\myreg.Reg[8][23] ), .B(\myreg.Reg[9][23] ), .S(fanout_net_34 ), .Z(_04788_ ) );
MUX2_X1 _12542_ ( .A(\myreg.Reg[10][23] ), .B(\myreg.Reg[11][23] ), .S(fanout_net_35 ), .Z(_04789_ ) );
MUX2_X1 _12543_ ( .A(_04788_ ), .B(_04789_ ), .S(fanout_net_38 ), .Z(_04790_ ) );
OAI211_X1 _12544_ ( .A(fanout_net_40 ), .B(_04787_ ), .C1(_04790_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04791_ ) );
NAND2_X1 _12545_ ( .A1(_04782_ ), .A2(_04791_ ), .ZN(_04792_ ) );
OAI21_X1 _12546_ ( .A(_04792_ ), .B1(_04253_ ), .B2(_04138_ ), .ZN(_04793_ ) );
INV_X1 _12547_ ( .A(\EX_LS_result_reg [23] ), .ZN(_04794_ ) );
OR3_X1 _12548_ ( .A1(_04253_ ), .A2(_04794_ ), .A3(_04103_ ), .ZN(_04795_ ) );
AND3_X1 _12549_ ( .A1(_02282_ ), .A2(_04793_ ), .A3(_04795_ ), .ZN(_04796_ ) );
AOI21_X1 _12550_ ( .A(_02282_ ), .B1(_04793_ ), .B2(_04795_ ), .ZN(_04797_ ) );
NOR2_X1 _12551_ ( .A1(_04796_ ), .A2(_04797_ ), .ZN(_04798_ ) );
AND2_X1 _12552_ ( .A1(_04773_ ), .A2(_04798_ ), .ZN(_04799_ ) );
NOR2_X1 _12553_ ( .A1(_04400_ ), .A2(\myreg.Reg[11][20] ), .ZN(_04800_ ) );
OAI21_X1 _12554_ ( .A(fanout_net_38 ), .B1(fanout_net_35 ), .B2(\myreg.Reg[10][20] ), .ZN(_04801_ ) );
NOR2_X1 _12555_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[8][20] ), .ZN(_04802_ ) );
OAI21_X1 _12556_ ( .A(_04150_ ), .B1(_04400_ ), .B2(\myreg.Reg[9][20] ), .ZN(_04803_ ) );
OAI221_X1 _12557_ ( .A(_04265_ ), .B1(_04800_ ), .B2(_04801_ ), .C1(_04802_ ), .C2(_04803_ ), .ZN(_04804_ ) );
MUX2_X1 _12558_ ( .A(\myreg.Reg[12][20] ), .B(\myreg.Reg[13][20] ), .S(fanout_net_35 ), .Z(_04805_ ) );
MUX2_X1 _12559_ ( .A(\myreg.Reg[14][20] ), .B(\myreg.Reg[15][20] ), .S(fanout_net_35 ), .Z(_04806_ ) );
MUX2_X1 _12560_ ( .A(_04805_ ), .B(_04806_ ), .S(fanout_net_38 ), .Z(_04807_ ) );
OAI211_X1 _12561_ ( .A(fanout_net_40 ), .B(_04804_ ), .C1(_04807_ ), .C2(_04157_ ), .ZN(_04808_ ) );
OR2_X1 _12562_ ( .A1(_04352_ ), .A2(\myreg.Reg[5][20] ), .ZN(_04809_ ) );
OAI211_X1 _12563_ ( .A(_04809_ ), .B(_04150_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[4][20] ), .ZN(_04810_ ) );
OR2_X1 _12564_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[6][20] ), .ZN(_04811_ ) );
OAI211_X1 _12565_ ( .A(_04811_ ), .B(fanout_net_38 ), .C1(_04153_ ), .C2(\myreg.Reg[7][20] ), .ZN(_04812_ ) );
NAND3_X1 _12566_ ( .A1(_04810_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04812_ ), .ZN(_04813_ ) );
MUX2_X1 _12567_ ( .A(\myreg.Reg[2][20] ), .B(\myreg.Reg[3][20] ), .S(fanout_net_35 ), .Z(_04814_ ) );
MUX2_X1 _12568_ ( .A(\myreg.Reg[0][20] ), .B(\myreg.Reg[1][20] ), .S(fanout_net_35 ), .Z(_04815_ ) );
MUX2_X1 _12569_ ( .A(_04814_ ), .B(_04815_ ), .S(_04150_ ), .Z(_04816_ ) );
OAI211_X1 _12570_ ( .A(_04148_ ), .B(_04813_ ), .C1(_04816_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04817_ ) );
NAND2_X1 _12571_ ( .A1(_04808_ ), .A2(_04817_ ), .ZN(_04818_ ) );
OAI21_X1 _12572_ ( .A(_04818_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04819_ ) );
NAND4_X1 _12573_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [20] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04820_ ) );
AND2_X1 _12574_ ( .A1(_04819_ ), .A2(_04820_ ), .ZN(_04821_ ) );
XOR2_X1 _12575_ ( .A(_02329_ ), .B(_04821_ ), .Z(_04822_ ) );
NAND2_X1 _12576_ ( .A1(_02332_ ), .A2(_02352_ ), .ZN(_04823_ ) );
NOR2_X1 _12577_ ( .A1(_04352_ ), .A2(\myreg.Reg[11][21] ), .ZN(_04824_ ) );
OAI21_X1 _12578_ ( .A(fanout_net_38 ), .B1(fanout_net_35 ), .B2(\myreg.Reg[10][21] ), .ZN(_04825_ ) );
NOR2_X1 _12579_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[8][21] ), .ZN(_04826_ ) );
OAI21_X1 _12580_ ( .A(_04268_ ), .B1(_04352_ ), .B2(\myreg.Reg[9][21] ), .ZN(_04827_ ) );
OAI221_X1 _12581_ ( .A(_04115_ ), .B1(_04824_ ), .B2(_04825_ ), .C1(_04826_ ), .C2(_04827_ ), .ZN(_04828_ ) );
MUX2_X1 _12582_ ( .A(\myreg.Reg[12][21] ), .B(\myreg.Reg[13][21] ), .S(fanout_net_35 ), .Z(_04829_ ) );
MUX2_X1 _12583_ ( .A(\myreg.Reg[14][21] ), .B(\myreg.Reg[15][21] ), .S(fanout_net_35 ), .Z(_04830_ ) );
MUX2_X1 _12584_ ( .A(_04829_ ), .B(_04830_ ), .S(fanout_net_38 ), .Z(_04831_ ) );
OAI211_X1 _12585_ ( .A(fanout_net_40 ), .B(_04828_ ), .C1(_04831_ ), .C2(_04265_ ), .ZN(_04832_ ) );
OR2_X1 _12586_ ( .A1(_04309_ ), .A2(\myreg.Reg[7][21] ), .ZN(_04833_ ) );
OAI211_X1 _12587_ ( .A(_04833_ ), .B(fanout_net_38 ), .C1(fanout_net_35 ), .C2(\myreg.Reg[6][21] ), .ZN(_04834_ ) );
OR2_X1 _12588_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[4][21] ), .ZN(_04835_ ) );
OAI211_X1 _12589_ ( .A(_04835_ ), .B(_04218_ ), .C1(_04352_ ), .C2(\myreg.Reg[5][21] ), .ZN(_04836_ ) );
NAND3_X1 _12590_ ( .A1(_04834_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04836_ ), .ZN(_04837_ ) );
MUX2_X1 _12591_ ( .A(\myreg.Reg[2][21] ), .B(\myreg.Reg[3][21] ), .S(fanout_net_35 ), .Z(_04838_ ) );
MUX2_X1 _12592_ ( .A(\myreg.Reg[0][21] ), .B(\myreg.Reg[1][21] ), .S(fanout_net_35 ), .Z(_04839_ ) );
MUX2_X1 _12593_ ( .A(_04838_ ), .B(_04839_ ), .S(_04268_ ), .Z(_04840_ ) );
OAI211_X1 _12594_ ( .A(_04148_ ), .B(_04837_ ), .C1(_04840_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04841_ ) );
NAND2_X1 _12595_ ( .A1(_04832_ ), .A2(_04841_ ), .ZN(_04842_ ) );
OAI21_X1 _12596_ ( .A(_04842_ ), .B1(_04145_ ), .B2(_04173_ ), .ZN(_04843_ ) );
NAND4_X1 _12597_ ( .A1(_04198_ ), .A2(\EX_LS_result_reg [21] ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04844_ ) );
AND2_X1 _12598_ ( .A1(_04843_ ), .A2(_04844_ ), .ZN(_04845_ ) );
AND2_X1 _12599_ ( .A1(_04823_ ), .A2(_04845_ ), .ZN(_04846_ ) );
NOR2_X1 _12600_ ( .A1(_04823_ ), .A2(_04845_ ), .ZN(_04847_ ) );
NOR2_X1 _12601_ ( .A1(_04846_ ), .A2(_04847_ ), .ZN(_04848_ ) );
AND3_X1 _12602_ ( .A1(_04799_ ), .A2(_04822_ ), .A3(_04848_ ), .ZN(_04849_ ) );
AND2_X1 _12603_ ( .A1(_04748_ ), .A2(_04849_ ), .ZN(_04850_ ) );
AND2_X1 _12604_ ( .A1(_04650_ ), .A2(_04850_ ), .ZN(_04851_ ) );
AND2_X1 _12605_ ( .A1(_04446_ ), .A2(_04851_ ), .ZN(_04852_ ) );
NAND2_X1 _12606_ ( .A1(_02502_ ), .A2(_04386_ ), .ZN(_04853_ ) );
OR2_X1 _12607_ ( .A1(_04151_ ), .A2(\myreg.Reg[9][4] ), .ZN(_04854_ ) );
OAI211_X1 _12608_ ( .A(_04854_ ), .B(_04268_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[8][4] ), .ZN(_04855_ ) );
OR2_X1 _12609_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[10][4] ), .ZN(_04856_ ) );
OAI211_X1 _12610_ ( .A(_04856_ ), .B(fanout_net_38 ), .C1(_04352_ ), .C2(\myreg.Reg[11][4] ), .ZN(_04857_ ) );
NAND3_X1 _12611_ ( .A1(_04855_ ), .A2(_04115_ ), .A3(_04857_ ), .ZN(_04858_ ) );
MUX2_X1 _12612_ ( .A(\myreg.Reg[14][4] ), .B(\myreg.Reg[15][4] ), .S(fanout_net_35 ), .Z(_04859_ ) );
MUX2_X1 _12613_ ( .A(\myreg.Reg[12][4] ), .B(\myreg.Reg[13][4] ), .S(fanout_net_35 ), .Z(_04860_ ) );
MUX2_X1 _12614_ ( .A(_04859_ ), .B(_04860_ ), .S(_04112_ ), .Z(_04861_ ) );
OAI211_X1 _12615_ ( .A(fanout_net_40 ), .B(_04858_ ), .C1(_04861_ ), .C2(_04265_ ), .ZN(_04862_ ) );
MUX2_X1 _12616_ ( .A(\myreg.Reg[2][4] ), .B(\myreg.Reg[3][4] ), .S(fanout_net_35 ), .Z(_04863_ ) );
AND2_X1 _12617_ ( .A1(_04863_ ), .A2(fanout_net_38 ), .ZN(_04864_ ) );
MUX2_X1 _12618_ ( .A(\myreg.Reg[0][4] ), .B(\myreg.Reg[1][4] ), .S(fanout_net_35 ), .Z(_04865_ ) );
AOI211_X1 _12619_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_04864_ ), .C1(_04150_ ), .C2(_04865_ ), .ZN(_04866_ ) );
MUX2_X1 _12620_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_35 ), .Z(_04867_ ) );
MUX2_X1 _12621_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_35 ), .Z(_04868_ ) );
MUX2_X1 _12622_ ( .A(_04867_ ), .B(_04868_ ), .S(_04207_ ), .Z(_04869_ ) );
OAI21_X1 _12623_ ( .A(_04106_ ), .B1(_04869_ ), .B2(_04115_ ), .ZN(_04870_ ) );
OAI221_X1 _12624_ ( .A(_04862_ ), .B1(_04866_ ), .B2(_04870_ ), .C1(_04394_ ), .C2(_04395_ ), .ZN(_04871_ ) );
OR3_X4 _12625_ ( .A1(_04394_ ), .A2(\EX_LS_result_reg [4] ), .A3(_04395_ ), .ZN(_04872_ ) );
NAND2_X2 _12626_ ( .A1(_04871_ ), .A2(_04872_ ), .ZN(_04873_ ) );
XNOR2_X1 _12627_ ( .A(_02656_ ), .B(_04873_ ), .ZN(_04874_ ) );
NAND2_X1 _12628_ ( .A1(_04447_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04875_ ) );
OR2_X1 _12629_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04876_ ) );
OAI211_X1 _12630_ ( .A(_04876_ ), .B(_04123_ ), .C1(_04152_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04877_ ) );
OR2_X1 _12631_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04878_ ) );
OAI211_X1 _12632_ ( .A(_04878_ ), .B(fanout_net_38 ), .C1(_04118_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04879_ ) );
NAND3_X1 _12633_ ( .A1(_04877_ ), .A2(_04879_ ), .A3(_04125_ ), .ZN(_04880_ ) );
MUX2_X1 _12634_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04881_ ) );
MUX2_X1 _12635_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04882_ ) );
MUX2_X1 _12636_ ( .A(_04881_ ), .B(_04882_ ), .S(_04207_ ), .Z(_04883_ ) );
OAI211_X1 _12637_ ( .A(_04106_ ), .B(_04880_ ), .C1(_04883_ ), .C2(_04126_ ), .ZN(_04884_ ) );
OR2_X1 _12638_ ( .A1(_04108_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04885_ ) );
OAI211_X1 _12639_ ( .A(_04885_ ), .B(_04123_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04886_ ) );
OR2_X1 _12640_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04887_ ) );
OAI211_X1 _12641_ ( .A(_04887_ ), .B(fanout_net_38 ), .C1(_04118_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04888_ ) );
NAND3_X1 _12642_ ( .A1(_04886_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04888_ ), .ZN(_04889_ ) );
MUX2_X1 _12643_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04890_ ) );
MUX2_X1 _12644_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04891_ ) );
MUX2_X1 _12645_ ( .A(_04890_ ), .B(_04891_ ), .S(fanout_net_38 ), .Z(_04892_ ) );
OAI211_X1 _12646_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04889_ ), .C1(_04892_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04893_ ) );
NAND2_X1 _12647_ ( .A1(_04884_ ), .A2(_04893_ ), .ZN(_04894_ ) );
OAI21_X1 _12648_ ( .A(_04894_ ), .B1(_04253_ ), .B2(_04138_ ), .ZN(_04895_ ) );
AND2_X1 _12649_ ( .A1(_04875_ ), .A2(_04895_ ), .ZN(_04896_ ) );
XNOR2_X1 _12650_ ( .A(_04896_ ), .B(_02579_ ), .ZN(_04897_ ) );
AND2_X2 _12651_ ( .A1(_04874_ ), .A2(_04897_ ), .ZN(_04898_ ) );
INV_X1 _12652_ ( .A(_02626_ ), .ZN(_04899_ ) );
OR3_X1 _12653_ ( .A1(_04394_ ), .A2(\EX_LS_result_reg [6] ), .A3(_04395_ ), .ZN(_04900_ ) );
OR2_X1 _12654_ ( .A1(_04108_ ), .A2(\myreg.Reg[5][6] ), .ZN(_04901_ ) );
OAI211_X1 _12655_ ( .A(_04901_ ), .B(_04112_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[4][6] ), .ZN(_04902_ ) );
OR2_X1 _12656_ ( .A1(_04108_ ), .A2(\myreg.Reg[7][6] ), .ZN(_04903_ ) );
OAI211_X1 _12657_ ( .A(_04903_ ), .B(fanout_net_38 ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[6][6] ), .ZN(_04904_ ) );
NAND3_X1 _12658_ ( .A1(_04902_ ), .A2(_04904_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04905_ ) );
MUX2_X1 _12659_ ( .A(\myreg.Reg[2][6] ), .B(\myreg.Reg[3][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04906_ ) );
MUX2_X1 _12660_ ( .A(\myreg.Reg[0][6] ), .B(\myreg.Reg[1][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04907_ ) );
MUX2_X1 _12661_ ( .A(_04906_ ), .B(_04907_ ), .S(_04123_ ), .Z(_04908_ ) );
OAI211_X1 _12662_ ( .A(_04106_ ), .B(_04905_ ), .C1(_04908_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04909_ ) );
NOR2_X1 _12663_ ( .A1(_04309_ ), .A2(\myreg.Reg[11][6] ), .ZN(_04910_ ) );
OAI21_X1 _12664_ ( .A(fanout_net_38 ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myreg.Reg[10][6] ), .ZN(_04911_ ) );
NOR2_X1 _12665_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[8][6] ), .ZN(_04912_ ) );
OAI21_X1 _12666_ ( .A(_04123_ ), .B1(_04118_ ), .B2(\myreg.Reg[9][6] ), .ZN(_04913_ ) );
OAI221_X1 _12667_ ( .A(_04125_ ), .B1(_04910_ ), .B2(_04911_ ), .C1(_04912_ ), .C2(_04913_ ), .ZN(_04914_ ) );
MUX2_X1 _12668_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04915_ ) );
MUX2_X1 _12669_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04916_ ) );
MUX2_X1 _12670_ ( .A(_04915_ ), .B(_04916_ ), .S(fanout_net_38 ), .Z(_04917_ ) );
OAI211_X1 _12671_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04914_ ), .C1(_04917_ ), .C2(_04126_ ), .ZN(_04918_ ) );
OAI211_X1 _12672_ ( .A(_04909_ ), .B(_04918_ ), .C1(_04394_ ), .C2(_04395_ ), .ZN(_04919_ ) );
NAND2_X2 _12673_ ( .A1(_04900_ ), .A2(_04919_ ), .ZN(_04920_ ) );
XNOR2_X1 _12674_ ( .A(_04899_ ), .B(_04920_ ), .ZN(_04921_ ) );
INV_X1 _12675_ ( .A(_02651_ ), .ZN(_04922_ ) );
INV_X1 _12676_ ( .A(\EX_LS_result_reg [7] ), .ZN(_04923_ ) );
OR3_X1 _12677_ ( .A1(_04100_ ), .A2(_04923_ ), .A3(_04103_ ), .ZN(_04924_ ) );
OR2_X1 _12678_ ( .A1(_04309_ ), .A2(\myreg.Reg[1][7] ), .ZN(_04925_ ) );
OAI211_X1 _12679_ ( .A(_04925_ ), .B(_04218_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[0][7] ), .ZN(_04926_ ) );
OR2_X1 _12680_ ( .A1(_04309_ ), .A2(\myreg.Reg[3][7] ), .ZN(_04927_ ) );
OAI211_X1 _12681_ ( .A(_04927_ ), .B(fanout_net_38 ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[2][7] ), .ZN(_04928_ ) );
NAND3_X1 _12682_ ( .A1(_04926_ ), .A2(_04928_ ), .A3(_04126_ ), .ZN(_04929_ ) );
MUX2_X1 _12683_ ( .A(\myreg.Reg[6][7] ), .B(\myreg.Reg[7][7] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04930_ ) );
MUX2_X1 _12684_ ( .A(\myreg.Reg[4][7] ), .B(\myreg.Reg[5][7] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04931_ ) );
MUX2_X1 _12685_ ( .A(_04930_ ), .B(_04931_ ), .S(_04268_ ), .Z(_04932_ ) );
OAI211_X1 _12686_ ( .A(_04148_ ), .B(_04929_ ), .C1(_04932_ ), .C2(_04265_ ), .ZN(_04933_ ) );
OR2_X1 _12687_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[14][7] ), .ZN(_04934_ ) );
OAI211_X1 _12688_ ( .A(_04934_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04310_ ), .C2(\myreg.Reg[15][7] ), .ZN(_04935_ ) );
OR2_X1 _12689_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[12][7] ), .ZN(_04936_ ) );
OAI211_X1 _12690_ ( .A(_04936_ ), .B(_04218_ ), .C1(_04352_ ), .C2(\myreg.Reg[13][7] ), .ZN(_04937_ ) );
NAND3_X1 _12691_ ( .A1(_04935_ ), .A2(_04937_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04938_ ) );
MUX2_X1 _12692_ ( .A(\myreg.Reg[8][7] ), .B(\myreg.Reg[9][7] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04939_ ) );
MUX2_X1 _12693_ ( .A(\myreg.Reg[10][7] ), .B(\myreg.Reg[11][7] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04940_ ) );
MUX2_X1 _12694_ ( .A(_04939_ ), .B(_04940_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04941_ ) );
OAI211_X1 _12695_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04938_ ), .C1(_04941_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04942_ ) );
NAND2_X1 _12696_ ( .A1(_04933_ ), .A2(_04942_ ), .ZN(_04943_ ) );
OAI21_X1 _12697_ ( .A(_04943_ ), .B1(_04253_ ), .B2(_04173_ ), .ZN(_04944_ ) );
AND2_X1 _12698_ ( .A1(_04924_ ), .A2(_04944_ ), .ZN(_04945_ ) );
XNOR2_X1 _12699_ ( .A(_04922_ ), .B(_04945_ ), .ZN(_04946_ ) );
AND2_X1 _12700_ ( .A1(_04921_ ), .A2(_04946_ ), .ZN(_04947_ ) );
AND2_X1 _12701_ ( .A1(_04898_ ), .A2(_04947_ ), .ZN(_04948_ ) );
AND3_X1 _12702_ ( .A1(_04852_ ), .A2(_04853_ ), .A3(_04948_ ), .ZN(_04949_ ) );
INV_X1 _12703_ ( .A(fanout_net_4 ), .ZN(_04950_ ) );
NOR2_X1 _12704_ ( .A1(_04950_ ), .A2(\ID_EX_typ [1] ), .ZN(_04951_ ) );
AND2_X2 _12705_ ( .A1(_04951_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04952_ ) );
INV_X1 _12706_ ( .A(_04952_ ), .ZN(_04953_ ) );
INV_X1 _12707_ ( .A(fanout_net_6 ), .ZN(_04954_ ) );
BUF_X4 _12708_ ( .A(_04954_ ), .Z(_04955_ ) );
BUF_X4 _12709_ ( .A(_04955_ ), .Z(_04956_ ) );
BUF_X2 _12710_ ( .A(_04956_ ), .Z(_04957_ ) );
OAI21_X1 _12711_ ( .A(_04957_ ), .B1(_04497_ ), .B2(_04498_ ), .ZN(_04958_ ) );
INV_X1 _12712_ ( .A(\ID_EX_imm [31] ), .ZN(_04959_ ) );
NAND2_X1 _12713_ ( .A1(_04959_ ), .A2(fanout_net_6 ), .ZN(_04960_ ) );
NAND2_X1 _12714_ ( .A1(_04958_ ), .A2(_04960_ ), .ZN(_04961_ ) );
NOR2_X1 _12715_ ( .A1(_04961_ ), .A2(_03006_ ), .ZN(_04962_ ) );
INV_X1 _12716_ ( .A(_03006_ ), .ZN(_04963_ ) );
AOI21_X1 _12717_ ( .A(_04963_ ), .B1(_04958_ ), .B2(_04960_ ), .ZN(_04964_ ) );
NOR2_X1 _12718_ ( .A1(_04962_ ), .A2(_04964_ ), .ZN(_04965_ ) );
INV_X1 _12719_ ( .A(_04965_ ), .ZN(_04966_ ) );
NAND3_X1 _12720_ ( .A1(_04448_ ), .A2(_04957_ ), .A3(_04474_ ), .ZN(_04967_ ) );
OR2_X1 _12721_ ( .A1(_04957_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04968_ ) );
NAND2_X1 _12722_ ( .A1(_04967_ ), .A2(_04968_ ), .ZN(_04969_ ) );
XNOR2_X1 _12723_ ( .A(_02178_ ), .B(_04969_ ), .ZN(_04970_ ) );
NOR2_X1 _12724_ ( .A1(_04966_ ), .A2(_04970_ ), .ZN(_04971_ ) );
NAND3_X1 _12725_ ( .A1(_04523_ ), .A2(_04957_ ), .A3(_04543_ ), .ZN(_04972_ ) );
NAND2_X1 _12726_ ( .A1(_02978_ ), .A2(fanout_net_6 ), .ZN(_04973_ ) );
NAND2_X1 _12727_ ( .A1(_04972_ ), .A2(_04973_ ), .ZN(_04974_ ) );
INV_X1 _12728_ ( .A(_02973_ ), .ZN(_04975_ ) );
XNOR2_X1 _12729_ ( .A(_04974_ ), .B(_04975_ ), .ZN(_04976_ ) );
INV_X1 _12730_ ( .A(_04976_ ), .ZN(_04977_ ) );
NAND3_X1 _12731_ ( .A1(_04501_ ), .A2(_04957_ ), .A3(_04520_ ), .ZN(_04978_ ) );
NAND2_X1 _12732_ ( .A1(fanout_net_6 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04979_ ) );
AND2_X2 _12733_ ( .A1(_04978_ ), .A2(_04979_ ), .ZN(_04980_ ) );
INV_X1 _12734_ ( .A(_02209_ ), .ZN(_04981_ ) );
XNOR2_X1 _12735_ ( .A(_04980_ ), .B(_04981_ ), .ZN(_04982_ ) );
INV_X1 _12736_ ( .A(_04982_ ), .ZN(_04983_ ) );
AND3_X1 _12737_ ( .A1(_04971_ ), .A2(_04977_ ), .A3(_04983_ ), .ZN(_04984_ ) );
NAND3_X1 _12738_ ( .A1(_04795_ ), .A2(_04955_ ), .A3(_04793_ ), .ZN(_04985_ ) );
NAND2_X1 _12739_ ( .A1(_02283_ ), .A2(fanout_net_6 ), .ZN(_04986_ ) );
NAND2_X1 _12740_ ( .A1(_04985_ ), .A2(_04986_ ), .ZN(_04987_ ) );
XNOR2_X1 _12741_ ( .A(_04987_ ), .B(_02282_ ), .ZN(_04988_ ) );
NAND3_X1 _12742_ ( .A1(_04751_ ), .A2(_04955_ ), .A3(_04771_ ), .ZN(_04989_ ) );
NAND2_X1 _12743_ ( .A1(_02306_ ), .A2(fanout_net_6 ), .ZN(_04990_ ) );
NAND2_X1 _12744_ ( .A1(_04989_ ), .A2(_04990_ ), .ZN(_04991_ ) );
INV_X1 _12745_ ( .A(_04991_ ), .ZN(_04992_ ) );
NOR3_X1 _12746_ ( .A1(_04988_ ), .A2(_04749_ ), .A3(_04992_ ), .ZN(_04993_ ) );
XNOR2_X1 _12747_ ( .A(_04991_ ), .B(_02305_ ), .ZN(_04994_ ) );
NOR2_X1 _12748_ ( .A1(_04988_ ), .A2(_04994_ ), .ZN(_04995_ ) );
AOI21_X1 _12749_ ( .A(fanout_net_6 ), .B1(_04843_ ), .B2(_04844_ ), .ZN(_04996_ ) );
AND2_X1 _12750_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [21] ), .ZN(_04997_ ) );
NOR2_X1 _12751_ ( .A1(_04996_ ), .A2(_04997_ ), .ZN(_04998_ ) );
XNOR2_X1 _12752_ ( .A(_04998_ ), .B(_04823_ ), .ZN(_04999_ ) );
INV_X1 _12753_ ( .A(_04999_ ), .ZN(_05000_ ) );
NAND3_X1 _12754_ ( .A1(_04819_ ), .A2(_04956_ ), .A3(_04820_ ), .ZN(_05001_ ) );
NAND2_X1 _12755_ ( .A1(_02330_ ), .A2(fanout_net_6 ), .ZN(_05002_ ) );
NAND2_X1 _12756_ ( .A1(_05001_ ), .A2(_05002_ ), .ZN(_05003_ ) );
XNOR2_X1 _12757_ ( .A(_05003_ ), .B(_02329_ ), .ZN(_05004_ ) );
INV_X1 _12758_ ( .A(_05004_ ), .ZN(_05005_ ) );
AND3_X1 _12759_ ( .A1(_04995_ ), .A2(_05000_ ), .A3(_05005_ ), .ZN(_05006_ ) );
AOI21_X1 _12760_ ( .A(fanout_net_6 ), .B1(_04653_ ), .B2(_04673_ ), .ZN(_05007_ ) );
AND2_X1 _12761_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [19] ), .ZN(_05008_ ) );
NOR2_X1 _12762_ ( .A1(_05007_ ), .A2(_05008_ ), .ZN(_05009_ ) );
XNOR2_X1 _12763_ ( .A(_05009_ ), .B(_02382_ ), .ZN(_05010_ ) );
NAND3_X1 _12764_ ( .A1(_04695_ ), .A2(_04956_ ), .A3(_04696_ ), .ZN(_05011_ ) );
NAND2_X1 _12765_ ( .A1(_02406_ ), .A2(fanout_net_6 ), .ZN(_05012_ ) );
NAND2_X1 _12766_ ( .A1(_05011_ ), .A2(_05012_ ), .ZN(_05013_ ) );
XNOR2_X1 _12767_ ( .A(_05013_ ), .B(_02405_ ), .ZN(_05014_ ) );
NOR2_X1 _12768_ ( .A1(_05010_ ), .A2(_05014_ ), .ZN(_05015_ ) );
NAND3_X1 _12769_ ( .A1(_04725_ ), .A2(_04955_ ), .A3(_04745_ ), .ZN(_05016_ ) );
NAND2_X1 _12770_ ( .A1(_02431_ ), .A2(fanout_net_6 ), .ZN(_05017_ ) );
NAND2_X1 _12771_ ( .A1(_05016_ ), .A2(_05017_ ), .ZN(_05018_ ) );
XNOR2_X1 _12772_ ( .A(_05018_ ), .B(_04723_ ), .ZN(_05019_ ) );
NAND3_X1 _12773_ ( .A1(_04719_ ), .A2(_04956_ ), .A3(_04720_ ), .ZN(_05020_ ) );
NAND2_X1 _12774_ ( .A1(_02455_ ), .A2(fanout_net_6 ), .ZN(_05021_ ) );
NAND2_X1 _12775_ ( .A1(_05020_ ), .A2(_05021_ ), .ZN(_05022_ ) );
AND3_X1 _12776_ ( .A1(_05019_ ), .A2(_02453_ ), .A3(_05022_ ), .ZN(_05023_ ) );
AOI22_X1 _12777_ ( .A1(_05016_ ), .A2(_05017_ ), .B1(_02429_ ), .B2(_02409_ ), .ZN(_05024_ ) );
OAI21_X1 _12778_ ( .A(_05015_ ), .B1(_05023_ ), .B2(_05024_ ), .ZN(_05025_ ) );
NAND2_X1 _12779_ ( .A1(_05009_ ), .A2(_02382_ ), .ZN(_05026_ ) );
NAND2_X1 _12780_ ( .A1(_05025_ ), .A2(_05026_ ), .ZN(_05027_ ) );
INV_X1 _12781_ ( .A(_05010_ ), .ZN(_05028_ ) );
AND3_X1 _12782_ ( .A1(_05028_ ), .A2(_02405_ ), .A3(_05013_ ), .ZN(_05029_ ) );
OAI21_X1 _12783_ ( .A(_05006_ ), .B1(_05027_ ), .B2(_05029_ ), .ZN(_05030_ ) );
AND3_X1 _12784_ ( .A1(_05000_ ), .A2(_02329_ ), .A3(_05003_ ), .ZN(_05031_ ) );
INV_X1 _12785_ ( .A(_04823_ ), .ZN(_05032_ ) );
NOR3_X1 _12786_ ( .A1(_05032_ ), .A2(_04997_ ), .A3(_04996_ ), .ZN(_05033_ ) );
OAI21_X1 _12787_ ( .A(_04995_ ), .B1(_05031_ ), .B2(_05033_ ), .ZN(_05034_ ) );
INV_X1 _12788_ ( .A(_02282_ ), .ZN(_05035_ ) );
INV_X1 _12789_ ( .A(_04987_ ), .ZN(_05036_ ) );
OAI211_X1 _12790_ ( .A(_05030_ ), .B(_05034_ ), .C1(_05035_ ), .C2(_05036_ ), .ZN(_05037_ ) );
INV_X1 _12791_ ( .A(_02731_ ), .ZN(_05038_ ) );
NAND3_X1 _12792_ ( .A1(_04331_ ), .A2(_04956_ ), .A3(_04332_ ), .ZN(_05039_ ) );
NAND2_X1 _12793_ ( .A1(_02732_ ), .A2(fanout_net_6 ), .ZN(_05040_ ) );
AOI21_X1 _12794_ ( .A(fanout_net_6 ), .B1(_04286_ ), .B2(_04306_ ), .ZN(_05041_ ) );
AND2_X1 _12795_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [13] ), .ZN(_05042_ ) );
NOR2_X1 _12796_ ( .A1(_05041_ ), .A2(_05042_ ), .ZN(_05043_ ) );
AND2_X1 _12797_ ( .A1(_05043_ ), .A2(_04284_ ), .ZN(_05044_ ) );
INV_X1 _12798_ ( .A(_05044_ ), .ZN(_05045_ ) );
NOR2_X1 _12799_ ( .A1(_05043_ ), .A2(_04284_ ), .ZN(_05046_ ) );
INV_X1 _12800_ ( .A(_05046_ ), .ZN(_05047_ ) );
AOI221_X4 _12801_ ( .A(_05038_ ), .B1(_05039_ ), .B2(_05040_ ), .C1(_05045_ ), .C2(_05047_ ), .ZN(_05048_ ) );
AOI21_X1 _12802_ ( .A(_05048_ ), .B1(_04283_ ), .B2(_05043_ ), .ZN(_05049_ ) );
NAND3_X1 _12803_ ( .A1(_04233_ ), .A2(_04955_ ), .A3(_04254_ ), .ZN(_05050_ ) );
NAND2_X1 _12804_ ( .A1(_02684_ ), .A2(fanout_net_6 ), .ZN(_05051_ ) );
NAND2_X1 _12805_ ( .A1(_05050_ ), .A2(_05051_ ), .ZN(_05052_ ) );
XNOR2_X1 _12806_ ( .A(_05052_ ), .B(_02683_ ), .ZN(_05053_ ) );
NAND3_X1 _12807_ ( .A1(_04278_ ), .A2(_04955_ ), .A3(_04279_ ), .ZN(_05054_ ) );
NAND2_X1 _12808_ ( .A1(_02708_ ), .A2(fanout_net_6 ), .ZN(_05055_ ) );
NAND2_X1 _12809_ ( .A1(_05054_ ), .A2(_05055_ ), .ZN(_05056_ ) );
XNOR2_X1 _12810_ ( .A(_05056_ ), .B(_02706_ ), .ZN(_05057_ ) );
NOR3_X1 _12811_ ( .A1(_05049_ ), .A2(_05053_ ), .A3(_05057_ ), .ZN(_05058_ ) );
XNOR2_X1 _12812_ ( .A(_05043_ ), .B(_04283_ ), .ZN(_05059_ ) );
NOR3_X1 _12813_ ( .A1(_05059_ ), .A2(_05053_ ), .A3(_05057_ ), .ZN(_05060_ ) );
NAND2_X1 _12814_ ( .A1(_05039_ ), .A2(_05040_ ), .ZN(_05061_ ) );
XNOR2_X1 _12815_ ( .A(_05061_ ), .B(_02731_ ), .ZN(_05062_ ) );
INV_X1 _12816_ ( .A(_05062_ ), .ZN(_05063_ ) );
NAND2_X1 _12817_ ( .A1(_05060_ ), .A2(_05063_ ), .ZN(_05064_ ) );
NAND3_X1 _12818_ ( .A1(_04226_ ), .A2(_04954_ ), .A3(_04227_ ), .ZN(_05065_ ) );
NAND2_X1 _12819_ ( .A1(_02829_ ), .A2(fanout_net_6 ), .ZN(_05066_ ) );
NAND2_X1 _12820_ ( .A1(_05065_ ), .A2(_05066_ ), .ZN(_05067_ ) );
XNOR2_X1 _12821_ ( .A(_05067_ ), .B(_02828_ ), .ZN(_05068_ ) );
NAND3_X1 _12822_ ( .A1(_04197_ ), .A2(_04954_ ), .A3(_04202_ ), .ZN(_05069_ ) );
NAND2_X1 _12823_ ( .A1(_02852_ ), .A2(fanout_net_6 ), .ZN(_05070_ ) );
NAND2_X1 _12824_ ( .A1(_05069_ ), .A2(_05070_ ), .ZN(_05071_ ) );
XNOR2_X1 _12825_ ( .A(_05071_ ), .B(_02851_ ), .ZN(_05072_ ) );
OR2_X1 _12826_ ( .A1(_05068_ ), .A2(_05072_ ), .ZN(_05073_ ) );
AOI21_X1 _12827_ ( .A(fanout_net_6 ), .B1(_04104_ ), .B2(_04139_ ), .ZN(_05074_ ) );
AND2_X1 _12828_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [9] ), .ZN(_05075_ ) );
NOR2_X1 _12829_ ( .A1(_05074_ ), .A2(_05075_ ), .ZN(_05076_ ) );
NAND2_X1 _12830_ ( .A1(_05076_ ), .A2(_02802_ ), .ZN(_05077_ ) );
NAND3_X1 _12831_ ( .A1(_04147_ ), .A2(_04956_ ), .A3(_04174_ ), .ZN(_05078_ ) );
NAND2_X1 _12832_ ( .A1(_02781_ ), .A2(fanout_net_6 ), .ZN(_05079_ ) );
NAND2_X1 _12833_ ( .A1(_05078_ ), .A2(_05079_ ), .ZN(_05080_ ) );
INV_X1 _12834_ ( .A(_02802_ ), .ZN(_05081_ ) );
AND2_X1 _12835_ ( .A1(_05076_ ), .A2(_05081_ ), .ZN(_05082_ ) );
NOR2_X1 _12836_ ( .A1(_05076_ ), .A2(_05081_ ), .ZN(_05083_ ) );
OAI211_X1 _12837_ ( .A(_02780_ ), .B(_05080_ ), .C1(_05082_ ), .C2(_05083_ ), .ZN(_05084_ ) );
AOI21_X1 _12838_ ( .A(_05073_ ), .B1(_05077_ ), .B2(_05084_ ), .ZN(_05085_ ) );
AOI21_X1 _12839_ ( .A(_05085_ ), .B1(_02851_ ), .B2(_05071_ ), .ZN(_05086_ ) );
INV_X1 _12840_ ( .A(_05072_ ), .ZN(_05087_ ) );
NAND3_X1 _12841_ ( .A1(_05087_ ), .A2(_02828_ ), .A3(_05067_ ), .ZN(_05088_ ) );
AOI21_X1 _12842_ ( .A(_05064_ ), .B1(_05086_ ), .B2(_05088_ ), .ZN(_05089_ ) );
AOI211_X1 _12843_ ( .A(_05058_ ), .B(_05089_ ), .C1(_02683_ ), .C2(_05052_ ), .ZN(_05090_ ) );
XNOR2_X1 _12844_ ( .A(_05076_ ), .B(_02802_ ), .ZN(_05091_ ) );
XNOR2_X1 _12845_ ( .A(_05080_ ), .B(_02780_ ), .ZN(_05092_ ) );
NOR4_X1 _12846_ ( .A1(_05064_ ), .A2(_05091_ ), .A3(_05073_ ), .A4(_05092_ ), .ZN(_05093_ ) );
NAND3_X1 _12847_ ( .A1(_04924_ ), .A2(_04956_ ), .A3(_04944_ ), .ZN(_05094_ ) );
NAND2_X1 _12848_ ( .A1(_02630_ ), .A2(fanout_net_6 ), .ZN(_05095_ ) );
NAND2_X1 _12849_ ( .A1(_05094_ ), .A2(_05095_ ), .ZN(_05096_ ) );
XNOR2_X1 _12850_ ( .A(_05096_ ), .B(_02651_ ), .ZN(_05097_ ) );
NAND2_X1 _12851_ ( .A1(_04873_ ), .A2(_04955_ ), .ZN(_05098_ ) );
NAND2_X1 _12852_ ( .A1(_02604_ ), .A2(fanout_net_6 ), .ZN(_05099_ ) );
NAND2_X2 _12853_ ( .A1(_05098_ ), .A2(_05099_ ), .ZN(_05100_ ) );
XNOR2_X1 _12854_ ( .A(_05100_ ), .B(_02603_ ), .ZN(_05101_ ) );
NAND2_X1 _12855_ ( .A1(_04920_ ), .A2(_04955_ ), .ZN(_05102_ ) );
NAND2_X1 _12856_ ( .A1(_02627_ ), .A2(fanout_net_6 ), .ZN(_05103_ ) );
NAND2_X2 _12857_ ( .A1(_05102_ ), .A2(_05103_ ), .ZN(_05104_ ) );
XNOR2_X1 _12858_ ( .A(_05104_ ), .B(_02626_ ), .ZN(_05105_ ) );
NAND3_X1 _12859_ ( .A1(_04875_ ), .A2(_04955_ ), .A3(_04895_ ), .ZN(_05106_ ) );
OR2_X1 _12860_ ( .A1(_04954_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05107_ ) );
NAND2_X1 _12861_ ( .A1(_05106_ ), .A2(_05107_ ), .ZN(_05108_ ) );
INV_X4 _12862_ ( .A(_02579_ ), .ZN(_05109_ ) );
XNOR2_X1 _12863_ ( .A(_05108_ ), .B(_05109_ ), .ZN(_05110_ ) );
OR4_X2 _12864_ ( .A1(_05097_ ), .A2(_05101_ ), .A3(_05105_ ), .A4(_05110_ ), .ZN(_05111_ ) );
NAND3_X1 _12865_ ( .A1(_04422_ ), .A2(_04956_ ), .A3(_04442_ ), .ZN(_05112_ ) );
NAND2_X1 _12866_ ( .A1(fanout_net_6 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_05113_ ) );
AND2_X2 _12867_ ( .A1(_05112_ ), .A2(_05113_ ), .ZN(_05114_ ) );
XNOR2_X1 _12868_ ( .A(_05114_ ), .B(_02555_ ), .ZN(_05115_ ) );
NAND2_X1 _12869_ ( .A1(_04419_ ), .A2(_04956_ ), .ZN(_05116_ ) );
INV_X1 _12870_ ( .A(\ID_EX_imm [2] ), .ZN(_05117_ ) );
NAND2_X1 _12871_ ( .A1(_05117_ ), .A2(fanout_net_6 ), .ZN(_05118_ ) );
NAND2_X2 _12872_ ( .A1(_05116_ ), .A2(_05118_ ), .ZN(_05119_ ) );
INV_X1 _12873_ ( .A(_05119_ ), .ZN(_05120_ ) );
NOR3_X1 _12874_ ( .A1(_05115_ ), .A2(_04390_ ), .A3(_05120_ ), .ZN(_05121_ ) );
INV_X1 _12875_ ( .A(_05114_ ), .ZN(_05122_ ) );
AOI21_X1 _12876_ ( .A(_05121_ ), .B1(_02527_ ), .B2(_05122_ ), .ZN(_05123_ ) );
XNOR2_X1 _12877_ ( .A(_05119_ ), .B(_02549_ ), .ZN(_05124_ ) );
INV_X1 _12878_ ( .A(_05124_ ), .ZN(_05125_ ) );
NAND3_X1 _12879_ ( .A1(_04341_ ), .A2(_04955_ ), .A3(_04362_ ), .ZN(_05126_ ) );
INV_X1 _12880_ ( .A(\ID_EX_imm [1] ), .ZN(_05127_ ) );
NAND2_X1 _12881_ ( .A1(_05127_ ), .A2(fanout_net_6 ), .ZN(_05128_ ) );
NAND2_X1 _12882_ ( .A1(_05126_ ), .A2(_05128_ ), .ZN(_05129_ ) );
NAND2_X1 _12883_ ( .A1(_05129_ ), .A2(_02478_ ), .ZN(_05130_ ) );
AND3_X1 _12884_ ( .A1(_05126_ ), .A2(_02478_ ), .A3(_05128_ ), .ZN(_05131_ ) );
AOI21_X1 _12885_ ( .A(_02478_ ), .B1(_05126_ ), .B2(_05128_ ), .ZN(_05132_ ) );
NOR2_X1 _12886_ ( .A1(_05131_ ), .A2(_05132_ ), .ZN(_05133_ ) );
NAND3_X1 _12887_ ( .A1(_04384_ ), .A2(_04954_ ), .A3(_04385_ ), .ZN(_05134_ ) );
NAND2_X1 _12888_ ( .A1(_02480_ ), .A2(\ID_EX_typ [4] ), .ZN(_05135_ ) );
NAND2_X2 _12889_ ( .A1(_05134_ ), .A2(_05135_ ), .ZN(_05136_ ) );
NOR2_X1 _12890_ ( .A1(_05136_ ), .A2(_02502_ ), .ZN(_05137_ ) );
OAI21_X1 _12891_ ( .A(_05130_ ), .B1(_05133_ ), .B2(_05137_ ), .ZN(_05138_ ) );
AND2_X1 _12892_ ( .A1(_05114_ ), .A2(_02527_ ), .ZN(_05139_ ) );
NOR2_X1 _12893_ ( .A1(_05114_ ), .A2(_02527_ ), .ZN(_05140_ ) );
OAI211_X1 _12894_ ( .A(_05125_ ), .B(_05138_ ), .C1(_05139_ ), .C2(_05140_ ), .ZN(_05141_ ) );
AOI21_X2 _12895_ ( .A(_05111_ ), .B1(_05123_ ), .B2(_05141_ ), .ZN(_05142_ ) );
INV_X1 _12896_ ( .A(_05105_ ), .ZN(_05143_ ) );
INV_X1 _12897_ ( .A(_05097_ ), .ZN(_05144_ ) );
AND3_X1 _12898_ ( .A1(_05106_ ), .A2(_02579_ ), .A3(_05107_ ), .ZN(_05145_ ) );
INV_X1 _12899_ ( .A(_05100_ ), .ZN(_05146_ ) );
NOR3_X1 _12900_ ( .A1(_05110_ ), .A2(_05146_ ), .A3(_02656_ ), .ZN(_05147_ ) );
OAI211_X1 _12901_ ( .A(_05143_ ), .B(_05144_ ), .C1(_05145_ ), .C2(_05147_ ), .ZN(_05148_ ) );
NAND2_X1 _12902_ ( .A1(_05096_ ), .A2(_02651_ ), .ZN(_05149_ ) );
NAND3_X1 _12903_ ( .A1(_05144_ ), .A2(_02626_ ), .A3(_05104_ ), .ZN(_05150_ ) );
NAND3_X1 _12904_ ( .A1(_05148_ ), .A2(_05149_ ), .A3(_05150_ ), .ZN(_05151_ ) );
OAI21_X1 _12905_ ( .A(_05093_ ), .B1(_05142_ ), .B2(_05151_ ), .ZN(_05152_ ) );
NAND2_X1 _12906_ ( .A1(_05056_ ), .A2(_02707_ ), .ZN(_05153_ ) );
OR2_X1 _12907_ ( .A1(_05053_ ), .A2(_05153_ ), .ZN(_05154_ ) );
NAND3_X1 _12908_ ( .A1(_05090_ ), .A2(_05152_ ), .A3(_05154_ ), .ZN(_05155_ ) );
AND4_X1 _12909_ ( .A1(_05000_ ), .A2(_05015_ ), .A3(_05005_ ), .A4(_04995_ ), .ZN(_05156_ ) );
XNOR2_X1 _12910_ ( .A(_05022_ ), .B(_02454_ ), .ZN(_05157_ ) );
INV_X1 _12911_ ( .A(_05157_ ), .ZN(_05158_ ) );
AND3_X1 _12912_ ( .A1(_05156_ ), .A2(_05019_ ), .A3(_05158_ ), .ZN(_05159_ ) );
AOI211_X1 _12913_ ( .A(_04993_ ), .B(_05037_ ), .C1(_05155_ ), .C2(_05159_ ), .ZN(_05160_ ) );
NAND3_X1 _12914_ ( .A1(_04568_ ), .A2(_04956_ ), .A3(_04570_ ), .ZN(_05161_ ) );
NAND2_X1 _12915_ ( .A1(_02257_ ), .A2(\ID_EX_typ [4] ), .ZN(_05162_ ) );
NAND2_X1 _12916_ ( .A1(_05161_ ), .A2(_05162_ ), .ZN(_05163_ ) );
INV_X1 _12917_ ( .A(_02256_ ), .ZN(_05164_ ) );
NOR2_X1 _12918_ ( .A1(_05163_ ), .A2(_05164_ ), .ZN(_05165_ ) );
AOI21_X1 _12919_ ( .A(_02256_ ), .B1(_05161_ ), .B2(_05162_ ), .ZN(_05166_ ) );
NOR2_X1 _12920_ ( .A1(_05165_ ), .A2(_05166_ ), .ZN(_05167_ ) );
NAND2_X1 _12921_ ( .A1(_04595_ ), .A2(_04957_ ), .ZN(_05168_ ) );
NAND2_X1 _12922_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [27] ), .ZN(_05169_ ) );
AND2_X1 _12923_ ( .A1(_05168_ ), .A2(_05169_ ), .ZN(_05170_ ) );
NOR2_X1 _12924_ ( .A1(_05170_ ), .A2(_04597_ ), .ZN(_05171_ ) );
INV_X1 _12925_ ( .A(_05171_ ), .ZN(_05172_ ) );
AND3_X1 _12926_ ( .A1(_05168_ ), .A2(_04597_ ), .A3(_05169_ ), .ZN(_05173_ ) );
INV_X1 _12927_ ( .A(_05173_ ), .ZN(_05174_ ) );
AOI21_X1 _12928_ ( .A(_05167_ ), .B1(_05172_ ), .B2(_05174_ ), .ZN(_05175_ ) );
INV_X1 _12929_ ( .A(_05175_ ), .ZN(_05176_ ) );
NAND3_X1 _12930_ ( .A1(_04618_ ), .A2(_04957_ ), .A3(_04620_ ), .ZN(_05177_ ) );
NAND2_X1 _12931_ ( .A1(_02916_ ), .A2(\ID_EX_typ [4] ), .ZN(_05178_ ) );
NAND2_X1 _12932_ ( .A1(_05177_ ), .A2(_05178_ ), .ZN(_05179_ ) );
NOR2_X1 _12933_ ( .A1(_05179_ ), .A2(_04622_ ), .ZN(_05180_ ) );
AOI21_X1 _12934_ ( .A(_02915_ ), .B1(_05177_ ), .B2(_05178_ ), .ZN(_05181_ ) );
NOR2_X1 _12935_ ( .A1(_05180_ ), .A2(_05181_ ), .ZN(_05182_ ) );
NAND3_X1 _12936_ ( .A1(_04642_ ), .A2(_04957_ ), .A3(_04644_ ), .ZN(_05183_ ) );
NAND2_X1 _12937_ ( .A1(_02939_ ), .A2(\ID_EX_typ [4] ), .ZN(_05184_ ) );
NAND2_X1 _12938_ ( .A1(_05183_ ), .A2(_05184_ ), .ZN(_05185_ ) );
NOR2_X1 _12939_ ( .A1(_05185_ ), .A2(_02946_ ), .ZN(_05186_ ) );
AOI21_X1 _12940_ ( .A(_02938_ ), .B1(_05183_ ), .B2(_05184_ ), .ZN(_05187_ ) );
NOR2_X1 _12941_ ( .A1(_05186_ ), .A2(_05187_ ), .ZN(_05188_ ) );
NOR4_X2 _12942_ ( .A1(_05160_ ), .A2(_05176_ ), .A3(_05182_ ), .A4(_05188_ ), .ZN(_05189_ ) );
NAND2_X1 _12943_ ( .A1(_05185_ ), .A2(_02938_ ), .ZN(_05190_ ) );
OAI211_X1 _12944_ ( .A(_02915_ ), .B(_05179_ ), .C1(_05186_ ), .C2(_05187_ ), .ZN(_05191_ ) );
AOI21_X1 _12945_ ( .A(_05176_ ), .B1(_05190_ ), .B2(_05191_ ), .ZN(_05192_ ) );
NAND2_X1 _12946_ ( .A1(_05163_ ), .A2(_02256_ ), .ZN(_05193_ ) );
AOI21_X1 _12947_ ( .A(_05193_ ), .B1(_05172_ ), .B2(_05174_ ), .ZN(_05194_ ) );
AND3_X1 _12948_ ( .A1(_05168_ ), .A2(_04596_ ), .A3(_05169_ ), .ZN(_05195_ ) );
OR3_X1 _12949_ ( .A1(_05192_ ), .A2(_05194_ ), .A3(_05195_ ), .ZN(_05196_ ) );
OAI21_X2 _12950_ ( .A(_04984_ ), .B1(_05189_ ), .B2(_05196_ ), .ZN(_05197_ ) );
AOI21_X1 _12951_ ( .A(_04969_ ), .B1(_02173_ ), .B2(_02177_ ), .ZN(_05198_ ) );
AND2_X1 _12952_ ( .A1(_04965_ ), .A2(_05198_ ), .ZN(_05199_ ) );
OR3_X1 _12953_ ( .A1(_04976_ ), .A2(_04981_ ), .A3(_04980_ ), .ZN(_05200_ ) );
OAI21_X1 _12954_ ( .A(_05200_ ), .B1(_04975_ ), .B2(_04974_ ), .ZN(_05201_ ) );
AOI211_X1 _12955_ ( .A(_04962_ ), .B(_05199_ ), .C1(_05201_ ), .C2(_04971_ ), .ZN(_05202_ ) );
AND2_X1 _12956_ ( .A1(_05197_ ), .A2(_05202_ ), .ZN(_05203_ ) );
AND3_X2 _12957_ ( .A1(_05203_ ), .A2(fanout_net_5 ), .A3(_04089_ ), .ZN(_05204_ ) );
AND2_X1 _12958_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_4 ), .ZN(_05205_ ) );
AND2_X1 _12959_ ( .A1(_05205_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05206_ ) );
INV_X1 _12960_ ( .A(_05206_ ), .ZN(_05207_ ) );
AND2_X1 _12961_ ( .A1(_02707_ ), .A2(_04280_ ), .ZN(_05208_ ) );
AND2_X1 _12962_ ( .A1(_04256_ ), .A2(_05208_ ), .ZN(_05209_ ) );
NOR2_X1 _12963_ ( .A1(_04307_ ), .A2(_04283_ ), .ZN(_05210_ ) );
AND2_X1 _12964_ ( .A1(_04307_ ), .A2(_04283_ ), .ZN(_05211_ ) );
INV_X1 _12965_ ( .A(_05211_ ), .ZN(_05212_ ) );
NAND2_X1 _12966_ ( .A1(_02731_ ), .A2(_04333_ ), .ZN(_05213_ ) );
AOI21_X1 _12967_ ( .A(_05210_ ), .B1(_05212_ ), .B2(_05213_ ), .ZN(_05214_ ) );
NAND3_X1 _12968_ ( .A1(_05214_ ), .A2(_04256_ ), .A3(_04281_ ), .ZN(_05215_ ) );
AND2_X1 _12969_ ( .A1(_04175_ ), .A2(_02780_ ), .ZN(_05216_ ) );
NAND2_X1 _12970_ ( .A1(_04143_ ), .A2(_05216_ ), .ZN(_05217_ ) );
INV_X1 _12971_ ( .A(_04141_ ), .ZN(_05218_ ) );
NAND2_X1 _12972_ ( .A1(_05217_ ), .A2(_05218_ ), .ZN(_05219_ ) );
AND3_X1 _12973_ ( .A1(_05219_ ), .A2(_04204_ ), .A3(_04229_ ), .ZN(_05220_ ) );
AND2_X1 _12974_ ( .A1(_02851_ ), .A2(_04203_ ), .ZN(_05221_ ) );
AND3_X1 _12975_ ( .A1(_04204_ ), .A2(_02828_ ), .A3(_04228_ ), .ZN(_05222_ ) );
NOR3_X1 _12976_ ( .A1(_05220_ ), .A2(_05221_ ), .A3(_05222_ ), .ZN(_05223_ ) );
INV_X1 _12977_ ( .A(_04336_ ), .ZN(_05224_ ) );
OAI21_X1 _12978_ ( .A(_05215_ ), .B1(_05223_ ), .B2(_05224_ ), .ZN(_05225_ ) );
AOI211_X1 _12979_ ( .A(_05209_ ), .B(_05225_ ), .C1(_02683_ ), .C2(_04255_ ), .ZN(_05226_ ) );
AND2_X1 _12980_ ( .A1(_04419_ ), .A2(_02549_ ), .ZN(_05227_ ) );
INV_X1 _12981_ ( .A(_05227_ ), .ZN(_05228_ ) );
NAND3_X1 _12982_ ( .A1(_02478_ ), .A2(_04362_ ), .A3(_04341_ ), .ZN(_05229_ ) );
AND2_X1 _12983_ ( .A1(_04389_ ), .A2(_05229_ ), .ZN(_05230_ ) );
OAI221_X1 _12984_ ( .A(_05228_ ), .B1(_02555_ ), .B2(_04443_ ), .C1(_05230_ ), .C2(_04421_ ), .ZN(_05231_ ) );
NAND2_X1 _12985_ ( .A1(_02555_ ), .A2(_04443_ ), .ZN(_05232_ ) );
NAND3_X1 _12986_ ( .A1(_05231_ ), .A2(_05232_ ), .A3(_04948_ ), .ZN(_05233_ ) );
AND3_X1 _12987_ ( .A1(_04946_ ), .A2(_02626_ ), .A3(_04920_ ), .ZN(_05234_ ) );
AND2_X1 _12988_ ( .A1(_04873_ ), .A2(_02603_ ), .ZN(_05235_ ) );
NAND2_X1 _12989_ ( .A1(_04897_ ), .A2(_05235_ ), .ZN(_05236_ ) );
OAI21_X1 _12990_ ( .A(_05236_ ), .B1(_05109_ ), .B2(_04896_ ), .ZN(_05237_ ) );
AOI221_X4 _12991_ ( .A(_05234_ ), .B1(_02651_ ), .B2(_04945_ ), .C1(_04947_ ), .C2(_05237_ ), .ZN(_05238_ ) );
AND2_X1 _12992_ ( .A1(_05233_ ), .A2(_05238_ ), .ZN(_05239_ ) );
OR2_X2 _12993_ ( .A1(_05239_ ), .A2(_04338_ ), .ZN(_05240_ ) );
AND2_X1 _12994_ ( .A1(_05226_ ), .A2(_05240_ ), .ZN(_05241_ ) );
INV_X1 _12995_ ( .A(_04851_ ), .ZN(_05242_ ) );
OR2_X4 _12996_ ( .A1(_05241_ ), .A2(_05242_ ), .ZN(_05243_ ) );
NAND2_X1 _12997_ ( .A1(_02329_ ), .A2(_04821_ ), .ZN(_05244_ ) );
NOR3_X1 _12998_ ( .A1(_04846_ ), .A2(_04847_ ), .A3(_05244_ ), .ZN(_05245_ ) );
OR2_X1 _12999_ ( .A1(_05245_ ), .A2(_04846_ ), .ZN(_05246_ ) );
NAND2_X1 _13000_ ( .A1(_05246_ ), .A2(_04799_ ), .ZN(_05247_ ) );
NOR2_X1 _13001_ ( .A1(_04746_ ), .A2(_02430_ ), .ZN(_05248_ ) );
AND2_X1 _13002_ ( .A1(_04746_ ), .A2(_02430_ ), .ZN(_05249_ ) );
INV_X1 _13003_ ( .A(_05249_ ), .ZN(_05250_ ) );
NAND2_X1 _13004_ ( .A1(_02454_ ), .A2(_04721_ ), .ZN(_05251_ ) );
AOI21_X1 _13005_ ( .A(_05248_ ), .B1(_05250_ ), .B2(_05251_ ), .ZN(_05252_ ) );
AND3_X1 _13006_ ( .A1(_05252_ ), .A2(_04675_ ), .A3(_04698_ ), .ZN(_05253_ ) );
AND3_X1 _13007_ ( .A1(_02382_ ), .A2(_04673_ ), .A3(_04653_ ), .ZN(_05254_ ) );
AND3_X1 _13008_ ( .A1(_04675_ ), .A2(_02405_ ), .A3(_04697_ ), .ZN(_05255_ ) );
NOR3_X1 _13009_ ( .A1(_05253_ ), .A2(_05254_ ), .A3(_05255_ ), .ZN(_05256_ ) );
INV_X1 _13010_ ( .A(_04849_ ), .ZN(_05257_ ) );
OAI21_X1 _13011_ ( .A(_05247_ ), .B1(_05256_ ), .B2(_05257_ ), .ZN(_05258_ ) );
NAND2_X1 _13012_ ( .A1(_04772_ ), .A2(_02305_ ), .ZN(_05259_ ) );
NOR3_X1 _13013_ ( .A1(_04796_ ), .A2(_04797_ ), .A3(_05259_ ), .ZN(_05260_ ) );
NOR3_X1 _13014_ ( .A1(_05258_ ), .A2(_04796_ ), .A3(_05260_ ), .ZN(_05261_ ) );
INV_X1 _13015_ ( .A(_04650_ ), .ZN(_05262_ ) );
NOR2_X1 _13016_ ( .A1(_05261_ ), .A2(_05262_ ), .ZN(_05263_ ) );
INV_X1 _13017_ ( .A(_04477_ ), .ZN(_05264_ ) );
INV_X1 _13018_ ( .A(_04500_ ), .ZN(_05265_ ) );
NOR2_X1 _13019_ ( .A1(_04975_ ), .A2(_04544_ ), .ZN(_05266_ ) );
NOR2_X1 _13020_ ( .A1(_04981_ ), .A2(_04521_ ), .ZN(_05267_ ) );
AOI21_X1 _13021_ ( .A(_05266_ ), .B1(_04545_ ), .B2(_05267_ ), .ZN(_05268_ ) );
NOR3_X1 _13022_ ( .A1(_05264_ ), .A2(_05265_ ), .A3(_05268_ ), .ZN(_05269_ ) );
NOR2_X1 _13023_ ( .A1(_02178_ ), .A2(_04475_ ), .ZN(_05270_ ) );
NAND2_X1 _13024_ ( .A1(_05270_ ), .A2(_04500_ ), .ZN(_05271_ ) );
OR3_X1 _13025_ ( .A1(_04598_ ), .A2(_05164_ ), .A3(_04571_ ), .ZN(_05272_ ) );
OAI21_X1 _13026_ ( .A(_05272_ ), .B1(_04597_ ), .B2(_04595_ ), .ZN(_05273_ ) );
NAND4_X1 _13027_ ( .A1(_04646_ ), .A2(_02915_ ), .A3(_04647_ ), .A4(_04621_ ), .ZN(_05274_ ) );
NAND2_X1 _13028_ ( .A1(_05274_ ), .A2(_04647_ ), .ZN(_05275_ ) );
AOI21_X1 _13029_ ( .A(_05273_ ), .B1(_04599_ ), .B2(_05275_ ), .ZN(_05276_ ) );
INV_X1 _13030_ ( .A(_04547_ ), .ZN(_05277_ ) );
OAI221_X1 _13031_ ( .A(_05271_ ), .B1(_04963_ ), .B2(_04499_ ), .C1(_05276_ ), .C2(_05277_ ), .ZN(_05278_ ) );
NOR3_X1 _13032_ ( .A1(_05263_ ), .A2(_05269_ ), .A3(_05278_ ), .ZN(_05279_ ) );
AOI21_X1 _13033_ ( .A(_05207_ ), .B1(_05243_ ), .B2(_05279_ ), .ZN(_05280_ ) );
AND2_X1 _13034_ ( .A1(_04951_ ), .A2(fanout_net_5 ), .ZN(_05281_ ) );
AND3_X1 _13035_ ( .A1(_05243_ ), .A2(_05279_ ), .A3(_05281_ ), .ZN(_05282_ ) );
OR4_X2 _13036_ ( .A1(_05204_ ), .A2(_05280_ ), .A3(_04952_ ), .A4(_05282_ ), .ZN(_05283_ ) );
INV_X1 _13037_ ( .A(\ID_EX_typ [1] ), .ZN(_05284_ ) );
NOR2_X1 _13038_ ( .A1(_05284_ ), .A2(fanout_net_4 ), .ZN(_05285_ ) );
INV_X1 _13039_ ( .A(fanout_net_5 ), .ZN(_05286_ ) );
AND2_X1 _13040_ ( .A1(_05285_ ), .A2(_05286_ ), .ZN(_05287_ ) );
BUF_X4 _13041_ ( .A(_05287_ ), .Z(_05288_ ) );
INV_X1 _13042_ ( .A(_05288_ ), .ZN(_05289_ ) );
AOI21_X1 _13043_ ( .A(_05289_ ), .B1(_05197_ ), .B2(_05202_ ), .ZN(_05290_ ) );
OAI221_X2 _13044_ ( .A(_04091_ ), .B1(_04949_ ), .B2(_04953_ ), .C1(_05283_ ), .C2(_05290_ ), .ZN(_05291_ ) );
OR2_X2 _13045_ ( .A1(_04949_ ), .A2(_04091_ ), .ZN(_05292_ ) );
AND2_X4 _13046_ ( .A1(_05291_ ), .A2(_05292_ ), .ZN(_05293_ ) );
BUF_X8 _13047_ ( .A(_05293_ ), .Z(_05294_ ) );
MUX2_X1 _13048_ ( .A(_03973_ ), .B(_04088_ ), .S(_05294_ ), .Z(_05295_ ) );
INV_X2 _13049_ ( .A(\ID_EX_typ [3] ), .ZN(_05296_ ) );
BUF_X4 _13050_ ( .A(_05296_ ), .Z(_05297_ ) );
MUX2_X1 _13051_ ( .A(_03954_ ), .B(_05295_ ), .S(_05297_ ), .Z(_05298_ ) );
BUF_X4 _13052_ ( .A(_03879_ ), .Z(_05299_ ) );
NAND2_X1 _13053_ ( .A1(_05298_ ), .A2(_05299_ ), .ZN(_05300_ ) );
BUF_X4 _13054_ ( .A(_03877_ ), .Z(_05301_ ) );
OR2_X1 _13055_ ( .A1(_04088_ ), .A2(fanout_net_4 ), .ZN(_05302_ ) );
BUF_X4 _13056_ ( .A(_04950_ ), .Z(_05303_ ) );
BUF_X4 _13057_ ( .A(_05303_ ), .Z(_05304_ ) );
OAI211_X1 _13058_ ( .A(_05301_ ), .B(_05302_ ), .C1(_03012_ ), .C2(_05304_ ), .ZN(_05305_ ) );
AOI21_X1 _13059_ ( .A(_03891_ ), .B1(_05300_ ), .B2(_05305_ ), .ZN(_00121_ ) );
INV_X2 _13060_ ( .A(_05293_ ), .ZN(_05306_ ) );
BUF_X2 _13061_ ( .A(_05306_ ), .Z(_05307_ ) );
NAND3_X1 _13062_ ( .A1(_03962_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_05308_ ) );
NAND4_X1 _13063_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_05309_ ) );
NOR2_X1 _13064_ ( .A1(_05308_ ), .A2(_05309_ ), .ZN(_05310_ ) );
AND2_X2 _13065_ ( .A1(_03961_ ), .A2(_05310_ ), .ZN(_05311_ ) );
AND4_X1 _13066_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_05312_ ) );
AND2_X1 _13067_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_05313_ ) );
AND4_X1 _13068_ ( .A1(\ID_EX_pc [21] ), .A2(_05312_ ), .A3(\ID_EX_pc [20] ), .A4(_05313_ ), .ZN(_05314_ ) );
AND2_X1 _13069_ ( .A1(_05311_ ), .A2(_05314_ ), .ZN(_05315_ ) );
AND3_X1 _13070_ ( .A1(_05315_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_05316_ ) );
NAND2_X1 _13071_ ( .A1(_05316_ ), .A2(\ID_EX_pc [28] ), .ZN(_05317_ ) );
XNOR2_X1 _13072_ ( .A(_05317_ ), .B(\ID_EX_pc [29] ), .ZN(_05318_ ) );
NAND2_X1 _13073_ ( .A1(_05307_ ), .A2(_05318_ ), .ZN(_05319_ ) );
BUF_X4 _13074_ ( .A(_05296_ ), .Z(_05320_ ) );
NAND2_X1 _13075_ ( .A1(_04082_ ), .A2(_04083_ ), .ZN(_05321_ ) );
NOR2_X1 _13076_ ( .A1(_04085_ ), .A2(_03974_ ), .ZN(_05322_ ) );
XNOR2_X1 _13077_ ( .A(_05321_ ), .B(_05322_ ), .ZN(_05323_ ) );
OAI211_X1 _13078_ ( .A(_05319_ ), .B(_05320_ ), .C1(_05307_ ), .C2(_05323_ ), .ZN(_05324_ ) );
BUF_X4 _13079_ ( .A(_03879_ ), .Z(_05325_ ) );
BUF_X4 _13080_ ( .A(_05297_ ), .Z(_05326_ ) );
INV_X1 _13081_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_05327_ ) );
INV_X1 _13082_ ( .A(\EX_LS_dest_csreg_mem [7] ), .ZN(_05328_ ) );
AOI22_X1 _13083_ ( .A1(_05327_ ), .A2(\ID_EX_csr [9] ), .B1(_05328_ ), .B2(\ID_EX_csr [7] ), .ZN(_05329_ ) );
AOI22_X1 _13084_ ( .A1(fanout_net_3 ), .A2(_03935_ ), .B1(_03926_ ), .B2(\EX_LS_dest_csreg_mem [7] ), .ZN(_05330_ ) );
NAND4_X1 _13085_ ( .A1(_02128_ ), .A2(_05329_ ), .A3(_03904_ ), .A4(_05330_ ), .ZN(_05331_ ) );
NAND2_X1 _13086_ ( .A1(_03903_ ), .A2(_03911_ ), .ZN(_05332_ ) );
NOR3_X1 _13087_ ( .A1(_05331_ ), .A2(_03897_ ), .A3(_05332_ ), .ZN(_05333_ ) );
INV_X1 _13088_ ( .A(\EX_LS_dest_csreg_mem [5] ), .ZN(_05334_ ) );
AOI22_X1 _13089_ ( .A1(\EX_LS_dest_csreg_mem [1] ), .A2(_03915_ ), .B1(_05334_ ), .B2(\ID_EX_csr [5] ), .ZN(_05335_ ) );
OAI221_X1 _13090_ ( .A(_05335_ ), .B1(fanout_net_3 ), .B2(_03935_ ), .C1(_05334_ ), .C2(\ID_EX_csr [5] ), .ZN(_05336_ ) );
OAI211_X1 _13091_ ( .A(_03900_ ), .B(_03908_ ), .C1(_05327_ ), .C2(\ID_EX_csr [9] ), .ZN(_05337_ ) );
INV_X1 _13092_ ( .A(\EX_LS_dest_csreg_mem [1] ), .ZN(_05338_ ) );
INV_X1 _13093_ ( .A(\ID_EX_csr [4] ), .ZN(_05339_ ) );
AOI22_X1 _13094_ ( .A1(_05338_ ), .A2(\ID_EX_csr [1] ), .B1(_05339_ ), .B2(\EX_LS_dest_csreg_mem [4] ), .ZN(_05340_ ) );
OAI211_X1 _13095_ ( .A(_05340_ ), .B(_03910_ ), .C1(\EX_LS_dest_csreg_mem [4] ), .C2(_05339_ ), .ZN(_05341_ ) );
NOR3_X1 _13096_ ( .A1(_05336_ ), .A2(_05337_ ), .A3(_05341_ ), .ZN(_05342_ ) );
AND2_X1 _13097_ ( .A1(_05333_ ), .A2(_05342_ ), .ZN(_05343_ ) );
INV_X1 _13098_ ( .A(_05343_ ), .ZN(_05344_ ) );
NOR2_X1 _13099_ ( .A1(_05344_ ), .A2(\EX_LS_result_csreg_mem [29] ), .ZN(_05345_ ) );
AND4_X1 _13100_ ( .A1(\ID_EX_csr [10] ), .A2(_03948_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_05346_ ) );
AND3_X1 _13101_ ( .A1(_05346_ ), .A2(_03946_ ), .A3(_03916_ ), .ZN(_05347_ ) );
AND2_X2 _13102_ ( .A1(_05347_ ), .A2(_03931_ ), .ZN(_05348_ ) );
NAND3_X1 _13103_ ( .A1(_03928_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_03943_ ), .ZN(_05349_ ) );
NAND3_X1 _13104_ ( .A1(_03928_ ), .A2(\mepc [29] ), .A3(_03931_ ), .ZN(_05350_ ) );
NOR2_X1 _13105_ ( .A1(_03930_ ), .A2(_03941_ ), .ZN(_05351_ ) );
BUF_X4 _13106_ ( .A(_03923_ ), .Z(_05352_ ) );
NAND4_X1 _13107_ ( .A1(_05351_ ), .A2(_05352_ ), .A3(\mtvec [29] ), .A4(_03919_ ), .ZN(_05353_ ) );
NAND4_X1 _13108_ ( .A1(_03936_ ), .A2(_03923_ ), .A3(\mycsreg.CSReg[0][29] ), .A4(_03919_ ), .ZN(_05354_ ) );
NAND4_X1 _13109_ ( .A1(_05349_ ), .A2(_05350_ ), .A3(_05353_ ), .A4(_05354_ ), .ZN(_05355_ ) );
NOR3_X1 _13110_ ( .A1(_05343_ ), .A2(_05348_ ), .A3(_05355_ ), .ZN(_05356_ ) );
NOR2_X1 _13111_ ( .A1(_05345_ ), .A2(_05356_ ), .ZN(_05357_ ) );
OAI211_X1 _13112_ ( .A(_05324_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05357_ ), .ZN(_05358_ ) );
MUX2_X1 _13113_ ( .A(_05323_ ), .B(_03049_ ), .S(fanout_net_4 ), .Z(_05359_ ) );
BUF_X2 _13114_ ( .A(_03878_ ), .Z(_05360_ ) );
OR2_X1 _13115_ ( .A1(_05359_ ), .A2(_05360_ ), .ZN(_05361_ ) );
AOI21_X1 _13116_ ( .A(_03891_ ), .B1(_05358_ ), .B2(_05361_ ), .ZN(_00122_ ) );
BUF_X4 _13117_ ( .A(_03878_ ), .Z(_05362_ ) );
BUF_X4 _13118_ ( .A(_05362_ ), .Z(_05363_ ) );
BUF_X4 _13119_ ( .A(_05297_ ), .Z(_05364_ ) );
BUF_X4 _13120_ ( .A(_05344_ ), .Z(_05365_ ) );
NAND3_X1 _13121_ ( .A1(_03929_ ), .A2(\mepc [20] ), .A3(_03931_ ), .ZN(_05366_ ) );
BUF_X2 _13122_ ( .A(_05351_ ), .Z(_05367_ ) );
BUF_X2 _13123_ ( .A(_03919_ ), .Z(_05368_ ) );
NAND4_X1 _13124_ ( .A1(_05367_ ), .A2(_03924_ ), .A3(\mtvec [20] ), .A4(_05368_ ), .ZN(_05369_ ) );
BUF_X4 _13125_ ( .A(_03936_ ), .Z(_05370_ ) );
NAND4_X1 _13126_ ( .A1(_05370_ ), .A2(_05352_ ), .A3(\mycsreg.CSReg[0][20] ), .A4(_05368_ ), .ZN(_05371_ ) );
AND3_X1 _13127_ ( .A1(_05366_ ), .A2(_05369_ ), .A3(_05371_ ), .ZN(_05372_ ) );
INV_X1 _13128_ ( .A(_05348_ ), .ZN(_05373_ ) );
BUF_X4 _13129_ ( .A(_03928_ ), .Z(_05374_ ) );
BUF_X4 _13130_ ( .A(_03943_ ), .Z(_05375_ ) );
NAND3_X1 _13131_ ( .A1(_05374_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_05375_ ), .ZN(_05376_ ) );
NAND2_X1 _13132_ ( .A1(_05347_ ), .A2(_03943_ ), .ZN(_05377_ ) );
BUF_X2 _13133_ ( .A(_05377_ ), .Z(_05378_ ) );
NAND4_X1 _13134_ ( .A1(_05372_ ), .A2(_05373_ ), .A3(_05376_ ), .A4(_05378_ ), .ZN(_05379_ ) );
NAND2_X1 _13135_ ( .A1(_05365_ ), .A2(_05379_ ), .ZN(_05380_ ) );
BUF_X2 _13136_ ( .A(_05333_ ), .Z(_05381_ ) );
BUF_X4 _13137_ ( .A(_05342_ ), .Z(_05382_ ) );
NAND3_X1 _13138_ ( .A1(_05381_ ), .A2(_05382_ ), .A3(\EX_LS_result_csreg_mem [20] ), .ZN(_05383_ ) );
AND2_X1 _13139_ ( .A1(_05380_ ), .A2(_05383_ ), .ZN(_05384_ ) );
INV_X1 _13140_ ( .A(_05384_ ), .ZN(_05385_ ) );
BUF_X8 _13141_ ( .A(_05293_ ), .Z(_05386_ ) );
BUF_X4 _13142_ ( .A(_05386_ ), .Z(_05387_ ) );
NAND3_X1 _13143_ ( .A1(_03961_ ), .A2(_05310_ ), .A3(_05313_ ), .ZN(_05388_ ) );
INV_X1 _13144_ ( .A(\ID_EX_pc [20] ), .ZN(_05389_ ) );
XNOR2_X1 _13145_ ( .A(_05388_ ), .B(_05389_ ), .ZN(_05390_ ) );
OAI21_X1 _13146_ ( .A(_05320_ ), .B1(_05387_ ), .B2(_05390_ ), .ZN(_05391_ ) );
NOR2_X1 _13147_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_05392_ ) );
NOR3_X1 _13148_ ( .A1(_04039_ ), .A2(_04056_ ), .A3(_05392_ ), .ZN(_05393_ ) );
NAND3_X1 _13149_ ( .A1(_05393_ ), .A2(_04050_ ), .A3(_04051_ ), .ZN(_05394_ ) );
NAND2_X1 _13150_ ( .A1(_05394_ ), .A2(_04064_ ), .ZN(_05395_ ) );
XNOR2_X1 _13151_ ( .A(_05395_ ), .B(_04044_ ), .ZN(_05396_ ) );
AND3_X1 _13152_ ( .A1(_05291_ ), .A2(_05292_ ), .A3(_05396_ ), .ZN(_05397_ ) );
OAI221_X1 _13153_ ( .A(_05363_ ), .B1(_05364_ ), .B2(_05385_ ), .C1(_05391_ ), .C2(_05397_ ), .ZN(_05398_ ) );
AND2_X2 _13154_ ( .A1(_03877_ ), .A2(fanout_net_4 ), .ZN(_05399_ ) );
AND3_X1 _13155_ ( .A1(_03020_ ), .A2(_03017_ ), .A3(_05399_ ), .ZN(_05400_ ) );
AND2_X2 _13156_ ( .A1(_03876_ ), .A2(_04950_ ), .ZN(_05401_ ) );
BUF_X4 _13157_ ( .A(_05401_ ), .Z(_05402_ ) );
AOI21_X1 _13158_ ( .A(_05400_ ), .B1(_05402_ ), .B2(_05396_ ), .ZN(_05403_ ) );
AOI21_X1 _13159_ ( .A(_03891_ ), .B1(_05398_ ), .B2(_05403_ ), .ZN(_00123_ ) );
BUF_X4 _13160_ ( .A(_03928_ ), .Z(_05404_ ) );
BUF_X4 _13161_ ( .A(_03943_ ), .Z(_05405_ ) );
NAND3_X1 _13162_ ( .A1(_05404_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_05405_ ), .ZN(_05406_ ) );
NAND3_X1 _13163_ ( .A1(_05404_ ), .A2(\mepc [19] ), .A3(_03932_ ), .ZN(_05407_ ) );
BUF_X2 _13164_ ( .A(_03936_ ), .Z(_05408_ ) );
BUF_X2 _13165_ ( .A(_03919_ ), .Z(_05409_ ) );
NAND4_X1 _13166_ ( .A1(_05408_ ), .A2(_03938_ ), .A3(\mycsreg.CSReg[0][19] ), .A4(_05409_ ), .ZN(_05410_ ) );
AND3_X1 _13167_ ( .A1(_05406_ ), .A2(_05407_ ), .A3(_05410_ ), .ZN(_05411_ ) );
BUF_X2 _13168_ ( .A(_05351_ ), .Z(_05412_ ) );
BUF_X4 _13169_ ( .A(_05352_ ), .Z(_05413_ ) );
BUF_X4 _13170_ ( .A(_03919_ ), .Z(_05414_ ) );
NAND4_X1 _13171_ ( .A1(_05412_ ), .A2(_05413_ ), .A3(\mtvec [19] ), .A4(_05414_ ), .ZN(_05415_ ) );
AND2_X1 _13172_ ( .A1(_05378_ ), .A2(_05415_ ), .ZN(_05416_ ) );
AOI22_X1 _13173_ ( .A1(_05411_ ), .A2(_05416_ ), .B1(_05382_ ), .B2(_05381_ ), .ZN(_05417_ ) );
CLKBUF_X2 _13174_ ( .A(_05333_ ), .Z(_05418_ ) );
CLKBUF_X2 _13175_ ( .A(_05342_ ), .Z(_05419_ ) );
AND3_X1 _13176_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(\EX_LS_result_csreg_mem [19] ), .ZN(_05420_ ) );
NOR2_X1 _13177_ ( .A1(_05417_ ), .A2(_05420_ ), .ZN(_05421_ ) );
INV_X1 _13178_ ( .A(_05421_ ), .ZN(_05422_ ) );
NAND3_X1 _13179_ ( .A1(_03961_ ), .A2(\ID_EX_pc [18] ), .A3(_05310_ ), .ZN(_05423_ ) );
INV_X1 _13180_ ( .A(\ID_EX_pc [19] ), .ZN(_05424_ ) );
XNOR2_X1 _13181_ ( .A(_05423_ ), .B(_05424_ ), .ZN(_05425_ ) );
OAI21_X1 _13182_ ( .A(_05320_ ), .B1(_05387_ ), .B2(_05425_ ), .ZN(_05426_ ) );
AND2_X1 _13183_ ( .A1(_05393_ ), .A2(_04051_ ), .ZN(_05427_ ) );
OAI21_X1 _13184_ ( .A(_04049_ ), .B1(_05427_ ), .B2(_04059_ ), .ZN(_05428_ ) );
INV_X1 _13185_ ( .A(_04062_ ), .ZN(_05429_ ) );
AND2_X1 _13186_ ( .A1(_05428_ ), .A2(_05429_ ), .ZN(_05430_ ) );
XNOR2_X1 _13187_ ( .A(_05430_ ), .B(_04048_ ), .ZN(_05431_ ) );
AND3_X1 _13188_ ( .A1(_05291_ ), .A2(_05292_ ), .A3(_05431_ ), .ZN(_05432_ ) );
OAI221_X1 _13189_ ( .A(_05363_ ), .B1(_05364_ ), .B2(_05422_ ), .C1(_05426_ ), .C2(_05432_ ), .ZN(_05433_ ) );
BUF_X2 _13190_ ( .A(_05303_ ), .Z(_05434_ ) );
NOR3_X1 _13191_ ( .A1(_03027_ ), .A2(_05434_ ), .A3(_05362_ ), .ZN(_05435_ ) );
AOI21_X1 _13192_ ( .A(_05435_ ), .B1(_05402_ ), .B2(_05431_ ), .ZN(_05436_ ) );
AOI21_X1 _13193_ ( .A(_03891_ ), .B1(_05433_ ), .B2(_05436_ ), .ZN(_00124_ ) );
INV_X1 _13194_ ( .A(\ID_EX_pc [18] ), .ZN(_05437_ ) );
XNOR2_X1 _13195_ ( .A(_05311_ ), .B(_05437_ ), .ZN(_05438_ ) );
NOR2_X1 _13196_ ( .A1(_05427_ ), .A2(_04059_ ), .ZN(_05439_ ) );
XNOR2_X1 _13197_ ( .A(_05439_ ), .B(_04049_ ), .ZN(_05440_ ) );
MUX2_X1 _13198_ ( .A(_05438_ ), .B(_05440_ ), .S(_05386_ ), .Z(_05441_ ) );
OR2_X2 _13199_ ( .A1(_05441_ ), .A2(\ID_EX_typ [3] ), .ZN(_05442_ ) );
NAND3_X1 _13200_ ( .A1(_05404_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_05405_ ), .ZN(_05443_ ) );
NAND3_X1 _13201_ ( .A1(_05404_ ), .A2(\mepc [18] ), .A3(_03932_ ), .ZN(_05444_ ) );
NAND4_X1 _13202_ ( .A1(_05370_ ), .A2(_03938_ ), .A3(\mycsreg.CSReg[0][18] ), .A4(_05409_ ), .ZN(_05445_ ) );
AND3_X1 _13203_ ( .A1(_05443_ ), .A2(_05444_ ), .A3(_05445_ ), .ZN(_05446_ ) );
NAND4_X1 _13204_ ( .A1(_05367_ ), .A2(_05413_ ), .A3(\mtvec [18] ), .A4(_05414_ ), .ZN(_05447_ ) );
AND2_X1 _13205_ ( .A1(_05378_ ), .A2(_05447_ ), .ZN(_05448_ ) );
AOI22_X1 _13206_ ( .A1(_05446_ ), .A2(_05448_ ), .B1(_05382_ ), .B2(_05418_ ), .ZN(_05449_ ) );
AND3_X1 _13207_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(\EX_LS_result_csreg_mem [18] ), .ZN(_05450_ ) );
NOR2_X1 _13208_ ( .A1(_05449_ ), .A2(_05450_ ), .ZN(_05451_ ) );
INV_X1 _13209_ ( .A(_05451_ ), .ZN(_05452_ ) );
OAI211_X1 _13210_ ( .A(_05442_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05452_ ), .ZN(_05453_ ) );
BUF_X4 _13211_ ( .A(_05399_ ), .Z(_05454_ ) );
AOI22_X1 _13212_ ( .A1(_03029_ ), .A2(_05454_ ), .B1(_05402_ ), .B2(_05440_ ), .ZN(_05455_ ) );
AOI21_X1 _13213_ ( .A(_03891_ ), .B1(_05453_ ), .B2(_05455_ ), .ZN(_00125_ ) );
BUF_X4 _13214_ ( .A(_05333_ ), .Z(_05456_ ) );
BUF_X4 _13215_ ( .A(_05456_ ), .Z(_05457_ ) );
BUF_X4 _13216_ ( .A(_05382_ ), .Z(_05458_ ) );
NAND3_X1 _13217_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(\EX_LS_result_csreg_mem [17] ), .ZN(_05459_ ) );
BUF_X4 _13218_ ( .A(_03928_ ), .Z(_05460_ ) );
AND3_X1 _13219_ ( .A1(_05460_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_05405_ ), .ZN(_05461_ ) );
AND4_X1 _13220_ ( .A1(\mycsreg.CSReg[0][17] ), .A2(_05408_ ), .A3(_03938_ ), .A4(_05414_ ), .ZN(_05462_ ) );
AND4_X1 _13221_ ( .A1(\mtvec [17] ), .A2(_05367_ ), .A3(_03938_ ), .A4(_05409_ ), .ZN(_05463_ ) );
NOR3_X1 _13222_ ( .A1(_05461_ ), .A2(_05462_ ), .A3(_05463_ ), .ZN(_05464_ ) );
AND2_X1 _13223_ ( .A1(_05347_ ), .A2(_03943_ ), .ZN(_05465_ ) );
NOR2_X1 _13224_ ( .A1(_05348_ ), .A2(_05465_ ), .ZN(_05466_ ) );
BUF_X4 _13225_ ( .A(_05460_ ), .Z(_05467_ ) );
BUF_X4 _13226_ ( .A(_03932_ ), .Z(_05468_ ) );
NAND3_X1 _13227_ ( .A1(_05467_ ), .A2(\mepc [17] ), .A3(_05468_ ), .ZN(_05469_ ) );
AND3_X1 _13228_ ( .A1(_05464_ ), .A2(_05466_ ), .A3(_05469_ ), .ZN(_05470_ ) );
BUF_X2 _13229_ ( .A(_05343_ ), .Z(_05471_ ) );
OAI21_X1 _13230_ ( .A(_05459_ ), .B1(_05470_ ), .B2(_05471_ ), .ZN(_05472_ ) );
INV_X1 _13231_ ( .A(_03961_ ), .ZN(_05473_ ) );
NOR2_X1 _13232_ ( .A1(_05473_ ), .A2(_05308_ ), .ZN(_05474_ ) );
AND3_X1 _13233_ ( .A1(_05474_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05475_ ) );
NAND2_X1 _13234_ ( .A1(_05475_ ), .A2(\ID_EX_pc [16] ), .ZN(_05476_ ) );
XNOR2_X1 _13235_ ( .A(_05476_ ), .B(\ID_EX_pc [17] ), .ZN(_05477_ ) );
AND2_X1 _13236_ ( .A1(_05307_ ), .A2(_05477_ ), .ZN(_05478_ ) );
OR2_X1 _13237_ ( .A1(_05393_ ), .A2(_04056_ ), .ZN(_05479_ ) );
XNOR2_X1 _13238_ ( .A(_05479_ ), .B(_04051_ ), .ZN(_05480_ ) );
OAI21_X1 _13239_ ( .A(_05297_ ), .B1(_05307_ ), .B2(_05480_ ), .ZN(_05481_ ) );
OAI221_X1 _13240_ ( .A(_05363_ ), .B1(_05364_ ), .B2(_05472_ ), .C1(_05478_ ), .C2(_05481_ ), .ZN(_05482_ ) );
NOR3_X1 _13241_ ( .A1(_03031_ ), .A2(_05304_ ), .A3(_03879_ ), .ZN(_05483_ ) );
NOR3_X1 _13242_ ( .A1(_05480_ ), .A2(fanout_net_4 ), .A3(_03879_ ), .ZN(_05484_ ) );
NOR2_X1 _13243_ ( .A1(_05483_ ), .A2(_05484_ ), .ZN(_05485_ ) );
AOI21_X1 _13244_ ( .A(_03891_ ), .B1(_05482_ ), .B2(_05485_ ), .ZN(_00126_ ) );
NAND3_X1 _13245_ ( .A1(_03929_ ), .A2(\mepc [16] ), .A3(_03931_ ), .ZN(_05486_ ) );
NAND4_X1 _13246_ ( .A1(_05367_ ), .A2(_05352_ ), .A3(\mtvec [16] ), .A4(_05368_ ), .ZN(_05487_ ) );
NAND4_X1 _13247_ ( .A1(_05370_ ), .A2(_05352_ ), .A3(\mycsreg.CSReg[0][16] ), .A4(_03919_ ), .ZN(_05488_ ) );
AND3_X1 _13248_ ( .A1(_05486_ ), .A2(_05487_ ), .A3(_05488_ ), .ZN(_05489_ ) );
NAND3_X1 _13249_ ( .A1(_05374_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_05375_ ), .ZN(_05490_ ) );
NAND4_X1 _13250_ ( .A1(_05489_ ), .A2(_05373_ ), .A3(_05378_ ), .A4(_05490_ ), .ZN(_05491_ ) );
NAND2_X1 _13251_ ( .A1(_05365_ ), .A2(_05491_ ), .ZN(_05492_ ) );
NAND3_X1 _13252_ ( .A1(_05381_ ), .A2(_05382_ ), .A3(\EX_LS_result_csreg_mem [16] ), .ZN(_05493_ ) );
AND2_X1 _13253_ ( .A1(_05492_ ), .A2(_05493_ ), .ZN(_05494_ ) );
INV_X1 _13254_ ( .A(_05494_ ), .ZN(_05495_ ) );
NAND3_X1 _13255_ ( .A1(_05474_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05496_ ) );
INV_X1 _13256_ ( .A(\ID_EX_pc [16] ), .ZN(_05497_ ) );
XNOR2_X1 _13257_ ( .A(_05496_ ), .B(_05497_ ), .ZN(_05498_ ) );
OAI21_X1 _13258_ ( .A(_05320_ ), .B1(_05387_ ), .B2(_05498_ ), .ZN(_05499_ ) );
XNOR2_X1 _13259_ ( .A(_04039_ ), .B(_04052_ ), .ZN(_05500_ ) );
AND3_X1 _13260_ ( .A1(_05291_ ), .A2(_05292_ ), .A3(_05500_ ), .ZN(_05501_ ) );
OAI221_X1 _13261_ ( .A(_05363_ ), .B1(_05364_ ), .B2(_05495_ ), .C1(_05499_ ), .C2(_05501_ ), .ZN(_05502_ ) );
NOR4_X1 _13262_ ( .A1(_03032_ ), .A2(_03022_ ), .A3(_05303_ ), .A4(_03878_ ), .ZN(_05503_ ) );
AOI21_X1 _13263_ ( .A(_05503_ ), .B1(_05402_ ), .B2(_05500_ ), .ZN(_05504_ ) );
AOI21_X1 _13264_ ( .A(_03891_ ), .B1(_05502_ ), .B2(_05504_ ), .ZN(_00127_ ) );
INV_X1 _13265_ ( .A(_04008_ ), .ZN(_05505_ ) );
NOR2_X1 _13266_ ( .A1(_04011_ ), .A2(_04012_ ), .ZN(_05506_ ) );
AND2_X1 _13267_ ( .A1(_04006_ ), .A2(_04020_ ), .ZN(_05507_ ) );
OAI21_X1 _13268_ ( .A(_05506_ ), .B1(_05507_ ), .B2(_04029_ ), .ZN(_05508_ ) );
AOI21_X1 _13269_ ( .A(_05505_ ), .B1(_05508_ ), .B2(_04034_ ), .ZN(_05509_ ) );
NOR2_X1 _13270_ ( .A1(_05509_ ), .A2(_04036_ ), .ZN(_05510_ ) );
XNOR2_X1 _13271_ ( .A(_05510_ ), .B(_04007_ ), .ZN(_05511_ ) );
AOI21_X1 _13272_ ( .A(\ID_EX_typ [3] ), .B1(_05386_ ), .B2(_05511_ ), .ZN(_05512_ ) );
INV_X1 _13273_ ( .A(\ID_EX_pc [14] ), .ZN(_05513_ ) );
NOR3_X1 _13274_ ( .A1(_05473_ ), .A2(_05513_ ), .A3(_05308_ ), .ZN(_05514_ ) );
XNOR2_X1 _13275_ ( .A(_05514_ ), .B(\ID_EX_pc [15] ), .ZN(_05515_ ) );
OAI21_X1 _13276_ ( .A(_05512_ ), .B1(_05387_ ), .B2(_05515_ ), .ZN(_05516_ ) );
NAND3_X1 _13277_ ( .A1(_05404_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_05405_ ), .ZN(_05517_ ) );
NAND3_X1 _13278_ ( .A1(_05404_ ), .A2(\mepc [15] ), .A3(_03932_ ), .ZN(_05518_ ) );
NAND4_X1 _13279_ ( .A1(_05370_ ), .A2(_03938_ ), .A3(\mycsreg.CSReg[0][15] ), .A4(_05409_ ), .ZN(_05519_ ) );
AND3_X1 _13280_ ( .A1(_05517_ ), .A2(_05518_ ), .A3(_05519_ ), .ZN(_05520_ ) );
NAND4_X1 _13281_ ( .A1(_05367_ ), .A2(_03938_ ), .A3(\mtvec [15] ), .A4(_05409_ ), .ZN(_05521_ ) );
AND2_X1 _13282_ ( .A1(_05377_ ), .A2(_05521_ ), .ZN(_05522_ ) );
AOI22_X1 _13283_ ( .A1(_05520_ ), .A2(_05522_ ), .B1(_05419_ ), .B2(_05418_ ), .ZN(_05523_ ) );
AND3_X1 _13284_ ( .A1(_05333_ ), .A2(_05342_ ), .A3(\EX_LS_result_csreg_mem [15] ), .ZN(_05524_ ) );
NOR2_X1 _13285_ ( .A1(_05523_ ), .A2(_05524_ ), .ZN(_05525_ ) );
INV_X1 _13286_ ( .A(_05525_ ), .ZN(_05526_ ) );
OAI211_X1 _13287_ ( .A(_05516_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05526_ ), .ZN(_05527_ ) );
BUF_X4 _13288_ ( .A(_05303_ ), .Z(_05528_ ) );
NOR3_X1 _13289_ ( .A1(_03042_ ), .A2(_05528_ ), .A3(_05362_ ), .ZN(_05529_ ) );
AOI21_X1 _13290_ ( .A(_05529_ ), .B1(_05402_ ), .B2(_05511_ ), .ZN(_05530_ ) );
AOI21_X1 _13291_ ( .A(_03891_ ), .B1(_05527_ ), .B2(_05530_ ), .ZN(_00128_ ) );
XNOR2_X1 _13292_ ( .A(_05474_ ), .B(_05513_ ), .ZN(_05531_ ) );
AND3_X1 _13293_ ( .A1(_05508_ ), .A2(_05505_ ), .A3(_04034_ ), .ZN(_05532_ ) );
NOR2_X1 _13294_ ( .A1(_05532_ ), .A2(_05509_ ), .ZN(_05533_ ) );
MUX2_X1 _13295_ ( .A(_05531_ ), .B(_05533_ ), .S(_05294_ ), .Z(_05534_ ) );
OR2_X1 _13296_ ( .A1(_05534_ ), .A2(\ID_EX_typ [3] ), .ZN(_05535_ ) );
NAND3_X1 _13297_ ( .A1(_03928_ ), .A2(\mepc [14] ), .A3(_03931_ ), .ZN(_05536_ ) );
NAND4_X1 _13298_ ( .A1(_05367_ ), .A2(_05352_ ), .A3(\mtvec [14] ), .A4(_05368_ ), .ZN(_05537_ ) );
NAND4_X1 _13299_ ( .A1(_05370_ ), .A2(_05352_ ), .A3(\mycsreg.CSReg[0][14] ), .A4(_03919_ ), .ZN(_05538_ ) );
AND3_X1 _13300_ ( .A1(_05536_ ), .A2(_05537_ ), .A3(_05538_ ), .ZN(_05539_ ) );
NAND3_X1 _13301_ ( .A1(_05374_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_05375_ ), .ZN(_05540_ ) );
NAND4_X1 _13302_ ( .A1(_05539_ ), .A2(_05373_ ), .A3(_05378_ ), .A4(_05540_ ), .ZN(_05541_ ) );
NAND2_X1 _13303_ ( .A1(_05365_ ), .A2(_05541_ ), .ZN(_05542_ ) );
NAND3_X1 _13304_ ( .A1(_05381_ ), .A2(_05382_ ), .A3(\EX_LS_result_csreg_mem [14] ), .ZN(_05543_ ) );
AND2_X1 _13305_ ( .A1(_05542_ ), .A2(_05543_ ), .ZN(_05544_ ) );
INV_X1 _13306_ ( .A(_05544_ ), .ZN(_05545_ ) );
OAI211_X1 _13307_ ( .A(_05535_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05545_ ), .ZN(_05546_ ) );
BUF_X4 _13308_ ( .A(_05401_ ), .Z(_05547_ ) );
AOI22_X1 _13309_ ( .A1(_03043_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05533_ ), .ZN(_05548_ ) );
AOI21_X1 _13310_ ( .A(_03891_ ), .B1(_05546_ ), .B2(_05548_ ), .ZN(_00129_ ) );
AND2_X1 _13311_ ( .A1(_03963_ ), .A2(\ID_EX_pc [12] ), .ZN(_05549_ ) );
INV_X1 _13312_ ( .A(\ID_EX_pc [13] ), .ZN(_05550_ ) );
XNOR2_X1 _13313_ ( .A(_05549_ ), .B(_05550_ ), .ZN(_05551_ ) );
OAI21_X1 _13314_ ( .A(_04010_ ), .B1(_05507_ ), .B2(_04029_ ), .ZN(_05552_ ) );
NAND2_X1 _13315_ ( .A1(_05552_ ), .A2(_04032_ ), .ZN(_05553_ ) );
XNOR2_X1 _13316_ ( .A(_05553_ ), .B(_04012_ ), .ZN(_05554_ ) );
MUX2_X1 _13317_ ( .A(_05551_ ), .B(_05554_ ), .S(_05294_ ), .Z(_05555_ ) );
OR2_X2 _13318_ ( .A1(_05555_ ), .A2(\ID_EX_typ [3] ), .ZN(_05556_ ) );
INV_X1 _13319_ ( .A(\EX_LS_result_csreg_mem [13] ), .ZN(_05557_ ) );
AND3_X1 _13320_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(_05557_ ), .ZN(_05558_ ) );
NOR2_X1 _13321_ ( .A1(_05343_ ), .A2(_05348_ ), .ZN(_05559_ ) );
BUF_X4 _13322_ ( .A(_03929_ ), .Z(_05560_ ) );
BUF_X4 _13323_ ( .A(_05405_ ), .Z(_05561_ ) );
NAND3_X1 _13324_ ( .A1(_05560_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_05561_ ), .ZN(_05562_ ) );
NAND3_X1 _13325_ ( .A1(_05560_ ), .A2(\mepc [13] ), .A3(_05468_ ), .ZN(_05563_ ) );
BUF_X2 _13326_ ( .A(_05351_ ), .Z(_05564_ ) );
BUF_X4 _13327_ ( .A(_03924_ ), .Z(_05565_ ) );
BUF_X2 _13328_ ( .A(_05368_ ), .Z(_05566_ ) );
NAND4_X1 _13329_ ( .A1(_05564_ ), .A2(_05565_ ), .A3(\mtvec [13] ), .A4(_05566_ ), .ZN(_05567_ ) );
BUF_X4 _13330_ ( .A(_05370_ ), .Z(_05568_ ) );
NAND4_X1 _13331_ ( .A1(_05568_ ), .A2(_05565_ ), .A3(\mycsreg.CSReg[0][13] ), .A4(_05566_ ), .ZN(_05569_ ) );
AND4_X1 _13332_ ( .A1(_05562_ ), .A2(_05563_ ), .A3(_05567_ ), .A4(_05569_ ), .ZN(_05570_ ) );
AOI21_X1 _13333_ ( .A(_05558_ ), .B1(_05559_ ), .B2(_05570_ ), .ZN(_05571_ ) );
OAI211_X1 _13334_ ( .A(_05556_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05571_ ), .ZN(_05572_ ) );
NOR3_X1 _13335_ ( .A1(_03046_ ), .A2(_05528_ ), .A3(_05362_ ), .ZN(_05573_ ) );
AOI21_X1 _13336_ ( .A(_05573_ ), .B1(_05402_ ), .B2(_05554_ ), .ZN(_05574_ ) );
AOI21_X1 _13337_ ( .A(_03891_ ), .B1(_05572_ ), .B2(_05574_ ), .ZN(_00130_ ) );
BUF_X4 _13338_ ( .A(_03890_ ), .Z(_05575_ ) );
INV_X1 _13339_ ( .A(\ID_EX_pc [12] ), .ZN(_05576_ ) );
XNOR2_X1 _13340_ ( .A(_03963_ ), .B(_05576_ ), .ZN(_05577_ ) );
NAND2_X1 _13341_ ( .A1(_05307_ ), .A2(_05577_ ), .ZN(_05578_ ) );
OR3_X1 _13342_ ( .A1(_05507_ ), .A2(_04010_ ), .A3(_04029_ ), .ZN(_05579_ ) );
AND2_X1 _13343_ ( .A1(_05579_ ), .A2(_05552_ ), .ZN(_05580_ ) );
NAND3_X1 _13344_ ( .A1(_05291_ ), .A2(_05292_ ), .A3(_05580_ ), .ZN(_05581_ ) );
AOI21_X1 _13345_ ( .A(\ID_EX_typ [3] ), .B1(_05578_ ), .B2(_05581_ ), .ZN(_05582_ ) );
NAND3_X1 _13346_ ( .A1(_03929_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_03943_ ), .ZN(_05583_ ) );
NAND3_X1 _13347_ ( .A1(_03928_ ), .A2(\mepc [12] ), .A3(_03931_ ), .ZN(_05584_ ) );
NAND4_X1 _13348_ ( .A1(_05370_ ), .A2(_05352_ ), .A3(\mycsreg.CSReg[0][12] ), .A4(_05368_ ), .ZN(_05585_ ) );
AND3_X1 _13349_ ( .A1(_05583_ ), .A2(_05584_ ), .A3(_05585_ ), .ZN(_05586_ ) );
BUF_X4 _13350_ ( .A(_05352_ ), .Z(_05587_ ) );
BUF_X2 _13351_ ( .A(_03919_ ), .Z(_05588_ ) );
NAND4_X1 _13352_ ( .A1(_05412_ ), .A2(_05587_ ), .A3(\mtvec [12] ), .A4(_05588_ ), .ZN(_05589_ ) );
NAND4_X1 _13353_ ( .A1(_05586_ ), .A2(_05373_ ), .A3(_05378_ ), .A4(_05589_ ), .ZN(_05590_ ) );
NAND2_X1 _13354_ ( .A1(_05344_ ), .A2(_05590_ ), .ZN(_05591_ ) );
NAND3_X1 _13355_ ( .A1(_05381_ ), .A2(_05382_ ), .A3(\EX_LS_result_csreg_mem [12] ), .ZN(_05592_ ) );
AOI21_X1 _13356_ ( .A(_05297_ ), .B1(_05591_ ), .B2(_05592_ ), .ZN(_05593_ ) );
OAI21_X1 _13357_ ( .A(_05299_ ), .B1(_05582_ ), .B2(_05593_ ), .ZN(_05594_ ) );
AND3_X1 _13358_ ( .A1(_03047_ ), .A2(_03044_ ), .A3(_05399_ ), .ZN(_05595_ ) );
AOI21_X1 _13359_ ( .A(_05595_ ), .B1(_05402_ ), .B2(_05580_ ), .ZN(_05596_ ) );
AOI21_X1 _13360_ ( .A(_05575_ ), .B1(_05594_ ), .B2(_05596_ ), .ZN(_00131_ ) );
BUF_X4 _13361_ ( .A(_05362_ ), .Z(_05597_ ) );
NAND3_X1 _13362_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(\EX_LS_result_csreg_mem [11] ), .ZN(_05598_ ) );
NAND3_X1 _13363_ ( .A1(_05467_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_05561_ ), .ZN(_05599_ ) );
NAND3_X1 _13364_ ( .A1(_05560_ ), .A2(\mepc [11] ), .A3(_05468_ ), .ZN(_05600_ ) );
BUF_X2 _13365_ ( .A(_03924_ ), .Z(_05601_ ) );
NAND4_X1 _13366_ ( .A1(_05568_ ), .A2(_05601_ ), .A3(\mycsreg.CSReg[0][11] ), .A4(_05566_ ), .ZN(_05602_ ) );
NAND3_X1 _13367_ ( .A1(_05599_ ), .A2(_05600_ ), .A3(_05602_ ), .ZN(_05603_ ) );
AND4_X1 _13368_ ( .A1(\mtvec [11] ), .A2(_05412_ ), .A3(_05587_ ), .A4(_05588_ ), .ZN(_05604_ ) );
NOR4_X1 _13369_ ( .A1(_05603_ ), .A2(_05348_ ), .A3(_05465_ ), .A4(_05604_ ), .ZN(_05605_ ) );
OAI21_X1 _13370_ ( .A(_05598_ ), .B1(_05605_ ), .B2(_05471_ ), .ZN(_05606_ ) );
AND2_X1 _13371_ ( .A1(_03961_ ), .A2(\ID_EX_pc [10] ), .ZN(_05607_ ) );
XNOR2_X1 _13372_ ( .A(_05607_ ), .B(\ID_EX_pc [11] ), .ZN(_05608_ ) );
OAI21_X1 _13373_ ( .A(_05320_ ), .B1(_05387_ ), .B2(_05608_ ), .ZN(_05609_ ) );
INV_X1 _13374_ ( .A(_04015_ ), .ZN(_05610_ ) );
NAND2_X1 _13375_ ( .A1(_04006_ ), .A2(_04019_ ), .ZN(_05611_ ) );
AOI21_X1 _13376_ ( .A(_05610_ ), .B1(_05611_ ), .B2(_04027_ ), .ZN(_05612_ ) );
NOR2_X1 _13377_ ( .A1(_05612_ ), .A2(_04022_ ), .ZN(_05613_ ) );
XNOR2_X1 _13378_ ( .A(_05613_ ), .B(_04014_ ), .ZN(_05614_ ) );
AND3_X1 _13379_ ( .A1(_05291_ ), .A2(_05292_ ), .A3(_05614_ ), .ZN(_05615_ ) );
OAI221_X1 _13380_ ( .A(_05597_ ), .B1(_05364_ ), .B2(_05606_ ), .C1(_05609_ ), .C2(_05615_ ), .ZN(_05616_ ) );
AOI21_X1 _13381_ ( .A(_02860_ ), .B1(_02662_ ), .B2(_02807_ ), .ZN(_05617_ ) );
AND3_X1 _13382_ ( .A1(_02808_ ), .A2(_02829_ ), .A3(_02827_ ), .ZN(_05618_ ) );
NOR3_X1 _13383_ ( .A1(_05617_ ), .A2(_02863_ ), .A3(_05618_ ), .ZN(_05619_ ) );
NOR2_X1 _13384_ ( .A1(_05619_ ), .A2(_02863_ ), .ZN(_05620_ ) );
XNOR2_X1 _13385_ ( .A(_05620_ ), .B(_02853_ ), .ZN(_05621_ ) );
AOI22_X1 _13386_ ( .A1(_05621_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05614_ ), .ZN(_05622_ ) );
AOI21_X1 _13387_ ( .A(_05575_ ), .B1(_05616_ ), .B2(_05622_ ), .ZN(_00132_ ) );
INV_X1 _13388_ ( .A(\EX_LS_result_csreg_mem [28] ), .ZN(_05623_ ) );
AND3_X1 _13389_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(_05623_ ), .ZN(_05624_ ) );
NAND3_X1 _13390_ ( .A1(_05560_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_05375_ ), .ZN(_05625_ ) );
NAND3_X1 _13391_ ( .A1(_05374_ ), .A2(\mepc [28] ), .A3(_03945_ ), .ZN(_05626_ ) );
NAND4_X1 _13392_ ( .A1(_05408_ ), .A2(_05587_ ), .A3(\mycsreg.CSReg[0][28] ), .A4(_05588_ ), .ZN(_05627_ ) );
NAND4_X1 _13393_ ( .A1(_05564_ ), .A2(_05587_ ), .A3(\mtvec [28] ), .A4(_05588_ ), .ZN(_05628_ ) );
AND4_X1 _13394_ ( .A1(_05625_ ), .A2(_05626_ ), .A3(_05627_ ), .A4(_05628_ ), .ZN(_05629_ ) );
AOI21_X1 _13395_ ( .A(_05624_ ), .B1(_05559_ ), .B2(_05629_ ), .ZN(_05630_ ) );
NAND3_X1 _13396_ ( .A1(_05315_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_05631_ ) );
XNOR2_X1 _13397_ ( .A(_05631_ ), .B(\ID_EX_pc [28] ), .ZN(_05632_ ) );
XOR2_X1 _13398_ ( .A(_04080_ ), .B(_04081_ ), .Z(_05633_ ) );
MUX2_X1 _13399_ ( .A(_05632_ ), .B(_05633_ ), .S(_05294_ ), .Z(_05634_ ) );
MUX2_X1 _13400_ ( .A(_05630_ ), .B(_05634_ ), .S(_05297_ ), .Z(_05635_ ) );
NAND2_X1 _13401_ ( .A1(_05635_ ), .A2(_05299_ ), .ZN(_05636_ ) );
OAI21_X1 _13402_ ( .A(fanout_net_4 ), .B1(_03050_ ), .B2(_02952_ ), .ZN(_05637_ ) );
OAI211_X1 _13403_ ( .A(_05637_ ), .B(_05301_ ), .C1(fanout_net_4 ), .C2(_05633_ ), .ZN(_05638_ ) );
AOI21_X1 _13404_ ( .A(_05575_ ), .B1(_05636_ ), .B2(_05638_ ), .ZN(_00133_ ) );
AND3_X1 _13405_ ( .A1(_05611_ ), .A2(_05610_ ), .A3(_04027_ ), .ZN(_05639_ ) );
NOR2_X1 _13406_ ( .A1(_05639_ ), .A2(_05612_ ), .ZN(_05640_ ) );
AOI21_X1 _13407_ ( .A(\ID_EX_typ [3] ), .B1(_05386_ ), .B2(_05640_ ), .ZN(_05641_ ) );
XNOR2_X1 _13408_ ( .A(_03961_ ), .B(\ID_EX_pc [10] ), .ZN(_05642_ ) );
OAI21_X1 _13409_ ( .A(_05641_ ), .B1(_05387_ ), .B2(_05642_ ), .ZN(_05643_ ) );
NAND3_X1 _13410_ ( .A1(_05460_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_05405_ ), .ZN(_05644_ ) );
NAND4_X1 _13411_ ( .A1(_05408_ ), .A2(_05413_ ), .A3(\mycsreg.CSReg[0][10] ), .A4(_05414_ ), .ZN(_05645_ ) );
NAND4_X1 _13412_ ( .A1(_05412_ ), .A2(_05413_ ), .A3(\mtvec [10] ), .A4(_05414_ ), .ZN(_05646_ ) );
AND3_X1 _13413_ ( .A1(_05644_ ), .A2(_05645_ ), .A3(_05646_ ), .ZN(_05647_ ) );
NAND3_X1 _13414_ ( .A1(_05460_ ), .A2(\mepc [10] ), .A3(_03945_ ), .ZN(_05648_ ) );
AND2_X1 _13415_ ( .A1(_05378_ ), .A2(_05648_ ), .ZN(_05649_ ) );
BUF_X2 _13416_ ( .A(_05342_ ), .Z(_05650_ ) );
AOI22_X1 _13417_ ( .A1(_05647_ ), .A2(_05649_ ), .B1(_05650_ ), .B2(_05381_ ), .ZN(_05651_ ) );
AND3_X1 _13418_ ( .A1(_05381_ ), .A2(_05382_ ), .A3(\EX_LS_result_csreg_mem [10] ), .ZN(_05652_ ) );
NOR2_X1 _13419_ ( .A1(_05651_ ), .A2(_05652_ ), .ZN(_05653_ ) );
INV_X1 _13420_ ( .A(_05653_ ), .ZN(_05654_ ) );
OAI211_X1 _13421_ ( .A(_05643_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05654_ ), .ZN(_05655_ ) );
XNOR2_X1 _13422_ ( .A(_05617_ ), .B(_02830_ ), .ZN(_05656_ ) );
AOI22_X1 _13423_ ( .A1(_05656_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05640_ ), .ZN(_05657_ ) );
AOI21_X1 _13424_ ( .A(_05575_ ), .B1(_05655_ ), .B2(_05657_ ), .ZN(_00134_ ) );
AND2_X1 _13425_ ( .A1(_04006_ ), .A2(_04017_ ), .ZN(_05658_ ) );
NOR2_X1 _13426_ ( .A1(_05658_ ), .A2(_04025_ ), .ZN(_05659_ ) );
XNOR2_X1 _13427_ ( .A(_05659_ ), .B(_04018_ ), .ZN(_05660_ ) );
AOI21_X1 _13428_ ( .A(\ID_EX_typ [3] ), .B1(_05386_ ), .B2(_05660_ ), .ZN(_05661_ ) );
XNOR2_X1 _13429_ ( .A(_03960_ ), .B(\ID_EX_pc [9] ), .ZN(_05662_ ) );
OAI21_X1 _13430_ ( .A(_05661_ ), .B1(_05387_ ), .B2(_05662_ ), .ZN(_05663_ ) );
NAND3_X1 _13431_ ( .A1(_05460_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_05405_ ), .ZN(_05664_ ) );
NAND3_X1 _13432_ ( .A1(_05460_ ), .A2(\mepc [9] ), .A3(_03945_ ), .ZN(_05665_ ) );
NAND4_X1 _13433_ ( .A1(_05408_ ), .A2(_05413_ ), .A3(\mycsreg.CSReg[0][9] ), .A4(_05414_ ), .ZN(_05666_ ) );
AND3_X1 _13434_ ( .A1(_05664_ ), .A2(_05665_ ), .A3(_05666_ ), .ZN(_05667_ ) );
NAND4_X1 _13435_ ( .A1(_05412_ ), .A2(_05413_ ), .A3(\mtvec [9] ), .A4(_05414_ ), .ZN(_05668_ ) );
AND2_X1 _13436_ ( .A1(_05378_ ), .A2(_05668_ ), .ZN(_05669_ ) );
AOI22_X1 _13437_ ( .A1(_05667_ ), .A2(_05669_ ), .B1(_05382_ ), .B2(_05381_ ), .ZN(_05670_ ) );
AND3_X1 _13438_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(\EX_LS_result_csreg_mem [9] ), .ZN(_05671_ ) );
NOR2_X1 _13439_ ( .A1(_05670_ ), .A2(_05671_ ), .ZN(_05672_ ) );
INV_X1 _13440_ ( .A(_05672_ ), .ZN(_05673_ ) );
OAI211_X1 _13441_ ( .A(_05663_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05673_ ), .ZN(_05674_ ) );
NAND2_X1 _13442_ ( .A1(_02662_ ), .A2(_02782_ ), .ZN(_05675_ ) );
AND2_X1 _13443_ ( .A1(_05675_ ), .A2(_02859_ ), .ZN(_05676_ ) );
XNOR2_X1 _13444_ ( .A(_05676_ ), .B(_02858_ ), .ZN(_05677_ ) );
NOR3_X1 _13445_ ( .A1(_05677_ ), .A2(_05528_ ), .A3(_05362_ ), .ZN(_05678_ ) );
AOI21_X1 _13446_ ( .A(_05678_ ), .B1(_05402_ ), .B2(_05660_ ), .ZN(_05679_ ) );
AOI21_X1 _13447_ ( .A(_05575_ ), .B1(_05674_ ), .B2(_05679_ ), .ZN(_00135_ ) );
NAND3_X1 _13448_ ( .A1(_03929_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_03943_ ), .ZN(_05680_ ) );
NAND3_X1 _13449_ ( .A1(_03929_ ), .A2(\mepc [8] ), .A3(_03932_ ), .ZN(_05681_ ) );
NAND4_X1 _13450_ ( .A1(_05370_ ), .A2(_03924_ ), .A3(\mycsreg.CSReg[0][8] ), .A4(_05409_ ), .ZN(_05682_ ) );
AND3_X1 _13451_ ( .A1(_05680_ ), .A2(_05681_ ), .A3(_05682_ ), .ZN(_05683_ ) );
NAND4_X1 _13452_ ( .A1(_05412_ ), .A2(_05587_ ), .A3(\mtvec [8] ), .A4(_05588_ ), .ZN(_05684_ ) );
NAND4_X1 _13453_ ( .A1(_05683_ ), .A2(_05373_ ), .A3(_05378_ ), .A4(_05684_ ), .ZN(_05685_ ) );
NAND2_X1 _13454_ ( .A1(_05365_ ), .A2(_05685_ ), .ZN(_05686_ ) );
NAND3_X1 _13455_ ( .A1(_05456_ ), .A2(_05650_ ), .A3(\EX_LS_result_csreg_mem [8] ), .ZN(_05687_ ) );
AND2_X1 _13456_ ( .A1(_05686_ ), .A2(_05687_ ), .ZN(_05688_ ) );
INV_X1 _13457_ ( .A(_05688_ ), .ZN(_05689_ ) );
XNOR2_X1 _13458_ ( .A(_03959_ ), .B(\ID_EX_pc [8] ), .ZN(_05690_ ) );
OAI21_X1 _13459_ ( .A(_05320_ ), .B1(_05387_ ), .B2(_05690_ ), .ZN(_05691_ ) );
XOR2_X1 _13460_ ( .A(_04006_ ), .B(_04017_ ), .Z(_05692_ ) );
AND3_X1 _13461_ ( .A1(_05291_ ), .A2(_05292_ ), .A3(_05692_ ), .ZN(_05693_ ) );
OAI221_X1 _13462_ ( .A(_05597_ ), .B1(_05364_ ), .B2(_05689_ ), .C1(_05691_ ), .C2(_05693_ ), .ZN(_05694_ ) );
XOR2_X1 _13463_ ( .A(_02662_ ), .B(_02782_ ), .Z(_05695_ ) );
AOI22_X1 _13464_ ( .A1(_05695_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05692_ ), .ZN(_05696_ ) );
AOI21_X1 _13465_ ( .A(_05575_ ), .B1(_05694_ ), .B2(_05696_ ), .ZN(_00136_ ) );
XNOR2_X1 _13466_ ( .A(\ID_EX_pc [7] ), .B(\ID_EX_imm [7] ), .ZN(_05697_ ) );
XNOR2_X1 _13467_ ( .A(_04002_ ), .B(_05697_ ), .ZN(_05698_ ) );
AOI21_X1 _13468_ ( .A(\ID_EX_typ [3] ), .B1(_05386_ ), .B2(_05698_ ), .ZN(_05699_ ) );
XNOR2_X1 _13469_ ( .A(_03958_ ), .B(\ID_EX_pc [7] ), .ZN(_05700_ ) );
OAI21_X1 _13470_ ( .A(_05699_ ), .B1(_05387_ ), .B2(_05700_ ), .ZN(_05701_ ) );
NAND3_X1 _13471_ ( .A1(_05404_ ), .A2(\mepc [7] ), .A3(_03932_ ), .ZN(_05702_ ) );
NAND3_X1 _13472_ ( .A1(_03929_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_03943_ ), .ZN(_05703_ ) );
NAND4_X1 _13473_ ( .A1(_05367_ ), .A2(_03924_ ), .A3(\mtvec [7] ), .A4(_05409_ ), .ZN(_05704_ ) );
NAND4_X1 _13474_ ( .A1(_05370_ ), .A2(_03924_ ), .A3(\mycsreg.CSReg[0][7] ), .A4(_05409_ ), .ZN(_05705_ ) );
AND4_X1 _13475_ ( .A1(_05702_ ), .A2(_05703_ ), .A3(_05704_ ), .A4(_05705_ ), .ZN(_05706_ ) );
OR2_X1 _13476_ ( .A1(_05471_ ), .A2(_05706_ ), .ZN(_05707_ ) );
NAND3_X1 _13477_ ( .A1(_05456_ ), .A2(_05650_ ), .A3(\EX_LS_result_csreg_mem [7] ), .ZN(_05708_ ) );
AND2_X1 _13478_ ( .A1(_05707_ ), .A2(_05708_ ), .ZN(_05709_ ) );
INV_X1 _13479_ ( .A(_05709_ ), .ZN(_05710_ ) );
OAI211_X1 _13480_ ( .A(_05701_ ), .B(_05325_ ), .C1(_05326_ ), .C2(_05710_ ), .ZN(_05711_ ) );
AND3_X1 _13481_ ( .A1(_02558_ ), .A2(_02581_ ), .A3(_02605_ ), .ZN(_05712_ ) );
OAI21_X1 _13482_ ( .A(_02628_ ), .B1(_05712_ ), .B2(_02660_ ), .ZN(_05713_ ) );
AND2_X1 _13483_ ( .A1(_02626_ ), .A2(\ID_EX_imm [6] ), .ZN(_05714_ ) );
INV_X1 _13484_ ( .A(_05714_ ), .ZN(_05715_ ) );
NAND2_X1 _13485_ ( .A1(_05713_ ), .A2(_05715_ ), .ZN(_05716_ ) );
NAND2_X1 _13486_ ( .A1(_02652_ ), .A2(_02650_ ), .ZN(_05717_ ) );
XNOR2_X1 _13487_ ( .A(_05716_ ), .B(_05717_ ), .ZN(_05718_ ) );
AOI22_X1 _13488_ ( .A1(_05718_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05698_ ), .ZN(_05719_ ) );
AOI21_X1 _13489_ ( .A(_05575_ ), .B1(_05711_ ), .B2(_05719_ ), .ZN(_00137_ ) );
INV_X1 _13490_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_05720_ ) );
AND3_X1 _13491_ ( .A1(_05333_ ), .A2(_05342_ ), .A3(_05720_ ), .ZN(_05721_ ) );
NAND3_X1 _13492_ ( .A1(_05374_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_05375_ ), .ZN(_05722_ ) );
NAND3_X1 _13493_ ( .A1(_05460_ ), .A2(\mepc [6] ), .A3(_03945_ ), .ZN(_05723_ ) );
NAND4_X1 _13494_ ( .A1(_05412_ ), .A2(_05413_ ), .A3(\mtvec [6] ), .A4(_05414_ ), .ZN(_05724_ ) );
NAND4_X1 _13495_ ( .A1(_05408_ ), .A2(_05413_ ), .A3(\mycsreg.CSReg[0][6] ), .A4(_05414_ ), .ZN(_05725_ ) );
AND4_X1 _13496_ ( .A1(_05722_ ), .A2(_05723_ ), .A3(_05724_ ), .A4(_05725_ ), .ZN(_05726_ ) );
AOI21_X1 _13497_ ( .A(_05721_ ), .B1(_05559_ ), .B2(_05726_ ), .ZN(_05727_ ) );
INV_X1 _13498_ ( .A(\ID_EX_pc [6] ), .ZN(_05728_ ) );
XNOR2_X1 _13499_ ( .A(_03957_ ), .B(_05728_ ), .ZN(_05729_ ) );
XOR2_X1 _13500_ ( .A(_03998_ ), .B(_03999_ ), .Z(_05730_ ) );
MUX2_X1 _13501_ ( .A(_05729_ ), .B(_05730_ ), .S(_05294_ ), .Z(_05731_ ) );
MUX2_X1 _13502_ ( .A(_05727_ ), .B(_05731_ ), .S(_05297_ ), .Z(_05732_ ) );
NAND2_X1 _13503_ ( .A1(_05732_ ), .A2(_05299_ ), .ZN(_05733_ ) );
NOR2_X1 _13504_ ( .A1(_05712_ ), .A2(_02660_ ), .ZN(_05734_ ) );
XNOR2_X1 _13505_ ( .A(_05734_ ), .B(_02628_ ), .ZN(_05735_ ) );
AOI22_X1 _13506_ ( .A1(_05735_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05730_ ), .ZN(_05736_ ) );
AOI21_X1 _13507_ ( .A(_05575_ ), .B1(_05733_ ), .B2(_05736_ ), .ZN(_00138_ ) );
INV_X1 _13508_ ( .A(\ID_EX_pc [5] ), .ZN(_05737_ ) );
XNOR2_X1 _13509_ ( .A(_03956_ ), .B(_05737_ ), .ZN(_05738_ ) );
AND2_X1 _13510_ ( .A1(_03994_ ), .A2(_03995_ ), .ZN(_05739_ ) );
NOR2_X1 _13511_ ( .A1(_05739_ ), .A2(_03983_ ), .ZN(_05740_ ) );
XOR2_X1 _13512_ ( .A(\ID_EX_pc [5] ), .B(\ID_EX_imm [5] ), .Z(_05741_ ) );
XNOR2_X1 _13513_ ( .A(_05740_ ), .B(_05741_ ), .ZN(_05742_ ) );
MUX2_X1 _13514_ ( .A(_05738_ ), .B(_05742_ ), .S(_05294_ ), .Z(_05743_ ) );
OR2_X1 _13515_ ( .A1(_05743_ ), .A2(\ID_EX_typ [3] ), .ZN(_05744_ ) );
AND2_X1 _13516_ ( .A1(_03950_ ), .A2(_03931_ ), .ZN(_05745_ ) );
INV_X1 _13517_ ( .A(_05745_ ), .ZN(_05746_ ) );
NAND3_X1 _13518_ ( .A1(_05374_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_05375_ ), .ZN(_05747_ ) );
NAND3_X1 _13519_ ( .A1(_05460_ ), .A2(\mepc [5] ), .A3(_03945_ ), .ZN(_05748_ ) );
NAND4_X1 _13520_ ( .A1(_03920_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [5] ), .A4(_05587_ ), .ZN(_05749_ ) );
NAND4_X1 _13521_ ( .A1(_05746_ ), .A2(_05747_ ), .A3(_05748_ ), .A4(_05749_ ), .ZN(_05750_ ) );
NAND3_X1 _13522_ ( .A1(_03937_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_05565_ ), .ZN(_05751_ ) );
OAI21_X1 _13523_ ( .A(_05751_ ), .B1(_03902_ ), .B2(_03912_ ), .ZN(_05752_ ) );
NOR2_X1 _13524_ ( .A1(_05750_ ), .A2(_05752_ ), .ZN(_05753_ ) );
CLKBUF_X2 _13525_ ( .A(_03902_ ), .Z(_05754_ ) );
CLKBUF_X2 _13526_ ( .A(_03912_ ), .Z(_05755_ ) );
NOR3_X1 _13527_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [5] ), .ZN(_05756_ ) );
NOR2_X1 _13528_ ( .A1(_05753_ ), .A2(_05756_ ), .ZN(_05757_ ) );
OAI211_X1 _13529_ ( .A(_05744_ ), .B(_05363_ ), .C1(_05326_ ), .C2(_05757_ ), .ZN(_05758_ ) );
OAI21_X1 _13530_ ( .A(_02605_ ), .B1(_02551_ ), .B2(_02556_ ), .ZN(_05759_ ) );
OAI21_X1 _13531_ ( .A(_05759_ ), .B1(_02604_ ), .B2(_02656_ ), .ZN(_05760_ ) );
XNOR2_X1 _13532_ ( .A(_05760_ ), .B(_02580_ ), .ZN(_05761_ ) );
AOI22_X1 _13533_ ( .A1(_05761_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05742_ ), .ZN(_05762_ ) );
AOI21_X1 _13534_ ( .A(_05575_ ), .B1(_05758_ ), .B2(_05762_ ), .ZN(_00139_ ) );
XNOR2_X1 _13535_ ( .A(_03955_ ), .B(\ID_EX_pc [4] ), .ZN(_05763_ ) );
XOR2_X1 _13536_ ( .A(_03994_ ), .B(_03995_ ), .Z(_05764_ ) );
INV_X1 _13537_ ( .A(_05764_ ), .ZN(_05765_ ) );
MUX2_X1 _13538_ ( .A(_05763_ ), .B(_05765_ ), .S(_05386_ ), .Z(_05766_ ) );
NAND2_X1 _13539_ ( .A1(_05766_ ), .A2(_05320_ ), .ZN(_05767_ ) );
INV_X1 _13540_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_05768_ ) );
AND3_X1 _13541_ ( .A1(_05456_ ), .A2(_05650_ ), .A3(_05768_ ), .ZN(_05769_ ) );
BUF_X4 _13542_ ( .A(_05565_ ), .Z(_05770_ ) );
BUF_X4 _13543_ ( .A(_05414_ ), .Z(_05771_ ) );
NAND4_X1 _13544_ ( .A1(_05564_ ), .A2(_05770_ ), .A3(\mtvec [4] ), .A4(_05771_ ), .ZN(_05772_ ) );
NAND3_X1 _13545_ ( .A1(_05467_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_05561_ ), .ZN(_05773_ ) );
NAND3_X1 _13546_ ( .A1(_05467_ ), .A2(\mepc [4] ), .A3(_05468_ ), .ZN(_05774_ ) );
NAND4_X1 _13547_ ( .A1(_05568_ ), .A2(_05770_ ), .A3(\mycsreg.CSReg[0][4] ), .A4(_05771_ ), .ZN(_05775_ ) );
AND4_X1 _13548_ ( .A1(_05772_ ), .A2(_05773_ ), .A3(_05774_ ), .A4(_05775_ ), .ZN(_05776_ ) );
AOI21_X1 _13549_ ( .A(_05769_ ), .B1(_05559_ ), .B2(_05776_ ), .ZN(_05777_ ) );
OAI211_X1 _13550_ ( .A(_05767_ ), .B(_05363_ ), .C1(_05326_ ), .C2(_05777_ ), .ZN(_05778_ ) );
XNOR2_X1 _13551_ ( .A(_02557_ ), .B(_02605_ ), .ZN(_05779_ ) );
AOI22_X1 _13552_ ( .A1(_05779_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05764_ ), .ZN(_05780_ ) );
AOI21_X1 _13553_ ( .A(_05575_ ), .B1(_05778_ ), .B2(_05780_ ), .ZN(_00140_ ) );
BUF_X4 _13554_ ( .A(_03890_ ), .Z(_05781_ ) );
NAND2_X1 _13555_ ( .A1(_03990_ ), .A2(_03991_ ), .ZN(_05782_ ) );
NOR2_X1 _13556_ ( .A1(_03993_ ), .A2(_03984_ ), .ZN(_05783_ ) );
XOR2_X1 _13557_ ( .A(_05782_ ), .B(_05783_ ), .Z(_05784_ ) );
AOI21_X1 _13558_ ( .A(\ID_EX_typ [3] ), .B1(_05386_ ), .B2(_05784_ ), .ZN(_05785_ ) );
XNOR2_X1 _13559_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .ZN(_05786_ ) );
OAI21_X1 _13560_ ( .A(_05785_ ), .B1(_05387_ ), .B2(_05786_ ), .ZN(_05787_ ) );
INV_X1 _13561_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_05788_ ) );
AND3_X1 _13562_ ( .A1(_05381_ ), .A2(_05419_ ), .A3(_05788_ ), .ZN(_05789_ ) );
NAND3_X1 _13563_ ( .A1(_05560_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_05561_ ), .ZN(_05790_ ) );
NAND3_X1 _13564_ ( .A1(_05560_ ), .A2(\mepc [3] ), .A3(_05468_ ), .ZN(_05791_ ) );
NAND4_X1 _13565_ ( .A1(_05568_ ), .A2(_05601_ ), .A3(\mycsreg.CSReg[0][3] ), .A4(_05566_ ), .ZN(_05792_ ) );
NAND4_X1 _13566_ ( .A1(_05564_ ), .A2(_05601_ ), .A3(\mtvec [3] ), .A4(_05566_ ), .ZN(_05793_ ) );
AND4_X1 _13567_ ( .A1(_05790_ ), .A2(_05791_ ), .A3(_05792_ ), .A4(_05793_ ), .ZN(_05794_ ) );
AOI21_X1 _13568_ ( .A(_05789_ ), .B1(_05559_ ), .B2(_05794_ ), .ZN(_05795_ ) );
OAI211_X1 _13569_ ( .A(_05787_ ), .B(_05363_ ), .C1(_05364_ ), .C2(_05795_ ), .ZN(_05796_ ) );
NOR2_X1 _13570_ ( .A1(_02505_ ), .A2(_02550_ ), .ZN(_05797_ ) );
NOR2_X1 _13571_ ( .A1(_05797_ ), .A2(_02553_ ), .ZN(_05798_ ) );
XNOR2_X1 _13572_ ( .A(_05798_ ), .B(_02552_ ), .ZN(_05799_ ) );
AOI22_X1 _13573_ ( .A1(_05799_ ), .A2(_05454_ ), .B1(_05547_ ), .B2(_05784_ ), .ZN(_05800_ ) );
AOI21_X1 _13574_ ( .A(_05781_ ), .B1(_05796_ ), .B2(_05800_ ), .ZN(_00141_ ) );
AND3_X1 _13575_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(\EX_LS_result_csreg_mem [2] ), .ZN(_05801_ ) );
INV_X1 _13576_ ( .A(_05801_ ), .ZN(_05802_ ) );
NAND3_X1 _13577_ ( .A1(_05404_ ), .A2(\mycsreg.CSReg[3][2] ), .A3(_05405_ ), .ZN(_05803_ ) );
NAND4_X1 _13578_ ( .A1(_05408_ ), .A2(_03938_ ), .A3(\mycsreg.CSReg[0][2] ), .A4(_05409_ ), .ZN(_05804_ ) );
NAND4_X1 _13579_ ( .A1(_05367_ ), .A2(_03938_ ), .A3(\mtvec [2] ), .A4(_05409_ ), .ZN(_05805_ ) );
AND3_X1 _13580_ ( .A1(_05803_ ), .A2(_05804_ ), .A3(_05805_ ), .ZN(_05806_ ) );
NAND3_X1 _13581_ ( .A1(_05404_ ), .A2(\mepc [2] ), .A3(_03945_ ), .ZN(_05807_ ) );
AND2_X1 _13582_ ( .A1(_05378_ ), .A2(_05807_ ), .ZN(_05808_ ) );
AND2_X1 _13583_ ( .A1(_05806_ ), .A2(_05808_ ), .ZN(_05809_ ) );
OAI21_X1 _13584_ ( .A(_05802_ ), .B1(_05809_ ), .B2(_05471_ ), .ZN(_05810_ ) );
OR3_X1 _13585_ ( .A1(_03988_ ), .A2(_03989_ ), .A3(_03985_ ), .ZN(_05811_ ) );
AND2_X1 _13586_ ( .A1(_05811_ ), .A2(_03990_ ), .ZN(_05812_ ) );
MUX2_X1 _13587_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B(_05812_ ), .S(_05294_ ), .Z(_05813_ ) );
MUX2_X1 _13588_ ( .A(_05810_ ), .B(_05813_ ), .S(_05297_ ), .Z(_05814_ ) );
NAND2_X1 _13589_ ( .A1(_05814_ ), .A2(_05299_ ), .ZN(_05815_ ) );
XOR2_X1 _13590_ ( .A(_02505_ ), .B(_02550_ ), .Z(_05816_ ) );
AOI22_X1 _13591_ ( .A1(_05816_ ), .A2(_05399_ ), .B1(_05547_ ), .B2(_05812_ ), .ZN(_05817_ ) );
AOI21_X1 _13592_ ( .A(_05781_ ), .B1(_05815_ ), .B2(_05817_ ), .ZN(_00142_ ) );
NAND3_X1 _13593_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(\EX_LS_result_csreg_mem [1] ), .ZN(_05818_ ) );
NAND3_X1 _13594_ ( .A1(_05467_ ), .A2(\mepc [1] ), .A3(_05468_ ), .ZN(_05819_ ) );
NAND3_X1 _13595_ ( .A1(_05467_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_05561_ ), .ZN(_05820_ ) );
BUF_X4 _13596_ ( .A(_05413_ ), .Z(_05821_ ) );
NAND4_X1 _13597_ ( .A1(_05564_ ), .A2(_05821_ ), .A3(\mtvec [1] ), .A4(_05771_ ), .ZN(_05822_ ) );
NAND4_X1 _13598_ ( .A1(_05568_ ), .A2(_05601_ ), .A3(\mycsreg.CSReg[0][1] ), .A4(_05771_ ), .ZN(_05823_ ) );
AND4_X1 _13599_ ( .A1(_05819_ ), .A2(_05820_ ), .A3(_05822_ ), .A4(_05823_ ), .ZN(_05824_ ) );
OAI21_X1 _13600_ ( .A(_05818_ ), .B1(_05471_ ), .B2(_05824_ ), .ZN(_05825_ ) );
XOR2_X1 _13601_ ( .A(_03986_ ), .B(_03987_ ), .Z(_05826_ ) );
INV_X1 _13602_ ( .A(_05826_ ), .ZN(_05827_ ) );
OAI21_X1 _13603_ ( .A(_05320_ ), .B1(_05307_ ), .B2(_05827_ ), .ZN(_05828_ ) );
INV_X1 _13604_ ( .A(\ID_EX_pc [1] ), .ZN(_05829_ ) );
AOI21_X1 _13605_ ( .A(_05829_ ), .B1(_05291_ ), .B2(_05292_ ), .ZN(_05830_ ) );
OAI221_X1 _13606_ ( .A(_05597_ ), .B1(_05320_ ), .B2(_05825_ ), .C1(_05828_ ), .C2(_05830_ ), .ZN(_05831_ ) );
AOI21_X1 _13607_ ( .A(_02480_ ), .B1(_02481_ ), .B2(_02501_ ), .ZN(_05832_ ) );
XNOR2_X1 _13608_ ( .A(_02479_ ), .B(_05832_ ), .ZN(_05833_ ) );
AOI22_X1 _13609_ ( .A1(_05833_ ), .A2(_05399_ ), .B1(_05401_ ), .B2(_05826_ ), .ZN(_05834_ ) );
AOI21_X1 _13610_ ( .A(_05781_ ), .B1(_05831_ ), .B2(_05834_ ), .ZN(_00143_ ) );
NAND3_X1 _13611_ ( .A1(_05311_ ), .A2(\ID_EX_pc [26] ), .A3(_05314_ ), .ZN(_05835_ ) );
XNOR2_X1 _13612_ ( .A(_05835_ ), .B(\ID_EX_pc [27] ), .ZN(_05836_ ) );
NAND2_X1 _13613_ ( .A1(_05307_ ), .A2(_05836_ ), .ZN(_05837_ ) );
OR2_X1 _13614_ ( .A1(_04054_ ), .A2(_04072_ ), .ZN(_05838_ ) );
AND2_X1 _13615_ ( .A1(_05838_ ), .A2(_03982_ ), .ZN(_05839_ ) );
OAI21_X1 _13616_ ( .A(_03976_ ), .B1(_05839_ ), .B2(_04078_ ), .ZN(_05840_ ) );
NAND2_X1 _13617_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_05841_ ) );
NAND2_X1 _13618_ ( .A1(_05840_ ), .A2(_05841_ ), .ZN(_05842_ ) );
XNOR2_X1 _13619_ ( .A(_05842_ ), .B(_03975_ ), .ZN(_05843_ ) );
OAI211_X1 _13620_ ( .A(_05837_ ), .B(_05320_ ), .C1(_05307_ ), .C2(_05843_ ), .ZN(_05844_ ) );
NAND3_X1 _13621_ ( .A1(_05467_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_05561_ ), .ZN(_05845_ ) );
NAND3_X1 _13622_ ( .A1(_05374_ ), .A2(\mepc [27] ), .A3(_05468_ ), .ZN(_05846_ ) );
NAND4_X1 _13623_ ( .A1(_05412_ ), .A2(_05587_ ), .A3(\mtvec [27] ), .A4(_05588_ ), .ZN(_05847_ ) );
AND2_X1 _13624_ ( .A1(_05846_ ), .A2(_05847_ ), .ZN(_05848_ ) );
BUF_X4 _13625_ ( .A(_05587_ ), .Z(_05849_ ) );
NAND4_X1 _13626_ ( .A1(_05568_ ), .A2(_05849_ ), .A3(\mycsreg.CSReg[0][27] ), .A4(_05771_ ), .ZN(_05850_ ) );
NAND4_X1 _13627_ ( .A1(_05559_ ), .A2(_05845_ ), .A3(_05848_ ), .A4(_05850_ ), .ZN(_05851_ ) );
INV_X1 _13628_ ( .A(\EX_LS_result_csreg_mem [27] ), .ZN(_05852_ ) );
NAND3_X1 _13629_ ( .A1(_05456_ ), .A2(_05650_ ), .A3(_05852_ ), .ZN(_05853_ ) );
AND2_X1 _13630_ ( .A1(_05851_ ), .A2(_05853_ ), .ZN(_05854_ ) );
OAI211_X1 _13631_ ( .A(_05844_ ), .B(_05363_ ), .C1(_05364_ ), .C2(_05854_ ), .ZN(_05855_ ) );
MUX2_X1 _13632_ ( .A(_05843_ ), .B(_03053_ ), .S(fanout_net_4 ), .Z(_05856_ ) );
OR2_X1 _13633_ ( .A1(_05856_ ), .A2(_05360_ ), .ZN(_05857_ ) );
AOI21_X1 _13634_ ( .A(_05781_ ), .B1(_05855_ ), .B2(_05857_ ), .ZN(_00144_ ) );
XOR2_X1 _13635_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05858_ ) );
OAI21_X1 _13636_ ( .A(_05296_ ), .B1(_05307_ ), .B2(_05858_ ), .ZN(_05859_ ) );
INV_X1 _13637_ ( .A(\ID_EX_pc [0] ), .ZN(_05860_ ) );
AOI21_X1 _13638_ ( .A(_05859_ ), .B1(_05860_ ), .B2(_05307_ ), .ZN(_05861_ ) );
OR3_X1 _13639_ ( .A1(_03902_ ), .A2(_03912_ ), .A3(\EX_LS_result_csreg_mem [0] ), .ZN(_05862_ ) );
NAND3_X1 _13640_ ( .A1(_03937_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_05601_ ), .ZN(_05863_ ) );
NAND3_X1 _13641_ ( .A1(_05560_ ), .A2(\mepc [0] ), .A3(_05468_ ), .ZN(_05864_ ) );
AND2_X1 _13642_ ( .A1(_05863_ ), .A2(_05864_ ), .ZN(_05865_ ) );
AOI22_X1 _13643_ ( .A1(_03944_ ), .A2(\mycsreg.CSReg[3][0] ), .B1(_05561_ ), .B2(_03950_ ), .ZN(_05866_ ) );
NAND2_X1 _13644_ ( .A1(_05865_ ), .A2(_05866_ ), .ZN(_05867_ ) );
NAND4_X1 _13645_ ( .A1(_03920_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [0] ), .A4(_05821_ ), .ZN(_05868_ ) );
BUF_X2 _13646_ ( .A(_03902_ ), .Z(_05869_ ) );
BUF_X2 _13647_ ( .A(_03912_ ), .Z(_05870_ ) );
OAI21_X1 _13648_ ( .A(_05868_ ), .B1(_05869_ ), .B2(_05870_ ), .ZN(_05871_ ) );
OAI211_X1 _13649_ ( .A(_05862_ ), .B(\ID_EX_typ [3] ), .C1(_05867_ ), .C2(_05871_ ), .ZN(_05872_ ) );
INV_X1 _13650_ ( .A(_05872_ ), .ZN(_05873_ ) );
OAI21_X1 _13651_ ( .A(_05299_ ), .B1(_05861_ ), .B2(_05873_ ), .ZN(_05874_ ) );
NAND3_X1 _13652_ ( .A1(_05858_ ), .A2(_05304_ ), .A3(_05301_ ), .ZN(_05875_ ) );
AOI21_X1 _13653_ ( .A(_05781_ ), .B1(_05874_ ), .B2(_05875_ ), .ZN(_00145_ ) );
NOR3_X1 _13654_ ( .A1(_05869_ ), .A2(_05870_ ), .A3(\EX_LS_result_csreg_mem [26] ), .ZN(_05876_ ) );
NAND3_X1 _13655_ ( .A1(_05374_ ), .A2(\mepc [26] ), .A3(_03945_ ), .ZN(_05877_ ) );
NAND4_X1 _13656_ ( .A1(_03920_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [26] ), .A4(_05565_ ), .ZN(_05878_ ) );
NAND3_X1 _13657_ ( .A1(_05374_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_05375_ ), .ZN(_05879_ ) );
NAND3_X1 _13658_ ( .A1(_03937_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_05601_ ), .ZN(_05880_ ) );
AND4_X1 _13659_ ( .A1(_05877_ ), .A2(_05878_ ), .A3(_05879_ ), .A4(_05880_ ), .ZN(_05881_ ) );
AOI21_X1 _13660_ ( .A(_05876_ ), .B1(_05881_ ), .B2(_03914_ ), .ZN(_05882_ ) );
NAND2_X1 _13661_ ( .A1(_05311_ ), .A2(_05314_ ), .ZN(_05883_ ) );
XNOR2_X1 _13662_ ( .A(_05883_ ), .B(\ID_EX_pc [26] ), .ZN(_05884_ ) );
OR3_X1 _13663_ ( .A1(_05839_ ), .A2(_03976_ ), .A3(_04078_ ), .ZN(_05885_ ) );
AND2_X1 _13664_ ( .A1(_05885_ ), .A2(_05840_ ), .ZN(_05886_ ) );
MUX2_X1 _13665_ ( .A(_05884_ ), .B(_05886_ ), .S(_05294_ ), .Z(_05887_ ) );
MUX2_X1 _13666_ ( .A(_05882_ ), .B(_05887_ ), .S(_05297_ ), .Z(_05888_ ) );
NAND2_X1 _13667_ ( .A1(_05888_ ), .A2(_05299_ ), .ZN(_05889_ ) );
AOI21_X1 _13668_ ( .A(_05528_ ), .B1(_03054_ ), .B2(_03051_ ), .ZN(_05890_ ) );
BUF_X2 _13669_ ( .A(_03877_ ), .Z(_05891_ ) );
OAI21_X1 _13670_ ( .A(_05891_ ), .B1(_05886_ ), .B2(fanout_net_4 ), .ZN(_05892_ ) );
OR2_X1 _13671_ ( .A1(_05890_ ), .A2(_05892_ ), .ZN(_05893_ ) );
AOI21_X1 _13672_ ( .A(_05781_ ), .B1(_05889_ ), .B2(_05893_ ), .ZN(_00146_ ) );
AND3_X1 _13673_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(\EX_LS_result_csreg_mem [25] ), .ZN(_05894_ ) );
INV_X1 _13674_ ( .A(_05894_ ), .ZN(_05895_ ) );
NAND3_X1 _13675_ ( .A1(_05560_ ), .A2(\mepc [25] ), .A3(_05468_ ), .ZN(_05896_ ) );
NAND3_X1 _13676_ ( .A1(_05374_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_05375_ ), .ZN(_05897_ ) );
NAND4_X1 _13677_ ( .A1(_05564_ ), .A2(_05565_ ), .A3(\mtvec [25] ), .A4(_05566_ ), .ZN(_05898_ ) );
NAND4_X1 _13678_ ( .A1(_05408_ ), .A2(_05565_ ), .A3(\mycsreg.CSReg[0][25] ), .A4(_05588_ ), .ZN(_05899_ ) );
AND4_X1 _13679_ ( .A1(_05896_ ), .A2(_05897_ ), .A3(_05898_ ), .A4(_05899_ ), .ZN(_05900_ ) );
OAI21_X1 _13680_ ( .A(_05895_ ), .B1(_05471_ ), .B2(_05900_ ), .ZN(_05901_ ) );
AND3_X1 _13681_ ( .A1(_05313_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05902_ ) );
AND2_X1 _13682_ ( .A1(_05311_ ), .A2(_05902_ ), .ZN(_05903_ ) );
NAND3_X1 _13683_ ( .A1(_05903_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05904_ ) );
INV_X1 _13684_ ( .A(\ID_EX_pc [24] ), .ZN(_05905_ ) );
NOR2_X1 _13685_ ( .A1(_05904_ ), .A2(_05905_ ), .ZN(_05906_ ) );
XNOR2_X1 _13686_ ( .A(_05906_ ), .B(_04077_ ), .ZN(_05907_ ) );
OAI21_X1 _13687_ ( .A(_03978_ ), .B1(_04054_ ), .B2(_04072_ ), .ZN(_05908_ ) );
AND2_X1 _13688_ ( .A1(_05908_ ), .A2(_04075_ ), .ZN(_05909_ ) );
XNOR2_X1 _13689_ ( .A(_05909_ ), .B(_03981_ ), .ZN(_05910_ ) );
MUX2_X1 _13690_ ( .A(_05907_ ), .B(_05910_ ), .S(_05293_ ), .Z(_05911_ ) );
MUX2_X1 _13691_ ( .A(_05901_ ), .B(_05911_ ), .S(_05296_ ), .Z(_05912_ ) );
NAND2_X1 _13692_ ( .A1(_05912_ ), .A2(_05299_ ), .ZN(_05913_ ) );
NOR3_X1 _13693_ ( .A1(_03057_ ), .A2(_05528_ ), .A3(_05362_ ), .ZN(_05914_ ) );
AOI21_X1 _13694_ ( .A(_05914_ ), .B1(_05402_ ), .B2(_05910_ ), .ZN(_05915_ ) );
AOI21_X1 _13695_ ( .A(_05781_ ), .B1(_05913_ ), .B2(_05915_ ), .ZN(_00147_ ) );
XNOR2_X1 _13696_ ( .A(_05904_ ), .B(\ID_EX_pc [24] ), .ZN(_05916_ ) );
XOR2_X1 _13697_ ( .A(_05838_ ), .B(_03978_ ), .Z(_05917_ ) );
MUX2_X1 _13698_ ( .A(_05916_ ), .B(_05917_ ), .S(_05294_ ), .Z(_05918_ ) );
OR2_X1 _13699_ ( .A1(_05918_ ), .A2(\ID_EX_typ [3] ), .ZN(_05919_ ) );
NAND3_X1 _13700_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(\EX_LS_result_csreg_mem [24] ), .ZN(_05920_ ) );
NAND3_X1 _13701_ ( .A1(_05467_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_05561_ ), .ZN(_05921_ ) );
NAND3_X1 _13702_ ( .A1(_05467_ ), .A2(\mepc [24] ), .A3(_05468_ ), .ZN(_05922_ ) );
NAND4_X1 _13703_ ( .A1(_05568_ ), .A2(_05849_ ), .A3(\mycsreg.CSReg[0][24] ), .A4(_05771_ ), .ZN(_05923_ ) );
NAND3_X1 _13704_ ( .A1(_05921_ ), .A2(_05922_ ), .A3(_05923_ ), .ZN(_05924_ ) );
AND4_X1 _13705_ ( .A1(\mtvec [24] ), .A2(_05564_ ), .A3(_05601_ ), .A4(_05566_ ), .ZN(_05925_ ) );
NOR4_X1 _13706_ ( .A1(_05924_ ), .A2(_05348_ ), .A3(_05465_ ), .A4(_05925_ ), .ZN(_05926_ ) );
OAI21_X1 _13707_ ( .A(_05920_ ), .B1(_05926_ ), .B2(_05471_ ), .ZN(_05927_ ) );
OAI211_X1 _13708_ ( .A(_05919_ ), .B(_05363_ ), .C1(_05364_ ), .C2(_05927_ ), .ZN(_05928_ ) );
AOI22_X1 _13709_ ( .A1(_03058_ ), .A2(_05399_ ), .B1(_05401_ ), .B2(_05917_ ), .ZN(_05929_ ) );
AOI21_X1 _13710_ ( .A(_05781_ ), .B1(_05928_ ), .B2(_05929_ ), .ZN(_00148_ ) );
NAND3_X1 _13711_ ( .A1(_05311_ ), .A2(\ID_EX_pc [22] ), .A3(_05902_ ), .ZN(_05930_ ) );
XNOR2_X1 _13712_ ( .A(_05930_ ), .B(\ID_EX_pc [23] ), .ZN(_05931_ ) );
AOI21_X1 _13713_ ( .A(\ID_EX_typ [3] ), .B1(_05306_ ), .B2(_05931_ ), .ZN(_05932_ ) );
NAND3_X1 _13714_ ( .A1(_05460_ ), .A2(\mepc [23] ), .A3(_03945_ ), .ZN(_05933_ ) );
NAND4_X1 _13715_ ( .A1(_05412_ ), .A2(_05587_ ), .A3(\mtvec [23] ), .A4(_05588_ ), .ZN(_05934_ ) );
AND2_X1 _13716_ ( .A1(_05933_ ), .A2(_05934_ ), .ZN(_05935_ ) );
NAND3_X1 _13717_ ( .A1(_05460_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_05405_ ), .ZN(_05936_ ) );
NAND4_X1 _13718_ ( .A1(_05408_ ), .A2(_05413_ ), .A3(\mycsreg.CSReg[0][23] ), .A4(_05588_ ), .ZN(_05937_ ) );
AND2_X1 _13719_ ( .A1(_05936_ ), .A2(_05937_ ), .ZN(_05938_ ) );
AOI22_X1 _13720_ ( .A1(_05935_ ), .A2(_05938_ ), .B1(_05650_ ), .B2(_05456_ ), .ZN(_05939_ ) );
AND3_X1 _13721_ ( .A1(_05333_ ), .A2(_05342_ ), .A3(\EX_LS_result_csreg_mem [23] ), .ZN(_05940_ ) );
NOR2_X1 _13722_ ( .A1(_05939_ ), .A2(_05940_ ), .ZN(_05941_ ) );
AOI211_X1 _13723_ ( .A(_05891_ ), .B(_05932_ ), .C1(\ID_EX_typ [3] ), .C2(_05941_ ), .ZN(_05942_ ) );
INV_X1 _13724_ ( .A(_04041_ ), .ZN(_05943_ ) );
NAND2_X1 _13725_ ( .A1(_05395_ ), .A2(_04046_ ), .ZN(_05944_ ) );
AOI21_X1 _13726_ ( .A(_05943_ ), .B1(_05944_ ), .B2(_04068_ ), .ZN(_05945_ ) );
OR2_X1 _13727_ ( .A1(_05945_ ), .A2(_04070_ ), .ZN(_05946_ ) );
XNOR2_X1 _13728_ ( .A(_05946_ ), .B(_04040_ ), .ZN(_05947_ ) );
INV_X1 _13729_ ( .A(_05940_ ), .ZN(_05948_ ) );
AND4_X1 _13730_ ( .A1(_05933_ ), .A2(_05936_ ), .A3(_05934_ ), .A4(_05937_ ), .ZN(_05949_ ) );
OAI21_X1 _13731_ ( .A(_05948_ ), .B1(_05471_ ), .B2(_05949_ ), .ZN(_05950_ ) );
OAI211_X1 _13732_ ( .A(_05386_ ), .B(_03878_ ), .C1(_05297_ ), .C2(_05950_ ), .ZN(_05951_ ) );
INV_X1 _13733_ ( .A(_05401_ ), .ZN(_05952_ ) );
AOI21_X1 _13734_ ( .A(_05947_ ), .B1(_05951_ ), .B2(_05952_ ), .ZN(_05953_ ) );
NOR2_X1 _13735_ ( .A1(_05942_ ), .A2(_05953_ ), .ZN(_05954_ ) );
OR3_X1 _13736_ ( .A1(_03064_ ), .A2(_05434_ ), .A3(_05362_ ), .ZN(_05955_ ) );
AOI21_X1 _13737_ ( .A(_05781_ ), .B1(_05954_ ), .B2(_05955_ ), .ZN(_00149_ ) );
NAND3_X1 _13738_ ( .A1(_05456_ ), .A2(_05650_ ), .A3(\EX_LS_result_csreg_mem [22] ), .ZN(_05956_ ) );
AND3_X1 _13739_ ( .A1(_03929_ ), .A2(\mepc [22] ), .A3(_03932_ ), .ZN(_05957_ ) );
AND4_X1 _13740_ ( .A1(\mtvec [22] ), .A2(_05367_ ), .A3(_03924_ ), .A4(_05368_ ), .ZN(_05958_ ) );
AND4_X1 _13741_ ( .A1(\mycsreg.CSReg[0][22] ), .A2(_03936_ ), .A3(_05352_ ), .A4(_05368_ ), .ZN(_05959_ ) );
NOR3_X1 _13742_ ( .A1(_05957_ ), .A2(_05958_ ), .A3(_05959_ ), .ZN(_05960_ ) );
NAND3_X1 _13743_ ( .A1(_05560_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_05375_ ), .ZN(_05961_ ) );
AND3_X1 _13744_ ( .A1(_05960_ ), .A2(_05466_ ), .A3(_05961_ ), .ZN(_05962_ ) );
OAI21_X1 _13745_ ( .A(_05956_ ), .B1(_05962_ ), .B2(_05471_ ), .ZN(_05963_ ) );
INV_X1 _13746_ ( .A(\ID_EX_pc [22] ), .ZN(_05964_ ) );
XNOR2_X1 _13747_ ( .A(_05903_ ), .B(_05964_ ), .ZN(_05965_ ) );
AND3_X1 _13748_ ( .A1(_05944_ ), .A2(_05943_ ), .A3(_04068_ ), .ZN(_05966_ ) );
NOR2_X1 _13749_ ( .A1(_05966_ ), .A2(_05945_ ), .ZN(_05967_ ) );
MUX2_X1 _13750_ ( .A(_05965_ ), .B(_05967_ ), .S(_05293_ ), .Z(_05968_ ) );
MUX2_X1 _13751_ ( .A(_05963_ ), .B(_05968_ ), .S(_05296_ ), .Z(_05969_ ) );
NAND2_X1 _13752_ ( .A1(_05969_ ), .A2(_05299_ ), .ZN(_05970_ ) );
AOI22_X1 _13753_ ( .A1(_03065_ ), .A2(_05399_ ), .B1(_05401_ ), .B2(_05967_ ), .ZN(_05971_ ) );
AOI21_X1 _13754_ ( .A(_05781_ ), .B1(_05970_ ), .B2(_05971_ ), .ZN(_00150_ ) );
NOR2_X1 _13755_ ( .A1(_05388_ ), .A2(_05389_ ), .ZN(_05972_ ) );
INV_X1 _13756_ ( .A(\ID_EX_pc [21] ), .ZN(_05973_ ) );
XNOR2_X1 _13757_ ( .A(_05972_ ), .B(_05973_ ), .ZN(_05974_ ) );
NAND2_X1 _13758_ ( .A1(_05395_ ), .A2(_04043_ ), .ZN(_05975_ ) );
NAND2_X1 _13759_ ( .A1(_05975_ ), .A2(_04066_ ), .ZN(_05976_ ) );
XNOR2_X1 _13760_ ( .A(_05976_ ), .B(_04045_ ), .ZN(_05977_ ) );
MUX2_X1 _13761_ ( .A(_05974_ ), .B(_05977_ ), .S(_05294_ ), .Z(_05978_ ) );
OR2_X1 _13762_ ( .A1(_05978_ ), .A2(\ID_EX_typ [3] ), .ZN(_05979_ ) );
NAND3_X1 _13763_ ( .A1(_05404_ ), .A2(\mepc [21] ), .A3(_03932_ ), .ZN(_05980_ ) );
NAND3_X1 _13764_ ( .A1(_05560_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_05375_ ), .ZN(_05981_ ) );
NAND4_X1 _13765_ ( .A1(_05568_ ), .A2(_05601_ ), .A3(\mycsreg.CSReg[0][21] ), .A4(_05566_ ), .ZN(_05982_ ) );
NAND4_X1 _13766_ ( .A1(_05564_ ), .A2(_05565_ ), .A3(\mtvec [21] ), .A4(_05566_ ), .ZN(_05983_ ) );
AND4_X1 _13767_ ( .A1(_05980_ ), .A2(_05981_ ), .A3(_05982_ ), .A4(_05983_ ), .ZN(_05984_ ) );
NAND3_X1 _13768_ ( .A1(_05365_ ), .A2(_05373_ ), .A3(_05984_ ), .ZN(_05985_ ) );
INV_X1 _13769_ ( .A(\EX_LS_result_csreg_mem [21] ), .ZN(_05986_ ) );
NAND3_X1 _13770_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(_05986_ ), .ZN(_05987_ ) );
AND2_X1 _13771_ ( .A1(_05985_ ), .A2(_05987_ ), .ZN(_05988_ ) );
OAI211_X1 _13772_ ( .A(_05979_ ), .B(_05363_ ), .C1(_05364_ ), .C2(_05988_ ), .ZN(_05989_ ) );
NOR3_X1 _13773_ ( .A1(_03019_ ), .A2(_05528_ ), .A3(_05362_ ), .ZN(_05990_ ) );
AOI21_X1 _13774_ ( .A(_05990_ ), .B1(_05402_ ), .B2(_05977_ ), .ZN(_05991_ ) );
AOI21_X1 _13775_ ( .A(_03890_ ), .B1(_05989_ ), .B2(_05991_ ), .ZN(_00151_ ) );
INV_X1 _13776_ ( .A(\ID_EX_pc [30] ), .ZN(_05992_ ) );
NOR2_X1 _13777_ ( .A1(_03972_ ), .A2(_05992_ ), .ZN(_05993_ ) );
INV_X1 _13778_ ( .A(\ID_EX_pc [31] ), .ZN(_05994_ ) );
XNOR2_X1 _13779_ ( .A(_05993_ ), .B(_05994_ ), .ZN(_05995_ ) );
AOI21_X1 _13780_ ( .A(\ID_EX_typ [3] ), .B1(_05306_ ), .B2(_05995_ ), .ZN(_05996_ ) );
NAND3_X1 _13781_ ( .A1(_03929_ ), .A2(\mepc [31] ), .A3(_03932_ ), .ZN(_05997_ ) );
NAND4_X1 _13782_ ( .A1(_05370_ ), .A2(_03924_ ), .A3(\mycsreg.CSReg[0][31] ), .A4(_05368_ ), .ZN(_05998_ ) );
AND2_X1 _13783_ ( .A1(_05997_ ), .A2(_05998_ ), .ZN(_05999_ ) );
NAND3_X1 _13784_ ( .A1(_03928_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_03943_ ), .ZN(_06000_ ) );
NAND4_X1 _13785_ ( .A1(_05367_ ), .A2(_03924_ ), .A3(\mtvec [31] ), .A4(_05368_ ), .ZN(_06001_ ) );
AND2_X1 _13786_ ( .A1(_06000_ ), .A2(_06001_ ), .ZN(_06002_ ) );
AOI22_X1 _13787_ ( .A1(_05999_ ), .A2(_06002_ ), .B1(_05419_ ), .B2(_05418_ ), .ZN(_06003_ ) );
AND3_X1 _13788_ ( .A1(_05333_ ), .A2(_05342_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_06004_ ) );
NOR2_X1 _13789_ ( .A1(_06003_ ), .A2(_06004_ ), .ZN(_06005_ ) );
AOI211_X1 _13790_ ( .A(_03877_ ), .B(_05996_ ), .C1(\ID_EX_typ [3] ), .C2(_06005_ ), .ZN(_06006_ ) );
NOR3_X1 _13791_ ( .A1(_03008_ ), .A2(_05303_ ), .A3(_03878_ ), .ZN(_06007_ ) );
OAI21_X1 _13792_ ( .A(_04087_ ), .B1(_04084_ ), .B2(_04085_ ), .ZN(_06008_ ) );
NAND2_X1 _13793_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_06009_ ) );
NAND2_X1 _13794_ ( .A1(_06008_ ), .A2(_06009_ ), .ZN(_06010_ ) );
XNOR2_X1 _13795_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_06011_ ) );
XOR2_X1 _13796_ ( .A(_06010_ ), .B(_06011_ ), .Z(_06012_ ) );
NAND3_X1 _13797_ ( .A1(_05333_ ), .A2(_05342_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_06013_ ) );
AND4_X1 _13798_ ( .A1(_05997_ ), .A2(_06000_ ), .A3(_05998_ ), .A4(_06001_ ), .ZN(_06014_ ) );
OAI21_X1 _13799_ ( .A(_06013_ ), .B1(_05471_ ), .B2(_06014_ ), .ZN(_06015_ ) );
OAI211_X1 _13800_ ( .A(_05386_ ), .B(_03878_ ), .C1(_05296_ ), .C2(_06015_ ), .ZN(_06016_ ) );
AOI21_X1 _13801_ ( .A(_06012_ ), .B1(_06016_ ), .B2(_05952_ ), .ZN(_06017_ ) );
OR4_X2 _13802_ ( .A1(_03890_ ), .A2(_06006_ ), .A3(_06007_ ), .A4(_06017_ ), .ZN(_00152_ ) );
AND3_X1 _13803_ ( .A1(_03889_ ), .A2(\ID_EX_pc [31] ), .A3(_03100_ ), .ZN(_00153_ ) );
AND3_X1 _13804_ ( .A1(_03889_ ), .A2(\ID_EX_pc [30] ), .A3(_03100_ ), .ZN(_00154_ ) );
AND3_X1 _13805_ ( .A1(_03889_ ), .A2(\ID_EX_pc [21] ), .A3(_03100_ ), .ZN(_00155_ ) );
CLKBUF_X2 _13806_ ( .A(_03099_ ), .Z(_06018_ ) );
AND3_X1 _13807_ ( .A1(_03889_ ), .A2(\ID_EX_pc [20] ), .A3(_06018_ ), .ZN(_00156_ ) );
AND3_X1 _13808_ ( .A1(_03889_ ), .A2(\ID_EX_pc [19] ), .A3(_06018_ ), .ZN(_00157_ ) );
CLKBUF_X2 _13809_ ( .A(_03888_ ), .Z(_06019_ ) );
AND3_X1 _13810_ ( .A1(_06019_ ), .A2(\ID_EX_pc [18] ), .A3(_06018_ ), .ZN(_00158_ ) );
AND3_X1 _13811_ ( .A1(_06019_ ), .A2(\ID_EX_pc [17] ), .A3(_06018_ ), .ZN(_00159_ ) );
AND3_X1 _13812_ ( .A1(_06019_ ), .A2(\ID_EX_pc [16] ), .A3(_06018_ ), .ZN(_00160_ ) );
AND3_X1 _13813_ ( .A1(_06019_ ), .A2(\ID_EX_pc [15] ), .A3(_06018_ ), .ZN(_00161_ ) );
AND3_X1 _13814_ ( .A1(_06019_ ), .A2(\ID_EX_pc [14] ), .A3(_06018_ ), .ZN(_00162_ ) );
AND3_X1 _13815_ ( .A1(_06019_ ), .A2(\ID_EX_pc [13] ), .A3(_06018_ ), .ZN(_00163_ ) );
AND3_X1 _13816_ ( .A1(_06019_ ), .A2(\ID_EX_pc [12] ), .A3(_06018_ ), .ZN(_00164_ ) );
AND3_X1 _13817_ ( .A1(_06019_ ), .A2(\ID_EX_pc [29] ), .A3(_06018_ ), .ZN(_00165_ ) );
CLKBUF_X2 _13818_ ( .A(_03067_ ), .Z(_06020_ ) );
AND3_X1 _13819_ ( .A1(_06019_ ), .A2(\ID_EX_pc [11] ), .A3(_06020_ ), .ZN(_00166_ ) );
AND3_X1 _13820_ ( .A1(_06019_ ), .A2(\ID_EX_pc [10] ), .A3(_06020_ ), .ZN(_00167_ ) );
CLKBUF_X2 _13821_ ( .A(_03888_ ), .Z(_06021_ ) );
AND3_X1 _13822_ ( .A1(_06021_ ), .A2(\ID_EX_pc [9] ), .A3(_06020_ ), .ZN(_00168_ ) );
AND3_X1 _13823_ ( .A1(_06021_ ), .A2(\ID_EX_pc [8] ), .A3(_06020_ ), .ZN(_00169_ ) );
AND3_X1 _13824_ ( .A1(_06021_ ), .A2(\ID_EX_pc [7] ), .A3(_06020_ ), .ZN(_00170_ ) );
AND3_X1 _13825_ ( .A1(_06021_ ), .A2(\ID_EX_pc [6] ), .A3(_06020_ ), .ZN(_00171_ ) );
AND3_X1 _13826_ ( .A1(_06021_ ), .A2(\ID_EX_pc [5] ), .A3(_06020_ ), .ZN(_00172_ ) );
AND3_X1 _13827_ ( .A1(_06021_ ), .A2(\ID_EX_pc [4] ), .A3(_06020_ ), .ZN(_00173_ ) );
AND3_X1 _13828_ ( .A1(_06021_ ), .A2(\ID_EX_pc [3] ), .A3(_06020_ ), .ZN(_00174_ ) );
AND3_X1 _13829_ ( .A1(_06021_ ), .A2(\ID_EX_pc [2] ), .A3(_06020_ ), .ZN(_00175_ ) );
CLKBUF_X2 _13830_ ( .A(_03067_ ), .Z(_06022_ ) );
AND3_X1 _13831_ ( .A1(_06021_ ), .A2(\ID_EX_pc [28] ), .A3(_06022_ ), .ZN(_00176_ ) );
AND3_X1 _13832_ ( .A1(_06021_ ), .A2(\ID_EX_pc [1] ), .A3(_06022_ ), .ZN(_00177_ ) );
CLKBUF_X2 _13833_ ( .A(_03883_ ), .Z(_06023_ ) );
AND3_X1 _13834_ ( .A1(_06023_ ), .A2(\ID_EX_pc [0] ), .A3(_06022_ ), .ZN(_00178_ ) );
AND3_X1 _13835_ ( .A1(_06023_ ), .A2(\ID_EX_pc [27] ), .A3(_06022_ ), .ZN(_00179_ ) );
AND3_X1 _13836_ ( .A1(_06023_ ), .A2(\ID_EX_pc [26] ), .A3(_06022_ ), .ZN(_00180_ ) );
AND3_X1 _13837_ ( .A1(_06023_ ), .A2(\ID_EX_pc [25] ), .A3(_06022_ ), .ZN(_00181_ ) );
AND3_X1 _13838_ ( .A1(_06023_ ), .A2(\ID_EX_pc [24] ), .A3(_06022_ ), .ZN(_00182_ ) );
AND3_X1 _13839_ ( .A1(_06023_ ), .A2(\ID_EX_pc [23] ), .A3(_06022_ ), .ZN(_00183_ ) );
AND3_X1 _13840_ ( .A1(_06023_ ), .A2(\ID_EX_pc [22] ), .A3(_06022_ ), .ZN(_00184_ ) );
AND3_X1 _13841_ ( .A1(_06023_ ), .A2(\ID_EX_typ [7] ), .A3(_06022_ ), .ZN(_00185_ ) );
INV_X1 _13842_ ( .A(io_master_awready ), .ZN(_06024_ ) );
NAND3_X1 _13843_ ( .A1(_03837_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A3(_06024_ ), .ZN(_06025_ ) );
OAI21_X1 _13844_ ( .A(_06025_ ), .B1(\mylsu.state [4] ), .B2(\mylsu.state [0] ), .ZN(_06026_ ) );
OAI21_X1 _13845_ ( .A(_02081_ ), .B1(_03820_ ), .B2(io_master_arready ), .ZN(_06027_ ) );
BUF_X2 _13846_ ( .A(_01973_ ), .Z(_06028_ ) );
INV_X2 _13847_ ( .A(_06028_ ), .ZN(_06029_ ) );
BUF_X2 _13848_ ( .A(_06029_ ), .Z(_06030_ ) );
BUF_X2 _13849_ ( .A(_06030_ ), .Z(_06031_ ) );
BUF_X4 _13850_ ( .A(_06031_ ), .Z(_06032_ ) );
NOR2_X1 _13851_ ( .A1(_06027_ ), .A2(_06032_ ), .ZN(_06033_ ) );
INV_X1 _13852_ ( .A(_06033_ ), .ZN(_06034_ ) );
AOI21_X1 _13853_ ( .A(_06026_ ), .B1(_06034_ ), .B2(_02041_ ), .ZN(_06035_ ) );
AND2_X1 _13854_ ( .A1(_03884_ ), .A2(EXU_valid_LSU ), .ZN(_06036_ ) );
INV_X1 _13855_ ( .A(_06036_ ), .ZN(_06037_ ) );
OAI22_X1 _13856_ ( .A1(_06035_ ), .A2(_06037_ ), .B1(_03886_ ), .B2(_03890_ ), .ZN(_00186_ ) );
AND3_X1 _13857_ ( .A1(_06023_ ), .A2(\ID_EX_typ [6] ), .A3(_03099_ ), .ZN(_00187_ ) );
AND3_X1 _13858_ ( .A1(_06023_ ), .A2(\ID_EX_typ [5] ), .A3(_03099_ ), .ZN(_00188_ ) );
AND3_X1 _13859_ ( .A1(_03888_ ), .A2(\ID_EX_typ [4] ), .A3(_03099_ ), .ZN(_00189_ ) );
AND3_X1 _13860_ ( .A1(_03888_ ), .A2(\ID_EX_typ [3] ), .A3(_03099_ ), .ZN(_00190_ ) );
AND3_X1 _13861_ ( .A1(_03888_ ), .A2(fanout_net_5 ), .A3(_03099_ ), .ZN(_00191_ ) );
AND3_X1 _13862_ ( .A1(_03888_ ), .A2(\ID_EX_typ [1] ), .A3(_03099_ ), .ZN(_00192_ ) );
AND3_X1 _13863_ ( .A1(_03888_ ), .A2(fanout_net_4 ), .A3(_03099_ ), .ZN(_00193_ ) );
AND2_X1 _13864_ ( .A1(_02071_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_06038_ ) );
CLKBUF_X2 _13865_ ( .A(_06038_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _13866_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .ZN(_06039_ ) );
BUF_X2 _13867_ ( .A(_06039_ ), .Z(_06040_ ) );
AND3_X1 _13868_ ( .A1(_02071_ ), .A2(_06040_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00241_ ) );
INV_X1 _13869_ ( .A(fanout_net_11 ), .ZN(_06041_ ) );
BUF_X4 _13870_ ( .A(_06041_ ), .Z(_06042_ ) );
BUF_X4 _13871_ ( .A(_06042_ ), .Z(_06043_ ) );
BUF_X2 _13872_ ( .A(_06043_ ), .Z(_06044_ ) );
AND3_X1 _13873_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06044_ ), .A3(fanout_net_7 ), .ZN(_00242_ ) );
INV_X1 _13874_ ( .A(fanout_net_7 ), .ZN(_06045_ ) );
BUF_X4 _13875_ ( .A(_06045_ ), .Z(_06046_ ) );
BUF_X4 _13876_ ( .A(_06046_ ), .Z(_06047_ ) );
BUF_X2 _13877_ ( .A(_06047_ ), .Z(_06048_ ) );
AND3_X1 _13878_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_11 ), .A3(_06048_ ), .ZN(_00243_ ) );
AND3_X1 _13879_ ( .A1(_03888_ ), .A2(\EX_LS_pc [2] ), .A3(_03099_ ), .ZN(_00281_ ) );
AND2_X1 _13880_ ( .A1(_03885_ ), .A2(\mylsu.state [3] ), .ZN(_00282_ ) );
INV_X1 _13881_ ( .A(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06049_ ) );
AND3_X1 _13882_ ( .A1(_03883_ ), .A2(_06049_ ), .A3(_03067_ ), .ZN(_06050_ ) );
NOR2_X1 _13883_ ( .A1(\mylsu.state [3] ), .A2(\mylsu.state [1] ), .ZN(_06051_ ) );
NAND2_X1 _13884_ ( .A1(_06050_ ), .A2(_06051_ ), .ZN(_06052_ ) );
OAI211_X1 _13885_ ( .A(_02058_ ), .B(_02100_ ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_06053_ ) );
AND2_X1 _13886_ ( .A1(_06053_ ), .A2(\EX_LS_flag [2] ), .ZN(_06054_ ) );
NOR2_X1 _13887_ ( .A1(_02092_ ), .A2(_06054_ ), .ZN(_06055_ ) );
NOR2_X1 _13888_ ( .A1(_03832_ ), .A2(_03841_ ), .ZN(_06056_ ) );
AOI21_X1 _13889_ ( .A(_06052_ ), .B1(_06055_ ), .B2(_06056_ ), .ZN(_00295_ ) );
AOI21_X1 _13890_ ( .A(_02092_ ), .B1(_03898_ ), .B2(_06054_ ), .ZN(_06057_ ) );
AOI21_X1 _13891_ ( .A(_06052_ ), .B1(_06057_ ), .B2(_06056_ ), .ZN(_00296_ ) );
NOR2_X1 _13892_ ( .A1(_02099_ ), .A2(_02101_ ), .ZN(_06058_ ) );
NAND3_X1 _13893_ ( .A1(_06058_ ), .A2(\EX_LS_flag [2] ), .A3(_02001_ ), .ZN(_06059_ ) );
NOR2_X1 _13894_ ( .A1(_06059_ ), .A2(_06052_ ), .ZN(_00297_ ) );
AOI21_X1 _13895_ ( .A(_06052_ ), .B1(_03834_ ), .B2(_02057_ ), .ZN(_00298_ ) );
AOI21_X1 _13896_ ( .A(_06052_ ), .B1(_06056_ ), .B2(_06059_ ), .ZN(_00299_ ) );
NAND3_X1 _13897_ ( .A1(_03885_ ), .A2(EXU_valid_LSU ), .A3(_06051_ ), .ZN(_06060_ ) );
OR3_X1 _13898_ ( .A1(_02067_ ), .A2(_03841_ ), .A3(_06060_ ), .ZN(_06061_ ) );
NOR3_X1 _13899_ ( .A1(_02101_ ), .A2(_03837_ ), .A3(_02025_ ), .ZN(_06062_ ) );
OAI21_X1 _13900_ ( .A(_06062_ ), .B1(_02099_ ), .B2(\EX_LS_flag [1] ), .ZN(_06063_ ) );
NOR2_X1 _13901_ ( .A1(_06033_ ), .A2(_06063_ ), .ZN(_06064_ ) );
OAI211_X1 _13902_ ( .A(_02041_ ), .B(_02056_ ), .C1(_06064_ ), .C2(_02040_ ), .ZN(_06065_ ) );
INV_X1 _13903_ ( .A(_02061_ ), .ZN(_06066_ ) );
AND2_X1 _13904_ ( .A1(_06066_ ), .A2(_06063_ ), .ZN(_06067_ ) );
AOI21_X1 _13905_ ( .A(_06061_ ), .B1(_06065_ ), .B2(_06067_ ), .ZN(_00300_ ) );
INV_X1 _13906_ ( .A(_00282_ ), .ZN(_06068_ ) );
NAND3_X1 _13907_ ( .A1(_06066_ ), .A2(EXU_valid_LSU ), .A3(_06051_ ), .ZN(_06069_ ) );
OAI21_X1 _13908_ ( .A(_03885_ ), .B1(_03835_ ), .B2(_02125_ ), .ZN(_06070_ ) );
OAI21_X1 _13909_ ( .A(_06068_ ), .B1(_06069_ ), .B2(_06070_ ), .ZN(_00301_ ) );
BUF_X2 _13910_ ( .A(_02035_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _13911_ ( .A(_01975_ ), .Z(_06071_ ) );
NOR3_X1 _13912_ ( .A1(_06071_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06072_ ) );
BUF_X4 _13913_ ( .A(_06032_ ), .Z(_06073_ ) );
INV_X1 _13914_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06074_ ) );
INV_X1 _13915_ ( .A(_01978_ ), .ZN(_06075_ ) );
AOI211_X1 _13916_ ( .A(_06072_ ), .B(_06073_ ), .C1(_06074_ ), .C2(_06075_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _13917_ ( .A1(_06071_ ), .A2(fanout_net_3 ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06076_ ) );
INV_X1 _13918_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06077_ ) );
AOI211_X1 _13919_ ( .A(_06076_ ), .B(_06073_ ), .C1(_06077_ ), .C2(_06075_ ), .ZN(\io_master_araddr [0] ) );
OR3_X1 _13920_ ( .A1(_06071_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06078_ ) );
BUF_X4 _13921_ ( .A(_01978_ ), .Z(_06079_ ) );
OAI21_X1 _13922_ ( .A(_06078_ ), .B1(_06079_ ), .B2(\mylsu.araddr_tmp [15] ), .ZN(_06080_ ) );
BUF_X4 _13923_ ( .A(_01982_ ), .Z(_06081_ ) );
BUF_X4 _13924_ ( .A(_06081_ ), .Z(_06082_ ) );
BUF_X4 _13925_ ( .A(_06082_ ), .Z(_06083_ ) );
OAI22_X1 _13926_ ( .A1(_06073_ ), .A2(_06080_ ), .B1(_03479_ ), .B2(_06083_ ), .ZN(\io_master_araddr [15] ) );
OAI221_X1 _13927_ ( .A(\IF_ID_pc [14] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01962_ ), .C2(_01963_ ), .ZN(_06084_ ) );
INV_X1 _13928_ ( .A(_01971_ ), .ZN(_06085_ ) );
OR3_X1 _13929_ ( .A1(_06071_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06086_ ) );
OAI211_X1 _13930_ ( .A(_06085_ ), .B(_06086_ ), .C1(\mylsu.araddr_tmp [14] ), .C2(_06079_ ), .ZN(_06087_ ) );
OAI21_X1 _13931_ ( .A(_06084_ ), .B1(\io_master_arburst [0] ), .B2(_06087_ ), .ZN(\io_master_araddr [14] ) );
NOR3_X1 _13932_ ( .A1(_06071_ ), .A2(_05334_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06088_ ) );
AOI21_X1 _13933_ ( .A(_06088_ ), .B1(_06075_ ), .B2(\mylsu.araddr_tmp [5] ), .ZN(_06089_ ) );
BUF_X2 _13934_ ( .A(_06081_ ), .Z(_06090_ ) );
OAI22_X1 _13935_ ( .A1(_06073_ ), .A2(_06089_ ), .B1(_03527_ ), .B2(_06090_ ), .ZN(\io_master_araddr [5] ) );
OAI221_X1 _13936_ ( .A(fanout_net_11 ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01962_ ), .C2(_01963_ ), .ZN(_06091_ ) );
OR3_X1 _13937_ ( .A1(_06071_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06092_ ) );
OAI211_X1 _13938_ ( .A(_06085_ ), .B(_06092_ ), .C1(\mylsu.araddr_tmp [4] ), .C2(_06079_ ), .ZN(_06093_ ) );
OAI21_X1 _13939_ ( .A(_06091_ ), .B1(\io_master_arburst [0] ), .B2(_06093_ ), .ZN(\io_master_araddr [4] ) );
NAND4_X1 _13940_ ( .A1(_01999_ ), .A2(_03907_ ), .A3(_02001_ ), .A4(_02025_ ), .ZN(_06094_ ) );
OAI21_X1 _13941_ ( .A(_06094_ ), .B1(_06079_ ), .B2(\mylsu.araddr_tmp [3] ), .ZN(_06095_ ) );
OAI22_X1 _13942_ ( .A1(_06073_ ), .A2(_06095_ ), .B1(_06048_ ), .B2(_06090_ ), .ZN(\io_master_araddr [3] ) );
OAI221_X1 _13943_ ( .A(\IF_ID_pc [13] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01962_ ), .C2(_01963_ ), .ZN(_06096_ ) );
OR3_X1 _13944_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06097_ ) );
OAI211_X1 _13945_ ( .A(_06085_ ), .B(_06097_ ), .C1(\mylsu.araddr_tmp [13] ), .C2(_06079_ ), .ZN(_06098_ ) );
OAI21_X1 _13946_ ( .A(_06096_ ), .B1(\io_master_arburst [0] ), .B2(_06098_ ), .ZN(\io_master_araddr [13] ) );
OAI221_X1 _13947_ ( .A(\IF_ID_pc [12] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01962_ ), .C2(_01963_ ), .ZN(_06099_ ) );
OR3_X1 _13948_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06100_ ) );
OAI211_X1 _13949_ ( .A(_06085_ ), .B(_06100_ ), .C1(\mylsu.araddr_tmp [12] ), .C2(_01978_ ), .ZN(_06101_ ) );
OAI21_X1 _13950_ ( .A(_06099_ ), .B1(\io_master_arburst [0] ), .B2(_06101_ ), .ZN(\io_master_araddr [12] ) );
OR3_X1 _13951_ ( .A1(_06071_ ), .A2(\EX_LS_dest_csreg_mem [11] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06102_ ) );
OAI21_X1 _13952_ ( .A(_06102_ ), .B1(_06079_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_06103_ ) );
OAI22_X1 _13953_ ( .A1(_06073_ ), .A2(_06103_ ), .B1(_01923_ ), .B2(_06090_ ), .ZN(\io_master_araddr [11] ) );
OR3_X1 _13954_ ( .A1(_06071_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06104_ ) );
OAI21_X1 _13955_ ( .A(_06104_ ), .B1(_06079_ ), .B2(\mylsu.araddr_tmp [10] ), .ZN(_06105_ ) );
OAI22_X1 _13956_ ( .A1(_06073_ ), .A2(_06105_ ), .B1(_01863_ ), .B2(_06090_ ), .ZN(\io_master_araddr [10] ) );
NAND4_X1 _13957_ ( .A1(_01999_ ), .A2(_05327_ ), .A3(_02001_ ), .A4(_02025_ ), .ZN(_06106_ ) );
OAI21_X1 _13958_ ( .A(_06106_ ), .B1(_06079_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06107_ ) );
OAI22_X1 _13959_ ( .A1(_06073_ ), .A2(_06107_ ), .B1(_01870_ ), .B2(_06090_ ), .ZN(\io_master_araddr [9] ) );
OR3_X1 _13960_ ( .A1(_06071_ ), .A2(\EX_LS_dest_csreg_mem [8] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06108_ ) );
OAI21_X1 _13961_ ( .A(_06108_ ), .B1(_06079_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_06109_ ) );
OAI22_X1 _13962_ ( .A1(_06073_ ), .A2(_06109_ ), .B1(_01810_ ), .B2(_06090_ ), .ZN(\io_master_araddr [8] ) );
NOR3_X1 _13963_ ( .A1(_06071_ ), .A2(_05328_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06110_ ) );
AOI21_X1 _13964_ ( .A(_06110_ ), .B1(_06075_ ), .B2(\mylsu.araddr_tmp [7] ), .ZN(_06111_ ) );
OAI22_X1 _13965_ ( .A1(_06073_ ), .A2(_06111_ ), .B1(_01789_ ), .B2(_06090_ ), .ZN(\io_master_araddr [7] ) );
OAI221_X1 _13966_ ( .A(\IF_ID_pc [6] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01962_ ), .C2(_01963_ ), .ZN(_06112_ ) );
OR3_X1 _13967_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [6] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06113_ ) );
OAI211_X1 _13968_ ( .A(_06085_ ), .B(_06113_ ), .C1(\mylsu.araddr_tmp [6] ), .C2(_01978_ ), .ZN(_06114_ ) );
OAI21_X1 _13969_ ( .A(_06112_ ), .B1(\io_master_arburst [0] ), .B2(_06114_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _13970_ ( .A1(_01975_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06115_ ) );
OAI211_X1 _13971_ ( .A(_06085_ ), .B(_06115_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01978_ ), .ZN(_06116_ ) );
NOR2_X1 _13972_ ( .A1(_01966_ ), .A2(_06116_ ), .ZN(_06117_ ) );
BUF_X4 _13973_ ( .A(_06117_ ), .Z(_06118_ ) );
BUF_X4 _13974_ ( .A(_06118_ ), .Z(_06119_ ) );
BUF_X2 _13975_ ( .A(_06119_ ), .Z(\io_master_araddr [2] ) );
CLKBUF_X2 _13976_ ( .A(_06028_ ), .Z(\io_master_arid [1] ) );
AND3_X1 _13977_ ( .A1(_06090_ ), .A2(\EX_LS_typ [3] ), .A3(_06085_ ), .ZN(\io_master_arsize [2] ) );
INV_X1 _13978_ ( .A(\EX_LS_typ [1] ), .ZN(_06120_ ) );
NOR3_X1 _13979_ ( .A1(\io_master_arburst [0] ), .A2(_06120_ ), .A3(_01971_ ), .ZN(\io_master_arsize [0] ) );
OAI21_X1 _13980_ ( .A(\EX_LS_typ [2] ), .B1(_06079_ ), .B2(_01970_ ), .ZN(_06121_ ) );
OAI21_X1 _13981_ ( .A(_06121_ ), .B1(_01964_ ), .B2(_01965_ ), .ZN(\io_master_arsize [1] ) );
BUF_X2 _13982_ ( .A(_02077_ ), .Z(_06122_ ) );
BUF_X2 _13983_ ( .A(_02080_ ), .Z(_06123_ ) );
AOI211_X1 _13984_ ( .A(_02070_ ), .B(_02072_ ), .C1(_06122_ ), .C2(_06123_ ), .ZN(io_master_arvalid ) );
BUF_X2 _13985_ ( .A(_02060_ ), .Z(_06124_ ) );
AND2_X1 _13986_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ) );
AND2_X1 _13987_ ( .A1(_06124_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_06125_ ) );
BUF_X4 _13988_ ( .A(_06125_ ), .Z(_06126_ ) );
BUF_X4 _13989_ ( .A(_06126_ ), .Z(_06127_ ) );
MUX2_X1 _13990_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06127_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _13991_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06127_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _13992_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06127_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _13993_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06127_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _13994_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06127_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _13995_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06127_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _13996_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06127_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _13997_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06127_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _13998_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06127_ ), .Z(\io_master_awaddr [15] ) );
MUX2_X1 _13999_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06127_ ), .Z(\io_master_awaddr [14] ) );
BUF_X4 _14000_ ( .A(_06126_ ), .Z(_06128_ ) );
MUX2_X1 _14001_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06128_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _14002_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06128_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _14003_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06128_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _14004_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06128_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _14005_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06128_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _14006_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06128_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _14007_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06128_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _14008_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06128_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _14009_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06128_ ), .Z(\io_master_awaddr [6] ) );
MUX2_X1 _14010_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06128_ ), .Z(\io_master_awaddr [5] ) );
BUF_X4 _14011_ ( .A(_06126_ ), .Z(_06129_ ) );
MUX2_X1 _14012_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06129_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _14013_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06129_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _14014_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06129_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _14015_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06129_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _14016_ ( .A(\mylsu.awaddr_tmp [1] ), .B(\EX_LS_dest_csreg_mem [1] ), .S(_06129_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _14017_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_3 ), .S(_06129_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _14018_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06129_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _14019_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06129_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _14020_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06129_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _14021_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06129_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _14022_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06126_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _14023_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06126_ ), .Z(\io_master_awaddr [22] ) );
NOR4_X1 _14024_ ( .A1(_03898_ ), .A2(_02050_ ), .A3(_02062_ ), .A4(_06120_ ), .ZN(\io_master_awsize [0] ) );
NAND2_X1 _14025_ ( .A1(_02063_ ), .A2(_02049_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _14026_ ( .A1(_02057_ ), .A2(_02068_ ), .A3(_06126_ ), .ZN(_06130_ ) );
INV_X1 _14027_ ( .A(\mylsu.state [4] ), .ZN(_06131_ ) );
NAND2_X1 _14028_ ( .A1(_06130_ ), .A2(_06131_ ), .ZN(io_master_awvalid ) );
OR3_X1 _14029_ ( .A1(io_master_awvalid ), .A2(\mylsu.state [2] ), .A3(\mylsu.state [1] ), .ZN(io_master_bready ) );
NOR3_X1 _14030_ ( .A1(_01970_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_06132_ ) );
INV_X1 _14031_ ( .A(\io_master_bid [2] ), .ZN(_06133_ ) );
INV_X1 _14032_ ( .A(\io_master_bresp [0] ), .ZN(_06134_ ) );
AND4_X1 _14033_ ( .A1(\io_master_bid [1] ), .A2(_06133_ ), .A3(_06134_ ), .A4(io_master_bvalid ), .ZN(_06135_ ) );
INV_X1 _14034_ ( .A(\io_master_bid [0] ), .ZN(_06136_ ) );
NOR3_X1 _14035_ ( .A1(_06136_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bresp [1] ), .ZN(_06137_ ) );
NAND2_X1 _14036_ ( .A1(_06135_ ), .A2(_06137_ ), .ZN(_06138_ ) );
NOR3_X1 _14037_ ( .A1(_02006_ ), .A2(_06031_ ), .A3(_02031_ ), .ZN(_06139_ ) );
NOR2_X1 _14038_ ( .A1(_03814_ ), .A2(\io_master_rid [0] ), .ZN(_06140_ ) );
AND2_X1 _14039_ ( .A1(_06140_ ), .A2(io_master_rlast ), .ZN(_06141_ ) );
AND4_X1 _14040_ ( .A1(\io_master_arid [1] ), .A2(_03812_ ), .A3(_03813_ ), .A4(_06141_ ), .ZN(_06142_ ) );
OAI21_X1 _14041_ ( .A(_03825_ ), .B1(_06139_ ), .B2(_06142_ ), .ZN(_06143_ ) );
AOI221_X4 _14042_ ( .A(_06132_ ), .B1(\mylsu.state [1] ), .B2(_06138_ ), .C1(_06143_ ), .C2(\mylsu.state [3] ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _14043_ ( .A(_02082_ ), .B(_02084_ ), .C1(_06122_ ), .C2(_06123_ ), .ZN(io_master_rready ) );
MUX2_X1 _14044_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_3 ), .Z(_06144_ ) );
CLKBUF_X2 _14045_ ( .A(_05338_ ), .Z(_06145_ ) );
AND2_X1 _14046_ ( .A1(_06144_ ), .A2(_06145_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _14047_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_3 ), .Z(_06146_ ) );
AND2_X1 _14048_ ( .A1(_06146_ ), .A2(_06145_ ), .ZN(\io_master_wdata [14] ) );
INV_X1 _14049_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_06147_ ) );
NOR3_X1 _14050_ ( .A1(_06147_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _14051_ ( .A1(_05768_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [4] ) );
NOR3_X1 _14052_ ( .A1(_05788_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14053_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_06148_ ) );
NOR3_X1 _14054_ ( .A1(_06148_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14055_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06149_ ) );
NOR3_X1 _14056_ ( .A1(_06149_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14057_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06150_ ) );
NOR3_X1 _14058_ ( .A1(_06150_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14059_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_3 ), .Z(_06151_ ) );
AND2_X1 _14060_ ( .A1(_06151_ ), .A2(_06145_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14061_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_3 ), .Z(_06152_ ) );
AND2_X1 _14062_ ( .A1(_06152_ ), .A2(_06145_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14063_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_3 ), .Z(_06153_ ) );
AND2_X1 _14064_ ( .A1(_06153_ ), .A2(_06145_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14065_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_3 ), .Z(_06154_ ) );
AND2_X1 _14066_ ( .A1(_06154_ ), .A2(_06145_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14067_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_3 ), .Z(_06155_ ) );
AND2_X1 _14068_ ( .A1(_06155_ ), .A2(_06145_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14069_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_3 ), .Z(_06156_ ) );
AND2_X1 _14070_ ( .A1(_06156_ ), .A2(_06145_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14071_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06157_ ) );
NOR3_X1 _14072_ ( .A1(_06157_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [7] ) );
NOR3_X1 _14073_ ( .A1(_05720_ ), .A2(fanout_net_3 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14074_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_3 ), .Z(_06158_ ) );
MUX2_X1 _14075_ ( .A(_06158_ ), .B(_06144_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14076_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_3 ), .Z(_06159_ ) );
MUX2_X1 _14077_ ( .A(_06159_ ), .B(_06146_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [30] ) );
MUX2_X1 _14078_ ( .A(_05986_ ), .B(_05557_ ), .S(fanout_net_3 ), .Z(_06160_ ) );
NOR2_X1 _14079_ ( .A1(_05338_ ), .A2(fanout_net_3 ), .ZN(_06161_ ) );
INV_X1 _14080_ ( .A(_06161_ ), .ZN(_06162_ ) );
OAI22_X1 _14081_ ( .A1(_06160_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06162_ ), .B2(_06147_ ), .ZN(\io_master_wdata [21] ) );
INV_X1 _14082_ ( .A(\EX_LS_result_csreg_mem [20] ), .ZN(_06163_ ) );
INV_X1 _14083_ ( .A(\EX_LS_result_csreg_mem [12] ), .ZN(_06164_ ) );
MUX2_X1 _14084_ ( .A(_06163_ ), .B(_06164_ ), .S(fanout_net_3 ), .Z(_06165_ ) );
OAI22_X1 _14085_ ( .A1(_06165_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06162_ ), .B2(_05768_ ), .ZN(\io_master_wdata [20] ) );
INV_X1 _14086_ ( .A(fanout_net_3 ), .ZN(_06166_ ) );
OAI21_X1 _14087_ ( .A(_05338_ ), .B1(_06166_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_06167_ ) );
NOR2_X1 _14088_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_06168_ ) );
OAI22_X1 _14089_ ( .A1(_06162_ ), .A2(_05788_ ), .B1(_06167_ ), .B2(_06168_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _14090_ ( .A(_05338_ ), .B1(_06166_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_06169_ ) );
NOR2_X1 _14091_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_06170_ ) );
OAI22_X1 _14092_ ( .A1(_06162_ ), .A2(_06148_ ), .B1(_06169_ ), .B2(_06170_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _14093_ ( .A(_05338_ ), .B1(_06166_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_06171_ ) );
NOR2_X1 _14094_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_06172_ ) );
OAI22_X1 _14095_ ( .A1(_06162_ ), .A2(_06149_ ), .B1(_06171_ ), .B2(_06172_ ), .ZN(\io_master_wdata [17] ) );
OAI21_X1 _14096_ ( .A(_05338_ ), .B1(_06166_ ), .B2(\EX_LS_result_csreg_mem [8] ), .ZN(_06173_ ) );
NOR2_X1 _14097_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [16] ), .ZN(_06174_ ) );
OAI22_X1 _14098_ ( .A1(_06162_ ), .A2(_06150_ ), .B1(_06173_ ), .B2(_06174_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14099_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06175_ ) );
MUX2_X1 _14100_ ( .A(_06175_ ), .B(_06151_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14101_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06176_ ) );
MUX2_X1 _14102_ ( .A(_06176_ ), .B(_06152_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14103_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06177_ ) );
MUX2_X1 _14104_ ( .A(_06177_ ), .B(_06153_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14105_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06178_ ) );
MUX2_X1 _14106_ ( .A(_06178_ ), .B(_06154_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14107_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06179_ ) );
MUX2_X1 _14108_ ( .A(_06179_ ), .B(_06155_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14109_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06180_ ) );
MUX2_X1 _14110_ ( .A(_06180_ ), .B(_06156_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [24] ) );
OAI21_X1 _14111_ ( .A(_05338_ ), .B1(_06166_ ), .B2(\EX_LS_result_csreg_mem [15] ), .ZN(_06181_ ) );
NOR2_X1 _14112_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [23] ), .ZN(_06182_ ) );
OAI22_X1 _14113_ ( .A1(_06162_ ), .A2(_06157_ ), .B1(_06181_ ), .B2(_06182_ ), .ZN(\io_master_wdata [23] ) );
OAI21_X1 _14114_ ( .A(_05338_ ), .B1(_06166_ ), .B2(\EX_LS_result_csreg_mem [14] ), .ZN(_06183_ ) );
NOR2_X1 _14115_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [22] ), .ZN(_06184_ ) );
OAI22_X1 _14116_ ( .A1(_06162_ ), .A2(_05720_ ), .B1(_06183_ ), .B2(_06184_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14117_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06185_ ) );
AND2_X1 _14118_ ( .A1(_06185_ ), .A2(_06145_ ), .ZN(\io_master_wstrb [1] ) );
NOR3_X1 _14119_ ( .A1(_02046_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14120_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06186_ ) );
MUX2_X1 _14121_ ( .A(_06186_ ), .B(_06185_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14122_ ( .A1(_06166_ ), .A2(_06145_ ), .A3(\EX_LS_typ [2] ), .ZN(_06187_ ) );
OAI221_X1 _14123_ ( .A(_06187_ ), .B1(_02052_ ), .B2(\EX_LS_dest_csreg_mem [1] ), .C1(_06162_ ), .C2(_02046_ ), .ZN(\io_master_wstrb [2] ) );
INV_X1 _14124_ ( .A(\mylsu.state [2] ), .ZN(_06188_ ) );
NAND2_X1 _14125_ ( .A1(_06130_ ), .A2(_06188_ ), .ZN(io_master_wvalid ) );
NOR4_X1 _14126_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .A3(\LS_WB_waddr_csreg [5] ), .A4(\LS_WB_waddr_csreg [4] ), .ZN(_06189_ ) );
NOR2_X1 _14127_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06190_ ) );
AND2_X1 _14128_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06191_ ) );
NAND3_X1 _14129_ ( .A1(_06189_ ), .A2(_06190_ ), .A3(_06191_ ), .ZN(_06192_ ) );
NOR2_X1 _14130_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_06193_ ) );
NAND3_X1 _14131_ ( .A1(_06193_ ), .A2(_01559_ ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_06194_ ) );
NOR4_X1 _14132_ ( .A1(_06192_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(\LS_WB_waddr_csreg [1] ), .A4(_06194_ ), .ZN(\mycsreg.CSReg[0]_$_DFFE_PP__Q_E ) );
INV_X1 _14133_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_06195_ ) );
NOR2_X1 _14134_ ( .A1(_06195_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_06196_ ) );
INV_X1 _14135_ ( .A(_06196_ ), .ZN(_06197_ ) );
INV_X1 _14136_ ( .A(\LS_WB_waddr_csreg [3] ), .ZN(_06198_ ) );
NAND4_X1 _14137_ ( .A1(_01559_ ), .A2(_06198_ ), .A3(\LS_WB_waddr_csreg [2] ), .A4(\LS_WB_wen_csreg [7] ), .ZN(_06199_ ) );
NOR3_X1 _14138_ ( .A1(_06192_ ), .A2(_06197_ ), .A3(_06199_ ), .ZN(\mycsreg.CSReg[1]_$_DFFE_PP__Q_E ) );
NOR2_X1 _14139_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06200_ ) );
NAND2_X1 _14140_ ( .A1(_06200_ ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06201_ ) );
NOR2_X1 _14141_ ( .A1(_06201_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06202_ ) );
NAND3_X1 _14142_ ( .A1(_06202_ ), .A2(_06190_ ), .A3(_06191_ ), .ZN(_06203_ ) );
NOR3_X1 _14143_ ( .A1(_06203_ ), .A2(_06194_ ), .A3(_06197_ ), .ZN(\mycsreg.CSReg[2]_$_DFFE_PP__Q_E ) );
MUX2_X1 _14144_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14145_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14146_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14147_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
AND3_X1 _14148_ ( .A1(_06193_ ), .A2(_06195_ ), .A3(\LS_WB_waddr_csreg [1] ), .ZN(_06204_ ) );
NAND4_X1 _14149_ ( .A1(_06202_ ), .A2(_06190_ ), .A3(_06191_ ), .A4(_06204_ ), .ZN(_06205_ ) );
AOI21_X1 _14150_ ( .A(reset ), .B1(_06205_ ), .B2(_02087_ ), .ZN(_06206_ ) );
AND2_X1 _14151_ ( .A1(_06206_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(\mycsreg.CSReg[3]_$_DFFE_PP__Q_E ) );
AND2_X1 _14152_ ( .A1(\LS_WB_wen_csreg [6] ), .A2(\LS_WB_wen_csreg [7] ), .ZN(\mycsreg.excp_written_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14153_ ( .A(_02069_ ), .ZN(_06207_ ) );
NOR2_X1 _14154_ ( .A1(_06058_ ), .A2(exception_quest_IDU ), .ZN(_06208_ ) );
NOR2_X1 _14155_ ( .A1(_06207_ ), .A2(_06208_ ), .ZN(_06209_ ) );
BUF_X4 _14156_ ( .A(_06209_ ), .Z(_06210_ ) );
MUX2_X1 _14157_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14158_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14159_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14160_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14161_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14162_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14163_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14164_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14165_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14166_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_06210_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14167_ ( .A(_06209_ ), .Z(_06211_ ) );
MUX2_X1 _14168_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14169_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14170_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14171_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14172_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14173_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14174_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14175_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14176_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14177_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_06211_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14178_ ( .A(_06209_ ), .Z(_06212_ ) );
MUX2_X1 _14179_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14180_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14181_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14182_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14183_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14184_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14185_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14186_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14187_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14188_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_06212_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14189_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_06209_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14190_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_06209_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
INV_X1 _14191_ ( .A(_02094_ ), .ZN(_06213_ ) );
NOR4_X1 _14192_ ( .A1(_06207_ ), .A2(exception_quest_IDU ), .A3(_06213_ ), .A4(_06208_ ), .ZN(_06214_ ) );
XNOR2_X1 _14193_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06215_ ) );
XNOR2_X1 _14194_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06216_ ) );
XNOR2_X1 _14195_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06217_ ) );
XNOR2_X1 _14196_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06218_ ) );
NAND4_X1 _14197_ ( .A1(_06215_ ), .A2(_06216_ ), .A3(_06217_ ), .A4(_06218_ ), .ZN(_06219_ ) );
XNOR2_X1 _14198_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_06220_ ) );
XNOR2_X1 _14199_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_06221_ ) );
NAND2_X1 _14200_ ( .A1(_06220_ ), .A2(_06221_ ), .ZN(_06222_ ) );
XOR2_X1 _14201_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .Z(_06223_ ) );
XOR2_X1 _14202_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .Z(_06224_ ) );
NOR4_X1 _14203_ ( .A1(_06219_ ), .A2(_06222_ ), .A3(_06223_ ), .A4(_06224_ ), .ZN(_06225_ ) );
XNOR2_X1 _14204_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06226_ ) );
XNOR2_X1 _14205_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06227_ ) );
XNOR2_X1 _14206_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06228_ ) );
XNOR2_X1 _14207_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06229_ ) );
AND4_X1 _14208_ ( .A1(_06226_ ), .A2(_06227_ ), .A3(_06228_ ), .A4(_06229_ ), .ZN(_06230_ ) );
XNOR2_X1 _14209_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06231_ ) );
XNOR2_X1 _14210_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06232_ ) );
XNOR2_X1 _14211_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06233_ ) );
XNOR2_X1 _14212_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06234_ ) );
AND4_X1 _14213_ ( .A1(_06231_ ), .A2(_06232_ ), .A3(_06233_ ), .A4(_06234_ ), .ZN(_06235_ ) );
AND3_X1 _14214_ ( .A1(_06225_ ), .A2(_06230_ ), .A3(_06235_ ), .ZN(_06236_ ) );
XNOR2_X1 _14215_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06237_ ) );
XNOR2_X1 _14216_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06238_ ) );
XNOR2_X1 _14217_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06239_ ) );
XNOR2_X1 _14218_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06240_ ) );
NAND4_X1 _14219_ ( .A1(_06237_ ), .A2(_06238_ ), .A3(_06239_ ), .A4(_06240_ ), .ZN(_06241_ ) );
XNOR2_X1 _14220_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06242_ ) );
XNOR2_X1 _14221_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06243_ ) );
XNOR2_X1 _14222_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06244_ ) );
XNOR2_X1 _14223_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06245_ ) );
NAND4_X1 _14224_ ( .A1(_06242_ ), .A2(_06243_ ), .A3(_06244_ ), .A4(_06245_ ), .ZN(_06246_ ) );
XNOR2_X1 _14225_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06247_ ) );
XNOR2_X1 _14226_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06248_ ) );
XNOR2_X1 _14227_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06249_ ) );
XNOR2_X1 _14228_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06250_ ) );
NAND4_X1 _14229_ ( .A1(_06247_ ), .A2(_06248_ ), .A3(_06249_ ), .A4(_06250_ ), .ZN(_06251_ ) );
XNOR2_X1 _14230_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06252_ ) );
XNOR2_X1 _14231_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06253_ ) );
XNOR2_X1 _14232_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06254_ ) );
XNOR2_X1 _14233_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06255_ ) );
NAND4_X1 _14234_ ( .A1(_06252_ ), .A2(_06253_ ), .A3(_06254_ ), .A4(_06255_ ), .ZN(_06256_ ) );
NOR4_X1 _14235_ ( .A1(_06241_ ), .A2(_06246_ ), .A3(_06251_ ), .A4(_06256_ ), .ZN(_06257_ ) );
NAND3_X1 _14236_ ( .A1(_06236_ ), .A2(excp_written ), .A3(_06257_ ), .ZN(_06258_ ) );
AOI21_X1 _14237_ ( .A(_06214_ ), .B1(_06213_ ), .B2(_06258_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _14238_ ( .A1(\ID_EX_typ [7] ), .A2(_03872_ ), .A3(_01998_ ), .A4(IDU_valid_EXU ), .ZN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _14239_ ( .A1(_05833_ ), .A2(_03013_ ), .ZN(_06259_ ) );
AND2_X2 _14240_ ( .A1(_03009_ ), .A2(_03875_ ), .ZN(_06260_ ) );
INV_X1 _14241_ ( .A(_06260_ ), .ZN(_06261_ ) );
BUF_X2 _14242_ ( .A(_06261_ ), .Z(_06262_ ) );
BUF_X4 _14243_ ( .A(_06262_ ), .Z(_06263_ ) );
OAI21_X1 _14244_ ( .A(_06259_ ), .B1(_03915_ ), .B2(_06263_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _14245_ ( .A(_02502_ ), .B(\ID_EX_imm [0] ), .ZN(_06264_ ) );
BUF_X4 _14246_ ( .A(_06260_ ), .Z(_06265_ ) );
BUF_X4 _14247_ ( .A(_06265_ ), .Z(_06266_ ) );
AOI22_X1 _14248_ ( .A1(_06264_ ), .A2(_03014_ ), .B1(_03935_ ), .B2(_06266_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND2_X1 _14249_ ( .A1(_03353_ ), .A2(\ID_EX_typ [7] ), .ZN(_06267_ ) );
BUF_X4 _14250_ ( .A(_06267_ ), .Z(_06268_ ) );
INV_X1 _14251_ ( .A(_06268_ ), .ZN(_06269_ ) );
BUF_X4 _14252_ ( .A(_06269_ ), .Z(_06270_ ) );
AND2_X1 _14253_ ( .A1(_05656_ ), .A2(_06270_ ), .ZN(_06271_ ) );
BUF_X4 _14254_ ( .A(_06261_ ), .Z(_06272_ ) );
MUX2_X1 _14255_ ( .A(\ID_EX_csr [10] ), .B(_06271_ ), .S(_06272_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
NOR4_X1 _14256_ ( .A1(_03348_ ), .A2(_03872_ ), .A3(\ID_EX_typ [5] ), .A4(\ID_EX_csr [9] ), .ZN(_06273_ ) );
AOI21_X1 _14257_ ( .A(_06273_ ), .B1(_05677_ ), .B2(_03014_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR2_X1 _14258_ ( .A1(_05695_ ), .A2(_06268_ ), .ZN(_06274_ ) );
MUX2_X1 _14259_ ( .A(\ID_EX_csr [8] ), .B(_06274_ ), .S(_06272_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _14260_ ( .A1(_05718_ ), .A2(_03013_ ), .ZN(_06275_ ) );
OAI21_X1 _14261_ ( .A(_06275_ ), .B1(_03926_ ), .B2(_06263_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
OR2_X1 _14262_ ( .A1(_05735_ ), .A2(_06268_ ), .ZN(_06276_ ) );
MUX2_X1 _14263_ ( .A(\ID_EX_csr [6] ), .B(_06276_ ), .S(_06262_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14264_ ( .A1(_05761_ ), .A2(_03013_ ), .ZN(_06277_ ) );
OAI21_X1 _14265_ ( .A(_06277_ ), .B1(_03948_ ), .B2(_06263_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _14266_ ( .A1(_05779_ ), .A2(_03013_ ), .ZN(_06278_ ) );
BUF_X4 _14267_ ( .A(_06261_ ), .Z(_06279_ ) );
BUF_X4 _14268_ ( .A(_06279_ ), .Z(_06280_ ) );
OAI21_X1 _14269_ ( .A(_06278_ ), .B1(_05339_ ), .B2(_06280_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _14270_ ( .A1(_05799_ ), .A2(_03013_ ), .ZN(_06281_ ) );
OAI21_X1 _14271_ ( .A(_06281_ ), .B1(_03909_ ), .B2(_06280_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _14272_ ( .A1(_05816_ ), .A2(_03013_ ), .ZN(_06282_ ) );
OAI21_X1 _14273_ ( .A(_06282_ ), .B1(_03941_ ), .B2(_06280_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
NAND2_X1 _14274_ ( .A1(_05621_ ), .A2(_03013_ ), .ZN(_06283_ ) );
OAI21_X1 _14275_ ( .A(_06283_ ), .B1(_03921_ ), .B2(_06280_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X2 _14276_ ( .A(_06261_ ), .Z(_06284_ ) );
NAND4_X1 _14277_ ( .A1(_03920_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [21] ), .A4(_05601_ ), .ZN(_06285_ ) );
AOI22_X1 _14278_ ( .A1(_03944_ ), .A2(\mycsreg.CSReg[3][21] ), .B1(_03945_ ), .B2(_03950_ ), .ZN(_06286_ ) );
NAND3_X1 _14279_ ( .A1(_03937_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_03938_ ), .ZN(_06287_ ) );
AND2_X1 _14280_ ( .A1(_06287_ ), .A2(_05980_ ), .ZN(_06288_ ) );
NAND4_X1 _14281_ ( .A1(_03914_ ), .A2(_06285_ ), .A3(_06286_ ), .A4(_06288_ ), .ZN(_06289_ ) );
OR3_X1 _14282_ ( .A1(_03902_ ), .A2(_03912_ ), .A3(\EX_LS_result_csreg_mem [21] ), .ZN(_06290_ ) );
NAND2_X1 _14283_ ( .A1(_06289_ ), .A2(_06290_ ), .ZN(_06291_ ) );
AOI22_X1 _14284_ ( .A1(_06291_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02333_ ), .ZN(_06292_ ) );
OAI21_X1 _14285_ ( .A(_06292_ ), .B1(fanout_net_4 ), .B2(_04823_ ), .ZN(_06293_ ) );
NOR2_X1 _14286_ ( .A1(_05284_ ), .A2(fanout_net_5 ), .ZN(_06294_ ) );
NAND3_X1 _14287_ ( .A1(_06289_ ), .A2(_06294_ ), .A3(_06290_ ), .ZN(_06295_ ) );
AOI21_X1 _14288_ ( .A(_06284_ ), .B1(_06293_ ), .B2(_06295_ ), .ZN(_06296_ ) );
AND3_X1 _14289_ ( .A1(_03362_ ), .A2(_05973_ ), .A3(\ID_EX_typ [7] ), .ZN(_06297_ ) );
BUF_X4 _14290_ ( .A(_06269_ ), .Z(_06298_ ) );
AOI211_X1 _14291_ ( .A(_06265_ ), .B(_06297_ ), .C1(_04845_ ), .C2(_06298_ ), .ZN(_06299_ ) );
OR2_X1 _14292_ ( .A1(_06296_ ), .A2(_06299_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
INV_X1 _14293_ ( .A(_06294_ ), .ZN(_06300_ ) );
AOI21_X1 _14294_ ( .A(_06300_ ), .B1(_05380_ ), .B2(_05383_ ), .ZN(_06301_ ) );
AOI22_X1 _14295_ ( .A1(_05384_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02330_ ), .ZN(_06302_ ) );
NAND3_X1 _14296_ ( .A1(_02309_ ), .A2(_02328_ ), .A3(_05528_ ), .ZN(_06303_ ) );
AOI211_X1 _14297_ ( .A(_06284_ ), .B(_06301_ ), .C1(_06302_ ), .C2(_06303_ ), .ZN(_06304_ ) );
MUX2_X1 _14298_ ( .A(_05389_ ), .B(_04821_ ), .S(_06270_ ), .Z(_06305_ ) );
AOI21_X1 _14299_ ( .A(_06304_ ), .B1(_06263_ ), .B2(_06305_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
NAND2_X1 _14300_ ( .A1(_05411_ ), .A2(_05416_ ), .ZN(_06306_ ) );
NAND2_X1 _14301_ ( .A1(_05365_ ), .A2(_06306_ ), .ZN(_06307_ ) );
NAND3_X1 _14302_ ( .A1(_05456_ ), .A2(_05650_ ), .A3(\EX_LS_result_csreg_mem [19] ), .ZN(_06308_ ) );
AOI21_X1 _14303_ ( .A(_06300_ ), .B1(_06307_ ), .B2(_06308_ ), .ZN(_06309_ ) );
NAND3_X1 _14304_ ( .A1(_02380_ ), .A2(_02381_ ), .A3(_05434_ ), .ZN(_06310_ ) );
AOI22_X1 _14305_ ( .A1(_05421_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02383_ ), .ZN(_06311_ ) );
AOI211_X1 _14306_ ( .A(_06284_ ), .B(_06309_ ), .C1(_06310_ ), .C2(_06311_ ), .ZN(_06312_ ) );
MUX2_X1 _14307_ ( .A(_05424_ ), .B(_04674_ ), .S(_06298_ ), .Z(_06313_ ) );
AOI21_X1 _14308_ ( .A(_06312_ ), .B1(_06313_ ), .B2(_06263_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
NAND2_X1 _14309_ ( .A1(_05446_ ), .A2(_05448_ ), .ZN(_06314_ ) );
NAND2_X1 _14310_ ( .A1(_05365_ ), .A2(_06314_ ), .ZN(_06315_ ) );
NAND3_X1 _14311_ ( .A1(_05456_ ), .A2(_05650_ ), .A3(\EX_LS_result_csreg_mem [18] ), .ZN(_06316_ ) );
AOI21_X1 _14312_ ( .A(_06300_ ), .B1(_06315_ ), .B2(_06316_ ), .ZN(_06317_ ) );
NAND3_X1 _14313_ ( .A1(_02385_ ), .A2(_05434_ ), .A3(_02404_ ), .ZN(_06318_ ) );
AOI22_X1 _14314_ ( .A1(_05451_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02406_ ), .ZN(_06319_ ) );
AOI211_X1 _14315_ ( .A(_06284_ ), .B(_06317_ ), .C1(_06318_ ), .C2(_06319_ ), .ZN(_06320_ ) );
MUX2_X1 _14316_ ( .A(_05437_ ), .B(_04697_ ), .S(_06270_ ), .Z(_06321_ ) );
AOI21_X1 _14317_ ( .A(_06320_ ), .B1(_06263_ ), .B2(_06321_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
BUF_X2 _14318_ ( .A(_03937_ ), .Z(_06322_ ) );
AND3_X1 _14319_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_05601_ ), .ZN(_06323_ ) );
NOR2_X1 _14320_ ( .A1(_03913_ ), .A2(_06323_ ), .ZN(_06324_ ) );
BUF_X4 _14321_ ( .A(_03920_ ), .Z(_06325_ ) );
NAND4_X1 _14322_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [17] ), .A4(_05770_ ), .ZN(_06326_ ) );
AND2_X1 _14323_ ( .A1(_03950_ ), .A2(_05405_ ), .ZN(_06327_ ) );
NOR3_X1 _14324_ ( .A1(_05745_ ), .A2(_06327_ ), .A3(_05461_ ), .ZN(_06328_ ) );
NAND4_X1 _14325_ ( .A1(_06324_ ), .A2(_05469_ ), .A3(_06326_ ), .A4(_06328_ ), .ZN(_06329_ ) );
OR3_X1 _14326_ ( .A1(_05869_ ), .A2(_05870_ ), .A3(\EX_LS_result_csreg_mem [17] ), .ZN(_06330_ ) );
NAND2_X1 _14327_ ( .A1(_06329_ ), .A2(_06330_ ), .ZN(_06331_ ) );
AOI22_X1 _14328_ ( .A1(_06331_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02431_ ), .ZN(_06332_ ) );
BUF_X4 _14329_ ( .A(_06260_ ), .Z(_06333_ ) );
OAI211_X1 _14330_ ( .A(_06332_ ), .B(_06333_ ), .C1(fanout_net_4 ), .C2(_02430_ ), .ZN(_06334_ ) );
BUF_X4 _14331_ ( .A(_06279_ ), .Z(_06335_ ) );
AOI21_X1 _14332_ ( .A(_06268_ ), .B1(_04725_ ), .B2(_04745_ ), .ZN(_06336_ ) );
AND3_X1 _14333_ ( .A1(_03362_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_typ [7] ), .ZN(_06337_ ) );
OAI21_X1 _14334_ ( .A(_06335_ ), .B1(_06336_ ), .B2(_06337_ ), .ZN(_06338_ ) );
BUF_X4 _14335_ ( .A(_06294_ ), .Z(_06339_ ) );
BUF_X4 _14336_ ( .A(_06260_ ), .Z(_06340_ ) );
NAND4_X1 _14337_ ( .A1(_06329_ ), .A2(_06339_ ), .A3(_06330_ ), .A4(_06340_ ), .ZN(_06341_ ) );
NAND3_X1 _14338_ ( .A1(_06334_ ), .A2(_06338_ ), .A3(_06341_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _14339_ ( .A(_06300_ ), .B1(_05492_ ), .B2(_05493_ ), .ZN(_06342_ ) );
AOI22_X1 _14340_ ( .A1(_05494_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02455_ ), .ZN(_06343_ ) );
NAND3_X1 _14341_ ( .A1(_02433_ ), .A2(_02452_ ), .A3(_05528_ ), .ZN(_06344_ ) );
AOI211_X1 _14342_ ( .A(_06284_ ), .B(_06342_ ), .C1(_06343_ ), .C2(_06344_ ), .ZN(_06345_ ) );
MUX2_X1 _14343_ ( .A(_05497_ ), .B(_04721_ ), .S(_06270_ ), .Z(_06346_ ) );
AOI21_X1 _14344_ ( .A(_06345_ ), .B1(_06263_ ), .B2(_06346_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
BUF_X4 _14345_ ( .A(_06260_ ), .Z(_06347_ ) );
OAI21_X1 _14346_ ( .A(_06339_ ), .B1(_05523_ ), .B2(_05524_ ), .ZN(_06348_ ) );
BUF_X2 _14347_ ( .A(_05286_ ), .Z(_06349_ ) );
OAI22_X1 _14348_ ( .A1(_05526_ ), .A2(_06349_ ), .B1(_05528_ ), .B2(\ID_EX_imm [15] ), .ZN(_06350_ ) );
AND3_X1 _14349_ ( .A1(_02663_ ), .A2(_05303_ ), .A3(_02682_ ), .ZN(_06351_ ) );
OAI211_X1 _14350_ ( .A(_06347_ ), .B(_06348_ ), .C1(_06350_ ), .C2(_06351_ ), .ZN(_06352_ ) );
NAND4_X1 _14351_ ( .A1(\ID_EX_pc [15] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06353_ ) );
BUF_X4 _14352_ ( .A(_06268_ ), .Z(_06354_ ) );
OAI211_X1 _14353_ ( .A(_06262_ ), .B(_06353_ ), .C1(_04255_ ), .C2(_06354_ ), .ZN(_06355_ ) );
AND2_X1 _14354_ ( .A1(_06352_ ), .A2(_06355_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _14355_ ( .A(_06300_ ), .B1(_05542_ ), .B2(_05543_ ), .ZN(_06356_ ) );
AOI22_X1 _14356_ ( .A1(_05544_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02708_ ), .ZN(_06357_ ) );
NAND3_X1 _14357_ ( .A1(_02686_ ), .A2(_02705_ ), .A3(_05528_ ), .ZN(_06358_ ) );
AOI211_X1 _14358_ ( .A(_06284_ ), .B(_06356_ ), .C1(_06357_ ), .C2(_06358_ ), .ZN(_06359_ ) );
MUX2_X1 _14359_ ( .A(_05513_ ), .B(_04280_ ), .S(_06270_ ), .Z(_06360_ ) );
AOI21_X1 _14360_ ( .A(_06359_ ), .B1(_06263_ ), .B2(_06360_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
NAND3_X1 _14361_ ( .A1(_05571_ ), .A2(_06339_ ), .A3(_06333_ ), .ZN(_06361_ ) );
AND3_X1 _14362_ ( .A1(_02734_ ), .A2(_05434_ ), .A3(_02754_ ), .ZN(_06362_ ) );
OAI221_X1 _14363_ ( .A(_06265_ ), .B1(_05434_ ), .B2(\ID_EX_imm [13] ), .C1(_05571_ ), .C2(_06349_ ), .ZN(_06363_ ) );
MUX2_X1 _14364_ ( .A(_05550_ ), .B(_04307_ ), .S(_06269_ ), .Z(_06364_ ) );
OAI221_X1 _14365_ ( .A(_06361_ ), .B1(_06362_ ), .B2(_06363_ ), .C1(_06364_ ), .C2(_06266_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AOI21_X1 _14366_ ( .A(_06300_ ), .B1(_05591_ ), .B2(_05592_ ), .ZN(_06365_ ) );
AND2_X1 _14367_ ( .A1(_05591_ ), .A2(_05592_ ), .ZN(_06366_ ) );
AOI22_X1 _14368_ ( .A1(_06366_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02732_ ), .ZN(_06367_ ) );
NAND3_X1 _14369_ ( .A1(_02711_ ), .A2(_05434_ ), .A3(_02730_ ), .ZN(_06368_ ) );
AOI211_X1 _14370_ ( .A(_06279_ ), .B(_06365_ ), .C1(_06367_ ), .C2(_06368_ ), .ZN(_06369_ ) );
MUX2_X1 _14371_ ( .A(_05576_ ), .B(_04333_ ), .S(_06270_ ), .Z(_06370_ ) );
AOI21_X1 _14372_ ( .A(_06369_ ), .B1(_06263_ ), .B2(_06370_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
NAND3_X1 _14373_ ( .A1(_03952_ ), .A2(_06294_ ), .A3(_03953_ ), .ZN(_06371_ ) );
AND3_X1 _14374_ ( .A1(_02173_ ), .A2(_05303_ ), .A3(_02177_ ), .ZN(_06372_ ) );
OAI22_X1 _14375_ ( .A1(_03954_ ), .A2(_06349_ ), .B1(_05303_ ), .B2(\ID_EX_imm [30] ), .ZN(_06373_ ) );
OAI211_X1 _14376_ ( .A(_06265_ ), .B(_06371_ ), .C1(_06372_ ), .C2(_06373_ ), .ZN(_06374_ ) );
INV_X1 _14377_ ( .A(_06374_ ), .ZN(_06375_ ) );
MUX2_X1 _14378_ ( .A(_05992_ ), .B(_04476_ ), .S(_06270_ ), .Z(_06376_ ) );
AOI21_X1 _14379_ ( .A(_06375_ ), .B1(_06263_ ), .B2(_06376_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
OR3_X1 _14380_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [11] ), .ZN(_06377_ ) );
INV_X1 _14381_ ( .A(_06327_ ), .ZN(_06378_ ) );
NAND4_X1 _14382_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [11] ), .A4(_05821_ ), .ZN(_06379_ ) );
NAND4_X1 _14383_ ( .A1(_05746_ ), .A2(_06378_ ), .A3(_05599_ ), .A4(_06379_ ), .ZN(_06380_ ) );
NAND3_X1 _14384_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_05849_ ), .ZN(_06381_ ) );
OAI211_X1 _14385_ ( .A(_05600_ ), .B(_06381_ ), .C1(_05869_ ), .C2(_05870_ ), .ZN(_06382_ ) );
OAI21_X1 _14386_ ( .A(_06377_ ), .B1(_06380_ ), .B2(_06382_ ), .ZN(_06383_ ) );
AOI22_X1 _14387_ ( .A1(_06383_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02852_ ), .ZN(_06384_ ) );
OAI211_X1 _14388_ ( .A(_06384_ ), .B(_06340_ ), .C1(_02851_ ), .C2(fanout_net_4 ), .ZN(_06385_ ) );
CLKBUF_X2 _14389_ ( .A(_06300_ ), .Z(_06386_ ) );
OR3_X1 _14390_ ( .A1(_06383_ ), .A2(_06386_ ), .A3(_06279_ ), .ZN(_06387_ ) );
BUF_X4 _14391_ ( .A(_06347_ ), .Z(_06388_ ) );
AOI21_X1 _14392_ ( .A(_06268_ ), .B1(_04197_ ), .B2(_04202_ ), .ZN(_06389_ ) );
AOI21_X1 _14393_ ( .A(_06389_ ), .B1(\ID_EX_pc [11] ), .B2(_06354_ ), .ZN(_06390_ ) );
OAI211_X1 _14394_ ( .A(_06385_ ), .B(_06387_ ), .C1(_06388_ ), .C2(_06390_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _14395_ ( .A(_06268_ ), .B1(_04226_ ), .B2(_04227_ ), .ZN(_06391_ ) );
AOI211_X1 _14396_ ( .A(_06347_ ), .B(_06391_ ), .C1(\ID_EX_pc [10] ), .C2(_06354_ ), .ZN(_06392_ ) );
NAND2_X1 _14397_ ( .A1(_05647_ ), .A2(_05649_ ), .ZN(_06393_ ) );
NAND2_X1 _14398_ ( .A1(_05365_ ), .A2(_06393_ ), .ZN(_06394_ ) );
NAND3_X1 _14399_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(\EX_LS_result_csreg_mem [10] ), .ZN(_06395_ ) );
AOI21_X1 _14400_ ( .A(_06300_ ), .B1(_06394_ ), .B2(_06395_ ), .ZN(_06396_ ) );
NAND3_X1 _14401_ ( .A1(_02808_ ), .A2(_02827_ ), .A3(_05304_ ), .ZN(_06397_ ) );
AOI22_X1 _14402_ ( .A1(_05653_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02829_ ), .ZN(_06398_ ) );
AOI211_X1 _14403_ ( .A(_06284_ ), .B(_06396_ ), .C1(_06397_ ), .C2(_06398_ ), .ZN(_06399_ ) );
NOR2_X1 _14404_ ( .A1(_06392_ ), .A2(_06399_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
AOI21_X1 _14405_ ( .A(_06268_ ), .B1(_04104_ ), .B2(_04139_ ), .ZN(_06400_ ) );
AOI211_X1 _14406_ ( .A(_06265_ ), .B(_06400_ ), .C1(\ID_EX_pc [9] ), .C2(_06354_ ), .ZN(_06401_ ) );
INV_X1 _14407_ ( .A(_05670_ ), .ZN(_06402_ ) );
INV_X1 _14408_ ( .A(_05671_ ), .ZN(_06403_ ) );
AOI21_X1 _14409_ ( .A(_06300_ ), .B1(_06402_ ), .B2(_06403_ ), .ZN(_06404_ ) );
NAND3_X1 _14410_ ( .A1(_02800_ ), .A2(_02801_ ), .A3(_05304_ ), .ZN(_06405_ ) );
AOI22_X1 _14411_ ( .A1(_05672_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02805_ ), .ZN(_06406_ ) );
AOI211_X1 _14412_ ( .A(_06284_ ), .B(_06404_ ), .C1(_06405_ ), .C2(_06406_ ), .ZN(_06407_ ) );
NOR2_X1 _14413_ ( .A1(_06401_ ), .A2(_06407_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _14414_ ( .A(_06386_ ), .B1(_05686_ ), .B2(_05687_ ), .ZN(_06408_ ) );
AOI22_X1 _14415_ ( .A1(_05688_ ), .A2(fanout_net_5 ), .B1(fanout_net_4 ), .B2(_02781_ ), .ZN(_06409_ ) );
NAND3_X1 _14416_ ( .A1(_02760_ ), .A2(_02779_ ), .A3(_05304_ ), .ZN(_06410_ ) );
AOI211_X1 _14417_ ( .A(_06262_ ), .B(_06408_ ), .C1(_06409_ ), .C2(_06410_ ), .ZN(_06411_ ) );
AOI21_X1 _14418_ ( .A(_06268_ ), .B1(_04147_ ), .B2(_04174_ ), .ZN(_06412_ ) );
AOI211_X1 _14419_ ( .A(_06265_ ), .B(_06412_ ), .C1(\ID_EX_pc [8] ), .C2(_06354_ ), .ZN(_06413_ ) );
NOR2_X1 _14420_ ( .A1(_06411_ ), .A2(_06413_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
BUF_X4 _14421_ ( .A(_06265_ ), .Z(_06414_ ) );
OAI22_X1 _14422_ ( .A1(_05709_ ), .A2(_06386_ ), .B1(_05304_ ), .B2(_02630_ ), .ZN(_06415_ ) );
AOI21_X1 _14423_ ( .A(fanout_net_4 ), .B1(_02629_ ), .B2(_02649_ ), .ZN(_06416_ ) );
OAI221_X1 _14424_ ( .A(_06414_ ), .B1(_06349_ ), .B2(_05710_ ), .C1(_06415_ ), .C2(_06416_ ), .ZN(_06417_ ) );
NAND3_X1 _14425_ ( .A1(_04924_ ), .A2(_04944_ ), .A3(_06298_ ), .ZN(_06418_ ) );
OAI211_X1 _14426_ ( .A(_06418_ ), .B(_06335_ ), .C1(\ID_EX_pc [7] ), .C2(_06298_ ), .ZN(_06419_ ) );
NAND2_X1 _14427_ ( .A1(_06417_ ), .A2(_06419_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
NAND3_X1 _14428_ ( .A1(_05727_ ), .A2(_06339_ ), .A3(_06340_ ), .ZN(_06420_ ) );
AND3_X1 _14429_ ( .A1(_02606_ ), .A2(_05434_ ), .A3(_02625_ ), .ZN(_06421_ ) );
OAI221_X1 _14430_ ( .A(_06265_ ), .B1(_05434_ ), .B2(\ID_EX_imm [6] ), .C1(_05727_ ), .C2(_06349_ ), .ZN(_06422_ ) );
MUX2_X1 _14431_ ( .A(_05728_ ), .B(_04920_ ), .S(_06269_ ), .Z(_06423_ ) );
OAI221_X1 _14432_ ( .A(_06420_ ), .B1(_06421_ ), .B2(_06422_ ), .C1(_06423_ ), .C2(_06266_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
BUF_X4 _14433_ ( .A(_06265_ ), .Z(_06424_ ) );
OAI22_X1 _14434_ ( .A1(_05757_ ), .A2(_06349_ ), .B1(_05303_ ), .B2(\ID_EX_imm [5] ), .ZN(_06425_ ) );
AOI21_X1 _14435_ ( .A(_06425_ ), .B1(_05304_ ), .B2(_05109_ ), .ZN(_06426_ ) );
INV_X1 _14436_ ( .A(_05756_ ), .ZN(_06427_ ) );
OAI211_X1 _14437_ ( .A(_06427_ ), .B(_06294_ ), .C1(_05750_ ), .C2(_05752_ ), .ZN(_06428_ ) );
INV_X1 _14438_ ( .A(_06428_ ), .ZN(_06429_ ) );
OAI21_X1 _14439_ ( .A(_06424_ ), .B1(_06426_ ), .B2(_06429_ ), .ZN(_06430_ ) );
NAND3_X1 _14440_ ( .A1(_03362_ ), .A2(_05737_ ), .A3(\ID_EX_typ [7] ), .ZN(_06431_ ) );
OAI211_X1 _14441_ ( .A(_06335_ ), .B(_06431_ ), .C1(_04896_ ), .C2(_06354_ ), .ZN(_06432_ ) );
NAND2_X1 _14442_ ( .A1(_06430_ ), .A2(_06432_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
OR3_X1 _14443_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [4] ), .ZN(_06433_ ) );
NAND3_X1 _14444_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_05821_ ), .ZN(_06434_ ) );
NAND4_X1 _14445_ ( .A1(_05746_ ), .A2(_05773_ ), .A3(_05774_ ), .A4(_06434_ ), .ZN(_06435_ ) );
NAND4_X1 _14446_ ( .A1(_03920_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [4] ), .A4(_05821_ ), .ZN(_06436_ ) );
OAI21_X1 _14447_ ( .A(_06436_ ), .B1(_05869_ ), .B2(_05870_ ), .ZN(_06437_ ) );
OAI21_X1 _14448_ ( .A(_06433_ ), .B1(_06435_ ), .B2(_06437_ ), .ZN(_06438_ ) );
AOI22_X1 _14449_ ( .A1(_06438_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_02604_ ), .ZN(_06439_ ) );
OAI211_X1 _14450_ ( .A(_06439_ ), .B(_06340_ ), .C1(_02603_ ), .C2(\ID_EX_typ [0] ), .ZN(_06440_ ) );
OR3_X1 _14451_ ( .A1(_06438_ ), .A2(_06386_ ), .A3(_06279_ ), .ZN(_06441_ ) );
AND3_X1 _14452_ ( .A1(_04871_ ), .A2(_04872_ ), .A3(_06269_ ), .ZN(_06442_ ) );
AOI21_X1 _14453_ ( .A(_06442_ ), .B1(\ID_EX_pc [4] ), .B2(_06354_ ), .ZN(_06443_ ) );
OAI211_X1 _14454_ ( .A(_06440_ ), .B(_06441_ ), .C1(_06443_ ), .C2(_06388_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
NAND3_X1 _14455_ ( .A1(_05795_ ), .A2(_06339_ ), .A3(_06340_ ), .ZN(_06444_ ) );
OAI221_X1 _14456_ ( .A(_06265_ ), .B1(_05304_ ), .B2(\ID_EX_imm [3] ), .C1(_05795_ ), .C2(_06349_ ), .ZN(_06445_ ) );
AND3_X1 _14457_ ( .A1(_02506_ ), .A2(_05434_ ), .A3(_02526_ ), .ZN(_06446_ ) );
AND4_X1 _14458_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06447_ ) );
AOI21_X1 _14459_ ( .A(_06447_ ), .B1(_04443_ ), .B2(_06298_ ), .ZN(_06448_ ) );
OAI221_X1 _14460_ ( .A(_06444_ ), .B1(_06445_ ), .B2(_06446_ ), .C1(_06448_ ), .C2(_06266_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
AND3_X1 _14461_ ( .A1(_04396_ ), .A2(_04418_ ), .A3(_06269_ ), .ZN(_06449_ ) );
AND3_X1 _14462_ ( .A1(_03362_ ), .A2(\ID_EX_pc [2] ), .A3(\ID_EX_typ [7] ), .ZN(_06450_ ) );
OAI21_X1 _14463_ ( .A(_06280_ ), .B1(_06449_ ), .B2(_06450_ ), .ZN(_06451_ ) );
OR3_X1 _14464_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [2] ), .ZN(_06452_ ) );
NAND3_X1 _14465_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_05821_ ), .ZN(_06453_ ) );
AND2_X1 _14466_ ( .A1(_06453_ ), .A2(_05807_ ), .ZN(_06454_ ) );
AOI22_X1 _14467_ ( .A1(_03944_ ), .A2(\mycsreg.CSReg[3][2] ), .B1(_05561_ ), .B2(_03950_ ), .ZN(_06455_ ) );
NAND2_X1 _14468_ ( .A1(_06454_ ), .A2(_06455_ ), .ZN(_06456_ ) );
NAND4_X1 _14469_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [2] ), .A4(_05849_ ), .ZN(_06457_ ) );
OAI21_X1 _14470_ ( .A(_06457_ ), .B1(_05869_ ), .B2(_05870_ ), .ZN(_06458_ ) );
OAI21_X1 _14471_ ( .A(_06452_ ), .B1(_06456_ ), .B2(_06458_ ), .ZN(_06459_ ) );
AOI22_X1 _14472_ ( .A1(_06459_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_05117_ ), .ZN(_06460_ ) );
OAI211_X1 _14473_ ( .A(_06333_ ), .B(_06460_ ), .C1(_02549_ ), .C2(\ID_EX_typ [0] ), .ZN(_06461_ ) );
OR3_X1 _14474_ ( .A1(_06459_ ), .A2(_06386_ ), .A3(_06279_ ), .ZN(_06462_ ) );
NAND3_X1 _14475_ ( .A1(_06451_ ), .A2(_06461_ ), .A3(_06462_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
INV_X1 _14476_ ( .A(_05357_ ), .ZN(_06463_ ) );
AOI221_X4 _14477_ ( .A(_06261_ ), .B1(\ID_EX_typ [0] ), .B2(_02974_ ), .C1(_06463_ ), .C2(fanout_net_5 ), .ZN(_06464_ ) );
OAI21_X1 _14478_ ( .A(_06464_ ), .B1(\ID_EX_typ [0] ), .B2(_02973_ ), .ZN(_06465_ ) );
NAND3_X1 _14479_ ( .A1(_05357_ ), .A2(_06339_ ), .A3(_06333_ ), .ZN(_06466_ ) );
AND4_X1 _14480_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06467_ ) );
AOI21_X1 _14481_ ( .A(_06467_ ), .B1(_04544_ ), .B2(_06298_ ), .ZN(_06468_ ) );
OAI211_X1 _14482_ ( .A(_06465_ ), .B(_06466_ ), .C1(_06388_ ), .C2(_06468_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
AOI21_X1 _14483_ ( .A(_06354_ ), .B1(_04341_ ), .B2(_04362_ ), .ZN(_06469_ ) );
AND3_X1 _14484_ ( .A1(_03362_ ), .A2(\ID_EX_pc [1] ), .A3(\ID_EX_typ [7] ), .ZN(_06470_ ) );
OAI21_X1 _14485_ ( .A(_06280_ ), .B1(_06469_ ), .B2(_06470_ ), .ZN(_06471_ ) );
OR3_X1 _14486_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [1] ), .ZN(_06472_ ) );
NAND4_X1 _14487_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [1] ), .A4(_05849_ ), .ZN(_06473_ ) );
NAND3_X1 _14488_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_05849_ ), .ZN(_06474_ ) );
NAND4_X1 _14489_ ( .A1(_06473_ ), .A2(_06474_ ), .A3(_05819_ ), .A4(_05820_ ), .ZN(_06475_ ) );
OAI21_X1 _14490_ ( .A(_06472_ ), .B1(_03913_ ), .B2(_06475_ ), .ZN(_06476_ ) );
AOI22_X1 _14491_ ( .A1(_06476_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_05127_ ), .ZN(_06477_ ) );
OAI211_X1 _14492_ ( .A(_06333_ ), .B(_06477_ ), .C1(_02478_ ), .C2(\ID_EX_typ [0] ), .ZN(_06478_ ) );
OR3_X1 _14493_ ( .A1(_06476_ ), .A2(_06386_ ), .A3(_06279_ ), .ZN(_06479_ ) );
NAND3_X1 _14494_ ( .A1(_06471_ ), .A2(_06478_ ), .A3(_06479_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
OAI21_X1 _14495_ ( .A(_05862_ ), .B1(_05867_ ), .B2(_05871_ ), .ZN(_06480_ ) );
AOI22_X1 _14496_ ( .A1(_06480_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_02480_ ), .ZN(_06481_ ) );
OAI211_X1 _14497_ ( .A(_06481_ ), .B(_06347_ ), .C1(_02502_ ), .C2(\ID_EX_typ [0] ), .ZN(_06482_ ) );
OR3_X1 _14498_ ( .A1(_06480_ ), .A2(_06386_ ), .A3(_06279_ ), .ZN(_06483_ ) );
MUX2_X1 _14499_ ( .A(_05860_ ), .B(_04386_ ), .S(_06270_ ), .Z(_06484_ ) );
OAI211_X1 _14500_ ( .A(_06482_ ), .B(_06483_ ), .C1(_06484_ ), .C2(_06388_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
NAND3_X1 _14501_ ( .A1(_02182_ ), .A2(_05304_ ), .A3(_02208_ ), .ZN(_06485_ ) );
OR2_X1 _14502_ ( .A1(_05303_ ), .A2(\ID_EX_imm [28] ), .ZN(_06486_ ) );
OR3_X1 _14503_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [28] ), .ZN(_06487_ ) );
NAND4_X1 _14504_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [28] ), .A4(_05770_ ), .ZN(_06488_ ) );
NAND3_X1 _14505_ ( .A1(_05746_ ), .A2(_05625_ ), .A3(_06488_ ), .ZN(_06489_ ) );
NAND3_X1 _14506_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_05849_ ), .ZN(_06490_ ) );
OAI211_X1 _14507_ ( .A(_05626_ ), .B(_06490_ ), .C1(_05869_ ), .C2(_05870_ ), .ZN(_06491_ ) );
OAI21_X1 _14508_ ( .A(_06487_ ), .B1(_06489_ ), .B2(_06491_ ), .ZN(_06492_ ) );
NAND2_X1 _14509_ ( .A1(_06492_ ), .A2(fanout_net_5 ), .ZN(_06493_ ) );
NAND4_X1 _14510_ ( .A1(_06485_ ), .A2(_06340_ ), .A3(_06486_ ), .A4(_06493_ ), .ZN(_06494_ ) );
OR3_X1 _14511_ ( .A1(_06492_ ), .A2(_06386_ ), .A3(_06279_ ), .ZN(_06495_ ) );
AND3_X1 _14512_ ( .A1(_03362_ ), .A2(\ID_EX_pc [28] ), .A3(\ID_EX_typ [7] ), .ZN(_06496_ ) );
AOI21_X1 _14513_ ( .A(_06496_ ), .B1(_04521_ ), .B2(_06298_ ), .ZN(_06497_ ) );
OAI211_X1 _14514_ ( .A(_06494_ ), .B(_06495_ ), .C1(_06497_ ), .C2(_06388_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND3_X1 _14515_ ( .A1(_05851_ ), .A2(_06294_ ), .A3(_05853_ ), .ZN(_06498_ ) );
NAND2_X1 _14516_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [27] ), .ZN(_06499_ ) );
NAND2_X1 _14517_ ( .A1(_06498_ ), .A2(_06499_ ), .ZN(_06500_ ) );
AOI21_X1 _14518_ ( .A(\ID_EX_typ [0] ), .B1(_02211_ ), .B2(_02232_ ), .ZN(_06501_ ) );
OAI221_X1 _14519_ ( .A(_06414_ ), .B1(_06349_ ), .B2(_05854_ ), .C1(_06500_ ), .C2(_06501_ ), .ZN(_06502_ ) );
OR4_X1 _14520_ ( .A1(\ID_EX_pc [27] ), .A2(_03348_ ), .A3(_03872_ ), .A4(_03875_ ), .ZN(_06503_ ) );
OAI211_X1 _14521_ ( .A(_06335_ ), .B(_06503_ ), .C1(_04595_ ), .C2(_06354_ ), .ZN(_06504_ ) );
NAND2_X1 _14522_ ( .A1(_06502_ ), .A2(_06504_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
NAND4_X1 _14523_ ( .A1(_05408_ ), .A2(_05565_ ), .A3(\mycsreg.CSReg[0][26] ), .A4(_05566_ ), .ZN(_06505_ ) );
AND2_X1 _14524_ ( .A1(_05877_ ), .A2(_06505_ ), .ZN(_06506_ ) );
NAND4_X1 _14525_ ( .A1(_05412_ ), .A2(_05587_ ), .A3(\mtvec [26] ), .A4(_05588_ ), .ZN(_06507_ ) );
AND2_X1 _14526_ ( .A1(_05879_ ), .A2(_06507_ ), .ZN(_06508_ ) );
AOI22_X1 _14527_ ( .A1(_06506_ ), .A2(_06508_ ), .B1(_05650_ ), .B2(_05456_ ), .ZN(_06509_ ) );
AND3_X1 _14528_ ( .A1(_05381_ ), .A2(_05382_ ), .A3(\EX_LS_result_csreg_mem [26] ), .ZN(_06510_ ) );
NOR2_X1 _14529_ ( .A1(_06509_ ), .A2(_06510_ ), .ZN(_06511_ ) );
AOI22_X1 _14530_ ( .A1(_06511_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_02257_ ), .ZN(_06512_ ) );
OAI211_X1 _14531_ ( .A(_06340_ ), .B(_06512_ ), .C1(_02256_ ), .C2(\ID_EX_typ [0] ), .ZN(_06513_ ) );
AND2_X1 _14532_ ( .A1(_05877_ ), .A2(_05879_ ), .ZN(_06514_ ) );
AND2_X1 _14533_ ( .A1(_05878_ ), .A2(_05880_ ), .ZN(_06515_ ) );
NAND3_X1 _14534_ ( .A1(_03914_ ), .A2(_06514_ ), .A3(_06515_ ), .ZN(_06516_ ) );
INV_X1 _14535_ ( .A(_05876_ ), .ZN(_06517_ ) );
NAND4_X1 _14536_ ( .A1(_06516_ ), .A2(_06339_ ), .A3(_06517_ ), .A4(_06347_ ), .ZN(_06518_ ) );
AND3_X1 _14537_ ( .A1(_03362_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_06519_ ) );
AOI21_X1 _14538_ ( .A(_06519_ ), .B1(_04571_ ), .B2(_06298_ ), .ZN(_06520_ ) );
OAI211_X1 _14539_ ( .A(_06513_ ), .B(_06518_ ), .C1(_06520_ ), .C2(_06388_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
OR3_X1 _14540_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [25] ), .ZN(_06521_ ) );
NAND4_X1 _14541_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [25] ), .A4(_05821_ ), .ZN(_06522_ ) );
NAND3_X1 _14542_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_05849_ ), .ZN(_06523_ ) );
NAND4_X1 _14543_ ( .A1(_06522_ ), .A2(_06523_ ), .A3(_05896_ ), .A4(_05897_ ), .ZN(_06524_ ) );
OAI21_X1 _14544_ ( .A(_06521_ ), .B1(_03913_ ), .B2(_06524_ ), .ZN(_06525_ ) );
AOI22_X1 _14545_ ( .A1(_06525_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_02939_ ), .ZN(_06526_ ) );
OAI211_X1 _14546_ ( .A(_06340_ ), .B(_06526_ ), .C1(_02938_ ), .C2(\ID_EX_typ [0] ), .ZN(_06527_ ) );
AND2_X1 _14547_ ( .A1(_05896_ ), .A2(_05897_ ), .ZN(_06528_ ) );
AND2_X1 _14548_ ( .A1(_06522_ ), .A2(_06523_ ), .ZN(_06529_ ) );
NAND3_X1 _14549_ ( .A1(_03914_ ), .A2(_06528_ ), .A3(_06529_ ), .ZN(_06530_ ) );
NAND4_X1 _14550_ ( .A1(_06530_ ), .A2(_06339_ ), .A3(_06521_ ), .A4(_06347_ ), .ZN(_06531_ ) );
AND3_X1 _14551_ ( .A1(_03362_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06532_ ) );
AOI21_X1 _14552_ ( .A(_06532_ ), .B1(_04645_ ), .B2(_06298_ ), .ZN(_06533_ ) );
OAI211_X1 _14553_ ( .A(_06527_ ), .B(_06531_ ), .C1(_06533_ ), .C2(_06388_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
OR3_X1 _14554_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [24] ), .ZN(_06534_ ) );
NAND4_X1 _14555_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [24] ), .A4(_05821_ ), .ZN(_06535_ ) );
NAND4_X1 _14556_ ( .A1(_05746_ ), .A2(_06378_ ), .A3(_05921_ ), .A4(_06535_ ), .ZN(_06536_ ) );
NAND3_X1 _14557_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_05849_ ), .ZN(_06537_ ) );
OAI211_X1 _14558_ ( .A(_05922_ ), .B(_06537_ ), .C1(_05869_ ), .C2(_05870_ ), .ZN(_06538_ ) );
OAI21_X1 _14559_ ( .A(_06534_ ), .B1(_06536_ ), .B2(_06538_ ), .ZN(_06539_ ) );
AOI22_X1 _14560_ ( .A1(_06539_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_02916_ ), .ZN(_06540_ ) );
OAI211_X1 _14561_ ( .A(_06540_ ), .B(_06347_ ), .C1(_02915_ ), .C2(\ID_EX_typ [0] ), .ZN(_06541_ ) );
OR3_X1 _14562_ ( .A1(_06539_ ), .A2(_06386_ ), .A3(_06261_ ), .ZN(_06542_ ) );
MUX2_X1 _14563_ ( .A(_05905_ ), .B(_04621_ ), .S(_06270_ ), .Z(_06543_ ) );
OAI211_X1 _14564_ ( .A(_06541_ ), .B(_06542_ ), .C1(_06543_ ), .C2(_06266_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
OR3_X1 _14565_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [23] ), .ZN(_06544_ ) );
NAND4_X1 _14566_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [23] ), .A4(_05821_ ), .ZN(_06545_ ) );
NAND3_X1 _14567_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_05849_ ), .ZN(_06546_ ) );
NAND4_X1 _14568_ ( .A1(_06545_ ), .A2(_06546_ ), .A3(_05933_ ), .A4(_05936_ ), .ZN(_06547_ ) );
OAI21_X1 _14569_ ( .A(_06544_ ), .B1(_03913_ ), .B2(_06547_ ), .ZN(_06548_ ) );
AOI22_X1 _14570_ ( .A1(_06548_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_02283_ ), .ZN(_06549_ ) );
OAI211_X1 _14571_ ( .A(_06340_ ), .B(_06549_ ), .C1(_02282_ ), .C2(\ID_EX_typ [0] ), .ZN(_06550_ ) );
AND2_X1 _14572_ ( .A1(_05933_ ), .A2(_05936_ ), .ZN(_06551_ ) );
AND2_X1 _14573_ ( .A1(_06545_ ), .A2(_06546_ ), .ZN(_06552_ ) );
NAND3_X1 _14574_ ( .A1(_03914_ ), .A2(_06551_ ), .A3(_06552_ ), .ZN(_06553_ ) );
NAND4_X1 _14575_ ( .A1(_06553_ ), .A2(_06339_ ), .A3(_06544_ ), .A4(_06347_ ), .ZN(_06554_ ) );
AOI21_X1 _14576_ ( .A(_06268_ ), .B1(_04795_ ), .B2(_04793_ ), .ZN(_06555_ ) );
AOI21_X1 _14577_ ( .A(_06555_ ), .B1(\ID_EX_pc [23] ), .B2(_06354_ ), .ZN(_06556_ ) );
OAI211_X1 _14578_ ( .A(_06550_ ), .B(_06554_ ), .C1(_06556_ ), .C2(_06266_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
OR3_X1 _14579_ ( .A1(_05754_ ), .A2(_05755_ ), .A3(\EX_LS_result_csreg_mem [22] ), .ZN(_06557_ ) );
NOR2_X1 _14580_ ( .A1(_05745_ ), .A2(_06327_ ), .ZN(_06558_ ) );
AND3_X1 _14581_ ( .A1(_03937_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_05565_ ), .ZN(_06559_ ) );
NOR2_X1 _14582_ ( .A1(_06559_ ), .A2(_05957_ ), .ZN(_06560_ ) );
NAND3_X1 _14583_ ( .A1(_06558_ ), .A2(_05961_ ), .A3(_06560_ ), .ZN(_06561_ ) );
NAND4_X1 _14584_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [22] ), .A4(_05821_ ), .ZN(_06562_ ) );
OAI21_X1 _14585_ ( .A(_06562_ ), .B1(_05869_ ), .B2(_05870_ ), .ZN(_06563_ ) );
OAI21_X1 _14586_ ( .A(_06557_ ), .B1(_06561_ ), .B2(_06563_ ), .ZN(_06564_ ) );
AOI22_X1 _14587_ ( .A1(_06564_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_02306_ ), .ZN(_06565_ ) );
OAI211_X1 _14588_ ( .A(_06565_ ), .B(_06347_ ), .C1(\ID_EX_typ [0] ), .C2(_02305_ ), .ZN(_06566_ ) );
OR3_X1 _14589_ ( .A1(_06564_ ), .A2(_06386_ ), .A3(_06261_ ), .ZN(_06567_ ) );
MUX2_X1 _14590_ ( .A(_05964_ ), .B(_04772_ ), .S(_06270_ ), .Z(_06568_ ) );
OAI211_X1 _14591_ ( .A(_06566_ ), .B(_06567_ ), .C1(_06568_ ), .C2(_06266_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
AOI22_X1 _14592_ ( .A1(_06005_ ), .A2(fanout_net_5 ), .B1(\ID_EX_typ [0] ), .B2(_04959_ ), .ZN(_06569_ ) );
OAI211_X1 _14593_ ( .A(_06340_ ), .B(_06569_ ), .C1(_03006_ ), .C2(\ID_EX_typ [0] ), .ZN(_06570_ ) );
AND2_X1 _14594_ ( .A1(_05997_ ), .A2(_06000_ ), .ZN(_06571_ ) );
NAND4_X1 _14595_ ( .A1(_06325_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [31] ), .A4(_05770_ ), .ZN(_06572_ ) );
NAND3_X1 _14596_ ( .A1(_06322_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_05770_ ), .ZN(_06573_ ) );
AND2_X1 _14597_ ( .A1(_06572_ ), .A2(_06573_ ), .ZN(_06574_ ) );
NAND3_X1 _14598_ ( .A1(_03914_ ), .A2(_06571_ ), .A3(_06574_ ), .ZN(_06575_ ) );
NOR3_X1 _14599_ ( .A1(_05869_ ), .A2(_05870_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_06576_ ) );
INV_X1 _14600_ ( .A(_06576_ ), .ZN(_06577_ ) );
NAND4_X1 _14601_ ( .A1(_06575_ ), .A2(_06339_ ), .A3(_06577_ ), .A4(_06347_ ), .ZN(_06578_ ) );
AND3_X1 _14602_ ( .A1(_03362_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06579_ ) );
AOI21_X1 _14603_ ( .A(_06579_ ), .B1(_04499_ ), .B2(_06298_ ), .ZN(_06580_ ) );
OAI211_X1 _14604_ ( .A(_06570_ ), .B(_06578_ ), .C1(_06580_ ), .C2(_06266_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
NAND3_X1 _14605_ ( .A1(_05985_ ), .A2(_05987_ ), .A3(_06333_ ), .ZN(_06581_ ) );
NOR2_X1 _14606_ ( .A1(_03875_ ), .A2(\ID_EX_typ [6] ), .ZN(_06582_ ) );
AND2_X2 _14607_ ( .A1(_06582_ ), .A2(_03348_ ), .ZN(_06583_ ) );
INV_X2 _14608_ ( .A(_06583_ ), .ZN(_06584_ ) );
BUF_X4 _14609_ ( .A(_06584_ ), .Z(_06585_ ) );
INV_X1 _14610_ ( .A(_05241_ ), .ZN(_06586_ ) );
NAND2_X1 _14611_ ( .A1(_06586_ ), .A2(_04748_ ), .ZN(_06587_ ) );
AND2_X1 _14612_ ( .A1(_06587_ ), .A2(_05256_ ), .ZN(_06588_ ) );
INV_X1 _14613_ ( .A(_04822_ ), .ZN(_06589_ ) );
OR2_X1 _14614_ ( .A1(_06588_ ), .A2(_06589_ ), .ZN(_06590_ ) );
AND2_X1 _14615_ ( .A1(_06590_ ), .A2(_05244_ ), .ZN(_06591_ ) );
XNOR2_X1 _14616_ ( .A(_06591_ ), .B(_04848_ ), .ZN(_06592_ ) );
AND3_X1 _14617_ ( .A1(_04089_ ), .A2(\ID_EX_typ [3] ), .A3(_06349_ ), .ZN(_06593_ ) );
AND2_X1 _14618_ ( .A1(_06593_ ), .A2(_04957_ ), .ZN(_06594_ ) );
BUF_X2 _14619_ ( .A(_06594_ ), .Z(_06595_ ) );
NAND2_X1 _14620_ ( .A1(_06592_ ), .A2(_06595_ ), .ZN(_06596_ ) );
NOR3_X1 _14621_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06597_ ) );
AND2_X2 _14622_ ( .A1(\ID_EX_typ [3] ), .A2(fanout_net_5 ), .ZN(_06598_ ) );
AND2_X2 _14623_ ( .A1(_06597_ ), .A2(_06598_ ), .ZN(_06599_ ) );
BUF_X4 _14624_ ( .A(_06599_ ), .Z(_06600_ ) );
NOR3_X1 _14625_ ( .A1(_05284_ ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06601_ ) );
AND2_X1 _14626_ ( .A1(_06601_ ), .A2(_06598_ ), .ZN(_06602_ ) );
BUF_X4 _14627_ ( .A(_06602_ ), .Z(_06603_ ) );
BUF_X4 _14628_ ( .A(_06603_ ), .Z(_06604_ ) );
AOI22_X1 _14629_ ( .A1(_05977_ ), .A2(_06600_ ), .B1(\ID_EX_imm [21] ), .B2(_06604_ ), .ZN(_06605_ ) );
AOI21_X1 _14630_ ( .A(_06585_ ), .B1(_06596_ ), .B2(_06605_ ), .ZN(_06606_ ) );
CLKBUF_X2 _14631_ ( .A(_03877_ ), .Z(_06607_ ) );
OR2_X1 _14632_ ( .A1(_06606_ ), .A2(_06607_ ), .ZN(_06608_ ) );
NOR2_X1 _14633_ ( .A1(_05119_ ), .A2(_04390_ ), .ZN(_06609_ ) );
INV_X1 _14634_ ( .A(_06609_ ), .ZN(_06610_ ) );
NOR2_X1 _14635_ ( .A1(_02503_ ), .A2(_05136_ ), .ZN(_06611_ ) );
INV_X1 _14636_ ( .A(_06611_ ), .ZN(_06612_ ) );
NOR3_X4 _14637_ ( .A1(_06612_ ), .A2(_05131_ ), .A3(_05132_ ), .ZN(_06613_ ) );
NOR2_X2 _14638_ ( .A1(_06613_ ), .A2(_05131_ ), .ZN(_06614_ ) );
OAI221_X2 _14639_ ( .A(_06610_ ), .B1(_02555_ ), .B2(_05122_ ), .C1(_05125_ ), .C2(_06614_ ), .ZN(_06615_ ) );
INV_X1 _14640_ ( .A(_05140_ ), .ZN(_06616_ ) );
OR2_X1 _14641_ ( .A1(_05104_ ), .A2(_04899_ ), .ZN(_06617_ ) );
NAND2_X1 _14642_ ( .A1(_05104_ ), .A2(_04899_ ), .ZN(_06618_ ) );
AND3_X1 _14643_ ( .A1(_06617_ ), .A2(_05097_ ), .A3(_06618_ ), .ZN(_06619_ ) );
NOR2_X1 _14644_ ( .A1(_05100_ ), .A2(_02656_ ), .ZN(_06620_ ) );
INV_X1 _14645_ ( .A(_06620_ ), .ZN(_06621_ ) );
NAND2_X1 _14646_ ( .A1(_05100_ ), .A2(_02656_ ), .ZN(_06622_ ) );
AND3_X1 _14647_ ( .A1(_06621_ ), .A2(_05110_ ), .A3(_06622_ ), .ZN(_06623_ ) );
NAND4_X1 _14648_ ( .A1(_06615_ ), .A2(_06616_ ), .A3(_06619_ ), .A4(_06623_ ), .ZN(_06624_ ) );
NOR2_X1 _14649_ ( .A1(_05096_ ), .A2(_04922_ ), .ZN(_06625_ ) );
NOR2_X1 _14650_ ( .A1(_05144_ ), .A2(_06617_ ), .ZN(_06626_ ) );
NOR2_X1 _14651_ ( .A1(_05108_ ), .A2(_02579_ ), .ZN(_06627_ ) );
AND2_X1 _14652_ ( .A1(_05108_ ), .A2(_02579_ ), .ZN(_06628_ ) );
INV_X1 _14653_ ( .A(_06628_ ), .ZN(_06629_ ) );
AOI21_X1 _14654_ ( .A(_06627_ ), .B1(_06621_ ), .B2(_06629_ ), .ZN(_06630_ ) );
AOI211_X1 _14655_ ( .A(_06625_ ), .B(_06626_ ), .C1(_06630_ ), .C2(_06619_ ), .ZN(_06631_ ) );
AND2_X2 _14656_ ( .A1(_06624_ ), .A2(_06631_ ), .ZN(_06632_ ) );
INV_X2 _14657_ ( .A(_06632_ ), .ZN(_06633_ ) );
NOR3_X1 _14658_ ( .A1(_05063_ ), .A2(_05046_ ), .A3(_05044_ ), .ZN(_06634_ ) );
AND3_X1 _14659_ ( .A1(_06634_ ), .A2(_05053_ ), .A3(_05057_ ), .ZN(_06635_ ) );
AND2_X1 _14660_ ( .A1(_05068_ ), .A2(_05072_ ), .ZN(_06636_ ) );
AND3_X1 _14661_ ( .A1(_06636_ ), .A2(_05091_ ), .A3(_05092_ ), .ZN(_06637_ ) );
NAND3_X1 _14662_ ( .A1(_06633_ ), .A2(_06635_ ), .A3(_06637_ ), .ZN(_06638_ ) );
INV_X1 _14663_ ( .A(_05082_ ), .ZN(_06639_ ) );
NOR2_X1 _14664_ ( .A1(_05080_ ), .A2(_04144_ ), .ZN(_06640_ ) );
AOI21_X1 _14665_ ( .A(_05083_ ), .B1(_06639_ ), .B2(_06640_ ), .ZN(_06641_ ) );
INV_X1 _14666_ ( .A(_06641_ ), .ZN(_06642_ ) );
NAND2_X1 _14667_ ( .A1(_06642_ ), .A2(_06636_ ), .ZN(_06643_ ) );
INV_X1 _14668_ ( .A(_02851_ ), .ZN(_06644_ ) );
NOR2_X1 _14669_ ( .A1(_06644_ ), .A2(_05071_ ), .ZN(_06645_ ) );
AOI21_X1 _14670_ ( .A(_02851_ ), .B1(_05069_ ), .B2(_05070_ ), .ZN(_06646_ ) );
INV_X1 _14671_ ( .A(_06646_ ), .ZN(_06647_ ) );
NOR2_X1 _14672_ ( .A1(_05067_ ), .A2(_04205_ ), .ZN(_06648_ ) );
AOI21_X1 _14673_ ( .A(_06645_ ), .B1(_06647_ ), .B2(_06648_ ), .ZN(_06649_ ) );
AND2_X1 _14674_ ( .A1(_06643_ ), .A2(_06649_ ), .ZN(_06650_ ) );
INV_X1 _14675_ ( .A(_06650_ ), .ZN(_06651_ ) );
NAND2_X1 _14676_ ( .A1(_06651_ ), .A2(_06635_ ), .ZN(_06652_ ) );
NOR2_X1 _14677_ ( .A1(_05038_ ), .A2(_05061_ ), .ZN(_06653_ ) );
INV_X1 _14678_ ( .A(_06653_ ), .ZN(_06654_ ) );
AOI21_X1 _14679_ ( .A(_05044_ ), .B1(_05047_ ), .B2(_06654_ ), .ZN(_06655_ ) );
NAND3_X1 _14680_ ( .A1(_06655_ ), .A2(_05053_ ), .A3(_05057_ ), .ZN(_06656_ ) );
NOR2_X1 _14681_ ( .A1(_05052_ ), .A2(_04231_ ), .ZN(_06657_ ) );
NAND2_X1 _14682_ ( .A1(_05052_ ), .A2(_04231_ ), .ZN(_06658_ ) );
INV_X1 _14683_ ( .A(_02707_ ), .ZN(_06659_ ) );
NOR2_X1 _14684_ ( .A1(_06659_ ), .A2(_05056_ ), .ZN(_06660_ ) );
AOI21_X1 _14685_ ( .A(_06657_ ), .B1(_06658_ ), .B2(_06660_ ), .ZN(_06661_ ) );
AND3_X1 _14686_ ( .A1(_06652_ ), .A2(_06656_ ), .A3(_06661_ ), .ZN(_06662_ ) );
NAND2_X2 _14687_ ( .A1(_06638_ ), .A2(_06662_ ), .ZN(_06663_ ) );
NOR2_X1 _14688_ ( .A1(_05158_ ), .A2(_05019_ ), .ZN(_06664_ ) );
NAND4_X1 _14689_ ( .A1(_06663_ ), .A2(_05010_ ), .A3(_05014_ ), .A4(_06664_ ), .ZN(_06665_ ) );
AND2_X1 _14690_ ( .A1(_05018_ ), .A2(_04723_ ), .ZN(_06666_ ) );
OR2_X1 _14691_ ( .A1(_05018_ ), .A2(_04723_ ), .ZN(_06667_ ) );
INV_X1 _14692_ ( .A(_02454_ ), .ZN(_06668_ ) );
OR2_X1 _14693_ ( .A1(_06668_ ), .A2(_05022_ ), .ZN(_06669_ ) );
AOI21_X1 _14694_ ( .A(_06666_ ), .B1(_06667_ ), .B2(_06669_ ), .ZN(_06670_ ) );
NAND3_X1 _14695_ ( .A1(_06670_ ), .A2(_05010_ ), .A3(_05014_ ), .ZN(_06671_ ) );
OR2_X1 _14696_ ( .A1(_05009_ ), .A2(_04651_ ), .ZN(_06672_ ) );
INV_X1 _14697_ ( .A(_02405_ ), .ZN(_06673_ ) );
NOR2_X1 _14698_ ( .A1(_06673_ ), .A2(_05013_ ), .ZN(_06674_ ) );
NAND2_X1 _14699_ ( .A1(_05010_ ), .A2(_06674_ ), .ZN(_06675_ ) );
AND3_X1 _14700_ ( .A1(_06671_ ), .A2(_06672_ ), .A3(_06675_ ), .ZN(_06676_ ) );
AOI21_X1 _14701_ ( .A(_05005_ ), .B1(_06665_ ), .B2(_06676_ ), .ZN(_06677_ ) );
INV_X1 _14702_ ( .A(_02329_ ), .ZN(_06678_ ) );
NOR2_X1 _14703_ ( .A1(_06678_ ), .A2(_05003_ ), .ZN(_06679_ ) );
NOR2_X1 _14704_ ( .A1(_06677_ ), .A2(_06679_ ), .ZN(_06680_ ) );
XNOR2_X1 _14705_ ( .A(_06680_ ), .B(_04999_ ), .ZN(_06681_ ) );
NOR2_X1 _14706_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06682_ ) );
INV_X1 _14707_ ( .A(_06682_ ), .ZN(_06683_ ) );
NOR2_X1 _14708_ ( .A1(_04952_ ), .A2(_06683_ ), .ZN(_06684_ ) );
BUF_X2 _14709_ ( .A(_06684_ ), .Z(_06685_ ) );
NAND2_X1 _14710_ ( .A1(_06681_ ), .A2(_06685_ ), .ZN(_06686_ ) );
AND2_X1 _14711_ ( .A1(_05205_ ), .A2(\ID_EX_typ [2] ), .ZN(_06687_ ) );
BUF_X4 _14712_ ( .A(_06687_ ), .Z(_06688_ ) );
AND4_X1 _14713_ ( .A1(_05043_ ), .A2(_05067_ ), .A3(_05061_ ), .A4(_05071_ ), .ZN(_06689_ ) );
AND2_X1 _14714_ ( .A1(_05076_ ), .A2(_05080_ ), .ZN(_06690_ ) );
NAND4_X1 _14715_ ( .A1(_06689_ ), .A2(_05096_ ), .A3(_05104_ ), .A4(_06690_ ), .ZN(_06691_ ) );
AND4_X1 _14716_ ( .A1(_05052_ ), .A2(_05018_ ), .A3(_05056_ ), .A4(_05022_ ), .ZN(_06692_ ) );
AND2_X1 _14717_ ( .A1(_05009_ ), .A2(_05013_ ), .ZN(_06693_ ) );
NAND4_X1 _14718_ ( .A1(_06692_ ), .A2(_04998_ ), .A3(_05003_ ), .A4(_06693_ ), .ZN(_06694_ ) );
NOR2_X1 _14719_ ( .A1(_06691_ ), .A2(_06694_ ), .ZN(_06695_ ) );
AND2_X1 _14720_ ( .A1(_05129_ ), .A2(_05136_ ), .ZN(_06696_ ) );
AND2_X1 _14721_ ( .A1(_06696_ ), .A2(_05119_ ), .ZN(_06697_ ) );
AND2_X1 _14722_ ( .A1(_06697_ ), .A2(_05122_ ), .ZN(_06698_ ) );
AND2_X2 _14723_ ( .A1(_06698_ ), .A2(_05100_ ), .ZN(_06699_ ) );
INV_X1 _14724_ ( .A(_05108_ ), .ZN(_06700_ ) );
OAI21_X1 _14725_ ( .A(_06695_ ), .B1(_06699_ ), .B2(_06700_ ), .ZN(_06701_ ) );
NAND2_X1 _14726_ ( .A1(_04987_ ), .A2(_04991_ ), .ZN(_06702_ ) );
NOR2_X1 _14727_ ( .A1(_06701_ ), .A2(_06702_ ), .ZN(_06703_ ) );
INV_X1 _14728_ ( .A(_06703_ ), .ZN(_06704_ ) );
NAND3_X1 _14729_ ( .A1(_06701_ ), .A2(_05036_ ), .A3(_04992_ ), .ZN(_06705_ ) );
AND4_X1 _14730_ ( .A1(_05043_ ), .A2(_05061_ ), .A3(_04998_ ), .A4(_05003_ ), .ZN(_06706_ ) );
AND2_X1 _14731_ ( .A1(_05067_ ), .A2(_05071_ ), .ZN(_06707_ ) );
AND3_X1 _14732_ ( .A1(_06706_ ), .A2(_06690_ ), .A3(_06707_ ), .ZN(_06708_ ) );
AND4_X1 _14733_ ( .A1(_05018_ ), .A2(_06708_ ), .A3(_05022_ ), .A4(_06693_ ), .ZN(_06709_ ) );
AND3_X1 _14734_ ( .A1(_06709_ ), .A2(_05052_ ), .A3(_05056_ ), .ZN(_06710_ ) );
NOR2_X1 _14735_ ( .A1(_06699_ ), .A2(_06700_ ), .ZN(_06711_ ) );
INV_X1 _14736_ ( .A(_06711_ ), .ZN(_06712_ ) );
NAND4_X1 _14737_ ( .A1(_06710_ ), .A2(_06712_ ), .A3(_05096_ ), .A4(_05104_ ), .ZN(_06713_ ) );
NAND4_X1 _14738_ ( .A1(_05050_ ), .A2(_05051_ ), .A3(_05054_ ), .A4(_05055_ ), .ZN(_06714_ ) );
OR3_X1 _14739_ ( .A1(_06714_ ), .A2(_05018_ ), .A3(_05022_ ), .ZN(_06715_ ) );
OR3_X1 _14740_ ( .A1(_06715_ ), .A2(_04998_ ), .A3(_05013_ ), .ZN(_06716_ ) );
NOR3_X1 _14741_ ( .A1(_06716_ ), .A2(_05003_ ), .A3(_05009_ ), .ZN(_06717_ ) );
INV_X1 _14742_ ( .A(_06717_ ), .ZN(_06718_ ) );
NAND4_X1 _14743_ ( .A1(_05102_ ), .A2(_05094_ ), .A3(_05095_ ), .A4(_05103_ ), .ZN(_06719_ ) );
OR3_X1 _14744_ ( .A1(_06719_ ), .A2(_05076_ ), .A3(_05080_ ), .ZN(_06720_ ) );
OR4_X1 _14745_ ( .A1(_05061_ ), .A2(_06720_ ), .A3(_05071_ ), .A4(_05067_ ), .ZN(_06721_ ) );
NOR3_X1 _14746_ ( .A1(_06718_ ), .A2(_06721_ ), .A3(_05043_ ), .ZN(_06722_ ) );
NAND2_X1 _14747_ ( .A1(_06722_ ), .A2(_06711_ ), .ZN(_06723_ ) );
AOI221_X4 _14748_ ( .A(_04963_ ), .B1(_06704_ ), .B2(_06705_ ), .C1(_06713_ ), .C2(_06723_ ), .ZN(_06724_ ) );
INV_X1 _14749_ ( .A(_04961_ ), .ZN(_06725_ ) );
NOR4_X1 _14750_ ( .A1(_06725_ ), .A2(_04980_ ), .A3(_04974_ ), .A4(_04969_ ), .ZN(_06726_ ) );
AND2_X1 _14751_ ( .A1(_05179_ ), .A2(_05185_ ), .ZN(_06727_ ) );
NAND4_X1 _14752_ ( .A1(_06726_ ), .A2(_05170_ ), .A3(_05163_ ), .A4(_06727_ ), .ZN(_06728_ ) );
OR3_X1 _14753_ ( .A1(_06701_ ), .A2(_06702_ ), .A3(_06728_ ), .ZN(_06729_ ) );
NOR4_X1 _14754_ ( .A1(_05170_ ), .A2(_05163_ ), .A3(_05179_ ), .A4(_05185_ ), .ZN(_06730_ ) );
AND4_X1 _14755_ ( .A1(_04974_ ), .A2(_06725_ ), .A3(_04980_ ), .A4(_04969_ ), .ZN(_06731_ ) );
NAND2_X1 _14756_ ( .A1(_06730_ ), .A2(_06731_ ), .ZN(_06732_ ) );
OAI21_X1 _14757_ ( .A(_06729_ ), .B1(_06703_ ), .B2(_06732_ ), .ZN(_06733_ ) );
AND2_X2 _14758_ ( .A1(_06724_ ), .A2(_06733_ ), .ZN(_06734_ ) );
XNOR2_X1 _14759_ ( .A(_06697_ ), .B(_05114_ ), .ZN(_06735_ ) );
INV_X1 _14760_ ( .A(_06735_ ), .ZN(_06736_ ) );
AND2_X1 _14761_ ( .A1(_06734_ ), .A2(_06736_ ), .ZN(_06737_ ) );
BUF_X4 _14762_ ( .A(_05120_ ), .Z(_06738_ ) );
BUF_X4 _14763_ ( .A(_06738_ ), .Z(_06739_ ) );
BUF_X4 _14764_ ( .A(_06739_ ), .Z(_06740_ ) );
BUF_X4 _14765_ ( .A(_05129_ ), .Z(_06741_ ) );
BUF_X4 _14766_ ( .A(_06741_ ), .Z(_06742_ ) );
BUF_X4 _14767_ ( .A(_05136_ ), .Z(_06743_ ) );
BUF_X4 _14768_ ( .A(_06743_ ), .Z(_06744_ ) );
XNOR2_X1 _14769_ ( .A(_06742_ ), .B(_06744_ ), .ZN(_06745_ ) );
OAI21_X1 _14770_ ( .A(_06737_ ), .B1(_06740_ ), .B2(_06745_ ), .ZN(_06746_ ) );
XNOR2_X1 _14771_ ( .A(_06698_ ), .B(_05100_ ), .ZN(_06747_ ) );
INV_X1 _14772_ ( .A(_06747_ ), .ZN(_06748_ ) );
BUF_X2 _14773_ ( .A(_06734_ ), .Z(_06749_ ) );
XNOR2_X1 _14774_ ( .A(_06699_ ), .B(_05108_ ), .ZN(_06750_ ) );
NAND2_X1 _14775_ ( .A1(_06749_ ), .A2(_06750_ ), .ZN(_06751_ ) );
NOR2_X1 _14776_ ( .A1(_06747_ ), .A2(_05108_ ), .ZN(_06752_ ) );
INV_X1 _14777_ ( .A(_06752_ ), .ZN(_06753_ ) );
AOI22_X1 _14778_ ( .A1(_06746_ ), .A2(_06748_ ), .B1(_06751_ ), .B2(_06753_ ), .ZN(_06754_ ) );
BUF_X2 _14779_ ( .A(_05120_ ), .Z(_06755_ ) );
BUF_X4 _14780_ ( .A(_06755_ ), .Z(_06756_ ) );
INV_X1 _14781_ ( .A(_05129_ ), .ZN(_06757_ ) );
BUF_X4 _14782_ ( .A(_06757_ ), .Z(_06758_ ) );
BUF_X4 _14783_ ( .A(_06743_ ), .Z(_06759_ ) );
NOR2_X1 _14784_ ( .A1(_06759_ ), .A2(_02256_ ), .ZN(_06760_ ) );
BUF_X4 _14785_ ( .A(_05134_ ), .Z(_06761_ ) );
BUF_X4 _14786_ ( .A(_06761_ ), .Z(_06762_ ) );
BUF_X4 _14787_ ( .A(_05135_ ), .Z(_06763_ ) );
BUF_X4 _14788_ ( .A(_06763_ ), .Z(_06764_ ) );
AOI21_X1 _14789_ ( .A(_02938_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06765_ ) );
NOR3_X1 _14790_ ( .A1(_06758_ ), .A2(_06760_ ), .A3(_06765_ ), .ZN(_06766_ ) );
NOR2_X1 _14791_ ( .A1(_06743_ ), .A2(_02209_ ), .ZN(_06767_ ) );
AOI21_X1 _14792_ ( .A(_04596_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06768_ ) );
BUF_X2 _14793_ ( .A(_05129_ ), .Z(_06769_ ) );
NOR3_X1 _14794_ ( .A1(_06767_ ), .A2(_06768_ ), .A3(_06769_ ), .ZN(_06770_ ) );
OAI21_X1 _14795_ ( .A(_06756_ ), .B1(_06766_ ), .B2(_06770_ ), .ZN(_06771_ ) );
NOR2_X1 _14796_ ( .A1(_06759_ ), .A2(_02305_ ), .ZN(_06772_ ) );
BUF_X4 _14797_ ( .A(_06761_ ), .Z(_06773_ ) );
BUF_X4 _14798_ ( .A(_06763_ ), .Z(_06774_ ) );
AOI21_X1 _14799_ ( .A(_04823_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06775_ ) );
OAI21_X1 _14800_ ( .A(_06741_ ), .B1(_06772_ ), .B2(_06775_ ), .ZN(_06776_ ) );
NOR2_X1 _14801_ ( .A1(_06759_ ), .A2(_02915_ ), .ZN(_06777_ ) );
AOI21_X1 _14802_ ( .A(_02282_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06778_ ) );
OAI21_X1 _14803_ ( .A(_06758_ ), .B1(_06777_ ), .B2(_06778_ ), .ZN(_06779_ ) );
BUF_X4 _14804_ ( .A(_05119_ ), .Z(_06780_ ) );
NAND3_X1 _14805_ ( .A1(_06776_ ), .A2(_06779_ ), .A3(_06780_ ), .ZN(_06781_ ) );
NAND2_X1 _14806_ ( .A1(_06771_ ), .A2(_06781_ ), .ZN(_06782_ ) );
INV_X1 _14807_ ( .A(_06743_ ), .ZN(_06783_ ) );
NAND3_X1 _14808_ ( .A1(_06783_ ), .A2(_02173_ ), .A3(_02177_ ), .ZN(_06784_ ) );
BUF_X2 _14809_ ( .A(_06743_ ), .Z(_06785_ ) );
NAND2_X1 _14810_ ( .A1(_04975_ ), .A2(_06785_ ), .ZN(_06786_ ) );
AND3_X1 _14811_ ( .A1(_06784_ ), .A2(_06769_ ), .A3(_06786_ ), .ZN(_06787_ ) );
BUF_X4 _14812_ ( .A(_06757_ ), .Z(_06788_ ) );
BUF_X4 _14813_ ( .A(_06788_ ), .Z(_06789_ ) );
AND2_X1 _14814_ ( .A1(_03006_ ), .A2(_06744_ ), .ZN(_06790_ ) );
AOI21_X1 _14815_ ( .A(_06787_ ), .B1(_06789_ ), .B2(_06790_ ), .ZN(_06791_ ) );
NOR2_X1 _14816_ ( .A1(_06791_ ), .A2(_06756_ ), .ZN(_06792_ ) );
BUF_X2 _14817_ ( .A(_05114_ ), .Z(_06793_ ) );
BUF_X2 _14818_ ( .A(_06793_ ), .Z(_06794_ ) );
MUX2_X1 _14819_ ( .A(_06782_ ), .B(_06792_ ), .S(_06794_ ), .Z(_06795_ ) );
BUF_X2 _14820_ ( .A(_05100_ ), .Z(_06796_ ) );
BUF_X2 _14821_ ( .A(_06796_ ), .Z(_06797_ ) );
AND2_X1 _14822_ ( .A1(_06795_ ), .A2(_06797_ ), .ZN(_06798_ ) );
OAI21_X1 _14823_ ( .A(_06688_ ), .B1(_06754_ ), .B2(_06798_ ), .ZN(_06799_ ) );
BUF_X4 _14824_ ( .A(_05281_ ), .Z(_06800_ ) );
BUF_X4 _14825_ ( .A(_05146_ ), .Z(_06801_ ) );
NOR2_X1 _14826_ ( .A1(_06744_ ), .A2(_02731_ ), .ZN(_06802_ ) );
AOI21_X1 _14827_ ( .A(_04283_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06803_ ) );
OR3_X1 _14828_ ( .A1(_06789_ ), .A2(_06802_ ), .A3(_06803_ ), .ZN(_06804_ ) );
NOR2_X1 _14829_ ( .A1(_06744_ ), .A2(_02828_ ), .ZN(_06805_ ) );
AOI21_X1 _14830_ ( .A(_02851_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06806_ ) );
BUF_X2 _14831_ ( .A(_06769_ ), .Z(_06807_ ) );
OR3_X1 _14832_ ( .A1(_06805_ ), .A2(_06806_ ), .A3(_06807_ ), .ZN(_06808_ ) );
BUF_X2 _14833_ ( .A(_05119_ ), .Z(_06809_ ) );
BUF_X2 _14834_ ( .A(_06809_ ), .Z(_06810_ ) );
AND3_X1 _14835_ ( .A1(_06804_ ), .A2(_06808_ ), .A3(_06810_ ), .ZN(_06811_ ) );
AOI21_X1 _14836_ ( .A(_02802_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06812_ ) );
NOR2_X1 _14837_ ( .A1(_06785_ ), .A2(_02780_ ), .ZN(_06813_ ) );
NOR3_X1 _14838_ ( .A1(_06758_ ), .A2(_06812_ ), .A3(_06813_ ), .ZN(_06814_ ) );
NOR2_X1 _14839_ ( .A1(_06785_ ), .A2(_02626_ ), .ZN(_06815_ ) );
AOI21_X1 _14840_ ( .A(_02651_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06816_ ) );
NOR3_X1 _14841_ ( .A1(_06815_ ), .A2(_06816_ ), .A3(_06769_ ), .ZN(_06817_ ) );
NOR3_X1 _14842_ ( .A1(_06814_ ), .A2(_06817_ ), .A3(_06810_ ), .ZN(_06818_ ) );
BUF_X4 _14843_ ( .A(_05122_ ), .Z(_06819_ ) );
BUF_X4 _14844_ ( .A(_06819_ ), .Z(_06820_ ) );
OR3_X1 _14845_ ( .A1(_06811_ ), .A2(_06818_ ), .A3(_06820_ ), .ZN(_06821_ ) );
BUF_X4 _14846_ ( .A(_06820_ ), .Z(_06822_ ) );
BUF_X2 _14847_ ( .A(_06780_ ), .Z(_06823_ ) );
BUF_X4 _14848_ ( .A(_06788_ ), .Z(_06824_ ) );
BUF_X4 _14849_ ( .A(_06824_ ), .Z(_06825_ ) );
NOR2_X1 _14850_ ( .A1(_06759_ ), .A2(_02454_ ), .ZN(_06826_ ) );
AOI21_X1 _14851_ ( .A(_02430_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06827_ ) );
OR3_X1 _14852_ ( .A1(_06825_ ), .A2(_06826_ ), .A3(_06827_ ), .ZN(_06828_ ) );
AOI21_X1 _14853_ ( .A(_02683_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06829_ ) );
INV_X1 _14854_ ( .A(_06829_ ), .ZN(_06830_ ) );
BUF_X4 _14855_ ( .A(_06789_ ), .Z(_06831_ ) );
OAI211_X1 _14856_ ( .A(_06830_ ), .B(_06831_ ), .C1(_02707_ ), .C2(_06744_ ), .ZN(_06832_ ) );
AOI21_X1 _14857_ ( .A(_06823_ ), .B1(_06828_ ), .B2(_06832_ ), .ZN(_06833_ ) );
AOI21_X1 _14858_ ( .A(_02382_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06834_ ) );
NOR2_X1 _14859_ ( .A1(_06785_ ), .A2(_02405_ ), .ZN(_06835_ ) );
OAI21_X1 _14860_ ( .A(_06825_ ), .B1(_06834_ ), .B2(_06835_ ), .ZN(_06836_ ) );
BUF_X2 _14861_ ( .A(_06807_ ), .Z(_06837_ ) );
NOR2_X1 _14862_ ( .A1(_06743_ ), .A2(_02329_ ), .ZN(_06838_ ) );
OAI21_X1 _14863_ ( .A(_06837_ ), .B1(_06838_ ), .B2(_06775_ ), .ZN(_06839_ ) );
AND3_X1 _14864_ ( .A1(_06836_ ), .A2(_06839_ ), .A3(_06810_ ), .ZN(_06840_ ) );
OAI21_X1 _14865_ ( .A(_06822_ ), .B1(_06833_ ), .B2(_06840_ ), .ZN(_06841_ ) );
AOI21_X1 _14866_ ( .A(_06801_ ), .B1(_06821_ ), .B2(_06841_ ), .ZN(_06842_ ) );
BUF_X2 _14867_ ( .A(_05146_ ), .Z(_06843_ ) );
NOR2_X1 _14868_ ( .A1(_06759_ ), .A2(_02603_ ), .ZN(_06844_ ) );
AOI21_X1 _14869_ ( .A(_02579_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06845_ ) );
NOR3_X1 _14870_ ( .A1(_06824_ ), .A2(_06844_ ), .A3(_06845_ ), .ZN(_06846_ ) );
NOR2_X1 _14871_ ( .A1(_06744_ ), .A2(_02549_ ), .ZN(_06847_ ) );
AOI21_X1 _14872_ ( .A(_02527_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06848_ ) );
BUF_X2 _14873_ ( .A(_05129_ ), .Z(_06849_ ) );
NOR3_X1 _14874_ ( .A1(_06847_ ), .A2(_06848_ ), .A3(_06849_ ), .ZN(_06850_ ) );
NOR2_X1 _14875_ ( .A1(_06846_ ), .A2(_06850_ ), .ZN(_06851_ ) );
BUF_X4 _14876_ ( .A(_06780_ ), .Z(_06852_ ) );
NAND2_X1 _14877_ ( .A1(_06851_ ), .A2(_06852_ ), .ZN(_06853_ ) );
BUF_X2 _14878_ ( .A(_06819_ ), .Z(_06854_ ) );
AOI21_X1 _14879_ ( .A(_02478_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06855_ ) );
NOR3_X1 _14880_ ( .A1(_06825_ ), .A2(_05137_ ), .A3(_06855_ ), .ZN(_06856_ ) );
BUF_X4 _14881_ ( .A(_06809_ ), .Z(_06857_ ) );
OR2_X1 _14882_ ( .A1(_06856_ ), .A2(_06857_ ), .ZN(_06858_ ) );
AND4_X1 _14883_ ( .A1(_06843_ ), .A2(_06853_ ), .A3(_06854_ ), .A4(_06858_ ), .ZN(_06859_ ) );
OAI21_X1 _14884_ ( .A(_06800_ ), .B1(_06842_ ), .B2(_06859_ ), .ZN(_06860_ ) );
BUF_X2 _14885_ ( .A(_05206_ ), .Z(_06861_ ) );
BUF_X2 _14886_ ( .A(_06861_ ), .Z(_06862_ ) );
NOR2_X1 _14887_ ( .A1(_04998_ ), .A2(_05032_ ), .ZN(_06863_ ) );
BUF_X4 _14888_ ( .A(_04952_ ), .Z(_06864_ ) );
AOI22_X1 _14889_ ( .A1(_04999_ ), .A2(_06862_ ), .B1(_06863_ ), .B2(_06864_ ), .ZN(_06865_ ) );
NAND4_X1 _14890_ ( .A1(_06686_ ), .A2(_06799_ ), .A3(_06860_ ), .A4(_06865_ ), .ZN(_06866_ ) );
CLKBUF_X2 _14891_ ( .A(_06797_ ), .Z(_06867_ ) );
AND2_X1 _14892_ ( .A1(_05285_ ), .A2(\ID_EX_typ [2] ), .ZN(_06868_ ) );
BUF_X2 _14893_ ( .A(_06868_ ), .Z(_06869_ ) );
BUF_X2 _14894_ ( .A(_06869_ ), .Z(_06870_ ) );
AND3_X1 _14895_ ( .A1(_06795_ ), .A2(_06867_ ), .A3(_06870_ ), .ZN(_06871_ ) );
BUF_X4 _14896_ ( .A(_05289_ ), .Z(_06872_ ) );
BUF_X4 _14897_ ( .A(_06872_ ), .Z(_06873_ ) );
AOI21_X1 _14898_ ( .A(_06873_ ), .B1(_04998_ ), .B2(_05032_ ), .ZN(_06874_ ) );
OR3_X1 _14899_ ( .A1(_06866_ ), .A2(_06871_ ), .A3(_06874_ ), .ZN(_06875_ ) );
INV_X1 _14900_ ( .A(_06594_ ), .ZN(_06876_ ) );
OAI21_X1 _14901_ ( .A(_06598_ ), .B1(_06601_ ), .B2(_06597_ ), .ZN(_06877_ ) );
NAND2_X1 _14902_ ( .A1(_06876_ ), .A2(_06877_ ), .ZN(_06878_ ) );
NOR2_X1 _14903_ ( .A1(_05296_ ), .A2(\ID_EX_typ [2] ), .ZN(_06879_ ) );
NAND3_X1 _14904_ ( .A1(_04951_ ), .A2(_06879_ ), .A3(_04957_ ), .ZN(_06880_ ) );
NAND4_X1 _14905_ ( .A1(_04089_ ), .A2(\ID_EX_typ [4] ), .A3(\ID_EX_typ [3] ), .A4(_06349_ ), .ZN(_06881_ ) );
NAND2_X1 _14906_ ( .A1(_06880_ ), .A2(_06881_ ), .ZN(_06882_ ) );
NOR2_X1 _14907_ ( .A1(_06878_ ), .A2(_06882_ ), .ZN(_06883_ ) );
NOR2_X2 _14908_ ( .A1(_06883_ ), .A2(_06584_ ), .ZN(_06884_ ) );
INV_X1 _14909_ ( .A(_06884_ ), .ZN(_06885_ ) );
BUF_X4 _14910_ ( .A(_06885_ ), .Z(_06886_ ) );
AOI21_X1 _14911_ ( .A(_06608_ ), .B1(_06875_ ), .B2(_06886_ ), .ZN(_06887_ ) );
BUF_X4 _14912_ ( .A(_06279_ ), .Z(_06888_ ) );
OAI21_X1 _14913_ ( .A(_06888_ ), .B1(_05974_ ), .B2(_05597_ ), .ZN(_06889_ ) );
OAI21_X1 _14914_ ( .A(_06581_ ), .B1(_06887_ ), .B2(_06889_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
OR2_X1 _14915_ ( .A1(_05384_ ), .A2(_06262_ ), .ZN(_06890_ ) );
BUF_X2 _14916_ ( .A(_06594_ ), .Z(_06891_ ) );
NAND3_X1 _14917_ ( .A1(_06587_ ), .A2(_06589_ ), .A3(_05256_ ), .ZN(_06892_ ) );
NAND3_X1 _14918_ ( .A1(_06590_ ), .A2(_06891_ ), .A3(_06892_ ), .ZN(_06893_ ) );
AOI22_X1 _14919_ ( .A1(_05396_ ), .A2(_06600_ ), .B1(\ID_EX_imm [20] ), .B2(_06604_ ), .ZN(_06894_ ) );
AOI21_X1 _14920_ ( .A(_06585_ ), .B1(_06893_ ), .B2(_06894_ ), .ZN(_06895_ ) );
OR2_X1 _14921_ ( .A1(_06895_ ), .A2(_06607_ ), .ZN(_06896_ ) );
BUF_X2 _14922_ ( .A(_06843_ ), .Z(_06897_ ) );
BUF_X2 _14923_ ( .A(_06793_ ), .Z(_06898_ ) );
BUF_X2 _14924_ ( .A(_06898_ ), .Z(_06899_ ) );
AOI21_X1 _14925_ ( .A(_02828_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06900_ ) );
INV_X1 _14926_ ( .A(_06900_ ), .ZN(_06901_ ) );
OAI211_X1 _14927_ ( .A(_06901_ ), .B(_06789_ ), .C1(_02802_ ), .C2(_06744_ ), .ZN(_06902_ ) );
NOR2_X1 _14928_ ( .A1(_06759_ ), .A2(_02851_ ), .ZN(_06903_ ) );
INV_X1 _14929_ ( .A(_06903_ ), .ZN(_06904_ ) );
AOI21_X1 _14930_ ( .A(_02731_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06905_ ) );
INV_X1 _14931_ ( .A(_06905_ ), .ZN(_06906_ ) );
NAND3_X1 _14932_ ( .A1(_06904_ ), .A2(_06906_ ), .A3(_06742_ ), .ZN(_06907_ ) );
AND3_X1 _14933_ ( .A1(_06902_ ), .A2(_06907_ ), .A3(_06823_ ), .ZN(_06908_ ) );
NOR2_X1 _14934_ ( .A1(_06743_ ), .A2(_02651_ ), .ZN(_06909_ ) );
AOI21_X1 _14935_ ( .A(_02780_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06910_ ) );
NOR3_X1 _14936_ ( .A1(_06788_ ), .A2(_06909_ ), .A3(_06910_ ), .ZN(_06911_ ) );
NOR2_X1 _14937_ ( .A1(_06785_ ), .A2(_02579_ ), .ZN(_06912_ ) );
AOI21_X1 _14938_ ( .A(_02626_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06913_ ) );
NOR3_X1 _14939_ ( .A1(_06912_ ), .A2(_06913_ ), .A3(_06769_ ), .ZN(_06914_ ) );
NOR3_X1 _14940_ ( .A1(_06911_ ), .A2(_06914_ ), .A3(_06823_ ), .ZN(_06915_ ) );
OAI21_X1 _14941_ ( .A(_06899_ ), .B1(_06908_ ), .B2(_06915_ ), .ZN(_06916_ ) );
BUF_X2 _14942_ ( .A(_06819_ ), .Z(_06917_ ) );
BUF_X2 _14943_ ( .A(_06917_ ), .Z(_06918_ ) );
NOR2_X1 _14944_ ( .A1(_06785_ ), .A2(_04283_ ), .ZN(_06919_ ) );
INV_X1 _14945_ ( .A(_06919_ ), .ZN(_06920_ ) );
AOI21_X1 _14946_ ( .A(_02707_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06921_ ) );
INV_X1 _14947_ ( .A(_06921_ ), .ZN(_06922_ ) );
NAND3_X1 _14948_ ( .A1(_06920_ ), .A2(_06922_ ), .A3(_06789_ ), .ZN(_06923_ ) );
NOR2_X1 _14949_ ( .A1(_06785_ ), .A2(_02683_ ), .ZN(_06924_ ) );
INV_X1 _14950_ ( .A(_06924_ ), .ZN(_06925_ ) );
AOI21_X1 _14951_ ( .A(_02454_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_06926_ ) );
INV_X1 _14952_ ( .A(_06926_ ), .ZN(_06927_ ) );
NAND3_X1 _14953_ ( .A1(_06925_ ), .A2(_06927_ ), .A3(_06807_ ), .ZN(_06928_ ) );
BUF_X2 _14954_ ( .A(_06756_ ), .Z(_06929_ ) );
AND3_X1 _14955_ ( .A1(_06923_ ), .A2(_06928_ ), .A3(_06929_ ), .ZN(_06930_ ) );
BUF_X4 _14956_ ( .A(_06742_ ), .Z(_06931_ ) );
NOR2_X1 _14957_ ( .A1(_06743_ ), .A2(_02382_ ), .ZN(_06932_ ) );
AOI21_X1 _14958_ ( .A(_02329_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06933_ ) );
OAI21_X1 _14959_ ( .A(_06931_ ), .B1(_06932_ ), .B2(_06933_ ), .ZN(_06934_ ) );
NOR2_X1 _14960_ ( .A1(_06759_ ), .A2(_02430_ ), .ZN(_06935_ ) );
AOI21_X1 _14961_ ( .A(_02405_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06936_ ) );
OAI21_X1 _14962_ ( .A(_06831_ ), .B1(_06935_ ), .B2(_06936_ ), .ZN(_06937_ ) );
AOI21_X1 _14963_ ( .A(_06929_ ), .B1(_06934_ ), .B2(_06937_ ), .ZN(_06938_ ) );
OAI21_X1 _14964_ ( .A(_06918_ ), .B1(_06930_ ), .B2(_06938_ ), .ZN(_06939_ ) );
AOI21_X1 _14965_ ( .A(_06897_ ), .B1(_06916_ ), .B2(_06939_ ), .ZN(_06940_ ) );
AND2_X1 _14966_ ( .A1(_06785_ ), .A2(_02502_ ), .ZN(_06941_ ) );
AND2_X1 _14967_ ( .A1(_06941_ ), .A2(_06849_ ), .ZN(_06942_ ) );
INV_X1 _14968_ ( .A(_06942_ ), .ZN(_06943_ ) );
NOR2_X1 _14969_ ( .A1(_06785_ ), .A2(_02527_ ), .ZN(_06944_ ) );
AOI21_X1 _14970_ ( .A(_02603_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06945_ ) );
NOR3_X1 _14971_ ( .A1(_06788_ ), .A2(_06944_ ), .A3(_06945_ ), .ZN(_06946_ ) );
NOR2_X1 _14972_ ( .A1(_06759_ ), .A2(_02478_ ), .ZN(_06947_ ) );
AOI21_X1 _14973_ ( .A(_02549_ ), .B1(_06762_ ), .B2(_06764_ ), .ZN(_06948_ ) );
NOR3_X1 _14974_ ( .A1(_06947_ ), .A2(_06948_ ), .A3(_06769_ ), .ZN(_06949_ ) );
NOR2_X1 _14975_ ( .A1(_06946_ ), .A2(_06949_ ), .ZN(_06950_ ) );
MUX2_X1 _14976_ ( .A(_06943_ ), .B(_06950_ ), .S(_06852_ ), .Z(_06951_ ) );
BUF_X2 _14977_ ( .A(_06898_ ), .Z(_06952_ ) );
NOR2_X1 _14978_ ( .A1(_06951_ ), .A2(_06952_ ), .ZN(_06953_ ) );
BUF_X4 _14979_ ( .A(_06796_ ), .Z(_06954_ ) );
BUF_X2 _14980_ ( .A(_06954_ ), .Z(_06955_ ) );
OAI21_X1 _14981_ ( .A(_06800_ ), .B1(_06953_ ), .B2(_06955_ ), .ZN(_06956_ ) );
NOR2_X1 _14982_ ( .A1(_06940_ ), .A2(_06956_ ), .ZN(_06957_ ) );
NAND2_X1 _14983_ ( .A1(_06679_ ), .A2(_06864_ ), .ZN(_06958_ ) );
BUF_X4 _14984_ ( .A(_05207_ ), .Z(_06959_ ) );
OAI21_X1 _14985_ ( .A(_06958_ ), .B1(_05005_ ), .B2(_06959_ ), .ZN(_06960_ ) );
OR4_X1 _14986_ ( .A1(_05043_ ), .A2(_05067_ ), .A3(_05061_ ), .A4(_05071_ ), .ZN(_06961_ ) );
OR4_X1 _14987_ ( .A1(_06712_ ), .A2(_06718_ ), .A3(_06720_ ), .A4(_06961_ ), .ZN(_06962_ ) );
AOI221_X4 _14988_ ( .A(_04963_ ), .B1(_06704_ ), .B2(_06705_ ), .C1(_06962_ ), .C2(_06701_ ), .ZN(_06963_ ) );
AND2_X1 _14989_ ( .A1(_06963_ ), .A2(_06733_ ), .ZN(_06964_ ) );
BUF_X2 _14990_ ( .A(_06736_ ), .Z(_06965_ ) );
BUF_X4 _14991_ ( .A(_06852_ ), .Z(_06966_ ) );
OAI21_X1 _14992_ ( .A(_06966_ ), .B1(_06831_ ), .B2(_06783_ ), .ZN(_06967_ ) );
NAND3_X1 _14993_ ( .A1(_06964_ ), .A2(_06965_ ), .A3(_06967_ ), .ZN(_06968_ ) );
AOI22_X1 _14994_ ( .A1(_06968_ ), .A2(_06748_ ), .B1(_06751_ ), .B2(_06753_ ), .ZN(_06969_ ) );
NOR2_X1 _14995_ ( .A1(_06785_ ), .A2(_04823_ ), .ZN(_06970_ ) );
OAI21_X1 _14996_ ( .A(_06741_ ), .B1(_06970_ ), .B2(_06933_ ), .ZN(_06971_ ) );
NOR2_X1 _14997_ ( .A1(_06743_ ), .A2(_02282_ ), .ZN(_06972_ ) );
AOI21_X1 _14998_ ( .A(_02305_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06973_ ) );
OAI21_X1 _14999_ ( .A(_06758_ ), .B1(_06972_ ), .B2(_06973_ ), .ZN(_06974_ ) );
AOI21_X1 _15000_ ( .A(_06755_ ), .B1(_06971_ ), .B2(_06974_ ), .ZN(_06975_ ) );
NOR2_X1 _15001_ ( .A1(_06743_ ), .A2(_02938_ ), .ZN(_06976_ ) );
AOI21_X1 _15002_ ( .A(_02915_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06977_ ) );
OAI21_X1 _15003_ ( .A(_06741_ ), .B1(_06976_ ), .B2(_06977_ ), .ZN(_06978_ ) );
NOR2_X1 _15004_ ( .A1(_05136_ ), .A2(_04596_ ), .ZN(_06979_ ) );
AOI21_X1 _15005_ ( .A(_02256_ ), .B1(_05134_ ), .B2(_05135_ ), .ZN(_06980_ ) );
OAI21_X1 _15006_ ( .A(_06758_ ), .B1(_06979_ ), .B2(_06980_ ), .ZN(_06981_ ) );
AOI21_X1 _15007_ ( .A(_06809_ ), .B1(_06978_ ), .B2(_06981_ ), .ZN(_06982_ ) );
NOR2_X1 _15008_ ( .A1(_06975_ ), .A2(_06982_ ), .ZN(_06983_ ) );
NOR2_X1 _15009_ ( .A1(_05136_ ), .A2(_02973_ ), .ZN(_06984_ ) );
AOI21_X1 _15010_ ( .A(_02209_ ), .B1(_06761_ ), .B2(_06763_ ), .ZN(_06985_ ) );
NOR3_X1 _15011_ ( .A1(_06788_ ), .A2(_06984_ ), .A3(_06985_ ), .ZN(_06986_ ) );
AND3_X1 _15012_ ( .A1(_02173_ ), .A2(_02177_ ), .A3(_05136_ ), .ZN(_06987_ ) );
AOI21_X1 _15013_ ( .A(_06987_ ), .B1(_04963_ ), .B2(_06783_ ), .ZN(_06988_ ) );
AOI21_X1 _15014_ ( .A(_06986_ ), .B1(_06988_ ), .B2(_06824_ ), .ZN(_06989_ ) );
NOR2_X1 _15015_ ( .A1(_06989_ ), .A2(_06738_ ), .ZN(_06990_ ) );
MUX2_X1 _15016_ ( .A(_06983_ ), .B(_06990_ ), .S(_06793_ ), .Z(_06991_ ) );
BUF_X2 _15017_ ( .A(_06796_ ), .Z(_06992_ ) );
AND2_X1 _15018_ ( .A1(_06991_ ), .A2(_06992_ ), .ZN(_06993_ ) );
OR2_X1 _15019_ ( .A1(_06969_ ), .A2(_06993_ ), .ZN(_06994_ ) );
BUF_X4 _15020_ ( .A(_06688_ ), .Z(_06995_ ) );
AOI211_X1 _15021_ ( .A(_06957_ ), .B(_06960_ ), .C1(_06994_ ), .C2(_06995_ ), .ZN(_06996_ ) );
INV_X1 _15022_ ( .A(_06684_ ), .ZN(_06997_ ) );
BUF_X2 _15023_ ( .A(_06997_ ), .Z(_06998_ ) );
NOR2_X1 _15024_ ( .A1(_06677_ ), .A2(_06998_ ), .ZN(_06999_ ) );
AND2_X1 _15025_ ( .A1(_06665_ ), .A2(_06676_ ), .ZN(_07000_ ) );
INV_X1 _15026_ ( .A(_07000_ ), .ZN(_07001_ ) );
OAI21_X1 _15027_ ( .A(_06999_ ), .B1(_05004_ ), .B2(_07001_ ), .ZN(_07002_ ) );
AOI21_X1 _15028_ ( .A(_06873_ ), .B1(_06678_ ), .B2(_05003_ ), .ZN(_07003_ ) );
AOI21_X1 _15029_ ( .A(_07003_ ), .B1(_06993_ ), .B2(_06870_ ), .ZN(_07004_ ) );
NAND3_X1 _15030_ ( .A1(_06996_ ), .A2(_07002_ ), .A3(_07004_ ), .ZN(_07005_ ) );
AOI21_X1 _15031_ ( .A(_06896_ ), .B1(_07005_ ), .B2(_06886_ ), .ZN(_07006_ ) );
NAND2_X1 _15032_ ( .A1(_05390_ ), .A2(_05301_ ), .ZN(_07007_ ) );
NAND2_X1 _15033_ ( .A1(_07007_ ), .A2(_06335_ ), .ZN(_07008_ ) );
OAI21_X1 _15034_ ( .A(_06890_ ), .B1(_07006_ ), .B2(_07008_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OAI21_X1 _15035_ ( .A(_06414_ ), .B1(_05417_ ), .B2(_05420_ ), .ZN(_07009_ ) );
AND2_X1 _15036_ ( .A1(_02454_ ), .A2(_04721_ ), .ZN(_07010_ ) );
AOI21_X1 _15037_ ( .A(_07010_ ), .B1(_06586_ ), .B2(_04722_ ), .ZN(_07011_ ) );
OAI21_X1 _15038_ ( .A(_05250_ ), .B1(_07011_ ), .B2(_05248_ ), .ZN(_07012_ ) );
AND2_X1 _15039_ ( .A1(_07012_ ), .A2(_04698_ ), .ZN(_07013_ ) );
AOI21_X1 _15040_ ( .A(_07013_ ), .B1(_02405_ ), .B2(_04697_ ), .ZN(_07014_ ) );
XNOR2_X1 _15041_ ( .A(_07014_ ), .B(_04675_ ), .ZN(_07015_ ) );
NAND2_X1 _15042_ ( .A1(_07015_ ), .A2(_06595_ ), .ZN(_07016_ ) );
AOI22_X1 _15043_ ( .A1(_05431_ ), .A2(_06600_ ), .B1(\ID_EX_imm [19] ), .B2(_06604_ ), .ZN(_07017_ ) );
AOI21_X1 _15044_ ( .A(_06585_ ), .B1(_07016_ ), .B2(_07017_ ), .ZN(_07018_ ) );
OR2_X1 _15045_ ( .A1(_07018_ ), .A2(_06607_ ), .ZN(_07019_ ) );
AND2_X2 _15046_ ( .A1(_06750_ ), .A2(_06747_ ), .ZN(_07020_ ) );
AND2_X1 _15047_ ( .A1(_06734_ ), .A2(_07020_ ), .ZN(_07021_ ) );
INV_X1 _15048_ ( .A(_06767_ ), .ZN(_07022_ ) );
INV_X1 _15049_ ( .A(_06768_ ), .ZN(_07023_ ) );
NAND3_X1 _15050_ ( .A1(_07022_ ), .A2(_07023_ ), .A3(_06769_ ), .ZN(_07024_ ) );
NAND3_X1 _15051_ ( .A1(_06784_ ), .A2(_06788_ ), .A3(_06786_ ), .ZN(_07025_ ) );
AOI21_X1 _15052_ ( .A(_06738_ ), .B1(_07024_ ), .B2(_07025_ ), .ZN(_07026_ ) );
AND4_X1 _15053_ ( .A1(_05116_ ), .A2(_06790_ ), .A3(_05118_ ), .A4(_06807_ ), .ZN(_07027_ ) );
OAI21_X1 _15054_ ( .A(_06793_ ), .B1(_07026_ ), .B2(_07027_ ), .ZN(_07028_ ) );
NOR3_X1 _15055_ ( .A1(_06788_ ), .A2(_06777_ ), .A3(_06778_ ), .ZN(_07029_ ) );
NOR3_X1 _15056_ ( .A1(_06760_ ), .A2(_06765_ ), .A3(_06769_ ), .ZN(_07030_ ) );
OR3_X1 _15057_ ( .A1(_07029_ ), .A2(_07030_ ), .A3(_06809_ ), .ZN(_07031_ ) );
OR3_X1 _15058_ ( .A1(_06772_ ), .A2(_06775_ ), .A3(_06849_ ), .ZN(_07032_ ) );
NOR2_X1 _15059_ ( .A1(_06834_ ), .A2(_06838_ ), .ZN(_07033_ ) );
NAND2_X1 _15060_ ( .A1(_07033_ ), .A2(_06807_ ), .ZN(_07034_ ) );
NAND3_X1 _15061_ ( .A1(_07032_ ), .A2(_07034_ ), .A3(_06780_ ), .ZN(_07035_ ) );
NAND2_X1 _15062_ ( .A1(_07031_ ), .A2(_07035_ ), .ZN(_07036_ ) );
OAI21_X1 _15063_ ( .A(_07028_ ), .B1(_07036_ ), .B2(_06794_ ), .ZN(_07037_ ) );
AND2_X1 _15064_ ( .A1(_07037_ ), .A2(_06954_ ), .ZN(_07038_ ) );
OR2_X1 _15065_ ( .A1(_07021_ ), .A2(_07038_ ), .ZN(_07039_ ) );
XNOR2_X1 _15066_ ( .A(_06696_ ), .B(_05119_ ), .ZN(_07040_ ) );
BUF_X2 _15067_ ( .A(_07040_ ), .Z(_07041_ ) );
NAND3_X1 _15068_ ( .A1(_06964_ ), .A2(_06965_ ), .A3(_07041_ ), .ZN(_07042_ ) );
INV_X1 _15069_ ( .A(_06750_ ), .ZN(_07043_ ) );
NOR2_X1 _15070_ ( .A1(_07042_ ), .A2(_07043_ ), .ZN(_07044_ ) );
OAI21_X1 _15071_ ( .A(_06688_ ), .B1(_07039_ ), .B2(_07044_ ), .ZN(_07045_ ) );
INV_X1 _15072_ ( .A(_05014_ ), .ZN(_07046_ ) );
NAND2_X1 _15073_ ( .A1(_06663_ ), .A2(_06664_ ), .ZN(_07047_ ) );
INV_X1 _15074_ ( .A(_06670_ ), .ZN(_07048_ ) );
AOI21_X1 _15075_ ( .A(_07046_ ), .B1(_07047_ ), .B2(_07048_ ), .ZN(_07049_ ) );
OR3_X1 _15076_ ( .A1(_07049_ ), .A2(_05010_ ), .A3(_06674_ ), .ZN(_07050_ ) );
OAI21_X1 _15077_ ( .A(_05010_ ), .B1(_07049_ ), .B2(_06674_ ), .ZN(_07051_ ) );
NAND3_X1 _15078_ ( .A1(_07050_ ), .A2(_06684_ ), .A3(_07051_ ), .ZN(_07052_ ) );
INV_X1 _15079_ ( .A(_06800_ ), .ZN(_07053_ ) );
NOR2_X1 _15080_ ( .A1(_06847_ ), .A2(_06848_ ), .ZN(_07054_ ) );
NOR2_X1 _15081_ ( .A1(_05137_ ), .A2(_06855_ ), .ZN(_07055_ ) );
MUX2_X1 _15082_ ( .A(_07054_ ), .B(_07055_ ), .S(_06824_ ), .Z(_07056_ ) );
NAND3_X1 _15083_ ( .A1(_07056_ ), .A2(_06819_ ), .A3(_06810_ ), .ZN(_07057_ ) );
AOI21_X1 _15084_ ( .A(_07053_ ), .B1(_07057_ ), .B2(_06897_ ), .ZN(_07058_ ) );
NOR2_X1 _15085_ ( .A1(_06759_ ), .A2(_02707_ ), .ZN(_07059_ ) );
OAI21_X1 _15086_ ( .A(_06742_ ), .B1(_07059_ ), .B2(_06829_ ), .ZN(_07060_ ) );
OAI21_X1 _15087_ ( .A(_06789_ ), .B1(_06802_ ), .B2(_06803_ ), .ZN(_07061_ ) );
NAND2_X1 _15088_ ( .A1(_07060_ ), .A2(_07061_ ), .ZN(_07062_ ) );
NOR3_X1 _15089_ ( .A1(_06789_ ), .A2(_06834_ ), .A3(_06835_ ), .ZN(_07063_ ) );
NOR3_X1 _15090_ ( .A1(_06826_ ), .A2(_06827_ ), .A3(_06807_ ), .ZN(_07064_ ) );
NOR2_X1 _15091_ ( .A1(_07063_ ), .A2(_07064_ ), .ZN(_07065_ ) );
MUX2_X1 _15092_ ( .A(_07062_ ), .B(_07065_ ), .S(_06857_ ), .Z(_07066_ ) );
OAI21_X1 _15093_ ( .A(_06992_ ), .B1(_07066_ ), .B2(_06899_ ), .ZN(_07067_ ) );
OAI21_X1 _15094_ ( .A(_06825_ ), .B1(_06812_ ), .B2(_06813_ ), .ZN(_07068_ ) );
OAI21_X1 _15095_ ( .A(_06742_ ), .B1(_06805_ ), .B2(_06806_ ), .ZN(_07069_ ) );
NAND2_X1 _15096_ ( .A1(_07068_ ), .A2(_07069_ ), .ZN(_07070_ ) );
NAND2_X1 _15097_ ( .A1(_07070_ ), .A2(_06852_ ), .ZN(_07071_ ) );
OAI21_X1 _15098_ ( .A(_06742_ ), .B1(_06815_ ), .B2(_06816_ ), .ZN(_07072_ ) );
OAI21_X1 _15099_ ( .A(_06789_ ), .B1(_06844_ ), .B2(_06845_ ), .ZN(_07073_ ) );
NAND2_X1 _15100_ ( .A1(_07072_ ), .A2(_07073_ ), .ZN(_07074_ ) );
NAND2_X1 _15101_ ( .A1(_07074_ ), .A2(_06739_ ), .ZN(_07075_ ) );
AND3_X1 _15102_ ( .A1(_07071_ ), .A2(_07075_ ), .A3(_06952_ ), .ZN(_07076_ ) );
OAI21_X1 _15103_ ( .A(_07058_ ), .B1(_07067_ ), .B2(_07076_ ), .ZN(_07077_ ) );
BUF_X4 _15104_ ( .A(_04953_ ), .Z(_07078_ ) );
NOR3_X1 _15105_ ( .A1(_05009_ ), .A2(_04651_ ), .A3(_07078_ ), .ZN(_07079_ ) );
AOI21_X1 _15106_ ( .A(_07079_ ), .B1(_05010_ ), .B2(_06862_ ), .ZN(_07080_ ) );
NAND4_X1 _15107_ ( .A1(_07045_ ), .A2(_07052_ ), .A3(_07077_ ), .A4(_07080_ ), .ZN(_07081_ ) );
AND3_X1 _15108_ ( .A1(_07037_ ), .A2(_06867_ ), .A3(_06870_ ), .ZN(_07082_ ) );
AOI21_X1 _15109_ ( .A(_06873_ ), .B1(_05009_ ), .B2(_04651_ ), .ZN(_07083_ ) );
OR3_X1 _15110_ ( .A1(_07081_ ), .A2(_07082_ ), .A3(_07083_ ), .ZN(_07084_ ) );
AOI21_X1 _15111_ ( .A(_07019_ ), .B1(_07084_ ), .B2(_06886_ ), .ZN(_07085_ ) );
NAND2_X1 _15112_ ( .A1(_05425_ ), .A2(_05301_ ), .ZN(_07086_ ) );
NAND2_X1 _15113_ ( .A1(_07086_ ), .A2(_06335_ ), .ZN(_07087_ ) );
OAI21_X1 _15114_ ( .A(_07009_ ), .B1(_07085_ ), .B2(_07087_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
OAI21_X1 _15115_ ( .A(_06414_ ), .B1(_05449_ ), .B2(_05450_ ), .ZN(_07088_ ) );
BUF_X2 _15116_ ( .A(_06876_ ), .Z(_07089_ ) );
AOI21_X1 _15117_ ( .A(_07089_ ), .B1(_07012_ ), .B2(_04698_ ), .ZN(_07090_ ) );
OAI21_X1 _15118_ ( .A(_07090_ ), .B1(_04698_ ), .B2(_07012_ ), .ZN(_07091_ ) );
AOI22_X1 _15119_ ( .A1(_05440_ ), .A2(_06600_ ), .B1(\ID_EX_imm [18] ), .B2(_06604_ ), .ZN(_07092_ ) );
AOI21_X1 _15120_ ( .A(_06585_ ), .B1(_07091_ ), .B2(_07092_ ), .ZN(_07093_ ) );
OR2_X1 _15121_ ( .A1(_07093_ ), .A2(_06607_ ), .ZN(_07094_ ) );
AND3_X1 _15122_ ( .A1(_06734_ ), .A2(_06736_ ), .A3(_07041_ ), .ZN(_07095_ ) );
AND2_X1 _15123_ ( .A1(_06783_ ), .A2(_06849_ ), .ZN(_07096_ ) );
INV_X1 _15124_ ( .A(_07096_ ), .ZN(_07097_ ) );
NAND2_X1 _15125_ ( .A1(_07095_ ), .A2(_07097_ ), .ZN(_07098_ ) );
AOI22_X1 _15126_ ( .A1(_07098_ ), .A2(_06748_ ), .B1(_06753_ ), .B2(_06751_ ), .ZN(_07099_ ) );
NAND3_X1 _15127_ ( .A1(_06988_ ), .A2(_06756_ ), .A3(_06837_ ), .ZN(_07100_ ) );
NOR3_X1 _15128_ ( .A1(_06757_ ), .A2(_06979_ ), .A3(_06980_ ), .ZN(_07101_ ) );
NOR3_X1 _15129_ ( .A1(_06984_ ), .A2(_06985_ ), .A3(_05129_ ), .ZN(_07102_ ) );
OAI21_X1 _15130_ ( .A(_06780_ ), .B1(_07101_ ), .B2(_07102_ ), .ZN(_07103_ ) );
AND2_X1 _15131_ ( .A1(_07100_ ), .A2(_07103_ ), .ZN(_07104_ ) );
OR3_X1 _15132_ ( .A1(_06788_ ), .A2(_06932_ ), .A3(_06936_ ), .ZN(_07105_ ) );
OR3_X1 _15133_ ( .A1(_06970_ ), .A2(_06933_ ), .A3(_06769_ ), .ZN(_07106_ ) );
NAND2_X1 _15134_ ( .A1(_07105_ ), .A2(_07106_ ), .ZN(_07107_ ) );
NAND2_X1 _15135_ ( .A1(_07107_ ), .A2(_06857_ ), .ZN(_07108_ ) );
OAI21_X1 _15136_ ( .A(_05129_ ), .B1(_06972_ ), .B2(_06973_ ), .ZN(_07109_ ) );
OAI21_X1 _15137_ ( .A(_06757_ ), .B1(_06976_ ), .B2(_06977_ ), .ZN(_07110_ ) );
NAND3_X1 _15138_ ( .A1(_07109_ ), .A2(_07110_ ), .A3(_06738_ ), .ZN(_07111_ ) );
AND2_X1 _15139_ ( .A1(_07108_ ), .A2(_07111_ ), .ZN(_07112_ ) );
MUX2_X1 _15140_ ( .A(_07104_ ), .B(_07112_ ), .S(_06820_ ), .Z(_07113_ ) );
NOR2_X1 _15141_ ( .A1(_07113_ ), .A2(_06897_ ), .ZN(_07114_ ) );
OAI21_X1 _15142_ ( .A(_06688_ ), .B1(_07099_ ), .B2(_07114_ ), .ZN(_07115_ ) );
AND3_X1 _15143_ ( .A1(_07047_ ), .A2(_07046_ ), .A3(_07048_ ), .ZN(_07116_ ) );
OR3_X1 _15144_ ( .A1(_07116_ ), .A2(_07049_ ), .A3(_06997_ ), .ZN(_07117_ ) );
NOR3_X1 _15145_ ( .A1(_06824_ ), .A2(_06912_ ), .A3(_06913_ ), .ZN(_07118_ ) );
NOR3_X1 _15146_ ( .A1(_06944_ ), .A2(_06945_ ), .A3(_06849_ ), .ZN(_07119_ ) );
OAI21_X1 _15147_ ( .A(_06929_ ), .B1(_07118_ ), .B2(_07119_ ), .ZN(_07120_ ) );
NOR2_X1 _15148_ ( .A1(_06759_ ), .A2(_02802_ ), .ZN(_07121_ ) );
OAI21_X1 _15149_ ( .A(_06741_ ), .B1(_07121_ ), .B2(_06900_ ), .ZN(_07122_ ) );
OAI21_X1 _15150_ ( .A(_06758_ ), .B1(_06909_ ), .B2(_06910_ ), .ZN(_07123_ ) );
NAND3_X1 _15151_ ( .A1(_07122_ ), .A2(_07123_ ), .A3(_06852_ ), .ZN(_07124_ ) );
NAND2_X1 _15152_ ( .A1(_07120_ ), .A2(_07124_ ), .ZN(_07125_ ) );
NAND2_X1 _15153_ ( .A1(_07125_ ), .A2(_06952_ ), .ZN(_07126_ ) );
OR3_X1 _15154_ ( .A1(_06824_ ), .A2(_06935_ ), .A3(_06936_ ), .ZN(_07127_ ) );
NAND3_X1 _15155_ ( .A1(_06925_ ), .A2(_06927_ ), .A3(_06789_ ), .ZN(_07128_ ) );
NAND3_X1 _15156_ ( .A1(_07127_ ), .A2(_06823_ ), .A3(_07128_ ), .ZN(_07129_ ) );
NAND3_X1 _15157_ ( .A1(_06904_ ), .A2(_06906_ ), .A3(_06789_ ), .ZN(_07130_ ) );
NAND3_X1 _15158_ ( .A1(_06920_ ), .A2(_06922_ ), .A3(_06807_ ), .ZN(_07131_ ) );
NAND3_X1 _15159_ ( .A1(_07130_ ), .A2(_07131_ ), .A3(_06929_ ), .ZN(_07132_ ) );
NAND3_X1 _15160_ ( .A1(_07129_ ), .A2(_06822_ ), .A3(_07132_ ), .ZN(_07133_ ) );
AOI21_X1 _15161_ ( .A(_06801_ ), .B1(_07126_ ), .B2(_07133_ ), .ZN(_07134_ ) );
OAI21_X1 _15162_ ( .A(_06741_ ), .B1(_06947_ ), .B2(_06948_ ), .ZN(_07135_ ) );
OAI21_X1 _15163_ ( .A(_07135_ ), .B1(_06807_ ), .B2(_06941_ ), .ZN(_07136_ ) );
BUF_X2 _15164_ ( .A(_06794_ ), .Z(_07137_ ) );
NOR4_X1 _15165_ ( .A1(_07136_ ), .A2(_06797_ ), .A3(_07137_ ), .A4(_06740_ ), .ZN(_07138_ ) );
OAI21_X1 _15166_ ( .A(_06800_ ), .B1(_07134_ ), .B2(_07138_ ), .ZN(_07139_ ) );
AOI22_X1 _15167_ ( .A1(_05014_ ), .A2(_06862_ ), .B1(_06674_ ), .B2(_06864_ ), .ZN(_07140_ ) );
NAND4_X1 _15168_ ( .A1(_07115_ ), .A2(_07117_ ), .A3(_07139_ ), .A4(_07140_ ), .ZN(_07141_ ) );
INV_X2 _15169_ ( .A(_06868_ ), .ZN(_07142_ ) );
NOR3_X1 _15170_ ( .A1(_07113_ ), .A2(_06897_ ), .A3(_07142_ ), .ZN(_07143_ ) );
AOI21_X1 _15171_ ( .A(_06873_ ), .B1(_06673_ ), .B2(_05013_ ), .ZN(_07144_ ) );
OR3_X1 _15172_ ( .A1(_07141_ ), .A2(_07143_ ), .A3(_07144_ ), .ZN(_07145_ ) );
AOI21_X1 _15173_ ( .A(_07094_ ), .B1(_07145_ ), .B2(_06886_ ), .ZN(_07146_ ) );
OAI21_X1 _15174_ ( .A(_06888_ ), .B1(_05438_ ), .B2(_05597_ ), .ZN(_07147_ ) );
OAI21_X1 _15175_ ( .A(_07088_ ), .B1(_07146_ ), .B2(_07147_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
NAND2_X1 _15176_ ( .A1(_05472_ ), .A2(_06424_ ), .ZN(_07148_ ) );
INV_X1 _15177_ ( .A(_06599_ ), .ZN(_07149_ ) );
INV_X1 _15178_ ( .A(_06603_ ), .ZN(_07150_ ) );
OAI22_X1 _15179_ ( .A1(_05480_ ), .A2(_07149_ ), .B1(_02431_ ), .B2(_07150_ ), .ZN(_07151_ ) );
XNOR2_X1 _15180_ ( .A(_07011_ ), .B(_04747_ ), .ZN(_07152_ ) );
AOI21_X1 _15181_ ( .A(_07151_ ), .B1(_07152_ ), .B2(_06595_ ), .ZN(_07153_ ) );
BUF_X4 _15182_ ( .A(_06584_ ), .Z(_07154_ ) );
OAI21_X1 _15183_ ( .A(_05360_ ), .B1(_07153_ ), .B2(_07154_ ), .ZN(_07155_ ) );
NAND4_X1 _15184_ ( .A1(_06964_ ), .A2(_06745_ ), .A3(_06965_ ), .A4(_07041_ ), .ZN(_07156_ ) );
AOI22_X1 _15185_ ( .A1(_06751_ ), .A2(_06753_ ), .B1(_06748_ ), .B2(_07156_ ), .ZN(_07157_ ) );
NAND2_X1 _15186_ ( .A1(_06791_ ), .A2(_06738_ ), .ZN(_07158_ ) );
OR3_X1 _15187_ ( .A1(_06766_ ), .A2(_06770_ ), .A3(_06755_ ), .ZN(_07159_ ) );
AOI21_X1 _15188_ ( .A(_06819_ ), .B1(_07158_ ), .B2(_07159_ ), .ZN(_07160_ ) );
NAND2_X1 _15189_ ( .A1(_07033_ ), .A2(_06758_ ), .ZN(_07161_ ) );
NOR2_X1 _15190_ ( .A1(_06835_ ), .A2(_06827_ ), .ZN(_07162_ ) );
NAND2_X1 _15191_ ( .A1(_07162_ ), .A2(_06849_ ), .ZN(_07163_ ) );
NAND2_X1 _15192_ ( .A1(_07161_ ), .A2(_07163_ ), .ZN(_07164_ ) );
NAND2_X1 _15193_ ( .A1(_07164_ ), .A2(_06809_ ), .ZN(_07165_ ) );
NAND3_X1 _15194_ ( .A1(_06776_ ), .A2(_06779_ ), .A3(_06755_ ), .ZN(_07166_ ) );
AND3_X1 _15195_ ( .A1(_07165_ ), .A2(_05122_ ), .A3(_07166_ ), .ZN(_07167_ ) );
NOR3_X1 _15196_ ( .A1(_07160_ ), .A2(_06897_ ), .A3(_07167_ ), .ZN(_07168_ ) );
OAI21_X1 _15197_ ( .A(_06995_ ), .B1(_07157_ ), .B2(_07168_ ), .ZN(_07169_ ) );
AND2_X1 _15198_ ( .A1(_06663_ ), .A2(_05157_ ), .ZN(_07170_ ) );
INV_X1 _15199_ ( .A(_07170_ ), .ZN(_07171_ ) );
AND3_X1 _15200_ ( .A1(_07171_ ), .A2(_05019_ ), .A3(_06669_ ), .ZN(_07172_ ) );
AOI21_X1 _15201_ ( .A(_05019_ ), .B1(_07171_ ), .B2(_06669_ ), .ZN(_07173_ ) );
OR3_X1 _15202_ ( .A1(_07172_ ), .A2(_07173_ ), .A3(_06998_ ), .ZN(_07174_ ) );
NOR2_X1 _15203_ ( .A1(_07160_ ), .A2(_07167_ ), .ZN(_07175_ ) );
AND3_X1 _15204_ ( .A1(_07175_ ), .A2(_06867_ ), .A3(_06869_ ), .ZN(_07176_ ) );
AND3_X1 _15205_ ( .A1(_06856_ ), .A2(_06917_ ), .A3(_06823_ ), .ZN(_07177_ ) );
OAI21_X1 _15206_ ( .A(_06800_ ), .B1(_07177_ ), .B2(_06992_ ), .ZN(_07178_ ) );
OR3_X1 _15207_ ( .A1(_06814_ ), .A2(_06817_ ), .A3(_06755_ ), .ZN(_07179_ ) );
NAND2_X1 _15208_ ( .A1(_06851_ ), .A2(_06738_ ), .ZN(_07180_ ) );
NAND2_X1 _15209_ ( .A1(_07179_ ), .A2(_07180_ ), .ZN(_07181_ ) );
AOI21_X1 _15210_ ( .A(_06929_ ), .B1(_06828_ ), .B2(_06832_ ), .ZN(_07182_ ) );
AOI21_X1 _15211_ ( .A(_06852_ ), .B1(_06804_ ), .B2(_06808_ ), .ZN(_07183_ ) );
NOR2_X1 _15212_ ( .A1(_07182_ ), .A2(_07183_ ), .ZN(_07184_ ) );
MUX2_X1 _15213_ ( .A(_07181_ ), .B(_07184_ ), .S(_06822_ ), .Z(_07185_ ) );
AOI21_X1 _15214_ ( .A(_07178_ ), .B1(_07185_ ), .B2(_06867_ ), .ZN(_07186_ ) );
BUF_X4 _15215_ ( .A(_07078_ ), .Z(_07187_ ) );
NOR3_X1 _15216_ ( .A1(_05018_ ), .A2(_04723_ ), .A3(_07187_ ), .ZN(_07188_ ) );
OAI22_X1 _15217_ ( .A1(_05019_ ), .A2(_06959_ ), .B1(_06666_ ), .B2(_06872_ ), .ZN(_07189_ ) );
NOR4_X1 _15218_ ( .A1(_07176_ ), .A2(_07186_ ), .A3(_07188_ ), .A4(_07189_ ), .ZN(_07190_ ) );
NAND3_X1 _15219_ ( .A1(_07169_ ), .A2(_07174_ ), .A3(_07190_ ), .ZN(_07191_ ) );
AOI21_X1 _15220_ ( .A(_07155_ ), .B1(_07191_ ), .B2(_06886_ ), .ZN(_07192_ ) );
OAI21_X1 _15221_ ( .A(_06888_ ), .B1(_05477_ ), .B2(_05597_ ), .ZN(_07193_ ) );
OAI21_X1 _15222_ ( .A(_07148_ ), .B1(_07192_ ), .B2(_07193_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
OR2_X1 _15223_ ( .A1(_05494_ ), .A2(_06262_ ), .ZN(_07194_ ) );
AOI21_X1 _15224_ ( .A(_07089_ ), .B1(_06586_ ), .B2(_04722_ ), .ZN(_07195_ ) );
OAI21_X1 _15225_ ( .A(_07195_ ), .B1(_04722_ ), .B2(_06586_ ), .ZN(_07196_ ) );
BUF_X2 _15226_ ( .A(_06599_ ), .Z(_07197_ ) );
NAND2_X1 _15227_ ( .A1(_05500_ ), .A2(_07197_ ), .ZN(_07198_ ) );
NAND3_X1 _15228_ ( .A1(_06601_ ), .A2(\ID_EX_imm [16] ), .A3(_06598_ ), .ZN(_07199_ ) );
AND3_X1 _15229_ ( .A1(_07196_ ), .A2(_07198_ ), .A3(_07199_ ), .ZN(_07200_ ) );
OAI21_X1 _15230_ ( .A(_05360_ ), .B1(_07200_ ), .B2(_07154_ ), .ZN(_07201_ ) );
INV_X1 _15231_ ( .A(_06698_ ), .ZN(_07202_ ) );
AOI21_X1 _15232_ ( .A(_06751_ ), .B1(_06867_ ), .B2(_07202_ ), .ZN(_07203_ ) );
NAND2_X1 _15233_ ( .A1(_06989_ ), .A2(_06756_ ), .ZN(_07204_ ) );
NAND2_X1 _15234_ ( .A1(_06978_ ), .A2(_06981_ ), .ZN(_07205_ ) );
NAND2_X1 _15235_ ( .A1(_07205_ ), .A2(_06857_ ), .ZN(_07206_ ) );
NAND3_X1 _15236_ ( .A1(_07204_ ), .A2(_06794_ ), .A3(_07206_ ), .ZN(_07207_ ) );
NOR3_X1 _15237_ ( .A1(_06824_ ), .A2(_06935_ ), .A3(_06926_ ), .ZN(_07208_ ) );
NOR3_X1 _15238_ ( .A1(_06932_ ), .A2(_06936_ ), .A3(_06741_ ), .ZN(_07209_ ) );
NOR3_X1 _15239_ ( .A1(_07208_ ), .A2(_07209_ ), .A3(_06755_ ), .ZN(_07210_ ) );
AOI21_X1 _15240_ ( .A(_06809_ ), .B1(_06971_ ), .B2(_06974_ ), .ZN(_07211_ ) );
OR3_X1 _15241_ ( .A1(_07210_ ), .A2(_06793_ ), .A3(_07211_ ), .ZN(_07212_ ) );
NAND2_X1 _15242_ ( .A1(_07207_ ), .A2(_07212_ ), .ZN(_07213_ ) );
AND2_X1 _15243_ ( .A1(_07213_ ), .A2(_06867_ ), .ZN(_07214_ ) );
OAI21_X1 _15244_ ( .A(_06995_ ), .B1(_07203_ ), .B2(_07214_ ), .ZN(_07215_ ) );
AOI21_X1 _15245_ ( .A(_06998_ ), .B1(_06663_ ), .B2(_05157_ ), .ZN(_07216_ ) );
OAI21_X1 _15246_ ( .A(_07216_ ), .B1(_05157_ ), .B2(_06663_ ), .ZN(_07217_ ) );
AND3_X1 _15247_ ( .A1(_06923_ ), .A2(_06928_ ), .A3(_06780_ ), .ZN(_07218_ ) );
AND2_X1 _15248_ ( .A1(_06902_ ), .A2(_06907_ ), .ZN(_07219_ ) );
AOI21_X1 _15249_ ( .A(_07218_ ), .B1(_06739_ ), .B2(_07219_ ), .ZN(_07220_ ) );
NOR2_X1 _15250_ ( .A1(_07220_ ), .A2(_07137_ ), .ZN(_07221_ ) );
OAI21_X1 _15251_ ( .A(_06755_ ), .B1(_06946_ ), .B2(_06949_ ), .ZN(_07222_ ) );
OAI21_X1 _15252_ ( .A(_06809_ ), .B1(_06911_ ), .B2(_06914_ ), .ZN(_07223_ ) );
AND2_X1 _15253_ ( .A1(_07222_ ), .A2(_07223_ ), .ZN(_07224_ ) );
AOI211_X1 _15254_ ( .A(_06801_ ), .B(_07221_ ), .C1(_06899_ ), .C2(_07224_ ), .ZN(_07225_ ) );
AND4_X1 _15255_ ( .A1(_06843_ ), .A2(_06942_ ), .A3(_06854_ ), .A4(_06966_ ), .ZN(_07226_ ) );
OAI21_X1 _15256_ ( .A(_06800_ ), .B1(_07225_ ), .B2(_07226_ ), .ZN(_07227_ ) );
OAI221_X1 _15257_ ( .A(_07227_ ), .B1(_06669_ ), .B2(_07187_ ), .C1(_05158_ ), .C2(_06959_ ), .ZN(_07228_ ) );
AND3_X1 _15258_ ( .A1(_07213_ ), .A2(_06867_ ), .A3(_06869_ ), .ZN(_07229_ ) );
AOI21_X1 _15259_ ( .A(_06873_ ), .B1(_06668_ ), .B2(_05022_ ), .ZN(_07230_ ) );
NOR3_X1 _15260_ ( .A1(_07228_ ), .A2(_07229_ ), .A3(_07230_ ), .ZN(_07231_ ) );
NAND3_X1 _15261_ ( .A1(_07215_ ), .A2(_07217_ ), .A3(_07231_ ), .ZN(_07232_ ) );
AOI21_X1 _15262_ ( .A(_07201_ ), .B1(_07232_ ), .B2(_06886_ ), .ZN(_07233_ ) );
NAND2_X1 _15263_ ( .A1(_05498_ ), .A2(_05891_ ), .ZN(_07234_ ) );
NAND2_X1 _15264_ ( .A1(_07234_ ), .A2(_06335_ ), .ZN(_07235_ ) );
OAI21_X1 _15265_ ( .A(_07194_ ), .B1(_07233_ ), .B2(_07235_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OAI21_X1 _15266_ ( .A(_06414_ ), .B1(_05523_ ), .B2(_05524_ ), .ZN(_07236_ ) );
NAND2_X1 _15267_ ( .A1(_05515_ ), .A2(_05891_ ), .ZN(_07237_ ) );
INV_X1 _15268_ ( .A(_05239_ ), .ZN(_07238_ ) );
NAND2_X1 _15269_ ( .A1(_07238_ ), .A2(_04230_ ), .ZN(_07239_ ) );
AND2_X1 _15270_ ( .A1(_07239_ ), .A2(_05223_ ), .ZN(_07240_ ) );
INV_X1 _15271_ ( .A(_04334_ ), .ZN(_07241_ ) );
OR2_X1 _15272_ ( .A1(_07240_ ), .A2(_07241_ ), .ZN(_07242_ ) );
AND2_X1 _15273_ ( .A1(_07242_ ), .A2(_05213_ ), .ZN(_07243_ ) );
OAI21_X1 _15274_ ( .A(_05212_ ), .B1(_07243_ ), .B2(_05210_ ), .ZN(_07244_ ) );
AND2_X1 _15275_ ( .A1(_07244_ ), .A2(_04281_ ), .ZN(_07245_ ) );
OR3_X1 _15276_ ( .A1(_07245_ ), .A2(_04256_ ), .A3(_05208_ ), .ZN(_07246_ ) );
OAI21_X1 _15277_ ( .A(_04256_ ), .B1(_07245_ ), .B2(_05208_ ), .ZN(_07247_ ) );
NAND3_X1 _15278_ ( .A1(_07246_ ), .A2(_06595_ ), .A3(_07247_ ), .ZN(_07248_ ) );
AOI22_X1 _15279_ ( .A1(_05511_ ), .A2(_07197_ ), .B1(\ID_EX_imm [15] ), .B2(_06604_ ), .ZN(_07249_ ) );
AOI21_X1 _15280_ ( .A(_06585_ ), .B1(_07248_ ), .B2(_07249_ ), .ZN(_07250_ ) );
OR2_X1 _15281_ ( .A1(_07250_ ), .A2(_05891_ ), .ZN(_07251_ ) );
NAND2_X1 _15282_ ( .A1(_07074_ ), .A2(_06810_ ), .ZN(_07252_ ) );
OAI21_X1 _15283_ ( .A(_07252_ ), .B1(_07056_ ), .B2(_06852_ ), .ZN(_07253_ ) );
NAND2_X1 _15284_ ( .A1(_07253_ ), .A2(_06952_ ), .ZN(_07254_ ) );
NAND2_X1 _15285_ ( .A1(_07062_ ), .A2(_06810_ ), .ZN(_07255_ ) );
NAND2_X1 _15286_ ( .A1(_07070_ ), .A2(_06739_ ), .ZN(_07256_ ) );
NAND2_X1 _15287_ ( .A1(_07255_ ), .A2(_07256_ ), .ZN(_07257_ ) );
NAND2_X1 _15288_ ( .A1(_07257_ ), .A2(_06918_ ), .ZN(_07258_ ) );
AND2_X1 _15289_ ( .A1(_05100_ ), .A2(_05281_ ), .ZN(_07259_ ) );
BUF_X4 _15290_ ( .A(_07259_ ), .Z(_07260_ ) );
NAND3_X1 _15291_ ( .A1(_07254_ ), .A2(_07258_ ), .A3(_07260_ ), .ZN(_07261_ ) );
INV_X1 _15292_ ( .A(_06688_ ), .ZN(_07262_ ) );
NAND2_X1 _15293_ ( .A1(_06734_ ), .A2(_07020_ ), .ZN(_07263_ ) );
NOR3_X1 _15294_ ( .A1(_07029_ ), .A2(_07030_ ), .A3(_06755_ ), .ZN(_07264_ ) );
AND3_X1 _15295_ ( .A1(_07024_ ), .A2(_07025_ ), .A3(_05120_ ), .ZN(_07265_ ) );
NOR2_X1 _15296_ ( .A1(_07264_ ), .A2(_07265_ ), .ZN(_07266_ ) );
NAND2_X1 _15297_ ( .A1(_07266_ ), .A2(_06898_ ), .ZN(_07267_ ) );
NAND3_X1 _15298_ ( .A1(_07032_ ), .A2(_07034_ ), .A3(_06756_ ), .ZN(_07268_ ) );
NAND2_X1 _15299_ ( .A1(_07162_ ), .A2(_06825_ ), .ZN(_07269_ ) );
OAI211_X1 _15300_ ( .A(_06830_ ), .B(_06742_ ), .C1(_02454_ ), .C2(_06744_ ), .ZN(_07270_ ) );
NAND3_X1 _15301_ ( .A1(_07269_ ), .A2(_07270_ ), .A3(_06857_ ), .ZN(_07271_ ) );
NAND2_X1 _15302_ ( .A1(_07268_ ), .A2(_07271_ ), .ZN(_07272_ ) );
OAI211_X1 _15303_ ( .A(_07267_ ), .B(_06954_ ), .C1(_07137_ ), .C2(_07272_ ), .ZN(_07273_ ) );
OAI21_X1 _15304_ ( .A(_06843_ ), .B1(_07202_ ), .B2(_04963_ ), .ZN(_07274_ ) );
NAND2_X1 _15305_ ( .A1(_07273_ ), .A2(_07274_ ), .ZN(_07275_ ) );
AOI21_X1 _15306_ ( .A(_07262_ ), .B1(_07263_ ), .B2(_07275_ ), .ZN(_07276_ ) );
AND3_X1 _15307_ ( .A1(_07273_ ), .A2(_06868_ ), .A3(_07274_ ), .ZN(_07277_ ) );
NOR2_X1 _15308_ ( .A1(_07276_ ), .A2(_07277_ ), .ZN(_07278_ ) );
OR3_X1 _15309_ ( .A1(_05052_ ), .A2(_04231_ ), .A3(_07078_ ), .ZN(_07279_ ) );
AOI22_X1 _15310_ ( .A1(_05053_ ), .A2(_06862_ ), .B1(_06658_ ), .B2(_05288_ ), .ZN(_07280_ ) );
AND4_X1 _15311_ ( .A1(_07261_ ), .A2(_07278_ ), .A3(_07279_ ), .A4(_07280_ ), .ZN(_07281_ ) );
INV_X1 _15312_ ( .A(_05057_ ), .ZN(_07282_ ) );
NAND2_X1 _15313_ ( .A1(_06633_ ), .A2(_06637_ ), .ZN(_07283_ ) );
AND2_X1 _15314_ ( .A1(_07283_ ), .A2(_06650_ ), .ZN(_07284_ ) );
INV_X1 _15315_ ( .A(_05059_ ), .ZN(_07285_ ) );
OR3_X1 _15316_ ( .A1(_07284_ ), .A2(_07285_ ), .A3(_05063_ ), .ZN(_07286_ ) );
INV_X1 _15317_ ( .A(_06655_ ), .ZN(_07287_ ) );
AOI21_X1 _15318_ ( .A(_07282_ ), .B1(_07286_ ), .B2(_07287_ ), .ZN(_07288_ ) );
OR3_X1 _15319_ ( .A1(_07288_ ), .A2(_05053_ ), .A3(_06660_ ), .ZN(_07289_ ) );
OAI21_X1 _15320_ ( .A(_05053_ ), .B1(_07288_ ), .B2(_06660_ ), .ZN(_07290_ ) );
NAND3_X1 _15321_ ( .A1(_07289_ ), .A2(_06685_ ), .A3(_07290_ ), .ZN(_07291_ ) );
AOI21_X1 _15322_ ( .A(_06884_ ), .B1(_07281_ ), .B2(_07291_ ), .ZN(_07292_ ) );
OAI21_X1 _15323_ ( .A(_07237_ ), .B1(_07251_ ), .B2(_07292_ ), .ZN(_07293_ ) );
OAI21_X1 _15324_ ( .A(_07236_ ), .B1(_07293_ ), .B2(_06388_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
OR2_X1 _15325_ ( .A1(_05544_ ), .A2(_06262_ ), .ZN(_07294_ ) );
AOI21_X1 _15326_ ( .A(_07089_ ), .B1(_07244_ ), .B2(_04281_ ), .ZN(_07295_ ) );
OAI21_X1 _15327_ ( .A(_07295_ ), .B1(_04281_ ), .B2(_07244_ ), .ZN(_07296_ ) );
AOI22_X1 _15328_ ( .A1(_05533_ ), .A2(_06600_ ), .B1(\ID_EX_imm [14] ), .B2(_06604_ ), .ZN(_07297_ ) );
AOI21_X1 _15329_ ( .A(_06585_ ), .B1(_07296_ ), .B2(_07297_ ), .ZN(_07298_ ) );
OR2_X1 _15330_ ( .A1(_07298_ ), .A2(_06607_ ), .ZN(_07299_ ) );
OAI211_X1 _15331_ ( .A(_06724_ ), .B(_06733_ ), .C1(_06929_ ), .C2(_07097_ ), .ZN(_07300_ ) );
INV_X1 _15332_ ( .A(_06734_ ), .ZN(_07301_ ) );
OAI21_X1 _15333_ ( .A(_07300_ ), .B1(_07301_ ), .B2(_06735_ ), .ZN(_07302_ ) );
BUF_X4 _15334_ ( .A(_07020_ ), .Z(_07303_ ) );
NAND2_X1 _15335_ ( .A1(_07302_ ), .A2(_07303_ ), .ZN(_07304_ ) );
OAI21_X1 _15336_ ( .A(_06849_ ), .B1(_06924_ ), .B2(_06921_ ), .ZN(_07305_ ) );
OAI21_X1 _15337_ ( .A(_06788_ ), .B1(_06935_ ), .B2(_06926_ ), .ZN(_07306_ ) );
NAND2_X1 _15338_ ( .A1(_07305_ ), .A2(_07306_ ), .ZN(_07307_ ) );
INV_X1 _15339_ ( .A(_07307_ ), .ZN(_07308_ ) );
MUX2_X1 _15340_ ( .A(_07308_ ), .B(_07107_ ), .S(_06738_ ), .Z(_07309_ ) );
NOR2_X1 _15341_ ( .A1(_07309_ ), .A2(_06794_ ), .ZN(_07310_ ) );
OAI21_X1 _15342_ ( .A(_05120_ ), .B1(_07101_ ), .B2(_07102_ ), .ZN(_07311_ ) );
NAND3_X1 _15343_ ( .A1(_07109_ ), .A2(_07110_ ), .A3(_05119_ ), .ZN(_07312_ ) );
AND3_X1 _15344_ ( .A1(_07311_ ), .A2(_06793_ ), .A3(_07312_ ), .ZN(_07313_ ) );
OAI21_X1 _15345_ ( .A(_06954_ ), .B1(_07310_ ), .B2(_07313_ ), .ZN(_07314_ ) );
AND3_X1 _15346_ ( .A1(_06988_ ), .A2(_05119_ ), .A3(_06769_ ), .ZN(_07315_ ) );
NAND2_X1 _15347_ ( .A1(_07315_ ), .A2(_06820_ ), .ZN(_07316_ ) );
NAND2_X1 _15348_ ( .A1(_07316_ ), .A2(_06843_ ), .ZN(_07317_ ) );
NAND2_X1 _15349_ ( .A1(_07314_ ), .A2(_07317_ ), .ZN(_07318_ ) );
AOI21_X1 _15350_ ( .A(_07262_ ), .B1(_07304_ ), .B2(_07318_ ), .ZN(_07319_ ) );
AND3_X1 _15351_ ( .A1(_07314_ ), .A2(_06868_ ), .A3(_07317_ ), .ZN(_07320_ ) );
AOI21_X1 _15352_ ( .A(_06738_ ), .B1(_07130_ ), .B2(_07131_ ), .ZN(_07321_ ) );
AND3_X1 _15353_ ( .A1(_07122_ ), .A2(_07123_ ), .A3(_06755_ ), .ZN(_07322_ ) );
OR2_X1 _15354_ ( .A1(_07321_ ), .A2(_07322_ ), .ZN(_07323_ ) );
AND2_X1 _15355_ ( .A1(_07323_ ), .A2(_06820_ ), .ZN(_07324_ ) );
NOR2_X1 _15356_ ( .A1(_07118_ ), .A2(_07119_ ), .ZN(_07325_ ) );
MUX2_X1 _15357_ ( .A(_07136_ ), .B(_07325_ ), .S(_06780_ ), .Z(_07326_ ) );
NOR2_X1 _15358_ ( .A1(_07326_ ), .A2(_06917_ ), .ZN(_07327_ ) );
NOR2_X1 _15359_ ( .A1(_07324_ ), .A2(_07327_ ), .ZN(_07328_ ) );
INV_X1 _15360_ ( .A(_07260_ ), .ZN(_07329_ ) );
NOR2_X1 _15361_ ( .A1(_07328_ ), .A2(_07329_ ), .ZN(_07330_ ) );
OR3_X1 _15362_ ( .A1(_07319_ ), .A2(_07320_ ), .A3(_07330_ ), .ZN(_07331_ ) );
AND3_X1 _15363_ ( .A1(_07286_ ), .A2(_07282_ ), .A3(_07287_ ), .ZN(_07332_ ) );
NOR3_X1 _15364_ ( .A1(_07332_ ), .A2(_07288_ ), .A3(_06998_ ), .ZN(_07333_ ) );
AND2_X1 _15365_ ( .A1(_05057_ ), .A2(_06861_ ), .ZN(_07334_ ) );
NOR3_X1 _15366_ ( .A1(_06659_ ), .A2(_05056_ ), .A3(_07078_ ), .ZN(_07335_ ) );
AOI21_X1 _15367_ ( .A(_05289_ ), .B1(_06659_ ), .B2(_05056_ ), .ZN(_07336_ ) );
OR3_X1 _15368_ ( .A1(_07334_ ), .A2(_07335_ ), .A3(_07336_ ), .ZN(_07337_ ) );
OR3_X1 _15369_ ( .A1(_07331_ ), .A2(_07333_ ), .A3(_07337_ ), .ZN(_07338_ ) );
AOI21_X1 _15370_ ( .A(_07299_ ), .B1(_06886_ ), .B2(_07338_ ), .ZN(_07339_ ) );
OAI21_X1 _15371_ ( .A(_06888_ ), .B1(_05531_ ), .B2(_05597_ ), .ZN(_07340_ ) );
OAI21_X1 _15372_ ( .A(_07294_ ), .B1(_07339_ ), .B2(_07340_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
NAND2_X1 _15373_ ( .A1(_05571_ ), .A2(_06424_ ), .ZN(_07341_ ) );
XNOR2_X1 _15374_ ( .A(_07243_ ), .B(_04308_ ), .ZN(_07342_ ) );
NAND2_X1 _15375_ ( .A1(_07342_ ), .A2(_06595_ ), .ZN(_07343_ ) );
AOI22_X1 _15376_ ( .A1(_05554_ ), .A2(_06600_ ), .B1(\ID_EX_imm [13] ), .B2(_06603_ ), .ZN(_07344_ ) );
AOI21_X1 _15377_ ( .A(_06585_ ), .B1(_07343_ ), .B2(_07344_ ), .ZN(_07345_ ) );
OR2_X1 _15378_ ( .A1(_07345_ ), .A2(_06607_ ), .ZN(_07346_ ) );
OR2_X1 _15379_ ( .A1(_07284_ ), .A2(_05063_ ), .ZN(_07347_ ) );
AND3_X1 _15380_ ( .A1(_07347_ ), .A2(_07285_ ), .A3(_06654_ ), .ZN(_07348_ ) );
AOI21_X1 _15381_ ( .A(_07285_ ), .B1(_07347_ ), .B2(_06654_ ), .ZN(_07349_ ) );
NOR3_X1 _15382_ ( .A1(_07348_ ), .A2(_07349_ ), .A3(_06998_ ), .ZN(_07350_ ) );
BUF_X4 _15383_ ( .A(_07262_ ), .Z(_07351_ ) );
NOR2_X1 _15384_ ( .A1(_06745_ ), .A2(_06739_ ), .ZN(_07352_ ) );
AND2_X1 _15385_ ( .A1(_06735_ ), .A2(_07352_ ), .ZN(_07353_ ) );
INV_X1 _15386_ ( .A(_07353_ ), .ZN(_07354_ ) );
NAND4_X1 _15387_ ( .A1(_06724_ ), .A2(_06733_ ), .A3(_07303_ ), .A4(_07354_ ), .ZN(_07355_ ) );
OAI21_X1 _15388_ ( .A(_06849_ ), .B1(_07059_ ), .B2(_06803_ ), .ZN(_07356_ ) );
OAI21_X1 _15389_ ( .A(_06788_ ), .B1(_06826_ ), .B2(_06829_ ), .ZN(_07357_ ) );
NAND2_X1 _15390_ ( .A1(_07356_ ), .A2(_07357_ ), .ZN(_07358_ ) );
INV_X1 _15391_ ( .A(_07358_ ), .ZN(_07359_ ) );
MUX2_X1 _15392_ ( .A(_07164_ ), .B(_07359_ ), .S(_06780_ ), .Z(_07360_ ) );
OR2_X1 _15393_ ( .A1(_07360_ ), .A2(_06794_ ), .ZN(_07361_ ) );
OAI211_X1 _15394_ ( .A(_07361_ ), .B(_06954_ ), .C1(_06854_ ), .C2(_06782_ ), .ZN(_07362_ ) );
NAND3_X1 _15395_ ( .A1(_06792_ ), .A2(_06843_ ), .A3(_06822_ ), .ZN(_07363_ ) );
AND2_X1 _15396_ ( .A1(_07362_ ), .A2(_07363_ ), .ZN(_07364_ ) );
AOI21_X1 _15397_ ( .A(_07351_ ), .B1(_07355_ ), .B2(_07364_ ), .ZN(_07365_ ) );
AOI21_X1 _15398_ ( .A(_07142_ ), .B1(_07362_ ), .B2(_07363_ ), .ZN(_07366_ ) );
AND3_X1 _15399_ ( .A1(_06853_ ), .A2(_06898_ ), .A3(_06858_ ), .ZN(_07367_ ) );
NOR3_X1 _15400_ ( .A1(_06811_ ), .A2(_06818_ ), .A3(_06898_ ), .ZN(_07368_ ) );
OAI21_X1 _15401_ ( .A(_07260_ ), .B1(_07367_ ), .B2(_07368_ ), .ZN(_07369_ ) );
OAI221_X1 _15402_ ( .A(_07369_ ), .B1(_05047_ ), .B2(_07078_ ), .C1(_07285_ ), .C2(_05207_ ), .ZN(_07370_ ) );
NOR4_X1 _15403_ ( .A1(_07350_ ), .A2(_07365_ ), .A3(_07366_ ), .A4(_07370_ ), .ZN(_07371_ ) );
OAI21_X1 _15404_ ( .A(_07371_ ), .B1(_05044_ ), .B2(_06873_ ), .ZN(_07372_ ) );
AOI21_X1 _15405_ ( .A(_07346_ ), .B1(_07372_ ), .B2(_06886_ ), .ZN(_07373_ ) );
OAI21_X1 _15406_ ( .A(_06888_ ), .B1(_05551_ ), .B2(_05597_ ), .ZN(_07374_ ) );
OAI21_X1 _15407_ ( .A(_07341_ ), .B1(_07373_ ), .B2(_07374_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
OR2_X1 _15408_ ( .A1(_06366_ ), .A2(_06262_ ), .ZN(_07375_ ) );
NAND3_X1 _15409_ ( .A1(_07239_ ), .A2(_07241_ ), .A3(_05223_ ), .ZN(_07376_ ) );
NAND3_X1 _15410_ ( .A1(_07242_ ), .A2(_06891_ ), .A3(_07376_ ), .ZN(_07377_ ) );
NAND3_X1 _15411_ ( .A1(_05579_ ), .A2(_05552_ ), .A3(_07197_ ), .ZN(_07378_ ) );
NAND3_X1 _15412_ ( .A1(_06601_ ), .A2(\ID_EX_imm [12] ), .A3(_06598_ ), .ZN(_07379_ ) );
AND3_X1 _15413_ ( .A1(_07377_ ), .A2(_07378_ ), .A3(_07379_ ), .ZN(_07380_ ) );
OAI21_X1 _15414_ ( .A(_05360_ ), .B1(_07380_ ), .B2(_07154_ ), .ZN(_07381_ ) );
NOR3_X1 _15415_ ( .A1(_06929_ ), .A2(_06898_ ), .A3(_06696_ ), .ZN(_07382_ ) );
INV_X1 _15416_ ( .A(_07382_ ), .ZN(_07383_ ) );
AND4_X1 _15417_ ( .A1(_06747_ ), .A2(_06964_ ), .A3(_06750_ ), .A4(_07383_ ), .ZN(_07384_ ) );
OR3_X1 _15418_ ( .A1(_07208_ ), .A2(_07209_ ), .A3(_06780_ ), .ZN(_07385_ ) );
NAND3_X1 _15419_ ( .A1(_06925_ ), .A2(_06922_ ), .A3(_06758_ ), .ZN(_07386_ ) );
NAND3_X1 _15420_ ( .A1(_06920_ ), .A2(_06906_ ), .A3(_06849_ ), .ZN(_07387_ ) );
NAND3_X1 _15421_ ( .A1(_07386_ ), .A2(_07387_ ), .A3(_06810_ ), .ZN(_07388_ ) );
NAND2_X1 _15422_ ( .A1(_07385_ ), .A2(_07388_ ), .ZN(_07389_ ) );
NAND2_X1 _15423_ ( .A1(_07389_ ), .A2(_06854_ ), .ZN(_07390_ ) );
OAI211_X1 _15424_ ( .A(_07390_ ), .B(_06992_ ), .C1(_06918_ ), .C2(_06983_ ), .ZN(_07391_ ) );
NAND3_X1 _15425_ ( .A1(_06990_ ), .A2(_06801_ ), .A3(_06918_ ), .ZN(_07392_ ) );
NAND2_X1 _15426_ ( .A1(_07391_ ), .A2(_07392_ ), .ZN(_07393_ ) );
OAI21_X1 _15427_ ( .A(_06995_ ), .B1(_07384_ ), .B2(_07393_ ), .ZN(_07394_ ) );
NAND2_X1 _15428_ ( .A1(_07393_ ), .A2(_06870_ ), .ZN(_07395_ ) );
NOR2_X1 _15429_ ( .A1(_06951_ ), .A2(_06918_ ), .ZN(_07396_ ) );
NOR3_X1 _15430_ ( .A1(_06908_ ), .A2(_06915_ ), .A3(_06952_ ), .ZN(_07397_ ) );
OAI21_X1 _15431_ ( .A(_07260_ ), .B1(_07396_ ), .B2(_07397_ ), .ZN(_07398_ ) );
AND3_X1 _15432_ ( .A1(_07394_ ), .A2(_07395_ ), .A3(_07398_ ), .ZN(_07399_ ) );
NAND3_X1 _15433_ ( .A1(_07283_ ), .A2(_05063_ ), .A3(_06650_ ), .ZN(_07400_ ) );
NAND3_X1 _15434_ ( .A1(_07347_ ), .A2(_06685_ ), .A3(_07400_ ), .ZN(_07401_ ) );
AND2_X1 _15435_ ( .A1(_05062_ ), .A2(_06862_ ), .ZN(_07402_ ) );
NOR3_X1 _15436_ ( .A1(_05038_ ), .A2(_05061_ ), .A3(_07187_ ), .ZN(_07403_ ) );
AOI21_X1 _15437_ ( .A(_06873_ ), .B1(_05038_ ), .B2(_05061_ ), .ZN(_07404_ ) );
NOR3_X1 _15438_ ( .A1(_07402_ ), .A2(_07403_ ), .A3(_07404_ ), .ZN(_07405_ ) );
NAND3_X1 _15439_ ( .A1(_07399_ ), .A2(_07401_ ), .A3(_07405_ ), .ZN(_07406_ ) );
AOI21_X1 _15440_ ( .A(_07381_ ), .B1(_07406_ ), .B2(_06886_ ), .ZN(_07407_ ) );
OAI21_X1 _15441_ ( .A(_06888_ ), .B1(_05577_ ), .B2(_05597_ ), .ZN(_07408_ ) );
OAI21_X1 _15442_ ( .A(_07375_ ), .B1(_07407_ ), .B2(_07408_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
NAND3_X1 _15443_ ( .A1(_05467_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_05561_ ), .ZN(_07409_ ) );
NAND4_X1 _15444_ ( .A1(_05568_ ), .A2(_05770_ ), .A3(\mycsreg.CSReg[0][30] ), .A4(_05771_ ), .ZN(_07410_ ) );
NAND4_X1 _15445_ ( .A1(_05564_ ), .A2(_05770_ ), .A3(\mtvec [30] ), .A4(_05771_ ), .ZN(_07411_ ) );
AND4_X1 _15446_ ( .A1(_03933_ ), .A2(_07409_ ), .A3(_07410_ ), .A4(_07411_ ), .ZN(_07412_ ) );
NAND3_X1 _15447_ ( .A1(_05365_ ), .A2(_05373_ ), .A3(_07412_ ), .ZN(_07413_ ) );
INV_X1 _15448_ ( .A(\EX_LS_result_csreg_mem [30] ), .ZN(_07414_ ) );
NAND3_X1 _15449_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(_07414_ ), .ZN(_07415_ ) );
NAND3_X1 _15450_ ( .A1(_07413_ ), .A2(_07415_ ), .A3(_06333_ ), .ZN(_07416_ ) );
OR2_X1 _15451_ ( .A1(_03973_ ), .A2(_05362_ ), .ZN(_07417_ ) );
INV_X1 _15452_ ( .A(_04970_ ), .ZN(_07418_ ) );
NOR2_X1 _15453_ ( .A1(_05171_ ), .A2(_05173_ ), .ZN(_07419_ ) );
INV_X1 _15454_ ( .A(_07419_ ), .ZN(_07420_ ) );
INV_X1 _15455_ ( .A(_05167_ ), .ZN(_07421_ ) );
AND2_X1 _15456_ ( .A1(_04999_ ), .A2(_05004_ ), .ZN(_07422_ ) );
NAND4_X1 _15457_ ( .A1(_07001_ ), .A2(_04988_ ), .A3(_04994_ ), .A4(_07422_ ), .ZN(_07423_ ) );
AND2_X1 _15458_ ( .A1(_04999_ ), .A2(_06679_ ), .ZN(_07424_ ) );
OAI211_X1 _15459_ ( .A(_04988_ ), .B(_04994_ ), .C1(_07424_ ), .C2(_06863_ ), .ZN(_07425_ ) );
OR2_X1 _15460_ ( .A1(_04987_ ), .A2(_05035_ ), .ZN(_07426_ ) );
NAND3_X1 _15461_ ( .A1(_04988_ ), .A2(_02305_ ), .A3(_04992_ ), .ZN(_07427_ ) );
AND3_X1 _15462_ ( .A1(_07425_ ), .A2(_07426_ ), .A3(_07427_ ), .ZN(_07428_ ) );
AND2_X2 _15463_ ( .A1(_07423_ ), .A2(_07428_ ), .ZN(_07429_ ) );
INV_X1 _15464_ ( .A(_07429_ ), .ZN(_07430_ ) );
NAND3_X1 _15465_ ( .A1(_07430_ ), .A2(_05182_ ), .A3(_05188_ ), .ZN(_07431_ ) );
AOI21_X1 _15466_ ( .A(_05186_ ), .B1(_05188_ ), .B2(_05180_ ), .ZN(_07432_ ) );
AOI211_X2 _15467_ ( .A(_07420_ ), .B(_07421_ ), .C1(_07431_ ), .C2(_07432_ ), .ZN(_07433_ ) );
AOI21_X1 _15468_ ( .A(_05171_ ), .B1(_05174_ ), .B2(_05165_ ), .ZN(_07434_ ) );
INV_X1 _15469_ ( .A(_07434_ ), .ZN(_07435_ ) );
OAI211_X2 _15470_ ( .A(_04976_ ), .B(_04982_ ), .C1(_07433_ ), .C2(_07435_ ), .ZN(_07436_ ) );
AND2_X1 _15471_ ( .A1(_04980_ ), .A2(_02209_ ), .ZN(_07437_ ) );
AND2_X1 _15472_ ( .A1(_07437_ ), .A2(_04976_ ), .ZN(_07438_ ) );
AOI21_X1 _15473_ ( .A(_07438_ ), .B1(_02973_ ), .B2(_04974_ ), .ZN(_07439_ ) );
AOI21_X1 _15474_ ( .A(_07418_ ), .B1(_07436_ ), .B2(_07439_ ), .ZN(_07440_ ) );
INV_X1 _15475_ ( .A(_07440_ ), .ZN(_07441_ ) );
NAND3_X1 _15476_ ( .A1(_07436_ ), .A2(_07418_ ), .A3(_07439_ ), .ZN(_07442_ ) );
NAND3_X1 _15477_ ( .A1(_07441_ ), .A2(_06685_ ), .A3(_07442_ ), .ZN(_07443_ ) );
NOR2_X1 _15478_ ( .A1(_07316_ ), .A2(_06801_ ), .ZN(_07444_ ) );
AOI21_X1 _15479_ ( .A(_07444_ ), .B1(_07302_ ), .B2(_06752_ ), .ZN(_07445_ ) );
AOI21_X1 _15480_ ( .A(_07351_ ), .B1(_07445_ ), .B2(_07263_ ), .ZN(_07446_ ) );
AOI21_X1 _15481_ ( .A(_06780_ ), .B1(_07127_ ), .B2(_07128_ ), .ZN(_07447_ ) );
OAI21_X1 _15482_ ( .A(_06741_ ), .B1(_06970_ ), .B2(_06973_ ), .ZN(_07448_ ) );
OAI21_X1 _15483_ ( .A(_06824_ ), .B1(_06932_ ), .B2(_06933_ ), .ZN(_07449_ ) );
AND3_X1 _15484_ ( .A1(_07448_ ), .A2(_07449_ ), .A3(_06809_ ), .ZN(_07450_ ) );
OR3_X1 _15485_ ( .A1(_07447_ ), .A2(_06917_ ), .A3(_07450_ ), .ZN(_07451_ ) );
OAI21_X1 _15486_ ( .A(_06931_ ), .B1(_06976_ ), .B2(_06980_ ), .ZN(_07452_ ) );
OAI21_X1 _15487_ ( .A(_06831_ ), .B1(_06972_ ), .B2(_06977_ ), .ZN(_07453_ ) );
NAND3_X1 _15488_ ( .A1(_07452_ ), .A2(_07453_ ), .A3(_06740_ ), .ZN(_07454_ ) );
NOR3_X1 _15489_ ( .A1(_06987_ ), .A2(_06831_ ), .A3(_06984_ ), .ZN(_07455_ ) );
NOR2_X1 _15490_ ( .A1(_06979_ ), .A2(_06985_ ), .ZN(_07456_ ) );
AOI21_X1 _15491_ ( .A(_07455_ ), .B1(_06831_ ), .B2(_07456_ ), .ZN(_07457_ ) );
OAI21_X1 _15492_ ( .A(_07454_ ), .B1(_07457_ ), .B2(_06740_ ), .ZN(_07458_ ) );
OAI211_X1 _15493_ ( .A(_07451_ ), .B(_06955_ ), .C1(_07458_ ), .C2(_06899_ ), .ZN(_07459_ ) );
OAI21_X1 _15494_ ( .A(_06897_ ), .B1(_07324_ ), .B2(_07327_ ), .ZN(_07460_ ) );
AOI21_X1 _15495_ ( .A(_07053_ ), .B1(_07459_ ), .B2(_07460_ ), .ZN(_07461_ ) );
INV_X1 _15496_ ( .A(_04969_ ), .ZN(_07462_ ) );
AOI21_X1 _15497_ ( .A(_06872_ ), .B1(_02178_ ), .B2(_07462_ ), .ZN(_07463_ ) );
OR3_X1 _15498_ ( .A1(_07316_ ), .A2(_06843_ ), .A3(_07142_ ), .ZN(_07464_ ) );
AOI21_X1 _15499_ ( .A(_07462_ ), .B1(_02173_ ), .B2(_02177_ ), .ZN(_07465_ ) );
INV_X1 _15500_ ( .A(_07465_ ), .ZN(_07466_ ) );
OAI221_X1 _15501_ ( .A(_07464_ ), .B1(_07466_ ), .B2(_07078_ ), .C1(_07418_ ), .C2(_05207_ ), .ZN(_07467_ ) );
NOR4_X1 _15502_ ( .A1(_07446_ ), .A2(_07461_ ), .A3(_07463_ ), .A4(_07467_ ), .ZN(_07468_ ) );
AOI21_X1 _15503_ ( .A(_06884_ ), .B1(_07443_ ), .B2(_07468_ ), .ZN(_07469_ ) );
NAND2_X1 _15504_ ( .A1(_06586_ ), .A2(_04850_ ), .ZN(_07470_ ) );
AND2_X1 _15505_ ( .A1(_07470_ ), .A2(_05261_ ), .ZN(_07471_ ) );
INV_X1 _15506_ ( .A(_07471_ ), .ZN(_07472_ ) );
AOI21_X1 _15507_ ( .A(_05275_ ), .B1(_07472_ ), .B2(_04649_ ), .ZN(_07473_ ) );
NOR3_X1 _15508_ ( .A1(_07473_ ), .A2(_04598_ ), .A3(_04573_ ), .ZN(_07474_ ) );
OAI21_X1 _15509_ ( .A(_04546_ ), .B1(_07474_ ), .B2(_05273_ ), .ZN(_07475_ ) );
AND3_X1 _15510_ ( .A1(_07475_ ), .A2(_05264_ ), .A3(_05268_ ), .ZN(_07476_ ) );
AOI21_X1 _15511_ ( .A(_05264_ ), .B1(_07475_ ), .B2(_05268_ ), .ZN(_07477_ ) );
OR3_X1 _15512_ ( .A1(_07476_ ), .A2(_07477_ ), .A3(_07089_ ), .ZN(_07478_ ) );
AOI22_X1 _15513_ ( .A1(_04088_ ), .A2(_07197_ ), .B1(\ID_EX_imm [30] ), .B2(_06604_ ), .ZN(_07479_ ) );
AOI21_X1 _15514_ ( .A(_06585_ ), .B1(_07478_ ), .B2(_07479_ ), .ZN(_07480_ ) );
OR2_X1 _15515_ ( .A1(_07480_ ), .A2(_05891_ ), .ZN(_07481_ ) );
OAI21_X1 _15516_ ( .A(_07417_ ), .B1(_07469_ ), .B2(_07481_ ), .ZN(_07482_ ) );
OAI21_X1 _15517_ ( .A(_07416_ ), .B1(_07482_ ), .B2(_06388_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
AND2_X1 _15518_ ( .A1(_04228_ ), .A2(_02828_ ), .ZN(_07483_ ) );
AOI21_X1 _15519_ ( .A(_05216_ ), .B1(_07238_ ), .B2(_04176_ ), .ZN(_07484_ ) );
OAI21_X1 _15520_ ( .A(_05218_ ), .B1(_07484_ ), .B2(_04142_ ), .ZN(_07485_ ) );
AOI21_X1 _15521_ ( .A(_07483_ ), .B1(_07485_ ), .B2(_04229_ ), .ZN(_07486_ ) );
XNOR2_X1 _15522_ ( .A(_07486_ ), .B(_04204_ ), .ZN(_07487_ ) );
AND2_X1 _15523_ ( .A1(_07487_ ), .A2(_06595_ ), .ZN(_07488_ ) );
NAND2_X1 _15524_ ( .A1(_05614_ ), .A2(_07197_ ), .ZN(_07489_ ) );
OAI21_X1 _15525_ ( .A(_07489_ ), .B1(_02852_ ), .B2(_07150_ ), .ZN(_07490_ ) );
OAI21_X1 _15526_ ( .A(_06583_ ), .B1(_07488_ ), .B2(_07490_ ), .ZN(_07491_ ) );
BUF_X4 _15527_ ( .A(_03878_ ), .Z(_07492_ ) );
OAI211_X1 _15528_ ( .A(_06749_ ), .B(_07303_ ), .C1(_06965_ ), .C2(_07041_ ), .ZN(_07493_ ) );
OAI21_X1 _15529_ ( .A(_06807_ ), .B1(_06802_ ), .B2(_06806_ ), .ZN(_07494_ ) );
OAI21_X1 _15530_ ( .A(_06824_ ), .B1(_07059_ ), .B2(_06803_ ), .ZN(_07495_ ) );
NAND2_X1 _15531_ ( .A1(_07494_ ), .A2(_07495_ ), .ZN(_07496_ ) );
NAND2_X1 _15532_ ( .A1(_07496_ ), .A2(_06823_ ), .ZN(_07497_ ) );
NAND3_X1 _15533_ ( .A1(_07269_ ), .A2(_07270_ ), .A3(_06929_ ), .ZN(_07498_ ) );
NAND3_X1 _15534_ ( .A1(_07497_ ), .A2(_07498_ ), .A3(_06854_ ), .ZN(_07499_ ) );
OAI211_X1 _15535_ ( .A(_06992_ ), .B(_07499_ ), .C1(_07036_ ), .C2(_06822_ ), .ZN(_07500_ ) );
OAI21_X1 _15536_ ( .A(_06819_ ), .B1(_07026_ ), .B2(_07027_ ), .ZN(_07501_ ) );
NAND2_X1 _15537_ ( .A1(_07501_ ), .A2(_06897_ ), .ZN(_07502_ ) );
NAND2_X1 _15538_ ( .A1(_07500_ ), .A2(_07502_ ), .ZN(_07503_ ) );
AOI21_X1 _15539_ ( .A(_07351_ ), .B1(_07493_ ), .B2(_07503_ ), .ZN(_07504_ ) );
INV_X1 _15540_ ( .A(_05091_ ), .ZN(_07505_ ) );
INV_X1 _15541_ ( .A(_05092_ ), .ZN(_07506_ ) );
NOR3_X1 _15542_ ( .A1(_06632_ ), .A2(_07505_ ), .A3(_07506_ ), .ZN(_07507_ ) );
NOR2_X1 _15543_ ( .A1(_07507_ ), .A2(_06642_ ), .ZN(_07508_ ) );
INV_X1 _15544_ ( .A(_05068_ ), .ZN(_07509_ ) );
NOR2_X1 _15545_ ( .A1(_07508_ ), .A2(_07509_ ), .ZN(_07510_ ) );
OAI21_X1 _15546_ ( .A(_05072_ ), .B1(_07510_ ), .B2(_06648_ ), .ZN(_07511_ ) );
INV_X1 _15547_ ( .A(_06648_ ), .ZN(_07512_ ) );
OAI211_X1 _15548_ ( .A(_05087_ ), .B(_07512_ ), .C1(_07508_ ), .C2(_07509_ ), .ZN(_07513_ ) );
AND3_X1 _15549_ ( .A1(_07511_ ), .A2(_06684_ ), .A3(_07513_ ), .ZN(_07514_ ) );
NAND3_X1 _15550_ ( .A1(_07500_ ), .A2(_06869_ ), .A3(_07502_ ), .ZN(_07515_ ) );
NAND2_X1 _15551_ ( .A1(_06645_ ), .A2(_06864_ ), .ZN(_07516_ ) );
AOI22_X1 _15552_ ( .A1(_05072_ ), .A2(_06861_ ), .B1(_06647_ ), .B2(_05288_ ), .ZN(_07517_ ) );
NAND3_X1 _15553_ ( .A1(_07071_ ), .A2(_07075_ ), .A3(_06917_ ), .ZN(_07518_ ) );
NAND3_X1 _15554_ ( .A1(_07056_ ), .A2(_06898_ ), .A3(_06823_ ), .ZN(_07519_ ) );
NAND2_X1 _15555_ ( .A1(_07518_ ), .A2(_07519_ ), .ZN(_07520_ ) );
NAND2_X1 _15556_ ( .A1(_07520_ ), .A2(_07260_ ), .ZN(_07521_ ) );
NAND4_X1 _15557_ ( .A1(_07515_ ), .A2(_07516_ ), .A3(_07517_ ), .A4(_07521_ ), .ZN(_07522_ ) );
NOR3_X1 _15558_ ( .A1(_07504_ ), .A2(_07514_ ), .A3(_07522_ ), .ZN(_07523_ ) );
OAI211_X1 _15559_ ( .A(_07491_ ), .B(_07492_ ), .C1(_06884_ ), .C2(_07523_ ), .ZN(_07524_ ) );
NAND2_X1 _15560_ ( .A1(_05608_ ), .A2(_05301_ ), .ZN(_07525_ ) );
NAND3_X1 _15561_ ( .A1(_07524_ ), .A2(_06280_ ), .A3(_07525_ ), .ZN(_07526_ ) );
NAND2_X1 _15562_ ( .A1(_05606_ ), .A2(_06266_ ), .ZN(_07527_ ) );
NAND2_X1 _15563_ ( .A1(_07526_ ), .A2(_07527_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OAI21_X1 _15564_ ( .A(_06414_ ), .B1(_05651_ ), .B2(_05652_ ), .ZN(_07528_ ) );
AOI21_X1 _15565_ ( .A(_07089_ ), .B1(_07485_ ), .B2(_04229_ ), .ZN(_07529_ ) );
OAI21_X1 _15566_ ( .A(_07529_ ), .B1(_04229_ ), .B2(_07485_ ), .ZN(_07530_ ) );
AOI22_X1 _15567_ ( .A1(_05640_ ), .A2(_06600_ ), .B1(\ID_EX_imm [10] ), .B2(_06603_ ), .ZN(_07531_ ) );
AOI21_X1 _15568_ ( .A(_06584_ ), .B1(_07530_ ), .B2(_07531_ ), .ZN(_07532_ ) );
OR2_X1 _15569_ ( .A1(_07532_ ), .A2(_06607_ ), .ZN(_07533_ ) );
AND4_X1 _15570_ ( .A1(_07097_ ), .A2(_06724_ ), .A3(_06733_ ), .A4(_07041_ ), .ZN(_07534_ ) );
OAI21_X1 _15571_ ( .A(_07303_ ), .B1(_06737_ ), .B2(_07534_ ), .ZN(_07535_ ) );
NAND3_X1 _15572_ ( .A1(_07108_ ), .A2(_06794_ ), .A3(_07111_ ), .ZN(_07536_ ) );
NAND3_X1 _15573_ ( .A1(_07305_ ), .A2(_07306_ ), .A3(_06756_ ), .ZN(_07537_ ) );
OAI21_X1 _15574_ ( .A(_06742_ ), .B1(_06903_ ), .B2(_06900_ ), .ZN(_07538_ ) );
OAI21_X1 _15575_ ( .A(_06825_ ), .B1(_06919_ ), .B2(_06905_ ), .ZN(_07539_ ) );
NAND3_X1 _15576_ ( .A1(_07538_ ), .A2(_07539_ ), .A3(_06857_ ), .ZN(_07540_ ) );
NAND3_X1 _15577_ ( .A1(_07537_ ), .A2(_07540_ ), .A3(_06819_ ), .ZN(_07541_ ) );
NAND3_X1 _15578_ ( .A1(_07536_ ), .A2(_06796_ ), .A3(_07541_ ), .ZN(_07542_ ) );
AOI21_X1 _15579_ ( .A(_06794_ ), .B1(_07100_ ), .B2(_07103_ ), .ZN(_07543_ ) );
NAND2_X1 _15580_ ( .A1(_07543_ ), .A2(_05146_ ), .ZN(_07544_ ) );
AND2_X1 _15581_ ( .A1(_07542_ ), .A2(_07544_ ), .ZN(_07545_ ) );
AOI21_X1 _15582_ ( .A(_07262_ ), .B1(_07535_ ), .B2(_07545_ ), .ZN(_07546_ ) );
AOI21_X1 _15583_ ( .A(_07142_ ), .B1(_07542_ ), .B2(_07544_ ), .ZN(_07547_ ) );
NAND2_X1 _15584_ ( .A1(_07125_ ), .A2(_06822_ ), .ZN(_07548_ ) );
OR3_X1 _15585_ ( .A1(_07136_ ), .A2(_06820_ ), .A3(_06739_ ), .ZN(_07549_ ) );
AOI21_X1 _15586_ ( .A(_07329_ ), .B1(_07548_ ), .B2(_07549_ ), .ZN(_07550_ ) );
OR3_X1 _15587_ ( .A1(_07546_ ), .A2(_07547_ ), .A3(_07550_ ), .ZN(_07551_ ) );
OAI21_X1 _15588_ ( .A(_06684_ ), .B1(_07508_ ), .B2(_07509_ ), .ZN(_07552_ ) );
AOI21_X1 _15589_ ( .A(_07552_ ), .B1(_07509_ ), .B2(_07508_ ), .ZN(_07553_ ) );
AND2_X1 _15590_ ( .A1(_05068_ ), .A2(_06861_ ), .ZN(_07554_ ) );
AOI21_X1 _15591_ ( .A(_05289_ ), .B1(_05067_ ), .B2(_04205_ ), .ZN(_07555_ ) );
NOR3_X1 _15592_ ( .A1(_05067_ ), .A2(_04205_ ), .A3(_07078_ ), .ZN(_07556_ ) );
OR3_X1 _15593_ ( .A1(_07554_ ), .A2(_07555_ ), .A3(_07556_ ), .ZN(_07557_ ) );
OR3_X1 _15594_ ( .A1(_07551_ ), .A2(_07553_ ), .A3(_07557_ ), .ZN(_07558_ ) );
AOI21_X1 _15595_ ( .A(_07533_ ), .B1(_07558_ ), .B2(_06886_ ), .ZN(_07559_ ) );
NAND2_X1 _15596_ ( .A1(_05642_ ), .A2(_05891_ ), .ZN(_07560_ ) );
NAND2_X1 _15597_ ( .A1(_07560_ ), .A2(_06335_ ), .ZN(_07561_ ) );
OAI21_X1 _15598_ ( .A(_07528_ ), .B1(_07559_ ), .B2(_07561_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
OAI21_X1 _15599_ ( .A(_06414_ ), .B1(_05670_ ), .B2(_05671_ ), .ZN(_07562_ ) );
XNOR2_X1 _15600_ ( .A(_07484_ ), .B(_04143_ ), .ZN(_07563_ ) );
NAND2_X1 _15601_ ( .A1(_07563_ ), .A2(_06595_ ), .ZN(_07564_ ) );
AOI22_X1 _15602_ ( .A1(_05660_ ), .A2(_06600_ ), .B1(\ID_EX_imm [9] ), .B2(_06603_ ), .ZN(_07565_ ) );
AOI21_X1 _15603_ ( .A(_06584_ ), .B1(_07564_ ), .B2(_07565_ ), .ZN(_07566_ ) );
OR2_X1 _15604_ ( .A1(_07566_ ), .A2(_06607_ ), .ZN(_07567_ ) );
AND2_X1 _15605_ ( .A1(_06964_ ), .A2(_06965_ ), .ZN(_07568_ ) );
AND4_X1 _15606_ ( .A1(_06745_ ), .A2(_06963_ ), .A3(_06733_ ), .A4(_07041_ ), .ZN(_07569_ ) );
OAI21_X1 _15607_ ( .A(_07303_ ), .B1(_07568_ ), .B2(_07569_ ), .ZN(_07570_ ) );
NAND3_X1 _15608_ ( .A1(_07165_ ), .A2(_06898_ ), .A3(_07166_ ), .ZN(_07571_ ) );
OAI21_X1 _15609_ ( .A(_06742_ ), .B1(_06812_ ), .B2(_06805_ ), .ZN(_07572_ ) );
OAI21_X1 _15610_ ( .A(_06825_ ), .B1(_06802_ ), .B2(_06806_ ), .ZN(_07573_ ) );
AOI21_X1 _15611_ ( .A(_06756_ ), .B1(_07572_ ), .B2(_07573_ ), .ZN(_07574_ ) );
AOI21_X1 _15612_ ( .A(_07574_ ), .B1(_06739_ ), .B2(_07358_ ), .ZN(_07575_ ) );
OAI211_X1 _15613_ ( .A(_07571_ ), .B(_06954_ ), .C1(_07137_ ), .C2(_07575_ ), .ZN(_07576_ ) );
NAND4_X1 _15614_ ( .A1(_07158_ ), .A2(_06843_ ), .A3(_06854_ ), .A4(_07159_ ), .ZN(_07577_ ) );
AND2_X1 _15615_ ( .A1(_07576_ ), .A2(_07577_ ), .ZN(_07578_ ) );
AOI21_X1 _15616_ ( .A(_07351_ ), .B1(_07570_ ), .B2(_07578_ ), .ZN(_07579_ ) );
AOI21_X1 _15617_ ( .A(_07506_ ), .B1(_06624_ ), .B2(_06631_ ), .ZN(_07580_ ) );
OR3_X1 _15618_ ( .A1(_07580_ ), .A2(_05091_ ), .A3(_06640_ ), .ZN(_07581_ ) );
OAI21_X1 _15619_ ( .A(_05091_ ), .B1(_07580_ ), .B2(_06640_ ), .ZN(_07582_ ) );
AND3_X1 _15620_ ( .A1(_07581_ ), .A2(_06684_ ), .A3(_07582_ ), .ZN(_07583_ ) );
NAND3_X1 _15621_ ( .A1(_07179_ ), .A2(_07180_ ), .A3(_06819_ ), .ZN(_07584_ ) );
NAND4_X1 _15622_ ( .A1(_07055_ ), .A2(_06793_ ), .A3(_06857_ ), .A4(_06837_ ), .ZN(_07585_ ) );
AOI21_X1 _15623_ ( .A(_07329_ ), .B1(_07584_ ), .B2(_07585_ ), .ZN(_07586_ ) );
AOI221_X4 _15624_ ( .A(_07586_ ), .B1(_05083_ ), .B2(_04952_ ), .C1(_05091_ ), .C2(_06861_ ), .ZN(_07587_ ) );
OAI221_X1 _15625_ ( .A(_07587_ ), .B1(_05082_ ), .B2(_06872_ ), .C1(_07142_ ), .C2(_07578_ ), .ZN(_07588_ ) );
OR3_X1 _15626_ ( .A1(_07579_ ), .A2(_07583_ ), .A3(_07588_ ), .ZN(_07589_ ) );
BUF_X4 _15627_ ( .A(_06885_ ), .Z(_07590_ ) );
AOI21_X1 _15628_ ( .A(_07567_ ), .B1(_07589_ ), .B2(_07590_ ), .ZN(_07591_ ) );
NAND2_X1 _15629_ ( .A1(_05662_ ), .A2(_05891_ ), .ZN(_07592_ ) );
NAND2_X1 _15630_ ( .A1(_07592_ ), .A2(_06335_ ), .ZN(_07593_ ) );
OAI21_X1 _15631_ ( .A(_07562_ ), .B1(_07591_ ), .B2(_07593_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
AND2_X1 _15632_ ( .A1(_05690_ ), .A2(_03877_ ), .ZN(_07594_ ) );
NOR2_X1 _15633_ ( .A1(_06697_ ), .A2(_06898_ ), .ZN(_07595_ ) );
INV_X1 _15634_ ( .A(_07595_ ), .ZN(_07596_ ) );
NAND4_X1 _15635_ ( .A1(_06724_ ), .A2(_07596_ ), .A3(_06733_ ), .A4(_07303_ ), .ZN(_07597_ ) );
OAI21_X1 _15636_ ( .A(_06793_ ), .B1(_07210_ ), .B2(_07211_ ), .ZN(_07598_ ) );
AND3_X1 _15637_ ( .A1(_07386_ ), .A2(_07387_ ), .A3(_06755_ ), .ZN(_07599_ ) );
NOR3_X1 _15638_ ( .A1(_06758_ ), .A2(_07121_ ), .A3(_06910_ ), .ZN(_07600_ ) );
NOR3_X1 _15639_ ( .A1(_06903_ ), .A2(_06900_ ), .A3(_06849_ ), .ZN(_07601_ ) );
NOR2_X1 _15640_ ( .A1(_07600_ ), .A2(_07601_ ), .ZN(_07602_ ) );
AOI21_X1 _15641_ ( .A(_07599_ ), .B1(_06857_ ), .B2(_07602_ ), .ZN(_07603_ ) );
OAI211_X1 _15642_ ( .A(_06796_ ), .B(_07598_ ), .C1(_07603_ ), .C2(_06794_ ), .ZN(_07604_ ) );
NAND4_X1 _15643_ ( .A1(_07204_ ), .A2(_05146_ ), .A3(_06819_ ), .A4(_07206_ ), .ZN(_07605_ ) );
AND2_X1 _15644_ ( .A1(_07604_ ), .A2(_07605_ ), .ZN(_07606_ ) );
AOI21_X1 _15645_ ( .A(_07262_ ), .B1(_07597_ ), .B2(_07606_ ), .ZN(_07607_ ) );
NAND3_X1 _15646_ ( .A1(_07222_ ), .A2(_07223_ ), .A3(_05122_ ), .ZN(_07608_ ) );
OAI21_X1 _15647_ ( .A(_05114_ ), .B1(_06943_ ), .B2(_06738_ ), .ZN(_07609_ ) );
AND3_X1 _15648_ ( .A1(_07608_ ), .A2(_07260_ ), .A3(_07609_ ), .ZN(_07610_ ) );
AND2_X1 _15649_ ( .A1(_05092_ ), .A2(_06861_ ), .ZN(_07611_ ) );
NOR3_X1 _15650_ ( .A1(_05080_ ), .A2(_04144_ ), .A3(_04953_ ), .ZN(_07612_ ) );
OR3_X1 _15651_ ( .A1(_07610_ ), .A2(_07611_ ), .A3(_07612_ ), .ZN(_07613_ ) );
AOI21_X1 _15652_ ( .A(_07142_ ), .B1(_07604_ ), .B2(_07605_ ), .ZN(_07614_ ) );
AOI21_X1 _15653_ ( .A(_05289_ ), .B1(_05080_ ), .B2(_04144_ ), .ZN(_07615_ ) );
OR3_X1 _15654_ ( .A1(_07613_ ), .A2(_07614_ ), .A3(_07615_ ), .ZN(_07616_ ) );
OR2_X1 _15655_ ( .A1(_07607_ ), .A2(_07616_ ), .ZN(_07617_ ) );
OAI21_X1 _15656_ ( .A(_06684_ ), .B1(_06632_ ), .B2(_07506_ ), .ZN(_07618_ ) );
AOI21_X1 _15657_ ( .A(_07618_ ), .B1(_07506_ ), .B2(_06632_ ), .ZN(_07619_ ) );
OAI21_X1 _15658_ ( .A(_06885_ ), .B1(_07617_ ), .B2(_07619_ ), .ZN(_07620_ ) );
AOI21_X1 _15659_ ( .A(_07089_ ), .B1(_07238_ ), .B2(_04176_ ), .ZN(_07621_ ) );
OAI21_X1 _15660_ ( .A(_07621_ ), .B1(_04176_ ), .B2(_07238_ ), .ZN(_07622_ ) );
AOI22_X1 _15661_ ( .A1(_05692_ ), .A2(_06599_ ), .B1(\ID_EX_imm [8] ), .B2(_06603_ ), .ZN(_07623_ ) );
AOI21_X1 _15662_ ( .A(_06584_ ), .B1(_07622_ ), .B2(_07623_ ), .ZN(_07624_ ) );
NOR2_X1 _15663_ ( .A1(_07624_ ), .A2(_03877_ ), .ZN(_07625_ ) );
AOI21_X1 _15664_ ( .A(_07594_ ), .B1(_07620_ ), .B2(_07625_ ), .ZN(_07626_ ) );
MUX2_X1 _15665_ ( .A(_05689_ ), .B(_07626_ ), .S(_06262_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
OR2_X1 _15666_ ( .A1(_05709_ ), .A2(_06284_ ), .ZN(_07627_ ) );
AND2_X1 _15667_ ( .A1(_05231_ ), .A2(_05232_ ), .ZN(_07628_ ) );
AOI21_X1 _15668_ ( .A(_05237_ ), .B1(_07628_ ), .B2(_04898_ ), .ZN(_07629_ ) );
INV_X1 _15669_ ( .A(_04921_ ), .ZN(_07630_ ) );
OR2_X1 _15670_ ( .A1(_07629_ ), .A2(_07630_ ), .ZN(_07631_ ) );
NAND2_X1 _15671_ ( .A1(_04920_ ), .A2(_02626_ ), .ZN(_07632_ ) );
AND2_X1 _15672_ ( .A1(_07631_ ), .A2(_07632_ ), .ZN(_07633_ ) );
XNOR2_X1 _15673_ ( .A(_07633_ ), .B(_04946_ ), .ZN(_07634_ ) );
NAND2_X1 _15674_ ( .A1(_07634_ ), .A2(_06891_ ), .ZN(_07635_ ) );
AOI22_X1 _15675_ ( .A1(_05698_ ), .A2(_06600_ ), .B1(\ID_EX_imm [7] ), .B2(_06603_ ), .ZN(_07636_ ) );
AOI21_X1 _15676_ ( .A(_06584_ ), .B1(_07635_ ), .B2(_07636_ ), .ZN(_07637_ ) );
OR2_X1 _15677_ ( .A1(_07637_ ), .A2(_06607_ ), .ZN(_07638_ ) );
AND4_X1 _15678_ ( .A1(_06965_ ), .A2(_06724_ ), .A3(_06733_ ), .A4(_07020_ ), .ZN(_07639_ ) );
AND3_X1 _15679_ ( .A1(_06809_ ), .A2(_06807_ ), .A3(_06790_ ), .ZN(_07640_ ) );
MUX2_X1 _15680_ ( .A(_07640_ ), .B(_07266_ ), .S(_05122_ ), .Z(_07641_ ) );
AND2_X1 _15681_ ( .A1(_07641_ ), .A2(_06843_ ), .ZN(_07642_ ) );
OR3_X1 _15682_ ( .A1(_06824_ ), .A2(_06813_ ), .A3(_06816_ ), .ZN(_07643_ ) );
OR3_X1 _15683_ ( .A1(_06812_ ), .A2(_06805_ ), .A3(_06741_ ), .ZN(_07644_ ) );
NAND3_X1 _15684_ ( .A1(_07643_ ), .A2(_07644_ ), .A3(_06857_ ), .ZN(_07645_ ) );
NAND2_X1 _15685_ ( .A1(_07496_ ), .A2(_06756_ ), .ZN(_07646_ ) );
AOI21_X1 _15686_ ( .A(_06793_ ), .B1(_07645_ ), .B2(_07646_ ), .ZN(_07647_ ) );
AOI211_X1 _15687_ ( .A(_05146_ ), .B(_07647_ ), .C1(_07137_ ), .C2(_07272_ ), .ZN(_07648_ ) );
OR2_X1 _15688_ ( .A1(_07642_ ), .A2(_07648_ ), .ZN(_07649_ ) );
OAI21_X1 _15689_ ( .A(_06995_ ), .B1(_07639_ ), .B2(_07649_ ), .ZN(_07650_ ) );
OAI21_X1 _15690_ ( .A(_06870_ ), .B1(_07642_ ), .B2(_07648_ ), .ZN(_07651_ ) );
OR3_X1 _15691_ ( .A1(_07253_ ), .A2(_06899_ ), .A3(_07329_ ), .ZN(_07652_ ) );
NAND3_X1 _15692_ ( .A1(_07650_ ), .A2(_07651_ ), .A3(_07652_ ), .ZN(_07653_ ) );
AND3_X1 _15693_ ( .A1(_06615_ ), .A2(_06616_ ), .A3(_06623_ ), .ZN(_07654_ ) );
OAI21_X1 _15694_ ( .A(_05105_ ), .B1(_07654_ ), .B2(_06630_ ), .ZN(_07655_ ) );
AND3_X1 _15695_ ( .A1(_07655_ ), .A2(_05144_ ), .A3(_06617_ ), .ZN(_07656_ ) );
AOI21_X1 _15696_ ( .A(_05144_ ), .B1(_07655_ ), .B2(_06617_ ), .ZN(_07657_ ) );
NOR3_X1 _15697_ ( .A1(_07656_ ), .A2(_07657_ ), .A3(_06998_ ), .ZN(_07658_ ) );
AOI21_X1 _15698_ ( .A(_05289_ ), .B1(_05096_ ), .B2(_04922_ ), .ZN(_07659_ ) );
AOI21_X1 _15699_ ( .A(_07659_ ), .B1(_06625_ ), .B2(_06864_ ), .ZN(_07660_ ) );
OAI21_X1 _15700_ ( .A(_07660_ ), .B1(_05144_ ), .B2(_06959_ ), .ZN(_07661_ ) );
OR3_X1 _15701_ ( .A1(_07653_ ), .A2(_07658_ ), .A3(_07661_ ), .ZN(_07662_ ) );
AOI21_X1 _15702_ ( .A(_07638_ ), .B1(_07662_ ), .B2(_07590_ ), .ZN(_07663_ ) );
NAND2_X1 _15703_ ( .A1(_05700_ ), .A2(_05891_ ), .ZN(_07664_ ) );
NAND2_X1 _15704_ ( .A1(_07664_ ), .A2(_06335_ ), .ZN(_07665_ ) );
OAI21_X1 _15705_ ( .A(_07627_ ), .B1(_07663_ ), .B2(_07665_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _15706_ ( .A1(_05727_ ), .A2(_06424_ ), .ZN(_07666_ ) );
NAND2_X1 _15707_ ( .A1(_07629_ ), .A2(_07630_ ), .ZN(_07667_ ) );
NAND3_X1 _15708_ ( .A1(_07631_ ), .A2(_06891_ ), .A3(_07667_ ), .ZN(_07668_ ) );
AOI22_X1 _15709_ ( .A1(_05730_ ), .A2(_06600_ ), .B1(\ID_EX_imm [6] ), .B2(_06603_ ), .ZN(_07669_ ) );
AOI21_X1 _15710_ ( .A(_06584_ ), .B1(_07668_ ), .B2(_07669_ ), .ZN(_07670_ ) );
OR2_X1 _15711_ ( .A1(_07670_ ), .A2(_06607_ ), .ZN(_07671_ ) );
INV_X1 _15712_ ( .A(_07020_ ), .ZN(_07672_ ) );
AND2_X1 _15713_ ( .A1(_07096_ ), .A2(_06809_ ), .ZN(_07673_ ) );
NOR4_X1 _15714_ ( .A1(_07301_ ), .A2(_06735_ ), .A3(_07672_ ), .A4(_07673_ ), .ZN(_07674_ ) );
NAND2_X1 _15715_ ( .A1(_07311_ ), .A2(_07312_ ), .ZN(_07675_ ) );
MUX2_X1 _15716_ ( .A(_07315_ ), .B(_07675_ ), .S(_05122_ ), .Z(_07676_ ) );
NAND2_X1 _15717_ ( .A1(_07676_ ), .A2(_06801_ ), .ZN(_07677_ ) );
OAI21_X1 _15718_ ( .A(_06837_ ), .B1(_06909_ ), .B2(_06913_ ), .ZN(_07678_ ) );
OAI21_X1 _15719_ ( .A(_06831_ ), .B1(_07121_ ), .B2(_06910_ ), .ZN(_07679_ ) );
AOI21_X1 _15720_ ( .A(_06739_ ), .B1(_07678_ ), .B2(_07679_ ), .ZN(_07680_ ) );
AOI21_X1 _15721_ ( .A(_06852_ ), .B1(_07538_ ), .B2(_07539_ ), .ZN(_07681_ ) );
OAI21_X1 _15722_ ( .A(_06917_ ), .B1(_07680_ ), .B2(_07681_ ), .ZN(_07682_ ) );
OAI211_X1 _15723_ ( .A(_06797_ ), .B(_07682_ ), .C1(_07309_ ), .C2(_06822_ ), .ZN(_07683_ ) );
NAND2_X1 _15724_ ( .A1(_07677_ ), .A2(_07683_ ), .ZN(_07684_ ) );
OAI21_X1 _15725_ ( .A(_06995_ ), .B1(_07674_ ), .B2(_07684_ ), .ZN(_07685_ ) );
NAND2_X1 _15726_ ( .A1(_07684_ ), .A2(_06870_ ), .ZN(_07686_ ) );
OR3_X1 _15727_ ( .A1(_07326_ ), .A2(_06899_ ), .A3(_07329_ ), .ZN(_07687_ ) );
NAND3_X1 _15728_ ( .A1(_07685_ ), .A2(_07686_ ), .A3(_07687_ ), .ZN(_07688_ ) );
OR3_X1 _15729_ ( .A1(_07654_ ), .A2(_05105_ ), .A3(_06630_ ), .ZN(_07689_ ) );
AND3_X1 _15730_ ( .A1(_07689_ ), .A2(_06684_ ), .A3(_07655_ ), .ZN(_07690_ ) );
NAND3_X1 _15731_ ( .A1(_06617_ ), .A2(_06618_ ), .A3(_06862_ ), .ZN(_07691_ ) );
OR3_X1 _15732_ ( .A1(_05104_ ), .A2(_04899_ ), .A3(_07078_ ), .ZN(_07692_ ) );
NAND2_X1 _15733_ ( .A1(_06618_ ), .A2(_05288_ ), .ZN(_07693_ ) );
NAND3_X1 _15734_ ( .A1(_07691_ ), .A2(_07692_ ), .A3(_07693_ ), .ZN(_07694_ ) );
OR3_X1 _15735_ ( .A1(_07688_ ), .A2(_07690_ ), .A3(_07694_ ), .ZN(_07695_ ) );
AOI21_X1 _15736_ ( .A(_07671_ ), .B1(_07695_ ), .B2(_07590_ ), .ZN(_07696_ ) );
OAI21_X1 _15737_ ( .A(_06888_ ), .B1(_05729_ ), .B2(_05597_ ), .ZN(_07697_ ) );
OAI21_X1 _15738_ ( .A(_07666_ ), .B1(_07696_ ), .B2(_07697_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
NAND4_X1 _15739_ ( .A1(_05564_ ), .A2(_05770_ ), .A3(\mtvec [5] ), .A4(_05771_ ), .ZN(_07698_ ) );
NAND4_X1 _15740_ ( .A1(_05568_ ), .A2(_05770_ ), .A3(\mycsreg.CSReg[0][5] ), .A4(_05771_ ), .ZN(_07699_ ) );
AND4_X1 _15741_ ( .A1(_05747_ ), .A2(_05748_ ), .A3(_07698_ ), .A4(_07699_ ), .ZN(_07700_ ) );
NAND3_X1 _15742_ ( .A1(_05365_ ), .A2(_05373_ ), .A3(_07700_ ), .ZN(_07701_ ) );
NAND3_X1 _15743_ ( .A1(_05457_ ), .A2(_05458_ ), .A3(_06147_ ), .ZN(_07702_ ) );
NAND3_X1 _15744_ ( .A1(_07701_ ), .A2(_07702_ ), .A3(_06333_ ), .ZN(_07703_ ) );
AND3_X1 _15745_ ( .A1(_05231_ ), .A2(_04874_ ), .A3(_05232_ ), .ZN(_07704_ ) );
OR3_X1 _15746_ ( .A1(_07704_ ), .A2(_04897_ ), .A3(_05235_ ), .ZN(_07705_ ) );
OAI21_X1 _15747_ ( .A(_04897_ ), .B1(_07704_ ), .B2(_05235_ ), .ZN(_07706_ ) );
NAND3_X1 _15748_ ( .A1(_07705_ ), .A2(_06891_ ), .A3(_07706_ ), .ZN(_07707_ ) );
AOI22_X1 _15749_ ( .A1(_05742_ ), .A2(_06599_ ), .B1(\ID_EX_imm [5] ), .B2(_06603_ ), .ZN(_07708_ ) );
AOI21_X1 _15750_ ( .A(_06584_ ), .B1(_07707_ ), .B2(_07708_ ), .ZN(_07709_ ) );
OR2_X1 _15751_ ( .A1(_07709_ ), .A2(_03877_ ), .ZN(_07710_ ) );
NOR4_X1 _15752_ ( .A1(_07301_ ), .A2(_07352_ ), .A3(_06735_ ), .A4(_07672_ ), .ZN(_07711_ ) );
NAND2_X1 _15753_ ( .A1(_06795_ ), .A2(_06801_ ), .ZN(_07712_ ) );
NAND3_X1 _15754_ ( .A1(_07572_ ), .A2(_07573_ ), .A3(_06929_ ), .ZN(_07713_ ) );
OAI21_X1 _15755_ ( .A(_06837_ ), .B1(_06815_ ), .B2(_06845_ ), .ZN(_07714_ ) );
OAI21_X1 _15756_ ( .A(_06825_ ), .B1(_06813_ ), .B2(_06816_ ), .ZN(_07715_ ) );
NAND2_X1 _15757_ ( .A1(_07714_ ), .A2(_07715_ ), .ZN(_07716_ ) );
OAI211_X1 _15758_ ( .A(_07713_ ), .B(_06917_ ), .C1(_07716_ ), .C2(_06929_ ), .ZN(_07717_ ) );
OAI211_X1 _15759_ ( .A(_06797_ ), .B(_07717_ ), .C1(_07360_ ), .C2(_06822_ ), .ZN(_07718_ ) );
NAND2_X1 _15760_ ( .A1(_07712_ ), .A2(_07718_ ), .ZN(_07719_ ) );
OAI21_X1 _15761_ ( .A(_06995_ ), .B1(_07711_ ), .B2(_07719_ ), .ZN(_07720_ ) );
OAI21_X1 _15762_ ( .A(_05288_ ), .B1(_05108_ ), .B2(_02579_ ), .ZN(_07721_ ) );
NAND3_X1 _15763_ ( .A1(_06615_ ), .A2(_06616_ ), .A3(_05101_ ), .ZN(_07722_ ) );
AND3_X1 _15764_ ( .A1(_07722_ ), .A2(_05110_ ), .A3(_06621_ ), .ZN(_07723_ ) );
AOI21_X1 _15765_ ( .A(_05110_ ), .B1(_07722_ ), .B2(_06621_ ), .ZN(_07724_ ) );
OAI21_X1 _15766_ ( .A(_06684_ ), .B1(_07723_ ), .B2(_07724_ ), .ZN(_07725_ ) );
NAND2_X1 _15767_ ( .A1(_07719_ ), .A2(_06870_ ), .ZN(_07726_ ) );
AND4_X1 _15768_ ( .A1(_06797_ ), .A2(_06853_ ), .A3(_06822_ ), .A4(_06858_ ), .ZN(_07727_ ) );
NAND2_X1 _15769_ ( .A1(_07727_ ), .A2(_06800_ ), .ZN(_07728_ ) );
AOI22_X1 _15770_ ( .A1(_05110_ ), .A2(_06862_ ), .B1(_06628_ ), .B2(_06864_ ), .ZN(_07729_ ) );
AND4_X1 _15771_ ( .A1(_07725_ ), .A2(_07726_ ), .A3(_07728_ ), .A4(_07729_ ), .ZN(_07730_ ) );
NAND3_X1 _15772_ ( .A1(_07720_ ), .A2(_07721_ ), .A3(_07730_ ), .ZN(_07731_ ) );
AOI21_X1 _15773_ ( .A(_07710_ ), .B1(_07731_ ), .B2(_07590_ ), .ZN(_07732_ ) );
OAI21_X1 _15774_ ( .A(_06888_ ), .B1(_05738_ ), .B2(_07492_ ), .ZN(_07733_ ) );
OAI21_X1 _15775_ ( .A(_07703_ ), .B1(_07732_ ), .B2(_07733_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
AOI21_X1 _15776_ ( .A(_04874_ ), .B1(_05231_ ), .B2(_05232_ ), .ZN(_07734_ ) );
NOR3_X1 _15777_ ( .A1(_07704_ ), .A2(_07734_ ), .A3(_07089_ ), .ZN(_07735_ ) );
OAI22_X1 _15778_ ( .A1(_05765_ ), .A2(_07149_ ), .B1(_02604_ ), .B2(_07150_ ), .ZN(_07736_ ) );
OAI21_X1 _15779_ ( .A(_06583_ ), .B1(_07735_ ), .B2(_07736_ ), .ZN(_07737_ ) );
AND2_X1 _15780_ ( .A1(_07737_ ), .A2(_03878_ ), .ZN(_07738_ ) );
NAND4_X1 _15781_ ( .A1(_06964_ ), .A2(_06965_ ), .A3(_06967_ ), .A4(_07303_ ), .ZN(_07739_ ) );
OR2_X1 _15782_ ( .A1(_06991_ ), .A2(_06796_ ), .ZN(_07740_ ) );
OAI21_X1 _15783_ ( .A(_06741_ ), .B1(_06912_ ), .B2(_06945_ ), .ZN(_07741_ ) );
OAI21_X1 _15784_ ( .A(_06758_ ), .B1(_06909_ ), .B2(_06913_ ), .ZN(_07742_ ) );
NAND2_X1 _15785_ ( .A1(_07741_ ), .A2(_07742_ ), .ZN(_07743_ ) );
MUX2_X1 _15786_ ( .A(_07743_ ), .B(_07602_ ), .S(_06738_ ), .Z(_07744_ ) );
OR2_X1 _15787_ ( .A1(_07744_ ), .A2(_06794_ ), .ZN(_07745_ ) );
OAI211_X1 _15788_ ( .A(_07745_ ), .B(_06954_ ), .C1(_06854_ ), .C2(_07389_ ), .ZN(_07746_ ) );
NAND2_X1 _15789_ ( .A1(_07740_ ), .A2(_07746_ ), .ZN(_07747_ ) );
AOI21_X1 _15790_ ( .A(_07351_ ), .B1(_07739_ ), .B2(_07747_ ), .ZN(_07748_ ) );
AND3_X1 _15791_ ( .A1(_06621_ ), .A2(_06622_ ), .A3(_06861_ ), .ZN(_07749_ ) );
NOR3_X1 _15792_ ( .A1(_06992_ ), .A2(_02656_ ), .A3(_07078_ ), .ZN(_07750_ ) );
NOR3_X1 _15793_ ( .A1(_06951_ ), .A2(_06899_ ), .A3(_07329_ ), .ZN(_07751_ ) );
NOR4_X1 _15794_ ( .A1(_07748_ ), .A2(_07749_ ), .A3(_07750_ ), .A4(_07751_ ), .ZN(_07752_ ) );
NAND3_X1 _15795_ ( .A1(_07740_ ), .A2(_06870_ ), .A3(_07746_ ), .ZN(_07753_ ) );
AOI21_X1 _15796_ ( .A(_05101_ ), .B1(_06615_ ), .B2(_06616_ ), .ZN(_07754_ ) );
NOR2_X1 _15797_ ( .A1(_07754_ ), .A2(_06997_ ), .ZN(_07755_ ) );
AOI22_X1 _15798_ ( .A1(_07755_ ), .A2(_07722_ ), .B1(_06622_ ), .B2(_05288_ ), .ZN(_07756_ ) );
AND3_X1 _15799_ ( .A1(_07752_ ), .A2(_07753_ ), .A3(_07756_ ), .ZN(_07757_ ) );
OAI21_X1 _15800_ ( .A(_07738_ ), .B1(_07757_ ), .B2(_06884_ ), .ZN(_07758_ ) );
NAND2_X1 _15801_ ( .A1(_05763_ ), .A2(_05301_ ), .ZN(_07759_ ) );
NAND3_X1 _15802_ ( .A1(_07758_ ), .A2(_06280_ ), .A3(_07759_ ), .ZN(_07760_ ) );
OR2_X1 _15803_ ( .A1(_06438_ ), .A2(_06262_ ), .ZN(_07761_ ) );
NAND2_X1 _15804_ ( .A1(_07760_ ), .A2(_07761_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
OR2_X1 _15805_ ( .A1(_05230_ ), .A2(_04421_ ), .ZN(_07762_ ) );
AND3_X1 _15806_ ( .A1(_07762_ ), .A2(_05228_ ), .A3(_04445_ ), .ZN(_07763_ ) );
AOI21_X1 _15807_ ( .A(_04445_ ), .B1(_07762_ ), .B2(_05228_ ), .ZN(_07764_ ) );
OR3_X1 _15808_ ( .A1(_07763_ ), .A2(_07764_ ), .A3(_07089_ ), .ZN(_07765_ ) );
AOI22_X1 _15809_ ( .A1(_05784_ ), .A2(_07197_ ), .B1(\ID_EX_imm [3] ), .B2(_06604_ ), .ZN(_07766_ ) );
AOI21_X1 _15810_ ( .A(_06585_ ), .B1(_07765_ ), .B2(_07766_ ), .ZN(_07767_ ) );
NOR2_X1 _15811_ ( .A1(_07767_ ), .A2(_05891_ ), .ZN(_07768_ ) );
NAND4_X1 _15812_ ( .A1(_06749_ ), .A2(_06965_ ), .A3(_07041_ ), .A4(_07303_ ), .ZN(_07769_ ) );
AOI21_X1 _15813_ ( .A(_06852_ ), .B1(_07643_ ), .B2(_07644_ ), .ZN(_07770_ ) );
NOR2_X1 _15814_ ( .A1(_06844_ ), .A2(_06848_ ), .ZN(_07771_ ) );
NOR2_X1 _15815_ ( .A1(_06815_ ), .A2(_06845_ ), .ZN(_07772_ ) );
MUX2_X1 _15816_ ( .A(_07771_ ), .B(_07772_ ), .S(_06831_ ), .Z(_07773_ ) );
AOI211_X1 _15817_ ( .A(_07137_ ), .B(_07770_ ), .C1(_06966_ ), .C2(_07773_ ), .ZN(_07774_ ) );
AOI21_X1 _15818_ ( .A(_06854_ ), .B1(_07497_ ), .B2(_07498_ ), .ZN(_07775_ ) );
OAI21_X1 _15819_ ( .A(_06992_ ), .B1(_07774_ ), .B2(_07775_ ), .ZN(_07776_ ) );
OAI211_X1 _15820_ ( .A(_06801_ ), .B(_07028_ ), .C1(_07036_ ), .C2(_06952_ ), .ZN(_07777_ ) );
NAND2_X1 _15821_ ( .A1(_07776_ ), .A2(_07777_ ), .ZN(_07778_ ) );
AOI21_X1 _15822_ ( .A(_07351_ ), .B1(_07769_ ), .B2(_07778_ ), .ZN(_07779_ ) );
NOR2_X1 _15823_ ( .A1(_05125_ ), .A2(_06614_ ), .ZN(_07780_ ) );
OAI22_X1 _15824_ ( .A1(_07780_ ), .A2(_06609_ ), .B1(_05139_ ), .B2(_05140_ ), .ZN(_07781_ ) );
OAI211_X1 _15825_ ( .A(_05115_ ), .B(_06610_ ), .C1(_05125_ ), .C2(_06614_ ), .ZN(_07782_ ) );
AOI21_X1 _15826_ ( .A(_06998_ ), .B1(_07781_ ), .B2(_07782_ ), .ZN(_07783_ ) );
NOR2_X1 _15827_ ( .A1(_07057_ ), .A2(_07329_ ), .ZN(_07784_ ) );
AOI221_X4 _15828_ ( .A(_07784_ ), .B1(_05139_ ), .B2(_04952_ ), .C1(_05115_ ), .C2(_06861_ ), .ZN(_07785_ ) );
OAI221_X1 _15829_ ( .A(_07785_ ), .B1(_05140_ ), .B2(_06872_ ), .C1(_07778_ ), .C2(_07142_ ), .ZN(_07786_ ) );
NOR3_X1 _15830_ ( .A1(_07779_ ), .A2(_07783_ ), .A3(_07786_ ), .ZN(_07787_ ) );
OAI21_X1 _15831_ ( .A(_07768_ ), .B1(_07787_ ), .B2(_06884_ ), .ZN(_07788_ ) );
NAND2_X1 _15832_ ( .A1(_05301_ ), .A2(_05786_ ), .ZN(_07789_ ) );
NAND3_X1 _15833_ ( .A1(_07788_ ), .A2(_06280_ ), .A3(_07789_ ), .ZN(_07790_ ) );
NAND2_X1 _15834_ ( .A1(_05795_ ), .A2(_06266_ ), .ZN(_07791_ ) );
NAND2_X1 _15835_ ( .A1(_07790_ ), .A2(_07791_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
AOI22_X1 _15836_ ( .A1(_05806_ ), .A2(_05808_ ), .B1(_05458_ ), .B2(_05457_ ), .ZN(_07792_ ) );
OAI21_X1 _15837_ ( .A(_06414_ ), .B1(_07792_ ), .B2(_05801_ ), .ZN(_07793_ ) );
NAND3_X1 _15838_ ( .A1(_04389_ ), .A2(_04421_ ), .A3(_05229_ ), .ZN(_07794_ ) );
NAND3_X1 _15839_ ( .A1(_07762_ ), .A2(_06891_ ), .A3(_07794_ ), .ZN(_07795_ ) );
AOI22_X1 _15840_ ( .A1(_05812_ ), .A2(_06599_ ), .B1(\ID_EX_imm [2] ), .B2(_06603_ ), .ZN(_07796_ ) );
AOI21_X1 _15841_ ( .A(_06584_ ), .B1(_07795_ ), .B2(_07796_ ), .ZN(_07797_ ) );
OR2_X1 _15842_ ( .A1(_07797_ ), .A2(_03877_ ), .ZN(_07798_ ) );
NAND3_X1 _15843_ ( .A1(_06749_ ), .A2(_06965_ ), .A3(_07041_ ), .ZN(_07799_ ) );
NOR3_X1 _15844_ ( .A1(_07799_ ), .A2(_07096_ ), .A3(_07672_ ), .ZN(_07800_ ) );
OR2_X1 _15845_ ( .A1(_07113_ ), .A2(_06955_ ), .ZN(_07801_ ) );
AND3_X1 _15846_ ( .A1(_07678_ ), .A2(_07679_ ), .A3(_06739_ ), .ZN(_07802_ ) );
NOR2_X1 _15847_ ( .A1(_06944_ ), .A2(_06948_ ), .ZN(_07803_ ) );
NOR2_X1 _15848_ ( .A1(_06912_ ), .A2(_06945_ ), .ZN(_07804_ ) );
MUX2_X1 _15849_ ( .A(_07803_ ), .B(_07804_ ), .S(_06831_ ), .Z(_07805_ ) );
AOI211_X1 _15850_ ( .A(_07137_ ), .B(_07802_ ), .C1(_06966_ ), .C2(_07805_ ), .ZN(_07806_ ) );
AND3_X1 _15851_ ( .A1(_07537_ ), .A2(_07540_ ), .A3(_07137_ ), .ZN(_07807_ ) );
OR3_X1 _15852_ ( .A1(_07806_ ), .A2(_06897_ ), .A3(_07807_ ), .ZN(_07808_ ) );
NAND2_X1 _15853_ ( .A1(_07801_ ), .A2(_07808_ ), .ZN(_07809_ ) );
OAI21_X1 _15854_ ( .A(_06995_ ), .B1(_07800_ ), .B2(_07809_ ), .ZN(_07810_ ) );
NAND2_X1 _15855_ ( .A1(_07809_ ), .A2(_06870_ ), .ZN(_07811_ ) );
OAI21_X1 _15856_ ( .A(_06684_ ), .B1(_05125_ ), .B2(_06614_ ), .ZN(_07812_ ) );
AOI21_X1 _15857_ ( .A(_07812_ ), .B1(_05125_ ), .B2(_06614_ ), .ZN(_07813_ ) );
NOR4_X1 _15858_ ( .A1(_07136_ ), .A2(_06801_ ), .A3(_06952_ ), .A4(_06740_ ), .ZN(_07814_ ) );
AND2_X1 _15859_ ( .A1(_07814_ ), .A2(_06800_ ), .ZN(_07815_ ) );
AOI21_X1 _15860_ ( .A(_06872_ ), .B1(_06966_ ), .B2(_04390_ ), .ZN(_07816_ ) );
OAI22_X1 _15861_ ( .A1(_05125_ ), .A2(_06959_ ), .B1(_06610_ ), .B2(_07187_ ), .ZN(_07817_ ) );
NOR4_X1 _15862_ ( .A1(_07813_ ), .A2(_07815_ ), .A3(_07816_ ), .A4(_07817_ ), .ZN(_07818_ ) );
NAND3_X1 _15863_ ( .A1(_07810_ ), .A2(_07811_ ), .A3(_07818_ ), .ZN(_07819_ ) );
AOI21_X1 _15864_ ( .A(_07798_ ), .B1(_07819_ ), .B2(_07590_ ), .ZN(_07820_ ) );
OAI21_X1 _15865_ ( .A(_06888_ ), .B1(_05325_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07821_ ) );
OAI21_X1 _15866_ ( .A(_07793_ ), .B1(_07820_ ), .B2(_07821_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
NAND2_X1 _15867_ ( .A1(_05357_ ), .A2(_06424_ ), .ZN(_07822_ ) );
NAND3_X1 _15868_ ( .A1(_07472_ ), .A2(_04599_ ), .A3(_04649_ ), .ZN(_07823_ ) );
AND2_X1 _15869_ ( .A1(_07823_ ), .A2(_05276_ ), .ZN(_07824_ ) );
INV_X1 _15870_ ( .A(_04522_ ), .ZN(_07825_ ) );
NOR2_X1 _15871_ ( .A1(_07824_ ), .A2(_07825_ ), .ZN(_07826_ ) );
OR3_X1 _15872_ ( .A1(_07826_ ), .A2(_04545_ ), .A3(_05267_ ), .ZN(_07827_ ) );
OAI21_X1 _15873_ ( .A(_04545_ ), .B1(_07826_ ), .B2(_05267_ ), .ZN(_07828_ ) );
AND3_X1 _15874_ ( .A1(_07827_ ), .A2(_06891_ ), .A3(_07828_ ), .ZN(_07829_ ) );
OAI22_X1 _15875_ ( .A1(_05323_ ), .A2(_07149_ ), .B1(_02974_ ), .B2(_07150_ ), .ZN(_07830_ ) );
OAI21_X1 _15876_ ( .A(_06583_ ), .B1(_07829_ ), .B2(_07830_ ), .ZN(_07831_ ) );
NAND2_X1 _15877_ ( .A1(_07831_ ), .A2(_05360_ ), .ZN(_07832_ ) );
INV_X1 _15878_ ( .A(_07433_ ), .ZN(_07833_ ) );
AOI21_X1 _15879_ ( .A(_04983_ ), .B1(_07833_ ), .B2(_07434_ ), .ZN(_07834_ ) );
OR3_X1 _15880_ ( .A1(_07834_ ), .A2(_04976_ ), .A3(_07437_ ), .ZN(_07835_ ) );
OAI21_X1 _15881_ ( .A(_04976_ ), .B1(_07834_ ), .B2(_07437_ ), .ZN(_07836_ ) );
NAND3_X1 _15882_ ( .A1(_07835_ ), .A2(_06685_ ), .A3(_07836_ ), .ZN(_07837_ ) );
NAND2_X1 _15883_ ( .A1(_04976_ ), .A2(_06862_ ), .ZN(_07838_ ) );
NAND3_X1 _15884_ ( .A1(_04974_ ), .A2(_02973_ ), .A3(_06864_ ), .ZN(_07839_ ) );
OAI21_X1 _15885_ ( .A(_05288_ ), .B1(_04974_ ), .B2(_02973_ ), .ZN(_07840_ ) );
AND3_X1 _15886_ ( .A1(_07838_ ), .A2(_07839_ ), .A3(_07840_ ), .ZN(_07841_ ) );
OAI211_X1 _15887_ ( .A(_06749_ ), .B(_06750_ ), .C1(_06747_ ), .C2(_07354_ ), .ZN(_07842_ ) );
NOR3_X1 _15888_ ( .A1(_06791_ ), .A2(_06952_ ), .A3(_06740_ ), .ZN(_07843_ ) );
NAND2_X1 _15889_ ( .A1(_07843_ ), .A2(_06867_ ), .ZN(_07844_ ) );
AOI21_X1 _15890_ ( .A(_07351_ ), .B1(_07842_ ), .B2(_07844_ ), .ZN(_07845_ ) );
OR3_X1 _15891_ ( .A1(_06833_ ), .A2(_06840_ ), .A3(_06917_ ), .ZN(_07846_ ) );
OR3_X1 _15892_ ( .A1(_06772_ ), .A2(_06778_ ), .A3(_06837_ ), .ZN(_07847_ ) );
NOR2_X1 _15893_ ( .A1(_06777_ ), .A2(_06765_ ), .ZN(_07848_ ) );
NAND2_X1 _15894_ ( .A1(_07848_ ), .A2(_06931_ ), .ZN(_07849_ ) );
NAND2_X1 _15895_ ( .A1(_07847_ ), .A2(_07849_ ), .ZN(_07850_ ) );
NOR2_X1 _15896_ ( .A1(_06760_ ), .A2(_06768_ ), .ZN(_07851_ ) );
AND2_X1 _15897_ ( .A1(_07022_ ), .A2(_06786_ ), .ZN(_07852_ ) );
MUX2_X1 _15898_ ( .A(_07851_ ), .B(_07852_ ), .S(_06931_ ), .Z(_07853_ ) );
MUX2_X1 _15899_ ( .A(_07850_ ), .B(_07853_ ), .S(_06966_ ), .Z(_07854_ ) );
OAI211_X1 _15900_ ( .A(_06955_ ), .B(_07846_ ), .C1(_07854_ ), .C2(_06899_ ), .ZN(_07855_ ) );
OAI21_X1 _15901_ ( .A(_06897_ ), .B1(_07367_ ), .B2(_07368_ ), .ZN(_07856_ ) );
AOI21_X1 _15902_ ( .A(_07053_ ), .B1(_07855_ ), .B2(_07856_ ), .ZN(_07857_ ) );
AND3_X1 _15903_ ( .A1(_07843_ ), .A2(_06955_ ), .A3(_06869_ ), .ZN(_07858_ ) );
NOR3_X1 _15904_ ( .A1(_07845_ ), .A2(_07857_ ), .A3(_07858_ ), .ZN(_07859_ ) );
NAND3_X1 _15905_ ( .A1(_07837_ ), .A2(_07841_ ), .A3(_07859_ ), .ZN(_07860_ ) );
AOI21_X1 _15906_ ( .A(_07832_ ), .B1(_07860_ ), .B2(_07590_ ), .ZN(_07861_ ) );
OAI21_X1 _15907_ ( .A(_06888_ ), .B1(_05318_ ), .B2(_07492_ ), .ZN(_07862_ ) );
OAI21_X1 _15908_ ( .A(_07822_ ), .B1(_07861_ ), .B2(_07862_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
NAND2_X1 _15909_ ( .A1(_05825_ ), .A2(_06424_ ), .ZN(_07863_ ) );
OR2_X1 _15910_ ( .A1(_04364_ ), .A2(_04388_ ), .ZN(_07864_ ) );
AND3_X1 _15911_ ( .A1(_07864_ ), .A2(_04389_ ), .A3(_06891_ ), .ZN(_07865_ ) );
OAI22_X1 _15912_ ( .A1(_05827_ ), .A2(_07149_ ), .B1(_05127_ ), .B2(_07150_ ), .ZN(_07866_ ) );
OAI21_X1 _15913_ ( .A(_06583_ ), .B1(_07865_ ), .B2(_07866_ ), .ZN(_07867_ ) );
NAND2_X1 _15914_ ( .A1(_07867_ ), .A2(_05360_ ), .ZN(_07868_ ) );
OR3_X1 _15915_ ( .A1(_07160_ ), .A2(_06796_ ), .A3(_07167_ ), .ZN(_07869_ ) );
OAI21_X1 _15916_ ( .A(_06837_ ), .B1(_06847_ ), .B2(_06855_ ), .ZN(_07870_ ) );
OAI211_X1 _15917_ ( .A(_07870_ ), .B(_06857_ ), .C1(_07771_ ), .C2(_06837_ ), .ZN(_07871_ ) );
OAI211_X1 _15918_ ( .A(_07871_ ), .B(_06820_ ), .C1(_06823_ ), .C2(_07716_ ), .ZN(_07872_ ) );
OAI211_X1 _15919_ ( .A(_06954_ ), .B(_07872_ ), .C1(_07575_ ), .C2(_06917_ ), .ZN(_07873_ ) );
AOI21_X1 _15920_ ( .A(_07142_ ), .B1(_07869_ ), .B2(_07873_ ), .ZN(_07874_ ) );
AND2_X1 _15921_ ( .A1(_06749_ ), .A2(_07041_ ), .ZN(_07875_ ) );
NAND4_X1 _15922_ ( .A1(_07875_ ), .A2(_06745_ ), .A3(_06736_ ), .A4(_07020_ ), .ZN(_07876_ ) );
NAND3_X1 _15923_ ( .A1(_07876_ ), .A2(_07873_ ), .A3(_07869_ ), .ZN(_07877_ ) );
AOI221_X4 _15924_ ( .A(_07874_ ), .B1(_07177_ ), .B2(_07260_ ), .C1(_07877_ ), .C2(_06688_ ), .ZN(_07878_ ) );
OAI21_X1 _15925_ ( .A(_06685_ ), .B1(_05133_ ), .B2(_06611_ ), .ZN(_07879_ ) );
OR2_X1 _15926_ ( .A1(_07879_ ), .A2(_06613_ ), .ZN(_07880_ ) );
NOR3_X1 _15927_ ( .A1(_05131_ ), .A2(_05132_ ), .A3(_06959_ ), .ZN(_07881_ ) );
NOR3_X1 _15928_ ( .A1(_06931_ ), .A2(_04339_ ), .A3(_07187_ ), .ZN(_07882_ ) );
AOI21_X1 _15929_ ( .A(_06873_ ), .B1(_06931_ ), .B2(_04339_ ), .ZN(_07883_ ) );
NOR3_X1 _15930_ ( .A1(_07881_ ), .A2(_07882_ ), .A3(_07883_ ), .ZN(_07884_ ) );
NAND3_X1 _15931_ ( .A1(_07878_ ), .A2(_07880_ ), .A3(_07884_ ), .ZN(_07885_ ) );
AOI21_X1 _15932_ ( .A(_07868_ ), .B1(_07885_ ), .B2(_07590_ ), .ZN(_07886_ ) );
OAI21_X1 _15933_ ( .A(_06272_ ), .B1(_05325_ ), .B2(\ID_EX_pc [1] ), .ZN(_07887_ ) );
OAI21_X1 _15934_ ( .A(_07863_ ), .B1(_07886_ ), .B2(_07887_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
OR2_X1 _15935_ ( .A1(_06480_ ), .A2(_06284_ ), .ZN(_07888_ ) );
AND3_X1 _15936_ ( .A1(_05197_ ), .A2(_05202_ ), .A3(_06882_ ), .ZN(_07889_ ) );
NAND3_X1 _15937_ ( .A1(_05858_ ), .A2(_06598_ ), .A3(_06597_ ), .ZN(_07890_ ) );
OAI21_X1 _15938_ ( .A(_07890_ ), .B1(_07150_ ), .B2(_02480_ ), .ZN(_07891_ ) );
AOI21_X1 _15939_ ( .A(_07089_ ), .B1(_04388_ ), .B2(_04853_ ), .ZN(_07892_ ) );
NOR3_X1 _15940_ ( .A1(_07889_ ), .A2(_07891_ ), .A3(_07892_ ), .ZN(_07893_ ) );
INV_X1 _15941_ ( .A(_05199_ ), .ZN(_07894_ ) );
NAND3_X1 _15942_ ( .A1(_05284_ ), .A2(_04950_ ), .A3(\ID_EX_typ [2] ), .ZN(_07895_ ) );
AOI211_X1 _15943_ ( .A(_04964_ ), .B(_07895_ ), .C1(_05201_ ), .C2(_04971_ ), .ZN(_07896_ ) );
NAND3_X1 _15944_ ( .A1(_05197_ ), .A2(_07894_ ), .A3(_07896_ ), .ZN(_07897_ ) );
AND4_X1 _15945_ ( .A1(_05108_ ), .A2(_06724_ ), .A3(_06699_ ), .A4(_06733_ ), .ZN(_07898_ ) );
NAND2_X1 _15946_ ( .A1(_07213_ ), .A2(_06801_ ), .ZN(_07899_ ) );
AOI21_X1 _15947_ ( .A(_02502_ ), .B1(_06773_ ), .B2(_06774_ ), .ZN(_07900_ ) );
OAI21_X1 _15948_ ( .A(_06837_ ), .B1(_06947_ ), .B2(_07900_ ), .ZN(_07901_ ) );
OAI211_X1 _15949_ ( .A(_07901_ ), .B(_06810_ ), .C1(_07803_ ), .C2(_06931_ ), .ZN(_07902_ ) );
OAI211_X1 _15950_ ( .A(_07902_ ), .B(_06820_ ), .C1(_06823_ ), .C2(_07743_ ), .ZN(_07903_ ) );
OAI211_X1 _15951_ ( .A(_06954_ ), .B(_07903_ ), .C1(_07603_ ), .C2(_06854_ ), .ZN(_07904_ ) );
NAND2_X1 _15952_ ( .A1(_07899_ ), .A2(_07904_ ), .ZN(_07905_ ) );
OAI21_X1 _15953_ ( .A(_06688_ ), .B1(_07898_ ), .B2(_07905_ ), .ZN(_07906_ ) );
NAND2_X1 _15954_ ( .A1(_07905_ ), .A2(_06869_ ), .ZN(_07907_ ) );
NAND4_X1 _15955_ ( .A1(_06698_ ), .A2(_02502_ ), .A3(_06955_ ), .A4(_06800_ ), .ZN(_07908_ ) );
NAND4_X1 _15956_ ( .A1(_07897_ ), .A2(_07906_ ), .A3(_07907_ ), .A4(_07908_ ), .ZN(_07909_ ) );
NOR3_X1 _15957_ ( .A1(_06611_ ), .A2(_07900_ ), .A3(_06997_ ), .ZN(_07910_ ) );
OAI21_X1 _15958_ ( .A(_06861_ ), .B1(_06941_ ), .B2(_05137_ ), .ZN(_07911_ ) );
OAI221_X1 _15959_ ( .A(_07911_ ), .B1(_06872_ ), .B2(_07900_ ), .C1(_07187_ ), .C2(_06612_ ), .ZN(_07912_ ) );
NOR3_X1 _15960_ ( .A1(_07909_ ), .A2(_07910_ ), .A3(_07912_ ), .ZN(_07913_ ) );
OAI221_X1 _15961_ ( .A(_03879_ ), .B1(_06585_ ), .B2(_07893_ ), .C1(_07913_ ), .C2(_06884_ ), .ZN(_07914_ ) );
OAI21_X1 _15962_ ( .A(_07914_ ), .B1(\ID_EX_pc [0] ), .B2(_05299_ ), .ZN(_07915_ ) );
OAI21_X1 _15963_ ( .A(_07888_ ), .B1(_07915_ ), .B2(_06388_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
NAND2_X1 _15964_ ( .A1(_05630_ ), .A2(_06424_ ), .ZN(_07916_ ) );
OAI21_X1 _15965_ ( .A(_06891_ ), .B1(_07824_ ), .B2(_07825_ ), .ZN(_07917_ ) );
AOI21_X1 _15966_ ( .A(_07917_ ), .B1(_07825_ ), .B2(_07824_ ), .ZN(_07918_ ) );
AND2_X1 _15967_ ( .A1(_05633_ ), .A2(_07197_ ), .ZN(_07919_ ) );
AND3_X1 _15968_ ( .A1(_06601_ ), .A2(\ID_EX_imm [28] ), .A3(_06598_ ), .ZN(_07920_ ) );
NOR3_X1 _15969_ ( .A1(_07918_ ), .A2(_07919_ ), .A3(_07920_ ), .ZN(_07921_ ) );
OAI21_X1 _15970_ ( .A(_05360_ ), .B1(_07921_ ), .B2(_07154_ ), .ZN(_07922_ ) );
NOR3_X1 _15971_ ( .A1(_07433_ ), .A2(_04982_ ), .A3(_07435_ ), .ZN(_07923_ ) );
OR3_X1 _15972_ ( .A1(_07834_ ), .A2(_06998_ ), .A3(_07923_ ), .ZN(_07924_ ) );
NAND2_X1 _15973_ ( .A1(_04982_ ), .A2(_06862_ ), .ZN(_07925_ ) );
OAI21_X1 _15974_ ( .A(_05288_ ), .B1(_04980_ ), .B2(_02209_ ), .ZN(_07926_ ) );
NAND3_X1 _15975_ ( .A1(_04980_ ), .A2(_02209_ ), .A3(_06864_ ), .ZN(_07927_ ) );
AND3_X1 _15976_ ( .A1(_07925_ ), .A2(_07926_ ), .A3(_07927_ ), .ZN(_07928_ ) );
OAI211_X1 _15977_ ( .A(_06749_ ), .B(_06735_ ), .C1(_06696_ ), .C2(_07041_ ), .ZN(_07929_ ) );
INV_X1 _15978_ ( .A(_07929_ ), .ZN(_07930_ ) );
OAI21_X1 _15979_ ( .A(_06752_ ), .B1(_07930_ ), .B2(_06737_ ), .ZN(_07931_ ) );
NOR3_X1 _15980_ ( .A1(_06989_ ), .A2(_06952_ ), .A3(_06740_ ), .ZN(_07932_ ) );
AOI22_X1 _15981_ ( .A1(_06749_ ), .A2(_07303_ ), .B1(_06955_ ), .B2(_07932_ ), .ZN(_07933_ ) );
AOI21_X1 _15982_ ( .A(_07351_ ), .B1(_07931_ ), .B2(_07933_ ), .ZN(_07934_ ) );
OAI21_X1 _15983_ ( .A(_06897_ ), .B1(_07396_ ), .B2(_07397_ ), .ZN(_07935_ ) );
OAI21_X1 _15984_ ( .A(_06952_ ), .B1(_06930_ ), .B2(_06938_ ), .ZN(_07936_ ) );
OAI21_X1 _15985_ ( .A(_06931_ ), .B1(_06972_ ), .B2(_06977_ ), .ZN(_07937_ ) );
OAI21_X1 _15986_ ( .A(_06831_ ), .B1(_06970_ ), .B2(_06973_ ), .ZN(_07938_ ) );
AND2_X1 _15987_ ( .A1(_07937_ ), .A2(_07938_ ), .ZN(_07939_ ) );
NOR2_X1 _15988_ ( .A1(_06976_ ), .A2(_06980_ ), .ZN(_07940_ ) );
MUX2_X1 _15989_ ( .A(_07940_ ), .B(_07456_ ), .S(_06931_ ), .Z(_07941_ ) );
MUX2_X1 _15990_ ( .A(_07939_ ), .B(_07941_ ), .S(_06823_ ), .Z(_07942_ ) );
OAI211_X1 _15991_ ( .A(_06955_ ), .B(_07936_ ), .C1(_07942_ ), .C2(_06899_ ), .ZN(_07943_ ) );
AOI21_X1 _15992_ ( .A(_07053_ ), .B1(_07935_ ), .B2(_07943_ ), .ZN(_07944_ ) );
AND3_X1 _15993_ ( .A1(_07932_ ), .A2(_06955_ ), .A3(_06869_ ), .ZN(_07945_ ) );
NOR3_X1 _15994_ ( .A1(_07934_ ), .A2(_07944_ ), .A3(_07945_ ), .ZN(_07946_ ) );
NAND3_X1 _15995_ ( .A1(_07924_ ), .A2(_07928_ ), .A3(_07946_ ), .ZN(_07947_ ) );
AOI21_X1 _15996_ ( .A(_07922_ ), .B1(_07947_ ), .B2(_07590_ ), .ZN(_07948_ ) );
OAI21_X1 _15997_ ( .A(_06272_ ), .B1(_05632_ ), .B2(_07492_ ), .ZN(_07949_ ) );
OAI21_X1 _15998_ ( .A(_07916_ ), .B1(_07948_ ), .B2(_07949_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND3_X1 _15999_ ( .A1(_05851_ ), .A2(_05853_ ), .A3(_06333_ ), .ZN(_07950_ ) );
OAI22_X1 _16000_ ( .A1(_05843_ ), .A2(_07149_ ), .B1(_02212_ ), .B2(_07150_ ), .ZN(_07951_ ) );
NOR2_X1 _16001_ ( .A1(_07473_ ), .A2(_04573_ ), .ZN(_07952_ ) );
NOR2_X1 _16002_ ( .A1(_04571_ ), .A2(_05164_ ), .ZN(_07953_ ) );
NOR2_X1 _16003_ ( .A1(_07952_ ), .A2(_07953_ ), .ZN(_07954_ ) );
OR2_X1 _16004_ ( .A1(_07954_ ), .A2(_04598_ ), .ZN(_07955_ ) );
AOI21_X1 _16005_ ( .A(_07089_ ), .B1(_07954_ ), .B2(_04598_ ), .ZN(_07956_ ) );
AOI21_X1 _16006_ ( .A(_07951_ ), .B1(_07955_ ), .B2(_07956_ ), .ZN(_07957_ ) );
OAI21_X1 _16007_ ( .A(_05360_ ), .B1(_07957_ ), .B2(_07154_ ), .ZN(_07958_ ) );
AOI21_X1 _16008_ ( .A(_07421_ ), .B1(_07431_ ), .B2(_07432_ ), .ZN(_07959_ ) );
OR3_X1 _16009_ ( .A1(_07959_ ), .A2(_07419_ ), .A3(_05165_ ), .ZN(_07960_ ) );
OAI21_X1 _16010_ ( .A(_07419_ ), .B1(_07959_ ), .B2(_05165_ ), .ZN(_07961_ ) );
AND3_X1 _16011_ ( .A1(_07960_ ), .A2(_06685_ ), .A3(_07961_ ), .ZN(_07962_ ) );
AOI22_X1 _16012_ ( .A1(_05171_ ), .A2(_06864_ ), .B1(_05174_ ), .B2(_05288_ ), .ZN(_07963_ ) );
OAI21_X1 _16013_ ( .A(_07963_ ), .B1(_07420_ ), .B2(_06959_ ), .ZN(_07964_ ) );
OAI211_X1 _16014_ ( .A(_06734_ ), .B(_06752_ ), .C1(_06736_ ), .C2(_07040_ ), .ZN(_07965_ ) );
OAI211_X1 _16015_ ( .A(_07965_ ), .B(_07263_ ), .C1(_05146_ ), .C2(_07501_ ), .ZN(_07966_ ) );
AND2_X1 _16016_ ( .A1(_07966_ ), .A2(_06688_ ), .ZN(_07967_ ) );
NOR2_X1 _16017_ ( .A1(_06796_ ), .A2(_07053_ ), .ZN(_07968_ ) );
INV_X1 _16018_ ( .A(_07968_ ), .ZN(_07969_ ) );
AOI21_X1 _16019_ ( .A(_07969_ ), .B1(_07518_ ), .B2(_07519_ ), .ZN(_07970_ ) );
OAI21_X1 _16020_ ( .A(_06742_ ), .B1(_06772_ ), .B2(_06778_ ), .ZN(_07971_ ) );
OAI21_X1 _16021_ ( .A(_06825_ ), .B1(_06838_ ), .B2(_06775_ ), .ZN(_07972_ ) );
NAND2_X1 _16022_ ( .A1(_07971_ ), .A2(_07972_ ), .ZN(_07973_ ) );
OAI21_X1 _16023_ ( .A(_06819_ ), .B1(_07973_ ), .B2(_06810_ ), .ZN(_07974_ ) );
NAND2_X1 _16024_ ( .A1(_07848_ ), .A2(_06825_ ), .ZN(_07975_ ) );
OAI211_X1 _16025_ ( .A(_07023_ ), .B(_06837_ ), .C1(_02256_ ), .C2(_06744_ ), .ZN(_07976_ ) );
AOI21_X1 _16026_ ( .A(_06756_ ), .B1(_07975_ ), .B2(_07976_ ), .ZN(_07977_ ) );
OAI21_X1 _16027_ ( .A(_07260_ ), .B1(_07974_ ), .B2(_07977_ ), .ZN(_07978_ ) );
AOI21_X1 _16028_ ( .A(_07978_ ), .B1(_07137_ ), .B2(_07066_ ), .ZN(_07979_ ) );
NOR3_X1 _16029_ ( .A1(_07501_ ), .A2(_06843_ ), .A3(_07142_ ), .ZN(_07980_ ) );
OR4_X1 _16030_ ( .A1(_07967_ ), .A2(_07970_ ), .A3(_07979_ ), .A4(_07980_ ), .ZN(_07981_ ) );
OR3_X1 _16031_ ( .A1(_07962_ ), .A2(_07964_ ), .A3(_07981_ ), .ZN(_07982_ ) );
AOI21_X1 _16032_ ( .A(_07958_ ), .B1(_07982_ ), .B2(_07590_ ), .ZN(_07983_ ) );
OAI21_X1 _16033_ ( .A(_06272_ ), .B1(_05836_ ), .B2(_07492_ ), .ZN(_00303_ ) );
OAI21_X1 _16034_ ( .A(_07950_ ), .B1(_07983_ ), .B2(_00303_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
OAI21_X1 _16035_ ( .A(_06414_ ), .B1(_06509_ ), .B2(_06510_ ), .ZN(_00304_ ) );
OAI21_X1 _16036_ ( .A(_06891_ ), .B1(_07473_ ), .B2(_04573_ ), .ZN(_00305_ ) );
AOI21_X1 _16037_ ( .A(_00305_ ), .B1(_04573_ ), .B2(_07473_ ), .ZN(_00306_ ) );
AND3_X1 _16038_ ( .A1(_05885_ ), .A2(_05840_ ), .A3(_06599_ ), .ZN(_00307_ ) );
AND3_X1 _16039_ ( .A1(_06601_ ), .A2(\ID_EX_imm [26] ), .A3(_06598_ ), .ZN(_00308_ ) );
NOR3_X1 _16040_ ( .A1(_00306_ ), .A2(_00307_ ), .A3(_00308_ ), .ZN(_00309_ ) );
OAI21_X1 _16041_ ( .A(_03879_ ), .B1(_00309_ ), .B2(_07154_ ), .ZN(_00310_ ) );
AND3_X1 _16042_ ( .A1(_07431_ ), .A2(_07421_ ), .A3(_07432_ ), .ZN(_00311_ ) );
OR3_X1 _16043_ ( .A1(_00311_ ), .A2(_07959_ ), .A3(_06998_ ), .ZN(_00312_ ) );
NOR3_X1 _16044_ ( .A1(_05165_ ), .A2(_05166_ ), .A3(_06959_ ), .ZN(_00313_ ) );
NOR3_X1 _16045_ ( .A1(_05163_ ), .A2(_05164_ ), .A3(_07187_ ), .ZN(_00314_ ) );
AOI21_X1 _16046_ ( .A(_06873_ ), .B1(_05163_ ), .B2(_05164_ ), .ZN(_00315_ ) );
NOR3_X1 _16047_ ( .A1(_00313_ ), .A2(_00314_ ), .A3(_00315_ ), .ZN(_00316_ ) );
AOI21_X1 _16048_ ( .A(_07534_ ), .B1(_06965_ ), .B2(_06749_ ), .ZN(_00317_ ) );
NOR2_X1 _16049_ ( .A1(_00317_ ), .A2(_06753_ ), .ZN(_00318_ ) );
NAND2_X1 _16050_ ( .A1(_07543_ ), .A2(_06797_ ), .ZN(_00319_ ) );
NAND2_X1 _16051_ ( .A1(_07263_ ), .A2(_00319_ ), .ZN(_00320_ ) );
OAI21_X1 _16052_ ( .A(_06688_ ), .B1(_00318_ ), .B2(_00320_ ), .ZN(_00321_ ) );
OAI21_X1 _16053_ ( .A(_00321_ ), .B1(_07142_ ), .B2(_00319_ ), .ZN(_00322_ ) );
AOI21_X1 _16054_ ( .A(_06918_ ), .B1(_07129_ ), .B2(_07132_ ), .ZN(_00323_ ) );
NAND3_X1 _16055_ ( .A1(_07452_ ), .A2(_07453_ ), .A3(_06966_ ), .ZN(_00324_ ) );
NAND3_X1 _16056_ ( .A1(_07448_ ), .A2(_07449_ ), .A3(_06740_ ), .ZN(_00325_ ) );
AND3_X1 _16057_ ( .A1(_00324_ ), .A2(_00325_ ), .A3(_06918_ ), .ZN(_00326_ ) );
NOR3_X1 _16058_ ( .A1(_00323_ ), .A2(_00326_ ), .A3(_07329_ ), .ZN(_00327_ ) );
AOI21_X1 _16059_ ( .A(_07969_ ), .B1(_07548_ ), .B2(_07549_ ), .ZN(_00328_ ) );
NOR3_X1 _16060_ ( .A1(_00322_ ), .A2(_00327_ ), .A3(_00328_ ), .ZN(_00329_ ) );
NAND3_X1 _16061_ ( .A1(_00312_ ), .A2(_00316_ ), .A3(_00329_ ), .ZN(_00330_ ) );
AOI21_X1 _16062_ ( .A(_00310_ ), .B1(_00330_ ), .B2(_07590_ ), .ZN(_00331_ ) );
OAI21_X1 _16063_ ( .A(_06272_ ), .B1(_05884_ ), .B2(_07492_ ), .ZN(_00332_ ) );
OAI21_X1 _16064_ ( .A(_00304_ ), .B1(_00331_ ), .B2(_00332_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
AND2_X1 _16065_ ( .A1(_05896_ ), .A2(_05898_ ), .ZN(_00333_ ) );
AND2_X1 _16066_ ( .A1(_05897_ ), .A2(_05899_ ), .ZN(_00334_ ) );
AOI22_X1 _16067_ ( .A1(_00333_ ), .A2(_00334_ ), .B1(_05458_ ), .B2(_05457_ ), .ZN(_00335_ ) );
OAI21_X1 _16068_ ( .A(_06414_ ), .B1(_00335_ ), .B2(_05894_ ), .ZN(_00336_ ) );
NAND2_X1 _16069_ ( .A1(_04621_ ), .A2(_02915_ ), .ZN(_00337_ ) );
INV_X1 _16070_ ( .A(_04623_ ), .ZN(_00338_ ) );
OAI21_X1 _16071_ ( .A(_00337_ ), .B1(_07471_ ), .B2(_00338_ ), .ZN(_00339_ ) );
OAI21_X1 _16072_ ( .A(_06594_ ), .B1(_00339_ ), .B2(_04648_ ), .ZN(_00340_ ) );
AOI21_X1 _16073_ ( .A(_00340_ ), .B1(_04648_ ), .B2(_00339_ ), .ZN(_00341_ ) );
AND2_X1 _16074_ ( .A1(_05910_ ), .A2(_07197_ ), .ZN(_00342_ ) );
AND3_X1 _16075_ ( .A1(_06601_ ), .A2(\ID_EX_imm [25] ), .A3(_06598_ ), .ZN(_00343_ ) );
NOR3_X1 _16076_ ( .A1(_00341_ ), .A2(_00342_ ), .A3(_00343_ ), .ZN(_00344_ ) );
OAI21_X1 _16077_ ( .A(_03879_ ), .B1(_00344_ ), .B2(_07154_ ), .ZN(_00345_ ) );
NOR3_X1 _16078_ ( .A1(_07429_ ), .A2(_05181_ ), .A3(_05180_ ), .ZN(_00346_ ) );
OR3_X1 _16079_ ( .A1(_00346_ ), .A2(_05180_ ), .A3(_05188_ ), .ZN(_00347_ ) );
OAI21_X1 _16080_ ( .A(_05188_ ), .B1(_00346_ ), .B2(_05180_ ), .ZN(_00348_ ) );
NAND3_X1 _16081_ ( .A1(_00347_ ), .A2(_06685_ ), .A3(_00348_ ), .ZN(_00349_ ) );
AND3_X1 _16082_ ( .A1(_07158_ ), .A2(_06820_ ), .A3(_07159_ ), .ZN(_00350_ ) );
AND3_X1 _16083_ ( .A1(_00350_ ), .A2(_06867_ ), .A3(_06870_ ), .ZN(_00351_ ) );
NOR3_X1 _16084_ ( .A1(_05186_ ), .A2(_05187_ ), .A3(_06959_ ), .ZN(_00352_ ) );
NOR3_X1 _16085_ ( .A1(_05185_ ), .A2(_02946_ ), .A3(_07187_ ), .ZN(_00353_ ) );
AOI21_X1 _16086_ ( .A(_06872_ ), .B1(_05185_ ), .B2(_02946_ ), .ZN(_00354_ ) );
NOR4_X1 _16087_ ( .A1(_00351_ ), .A2(_00352_ ), .A3(_00353_ ), .A4(_00354_ ), .ZN(_00355_ ) );
OAI21_X1 _16088_ ( .A(_06752_ ), .B1(_07568_ ), .B2(_07569_ ), .ZN(_00356_ ) );
AND2_X1 _16089_ ( .A1(_00350_ ), .A2(_06797_ ), .ZN(_00357_ ) );
AOI21_X1 _16090_ ( .A(_00357_ ), .B1(_06749_ ), .B2(_07303_ ), .ZN(_00358_ ) );
AOI21_X1 _16091_ ( .A(_07351_ ), .B1(_00356_ ), .B2(_00358_ ), .ZN(_00359_ ) );
AOI21_X1 _16092_ ( .A(_07969_ ), .B1(_07584_ ), .B2(_07585_ ), .ZN(_00360_ ) );
NAND2_X1 _16093_ ( .A1(_07850_ ), .A2(_06966_ ), .ZN(_00361_ ) );
NAND3_X1 _16094_ ( .A1(_06836_ ), .A2(_06839_ ), .A3(_06740_ ), .ZN(_00362_ ) );
NAND3_X1 _16095_ ( .A1(_00361_ ), .A2(_00362_ ), .A3(_06918_ ), .ZN(_00363_ ) );
NAND2_X1 _16096_ ( .A1(_00363_ ), .A2(_07260_ ), .ZN(_00364_ ) );
AOI21_X1 _16097_ ( .A(_00364_ ), .B1(_06899_ ), .B2(_07184_ ), .ZN(_00365_ ) );
NOR3_X1 _16098_ ( .A1(_00359_ ), .A2(_00360_ ), .A3(_00365_ ), .ZN(_00366_ ) );
NAND3_X1 _16099_ ( .A1(_00349_ ), .A2(_00355_ ), .A3(_00366_ ), .ZN(_00367_ ) );
AOI21_X1 _16100_ ( .A(_00345_ ), .B1(_00367_ ), .B2(_06885_ ), .ZN(_00368_ ) );
OAI21_X1 _16101_ ( .A(_06272_ ), .B1(_05907_ ), .B2(_07492_ ), .ZN(_00369_ ) );
OAI21_X1 _16102_ ( .A(_00336_ ), .B1(_00368_ ), .B2(_00369_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _16103_ ( .A1(_05927_ ), .A2(_06424_ ), .ZN(_00370_ ) );
OAI21_X1 _16104_ ( .A(_06594_ ), .B1(_07471_ ), .B2(_00338_ ), .ZN(_00371_ ) );
AOI21_X1 _16105_ ( .A(_00371_ ), .B1(_00338_ ), .B2(_07471_ ), .ZN(_00372_ ) );
AND2_X1 _16106_ ( .A1(_05917_ ), .A2(_07197_ ), .ZN(_00373_ ) );
AND3_X1 _16107_ ( .A1(_06601_ ), .A2(\ID_EX_imm [24] ), .A3(_06598_ ), .ZN(_00374_ ) );
NOR3_X1 _16108_ ( .A1(_00372_ ), .A2(_00373_ ), .A3(_00374_ ), .ZN(_00375_ ) );
OAI21_X1 _16109_ ( .A(_03879_ ), .B1(_00375_ ), .B2(_07154_ ), .ZN(_00376_ ) );
AOI21_X1 _16110_ ( .A(_06998_ ), .B1(_07430_ ), .B2(_05182_ ), .ZN(_00377_ ) );
OAI21_X1 _16111_ ( .A(_00377_ ), .B1(_05182_ ), .B2(_07430_ ), .ZN(_00378_ ) );
NOR3_X1 _16112_ ( .A1(_05180_ ), .A2(_05181_ ), .A3(_06959_ ), .ZN(_00379_ ) );
NOR3_X1 _16113_ ( .A1(_05179_ ), .A2(_04622_ ), .A3(_07187_ ), .ZN(_00380_ ) );
AOI21_X1 _16114_ ( .A(_06873_ ), .B1(_05179_ ), .B2(_04622_ ), .ZN(_00381_ ) );
NOR3_X1 _16115_ ( .A1(_00379_ ), .A2(_00380_ ), .A3(_00381_ ), .ZN(_00382_ ) );
NAND4_X1 _16116_ ( .A1(_06724_ ), .A2(_07596_ ), .A3(_06733_ ), .A4(_06752_ ), .ZN(_00383_ ) );
AND3_X1 _16117_ ( .A1(_07204_ ), .A2(_06917_ ), .A3(_07206_ ), .ZN(_00384_ ) );
NAND2_X1 _16118_ ( .A1(_00384_ ), .A2(_06992_ ), .ZN(_00385_ ) );
NAND2_X1 _16119_ ( .A1(_00383_ ), .A2(_00385_ ), .ZN(_00386_ ) );
OAI21_X1 _16120_ ( .A(_06995_ ), .B1(_07021_ ), .B2(_00386_ ), .ZN(_00387_ ) );
NAND3_X1 _16121_ ( .A1(_07608_ ), .A2(_07609_ ), .A3(_07968_ ), .ZN(_00388_ ) );
NAND3_X1 _16122_ ( .A1(_06934_ ), .A2(_06937_ ), .A3(_06740_ ), .ZN(_00389_ ) );
NAND3_X1 _16123_ ( .A1(_07937_ ), .A2(_07938_ ), .A3(_06966_ ), .ZN(_00390_ ) );
NAND3_X1 _16124_ ( .A1(_00389_ ), .A2(_00390_ ), .A3(_06918_ ), .ZN(_00391_ ) );
OAI211_X1 _16125_ ( .A(_07260_ ), .B(_00391_ ), .C1(_07220_ ), .C2(_06918_ ), .ZN(_00392_ ) );
NAND3_X1 _16126_ ( .A1(_00384_ ), .A2(_06867_ ), .A3(_06869_ ), .ZN(_00393_ ) );
AND4_X1 _16127_ ( .A1(_00387_ ), .A2(_00388_ ), .A3(_00392_ ), .A4(_00393_ ), .ZN(_00394_ ) );
NAND3_X1 _16128_ ( .A1(_00378_ ), .A2(_00382_ ), .A3(_00394_ ), .ZN(_00395_ ) );
AOI21_X1 _16129_ ( .A(_00376_ ), .B1(_00395_ ), .B2(_06885_ ), .ZN(_00396_ ) );
OAI21_X1 _16130_ ( .A(_06272_ ), .B1(_05916_ ), .B2(_07492_ ), .ZN(_00397_ ) );
OAI21_X1 _16131_ ( .A(_00370_ ), .B1(_00396_ ), .B2(_00397_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
NOR4_X1 _16132_ ( .A1(_06588_ ), .A2(_06589_ ), .A3(_04846_ ), .A4(_04847_ ), .ZN(_00398_ ) );
OAI21_X1 _16133_ ( .A(_04773_ ), .B1(_00398_ ), .B2(_05246_ ), .ZN(_00399_ ) );
AND2_X1 _16134_ ( .A1(_00399_ ), .A2(_05259_ ), .ZN(_00400_ ) );
XNOR2_X1 _16135_ ( .A(_00400_ ), .B(_04798_ ), .ZN(_00401_ ) );
AND2_X1 _16136_ ( .A1(_00401_ ), .A2(_06595_ ), .ZN(_00402_ ) );
OAI22_X1 _16137_ ( .A1(_05947_ ), .A2(_07149_ ), .B1(_02283_ ), .B2(_07150_ ), .ZN(_00403_ ) );
OAI21_X1 _16138_ ( .A(_06583_ ), .B1(_00402_ ), .B2(_00403_ ), .ZN(_00404_ ) );
NAND2_X1 _16139_ ( .A1(_07001_ ), .A2(_07422_ ), .ZN(_00405_ ) );
AOI21_X1 _16140_ ( .A(_06863_ ), .B1(_04999_ ), .B2(_06679_ ), .ZN(_00406_ ) );
AND2_X1 _16141_ ( .A1(_00405_ ), .A2(_00406_ ), .ZN(_00407_ ) );
INV_X1 _16142_ ( .A(_04994_ ), .ZN(_00408_ ) );
OR2_X1 _16143_ ( .A1(_00407_ ), .A2(_00408_ ), .ZN(_00409_ ) );
INV_X1 _16144_ ( .A(_04988_ ), .ZN(_00410_ ) );
OR2_X1 _16145_ ( .A1(_04991_ ), .A2(_04749_ ), .ZN(_00411_ ) );
AND3_X1 _16146_ ( .A1(_00409_ ), .A2(_00410_ ), .A3(_00411_ ), .ZN(_00412_ ) );
AOI21_X1 _16147_ ( .A(_00410_ ), .B1(_00409_ ), .B2(_00411_ ), .ZN(_00413_ ) );
OR3_X1 _16148_ ( .A1(_00412_ ), .A2(_00413_ ), .A3(_06997_ ), .ZN(_00414_ ) );
AOI21_X1 _16149_ ( .A(_06751_ ), .B1(_06748_ ), .B2(_06735_ ), .ZN(_00415_ ) );
AND2_X1 _16150_ ( .A1(_07641_ ), .A2(_06992_ ), .ZN(_00416_ ) );
OAI21_X1 _16151_ ( .A(_06995_ ), .B1(_00415_ ), .B2(_00416_ ), .ZN(_00417_ ) );
NAND3_X1 _16152_ ( .A1(_07641_ ), .A2(_06992_ ), .A3(_06869_ ), .ZN(_00418_ ) );
AOI21_X1 _16153_ ( .A(_02282_ ), .B1(_04985_ ), .B2(_04986_ ), .ZN(_00419_ ) );
OAI21_X1 _16154_ ( .A(_00418_ ), .B1(_00419_ ), .B2(_06872_ ), .ZN(_00420_ ) );
NOR2_X1 _16155_ ( .A1(_07253_ ), .A2(_07137_ ), .ZN(_00421_ ) );
OAI21_X1 _16156_ ( .A(_06800_ ), .B1(_00421_ ), .B2(_06797_ ), .ZN(_00422_ ) );
NAND2_X1 _16157_ ( .A1(_07065_ ), .A2(_06739_ ), .ZN(_00423_ ) );
NAND2_X1 _16158_ ( .A1(_07973_ ), .A2(_06810_ ), .ZN(_00424_ ) );
NAND2_X1 _16159_ ( .A1(_00423_ ), .A2(_00424_ ), .ZN(_00425_ ) );
MUX2_X1 _16160_ ( .A(_07257_ ), .B(_00425_ ), .S(_06820_ ), .Z(_00426_ ) );
AOI21_X1 _16161_ ( .A(_00422_ ), .B1(_06955_ ), .B2(_00426_ ), .ZN(_00427_ ) );
OAI22_X1 _16162_ ( .A1(_00410_ ), .A2(_05207_ ), .B1(_07426_ ), .B2(_07078_ ), .ZN(_00428_ ) );
NOR3_X1 _16163_ ( .A1(_00420_ ), .A2(_00427_ ), .A3(_00428_ ), .ZN(_00429_ ) );
AND3_X1 _16164_ ( .A1(_00414_ ), .A2(_00417_ ), .A3(_00429_ ), .ZN(_00430_ ) );
OAI211_X1 _16165_ ( .A(_00404_ ), .B(_05360_ ), .C1(_06884_ ), .C2(_00430_ ), .ZN(_00431_ ) );
OR2_X1 _16166_ ( .A1(_05931_ ), .A2(_03879_ ), .ZN(_00432_ ) );
NAND3_X1 _16167_ ( .A1(_00431_ ), .A2(_06280_ ), .A3(_00432_ ), .ZN(_00433_ ) );
OAI21_X1 _16168_ ( .A(_06424_ ), .B1(_05939_ ), .B2(_05940_ ), .ZN(_00434_ ) );
NAND2_X1 _16169_ ( .A1(_00433_ ), .A2(_00434_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _16170_ ( .A1(_05963_ ), .A2(_06424_ ), .ZN(_00435_ ) );
NOR4_X1 _16171_ ( .A1(_07301_ ), .A2(_06735_ ), .A3(_06753_ ), .A4(_07673_ ), .ZN(_00436_ ) );
AND2_X1 _16172_ ( .A1(_07676_ ), .A2(_06796_ ), .ZN(_00437_ ) );
OR3_X1 _16173_ ( .A1(_00436_ ), .A2(_07021_ ), .A3(_00437_ ), .ZN(_00438_ ) );
AND2_X1 _16174_ ( .A1(_00438_ ), .A2(_06688_ ), .ZN(_00439_ ) );
OR3_X1 _16175_ ( .A1(_07326_ ), .A2(_06796_ ), .A3(_06898_ ), .ZN(_00440_ ) );
OR3_X1 _16176_ ( .A1(_07447_ ), .A2(_06793_ ), .A3(_07450_ ), .ZN(_00441_ ) );
OAI211_X1 _16177_ ( .A(_00441_ ), .B(_06954_ ), .C1(_06854_ ), .C2(_07323_ ), .ZN(_00442_ ) );
AOI21_X1 _16178_ ( .A(_07053_ ), .B1(_00440_ ), .B2(_00442_ ), .ZN(_00443_ ) );
AND3_X1 _16179_ ( .A1(_07676_ ), .A2(_06797_ ), .A3(_06868_ ), .ZN(_00444_ ) );
OR3_X1 _16180_ ( .A1(_00439_ ), .A2(_00443_ ), .A3(_00444_ ), .ZN(_00445_ ) );
AND2_X1 _16181_ ( .A1(_04994_ ), .A2(_06862_ ), .ZN(_00446_ ) );
NOR3_X1 _16182_ ( .A1(_04991_ ), .A2(_04749_ ), .A3(_07187_ ), .ZN(_00447_ ) );
AOI21_X1 _16183_ ( .A(_06872_ ), .B1(_04991_ ), .B2(_04749_ ), .ZN(_00448_ ) );
NOR4_X1 _16184_ ( .A1(_00445_ ), .A2(_00446_ ), .A3(_00447_ ), .A4(_00448_ ), .ZN(_00449_ ) );
NAND3_X1 _16185_ ( .A1(_00405_ ), .A2(_00408_ ), .A3(_00406_ ), .ZN(_00450_ ) );
NAND3_X1 _16186_ ( .A1(_00409_ ), .A2(_06685_ ), .A3(_00450_ ), .ZN(_00451_ ) );
AOI21_X1 _16187_ ( .A(_06884_ ), .B1(_00449_ ), .B2(_00451_ ), .ZN(_00452_ ) );
OR3_X1 _16188_ ( .A1(_00398_ ), .A2(_04773_ ), .A3(_05246_ ), .ZN(_00453_ ) );
NAND3_X1 _16189_ ( .A1(_00453_ ), .A2(_06595_ ), .A3(_00399_ ), .ZN(_00454_ ) );
AOI22_X1 _16190_ ( .A1(_05967_ ), .A2(_07197_ ), .B1(\ID_EX_imm [22] ), .B2(_06604_ ), .ZN(_00455_ ) );
AOI21_X1 _16191_ ( .A(_07154_ ), .B1(_00454_ ), .B2(_00455_ ), .ZN(_00456_ ) );
NOR3_X1 _16192_ ( .A1(_00452_ ), .A2(_05301_ ), .A3(_00456_ ), .ZN(_00457_ ) );
OAI21_X1 _16193_ ( .A(_06272_ ), .B1(_05965_ ), .B2(_07492_ ), .ZN(_00458_ ) );
OAI21_X1 _16194_ ( .A(_00435_ ), .B1(_00457_ ), .B2(_00458_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
OAI21_X1 _16195_ ( .A(_06333_ ), .B1(_06003_ ), .B2(_06004_ ), .ZN(_00459_ ) );
NAND3_X1 _16196_ ( .A1(_07441_ ), .A2(_04965_ ), .A3(_07466_ ), .ZN(_00460_ ) );
OAI21_X1 _16197_ ( .A(_04966_ ), .B1(_07440_ ), .B2(_07465_ ), .ZN(_00461_ ) );
NAND3_X1 _16198_ ( .A1(_00460_ ), .A2(_06685_ ), .A3(_00461_ ), .ZN(_00462_ ) );
NAND2_X1 _16199_ ( .A1(_06699_ ), .A2(_03006_ ), .ZN(_00463_ ) );
AOI21_X1 _16200_ ( .A(_07351_ ), .B1(_06751_ ), .B2(_00463_ ), .ZN(_00464_ ) );
AOI21_X1 _16201_ ( .A(_06852_ ), .B1(_07975_ ), .B2(_07976_ ), .ZN(_00465_ ) );
AOI21_X1 _16202_ ( .A(_06744_ ), .B1(_02173_ ), .B2(_02177_ ), .ZN(_00466_ ) );
OR2_X1 _16203_ ( .A1(_00466_ ), .A2(_06790_ ), .ZN(_00467_ ) );
MUX2_X1 _16204_ ( .A(_07852_ ), .B(_00467_ ), .S(_06931_ ), .Z(_00468_ ) );
AOI21_X1 _16205_ ( .A(_00465_ ), .B1(_00468_ ), .B2(_06966_ ), .ZN(_00469_ ) );
MUX2_X1 _16206_ ( .A(_00425_ ), .B(_00469_ ), .S(_06822_ ), .Z(_00470_ ) );
NOR2_X1 _16207_ ( .A1(_00470_ ), .A2(_07329_ ), .ZN(_00471_ ) );
AND3_X1 _16208_ ( .A1(_07254_ ), .A2(_07258_ ), .A3(_07968_ ), .ZN(_00472_ ) );
NAND3_X1 _16209_ ( .A1(_06699_ ), .A2(_03006_ ), .A3(_06869_ ), .ZN(_00473_ ) );
OAI21_X1 _16210_ ( .A(_06861_ ), .B1(_04962_ ), .B2(_04964_ ), .ZN(_00474_ ) );
NAND3_X1 _16211_ ( .A1(_06725_ ), .A2(_03006_ ), .A3(_06864_ ), .ZN(_00475_ ) );
OAI21_X1 _16212_ ( .A(_05288_ ), .B1(_06725_ ), .B2(_03006_ ), .ZN(_00476_ ) );
NAND4_X1 _16213_ ( .A1(_00473_ ), .A2(_00474_ ), .A3(_00475_ ), .A4(_00476_ ), .ZN(_00477_ ) );
NOR4_X1 _16214_ ( .A1(_00464_ ), .A2(_00471_ ), .A3(_00472_ ), .A4(_00477_ ), .ZN(_00478_ ) );
AOI21_X1 _16215_ ( .A(_06884_ ), .B1(_00462_ ), .B2(_00478_ ), .ZN(_00479_ ) );
OR3_X1 _16216_ ( .A1(_07477_ ), .A2(_04500_ ), .A3(_05270_ ), .ZN(_00480_ ) );
OAI21_X1 _16217_ ( .A(_04500_ ), .B1(_07477_ ), .B2(_05270_ ), .ZN(_00481_ ) );
NAND3_X1 _16218_ ( .A1(_00480_ ), .A2(_06595_ ), .A3(_00481_ ), .ZN(_00482_ ) );
NOR2_X1 _16219_ ( .A1(_06012_ ), .A2(_07149_ ), .ZN(_00483_ ) );
AOI21_X1 _16220_ ( .A(_00483_ ), .B1(\ID_EX_imm [31] ), .B2(_06604_ ), .ZN(_00484_ ) );
AOI21_X1 _16221_ ( .A(_07154_ ), .B1(_00482_ ), .B2(_00484_ ), .ZN(_00485_ ) );
NOR3_X1 _16222_ ( .A1(_00479_ ), .A2(_05301_ ), .A3(_00485_ ), .ZN(_00486_ ) );
OAI21_X1 _16223_ ( .A(_06272_ ), .B1(_05995_ ), .B2(_07492_ ), .ZN(_00487_ ) );
OAI21_X1 _16224_ ( .A(_00459_ ), .B1(_00486_ ), .B2(_00487_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
AND3_X1 _16225_ ( .A1(\myexu.state_$_ANDNOT__B_Y ), .A2(_03100_ ), .A3(_03888_ ), .ZN(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ) );
AOI21_X1 _16226_ ( .A(_02095_ ), .B1(_02069_ ), .B2(_02102_ ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16227_ ( .A(IDU_ready_IFU ), .ZN(_00488_ ) );
NAND2_X1 _16228_ ( .A1(_00488_ ), .A2(IDU_valid_EXU ), .ZN(_00489_ ) );
OAI21_X1 _16229_ ( .A(_00489_ ), .B1(_03340_ ), .B2(_03234_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16230_ ( .A1(_03307_ ), .A2(_03234_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16231_ ( .A1(_03307_ ), .A2(_03234_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16232_ ( .A(_03231_ ), .ZN(_00490_ ) );
NOR4_X1 _16233_ ( .A1(_03307_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03095_ ), .A4(_00490_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16234_ ( .A1(_03634_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03069_ ), .A4(_03230_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16235_ ( .A(_03829_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16236_ ( .A(_00489_ ), .B1(_00490_ ), .B2(_00488_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16237_ ( .A1(_03231_ ), .A2(_00488_ ), .B1(_01998_ ), .B2(_03345_ ), .ZN(_00491_ ) );
INV_X1 _16238_ ( .A(loaduse_clear ), .ZN(_00492_ ) );
AOI221_X4 _16239_ ( .A(_00491_ ), .B1(\myidu.state [2] ), .B2(_00492_ ), .C1(_03305_ ), .C2(_03829_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16240_ ( .A(_03360_ ), .B1(_03284_ ), .B2(_03370_ ), .ZN(_00493_ ) );
OAI211_X1 _16241_ ( .A(_03231_ ), .B(_03375_ ), .C1(_00493_ ), .C2(_03303_ ), .ZN(_00494_ ) );
NAND3_X1 _16242_ ( .A1(_03145_ ), .A2(IDU_valid_EXU ), .A3(_06049_ ), .ZN(_00495_ ) );
INV_X1 _16243_ ( .A(_00207_ ), .ZN(_00496_ ) );
OAI211_X1 _16244_ ( .A(_00494_ ), .B(_00495_ ), .C1(_00492_ ), .C2(_00496_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16245_ ( .A(_03145_ ), .B(_03886_ ), .C1(_03231_ ), .C2(_00488_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
AND3_X1 _16246_ ( .A1(_03355_ ), .A2(_03356_ ), .A3(_03357_ ), .ZN(_00497_ ) );
OAI21_X1 _16247_ ( .A(_00497_ ), .B1(_03359_ ), .B2(_03088_ ), .ZN(_00498_ ) );
AND2_X1 _16248_ ( .A1(_00498_ ), .A2(_03284_ ), .ZN(_00499_ ) );
NAND4_X1 _16249_ ( .A1(_03643_ ), .A2(_03229_ ), .A3(_03370_ ), .A4(_03375_ ), .ZN(_00500_ ) );
OAI22_X1 _16250_ ( .A1(_00499_ ), .A2(_00500_ ), .B1(loaduse_clear ), .B2(_00496_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16251_ ( .A1(_03228_ ), .A2(IDU_ready_IFU ), .ZN(_00501_ ) );
NOR2_X1 _16252_ ( .A1(_03228_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00502_ ) );
NOR2_X1 _16253_ ( .A1(\myifu.state [0] ), .A2(\myifu.state [1] ), .ZN(_00503_ ) );
NOR4_X1 _16254_ ( .A1(_00501_ ), .A2(_00502_ ), .A3(reset ), .A4(_00503_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
CLKBUF_X2 _16255_ ( .A(_06116_ ), .Z(_00504_ ) );
OR3_X1 _16256_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00505_ ) );
OAI21_X1 _16257_ ( .A(_00505_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06118_ ), .ZN(_00506_ ) );
MUX2_X1 _16258_ ( .A(\io_master_rdata [31] ), .B(_00506_ ), .S(_03818_ ), .Z(_00507_ ) );
AND2_X1 _16259_ ( .A1(_00507_ ), .A2(\io_master_arburst [0] ), .ZN(\myifu.data_in [31] ) );
BUF_X8 _16260_ ( .A(_03817_ ), .Z(_00508_ ) );
OR3_X1 _16261_ ( .A1(_01966_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00509_ ) );
OAI211_X1 _16262_ ( .A(_00508_ ), .B(_00509_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06117_ ), .ZN(_00510_ ) );
OAI21_X2 _16263_ ( .A(_00510_ ), .B1(_00508_ ), .B2(\io_master_rdata [30] ), .ZN(_00511_ ) );
NOR2_X1 _16264_ ( .A1(_00511_ ), .A2(_06082_ ), .ZN(\myifu.data_in [30] ) );
MUX2_X1 _16265_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06119_ ), .Z(_00512_ ) );
AND3_X1 _16266_ ( .A1(_06122_ ), .A2(_06123_ ), .A3(_00512_ ), .ZN(_00513_ ) );
AOI21_X1 _16267_ ( .A(\io_master_rdata [21] ), .B1(_06122_ ), .B2(_06123_ ), .ZN(_00514_ ) );
NOR3_X1 _16268_ ( .A1(_00513_ ), .A2(_00514_ ), .A3(_06081_ ), .ZN(\myifu.data_in [21] ) );
OR3_X1 _16269_ ( .A1(_01966_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00515_ ) );
OAI211_X1 _16270_ ( .A(_00508_ ), .B(_00515_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06117_ ), .ZN(_00516_ ) );
OAI21_X2 _16271_ ( .A(_00516_ ), .B1(\io_master_rdata [20] ), .B2(_00508_ ), .ZN(_00517_ ) );
NOR2_X1 _16272_ ( .A1(_00517_ ), .A2(_06083_ ), .ZN(\myifu.data_in [20] ) );
BUF_X2 _16273_ ( .A(_03818_ ), .Z(_00518_ ) );
OR2_X1 _16274_ ( .A1(_00518_ ), .A2(\io_master_rdata [19] ), .ZN(_00519_ ) );
CLKBUF_X2 _16275_ ( .A(_00504_ ), .Z(_00520_ ) );
OR3_X1 _16276_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00521_ ) );
OAI211_X1 _16277_ ( .A(_00518_ ), .B(_00521_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00522_ ) );
AND3_X1 _16278_ ( .A1(_00519_ ), .A2(_00522_ ), .A3(_02035_ ), .ZN(\myifu.data_in [19] ) );
OR2_X1 _16279_ ( .A1(_00518_ ), .A2(\io_master_rdata [18] ), .ZN(_00523_ ) );
OR3_X1 _16280_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00524_ ) );
OAI211_X1 _16281_ ( .A(_00518_ ), .B(_00524_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00525_ ) );
AND3_X1 _16282_ ( .A1(_00523_ ), .A2(_00525_ ), .A3(_02035_ ), .ZN(\myifu.data_in [18] ) );
MUX2_X1 _16283_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06119_ ), .Z(_00526_ ) );
AND3_X1 _16284_ ( .A1(_06122_ ), .A2(_06123_ ), .A3(_00526_ ), .ZN(_00527_ ) );
AOI21_X1 _16285_ ( .A(\io_master_rdata [17] ), .B1(_06122_ ), .B2(_06123_ ), .ZN(_00528_ ) );
NOR3_X1 _16286_ ( .A1(_00527_ ), .A2(_00528_ ), .A3(_01982_ ), .ZN(\myifu.data_in [17] ) );
MUX2_X1 _16287_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06119_ ), .Z(_00529_ ) );
AND3_X1 _16288_ ( .A1(_02077_ ), .A2(_02080_ ), .A3(_00529_ ), .ZN(_00530_ ) );
AOI21_X1 _16289_ ( .A(\io_master_rdata [16] ), .B1(_06122_ ), .B2(_06123_ ), .ZN(_00531_ ) );
NOR3_X1 _16290_ ( .A1(_00530_ ), .A2(_00531_ ), .A3(_01982_ ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16291_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00532_ ) );
OAI211_X1 _16292_ ( .A(_00508_ ), .B(_00532_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00533_ ) );
OAI21_X1 _16293_ ( .A(_00533_ ), .B1(_03818_ ), .B2(\io_master_rdata [15] ), .ZN(_00534_ ) );
NOR2_X1 _16294_ ( .A1(_00534_ ), .A2(_06083_ ), .ZN(\myifu.data_in [15] ) );
OR3_X1 _16295_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00535_ ) );
OAI211_X1 _16296_ ( .A(_03818_ ), .B(_00535_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00536_ ) );
OAI21_X1 _16297_ ( .A(_00536_ ), .B1(_03818_ ), .B2(\io_master_rdata [14] ), .ZN(_00537_ ) );
NOR2_X1 _16298_ ( .A1(_00537_ ), .A2(_06083_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16299_ ( .A1(_03820_ ), .A2(\io_master_rdata [13] ), .ZN(_00538_ ) );
CLKBUF_X2 _16300_ ( .A(_00520_ ), .Z(_00539_ ) );
OR3_X1 _16301_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00540_ ) );
OAI211_X1 _16302_ ( .A(_03820_ ), .B(_00540_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00541_ ) );
AND3_X1 _16303_ ( .A1(_00538_ ), .A2(_00541_ ), .A3(_02034_ ), .ZN(\myifu.data_in [13] ) );
OR3_X1 _16304_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00542_ ) );
OAI211_X1 _16305_ ( .A(_00518_ ), .B(_00542_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00543_ ) );
OAI21_X1 _16306_ ( .A(_00543_ ), .B1(_00518_ ), .B2(\io_master_rdata [12] ), .ZN(_00544_ ) );
NOR2_X1 _16307_ ( .A1(_00544_ ), .A2(_06083_ ), .ZN(\myifu.data_in [12] ) );
MUX2_X1 _16308_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06119_ ), .Z(_00545_ ) );
OR3_X1 _16309_ ( .A1(_02006_ ), .A2(_02031_ ), .A3(_00545_ ), .ZN(_00546_ ) );
OAI21_X1 _16310_ ( .A(\io_master_rdata [29] ), .B1(_02006_ ), .B2(_02031_ ), .ZN(_00547_ ) );
AOI21_X1 _16311_ ( .A(_06081_ ), .B1(_00546_ ), .B2(_00547_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16312_ ( .A1(_03819_ ), .A2(\io_master_rdata [11] ), .ZN(_00548_ ) );
OR3_X1 _16313_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00549_ ) );
OAI211_X1 _16314_ ( .A(_03820_ ), .B(_00549_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00550_ ) );
AND3_X1 _16315_ ( .A1(_00548_ ), .A2(_00550_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16316_ ( .A1(_03819_ ), .A2(\io_master_rdata [10] ), .ZN(_00551_ ) );
OR3_X1 _16317_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00552_ ) );
OAI211_X1 _16318_ ( .A(_03819_ ), .B(_00552_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06119_ ), .ZN(_00553_ ) );
AND3_X1 _16319_ ( .A1(_00551_ ), .A2(_00553_ ), .A3(_02035_ ), .ZN(\myifu.data_in [10] ) );
BUF_X2 _16320_ ( .A(_03820_ ), .Z(_00554_ ) );
OR2_X1 _16321_ ( .A1(_00554_ ), .A2(\io_master_rdata [9] ), .ZN(_00555_ ) );
OR3_X1 _16322_ ( .A1(_02034_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00556_ ) );
OAI211_X1 _16323_ ( .A(_00554_ ), .B(_00556_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00557_ ) );
AND3_X1 _16324_ ( .A1(_00555_ ), .A2(_00557_ ), .A3(_02035_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16325_ ( .A1(_03820_ ), .A2(\io_master_rdata [8] ), .ZN(_00558_ ) );
OR3_X1 _16326_ ( .A1(_02034_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00559_ ) );
OAI211_X1 _16327_ ( .A(_00554_ ), .B(_00559_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00560_ ) );
AND3_X1 _16328_ ( .A1(_00558_ ), .A2(_00560_ ), .A3(_02035_ ), .ZN(\myifu.data_in [8] ) );
OR2_X1 _16329_ ( .A1(_03819_ ), .A2(\io_master_rdata [7] ), .ZN(_00561_ ) );
OR3_X1 _16330_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00562_ ) );
OAI211_X1 _16331_ ( .A(_03819_ ), .B(_00562_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06119_ ), .ZN(_00563_ ) );
AND3_X1 _16332_ ( .A1(_00561_ ), .A2(_00563_ ), .A3(_02034_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16333_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00564_ ) );
OAI211_X1 _16334_ ( .A(_00508_ ), .B(_00564_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06117_ ), .ZN(_00565_ ) );
OAI21_X2 _16335_ ( .A(_00565_ ), .B1(_03818_ ), .B2(\io_master_rdata [6] ), .ZN(_00566_ ) );
NOR2_X1 _16336_ ( .A1(_00566_ ), .A2(_06082_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16337_ ( .A1(_02034_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00567_ ) );
OAI211_X1 _16338_ ( .A(_00554_ ), .B(_00567_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00568_ ) );
OAI21_X1 _16339_ ( .A(_00568_ ), .B1(_00554_ ), .B2(\io_master_rdata [5] ), .ZN(_00569_ ) );
NOR2_X1 _16340_ ( .A1(_00569_ ), .A2(_06083_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16341_ ( .A1(_01966_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00570_ ) );
OAI211_X1 _16342_ ( .A(_00508_ ), .B(_00570_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06117_ ), .ZN(_00571_ ) );
OAI21_X2 _16343_ ( .A(_00571_ ), .B1(_00508_ ), .B2(\io_master_rdata [4] ), .ZN(_00572_ ) );
NOR2_X1 _16344_ ( .A1(_00572_ ), .A2(_06083_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16345_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00573_ ) );
OAI211_X1 _16346_ ( .A(_00518_ ), .B(_00573_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00574_ ) );
OAI21_X1 _16347_ ( .A(_00574_ ), .B1(_00518_ ), .B2(\io_master_rdata [3] ), .ZN(_00575_ ) );
NOR2_X1 _16348_ ( .A1(_00575_ ), .A2(_06083_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16349_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00576_ ) );
OAI211_X1 _16350_ ( .A(_03818_ ), .B(_00576_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00577_ ) );
OAI21_X1 _16351_ ( .A(_00577_ ), .B1(_00518_ ), .B2(\io_master_rdata [2] ), .ZN(_00578_ ) );
NOR2_X1 _16352_ ( .A1(_00578_ ), .A2(_06083_ ), .ZN(\myifu.data_in [2] ) );
OR3_X1 _16353_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00579_ ) );
OAI211_X1 _16354_ ( .A(_03818_ ), .B(_00579_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06118_ ), .ZN(_00580_ ) );
OAI21_X1 _16355_ ( .A(_00580_ ), .B1(_03818_ ), .B2(\io_master_rdata [28] ), .ZN(_00581_ ) );
NOR2_X1 _16356_ ( .A1(_00581_ ), .A2(_06081_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16357_ ( .A1(_02034_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00582_ ) );
OAI211_X1 _16358_ ( .A(_00554_ ), .B(_00582_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00583_ ) );
OAI21_X1 _16359_ ( .A(_00583_ ), .B1(_00554_ ), .B2(\io_master_rdata [1] ), .ZN(_00584_ ) );
NOR2_X1 _16360_ ( .A1(_00584_ ), .A2(_06083_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16361_ ( .A1(_02034_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00539_ ), .ZN(_00585_ ) );
OAI211_X1 _16362_ ( .A(_03820_ ), .B(_00585_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00586_ ) );
OAI21_X1 _16363_ ( .A(_00586_ ), .B1(\io_master_rdata [0] ), .B2(_03820_ ), .ZN(_00587_ ) );
NOR2_X1 _16364_ ( .A1(_00587_ ), .A2(_06081_ ), .ZN(\myifu.data_in [0] ) );
OR2_X1 _16365_ ( .A1(_03819_ ), .A2(\io_master_rdata [27] ), .ZN(_00588_ ) );
OR3_X1 _16366_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00589_ ) );
OAI211_X1 _16367_ ( .A(_03819_ ), .B(_00589_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06119_ ), .ZN(_00590_ ) );
AND3_X1 _16368_ ( .A1(_00588_ ), .A2(_00590_ ), .A3(_02035_ ), .ZN(\myifu.data_in [27] ) );
OR3_X1 _16369_ ( .A1(_02033_ ), .A2(_01693_ ), .A3(_00520_ ), .ZN(_00591_ ) );
OAI211_X1 _16370_ ( .A(_03819_ ), .B(_00591_ ), .C1(_01677_ ), .C2(_06119_ ), .ZN(_00592_ ) );
OAI21_X1 _16371_ ( .A(\io_master_rdata [26] ), .B1(_02006_ ), .B2(_02031_ ), .ZN(_00593_ ) );
AOI21_X1 _16372_ ( .A(_06081_ ), .B1(_00592_ ), .B2(_00593_ ), .ZN(\myifu.data_in [26] ) );
OR2_X1 _16373_ ( .A1(_00554_ ), .A2(\io_master_rdata [25] ), .ZN(_00594_ ) );
OR3_X1 _16374_ ( .A1(_02034_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00539_ ), .ZN(_00595_ ) );
OAI211_X1 _16375_ ( .A(_00554_ ), .B(_00595_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00596_ ) );
AND3_X1 _16376_ ( .A1(_00594_ ), .A2(_00596_ ), .A3(_02035_ ), .ZN(\myifu.data_in [25] ) );
OR3_X1 _16377_ ( .A1(_02034_ ), .A2(_01758_ ), .A3(_00539_ ), .ZN(_00597_ ) );
OAI211_X1 _16378_ ( .A(_03820_ ), .B(_00597_ ), .C1(_01683_ ), .C2(\io_master_araddr [2] ), .ZN(_00598_ ) );
OAI21_X1 _16379_ ( .A(\io_master_rdata [24] ), .B1(_02006_ ), .B2(_02031_ ), .ZN(_00599_ ) );
AOI21_X1 _16380_ ( .A(_06081_ ), .B1(_00598_ ), .B2(_00599_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16381_ ( .A1(_02033_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00520_ ), .ZN(_00600_ ) );
OAI211_X1 _16382_ ( .A(_00518_ ), .B(_00600_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06119_ ), .ZN(_00601_ ) );
OAI21_X1 _16383_ ( .A(_00601_ ), .B1(_03819_ ), .B2(\io_master_rdata [23] ), .ZN(_00602_ ) );
NOR2_X1 _16384_ ( .A1(_00602_ ), .A2(_06081_ ), .ZN(\myifu.data_in [23] ) );
OR3_X1 _16385_ ( .A1(_02032_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00504_ ), .ZN(_00603_ ) );
OAI211_X1 _16386_ ( .A(_00508_ ), .B(_00603_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06117_ ), .ZN(_00604_ ) );
OAI21_X2 _16387_ ( .A(_00604_ ), .B1(\io_master_rdata [22] ), .B2(_00508_ ), .ZN(_00605_ ) );
NOR2_X1 _16388_ ( .A1(_00605_ ), .A2(_06081_ ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16389_ ( .A(_00241_ ), .ZN(_00606_ ) );
NAND2_X1 _16390_ ( .A1(_00606_ ), .A2(_02071_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16391_ ( .A1(_06044_ ), .A2(fanout_net_7 ), .ZN(_00607_ ) );
INV_X1 _16392_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00608_ ) );
OAI21_X1 _16393_ ( .A(_02071_ ), .B1(_00607_ ), .B2(_00608_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16394_ ( .A1(_06048_ ), .A2(fanout_net_11 ), .ZN(_00609_ ) );
OAI21_X1 _16395_ ( .A(_02071_ ), .B1(_00609_ ), .B2(_00608_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16396_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .ZN(_00610_ ) );
OAI21_X1 _16397_ ( .A(_02071_ ), .B1(_00610_ ), .B2(_00608_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
OAI21_X1 _16398_ ( .A(\IF_ID_inst [8] ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_00611_ ) );
NOR2_X1 _16399_ ( .A1(_03264_ ), .A2(_03265_ ), .ZN(_00612_ ) );
INV_X1 _16400_ ( .A(_03167_ ), .ZN(_00613_ ) );
AND2_X1 _16401_ ( .A1(_00612_ ), .A2(_00613_ ), .ZN(_00614_ ) );
AND2_X1 _16402_ ( .A1(_03391_ ), .A2(_03398_ ), .ZN(_00615_ ) );
INV_X1 _16403_ ( .A(_03260_ ), .ZN(_00616_ ) );
NOR4_X1 _16404_ ( .A1(_03377_ ), .A2(_03162_ ), .A3(_00616_ ), .A4(_03316_ ), .ZN(_00617_ ) );
NAND3_X1 _16405_ ( .A1(_00614_ ), .A2(_00615_ ), .A3(_00617_ ), .ZN(_00618_ ) );
AND2_X1 _16406_ ( .A1(_00618_ ), .A2(_03557_ ), .ZN(_00619_ ) );
OAI221_X1 _16407_ ( .A(_00611_ ), .B1(_03309_ ), .B2(_03087_ ), .C1(_00619_ ), .C2(_03085_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
AND2_X1 _16408_ ( .A1(_03162_ ), .A2(\IF_ID_inst [31] ), .ZN(_00620_ ) );
INV_X1 _16409_ ( .A(_00620_ ), .ZN(_00621_ ) );
OAI221_X1 _16410_ ( .A(_00621_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_03302_ ), .C1(_00614_ ), .C2(_03066_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
NOR2_X1 _16411_ ( .A1(_03302_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_00622_ ) );
INV_X1 _16412_ ( .A(_00622_ ), .ZN(_00623_ ) );
OAI21_X1 _16413_ ( .A(\IF_ID_inst [31] ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_00624_ ) );
AND2_X1 _16414_ ( .A1(_00623_ ), .A2(_00624_ ), .ZN(_00625_ ) );
BUF_X4 _16415_ ( .A(_00625_ ), .Z(_00626_ ) );
BUF_X4 _16416_ ( .A(_00621_ ), .Z(_00627_ ) );
BUF_X4 _16417_ ( .A(_00613_ ), .Z(_00628_ ) );
OAI211_X1 _16418_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03084_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16419_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03085_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16420_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03089_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
BUF_X2 _16421_ ( .A(_03302_ ), .Z(_00629_ ) );
OAI221_X1 _16422_ ( .A(_00624_ ), .B1(_03170_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI221_X1 _16423_ ( .A(_00624_ ), .B1(_03181_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI221_X1 _16424_ ( .A(_00624_ ), .B1(_03182_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16425_ ( .A(_00624_ ), .B1(_03309_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _16426_ ( .A(_00624_ ), .B1(_03121_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16427_ ( .A(_00624_ ), .B1(_03118_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16428_ ( .A(_00624_ ), .B1(_03119_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16429_ ( .A(_00624_ ), .B1(_03106_ ), .B2(_03168_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16430_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03090_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
OR2_X1 _16431_ ( .A1(_03153_ ), .A2(_03066_ ), .ZN(_00630_ ) );
NAND3_X1 _16432_ ( .A1(_03262_ ), .A2(\IF_ID_inst [7] ), .A3(_03263_ ), .ZN(_00631_ ) );
NAND4_X1 _16433_ ( .A1(_00623_ ), .A2(_03496_ ), .A3(_00630_ ), .A4(_00631_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
OAI21_X1 _16434_ ( .A(\IF_ID_inst [30] ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_00632_ ) );
OAI221_X1 _16435_ ( .A(_00632_ ), .B1(_03084_ ), .B2(_03557_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
INV_X1 _16436_ ( .A(_03505_ ), .ZN(_00633_ ) );
OAI221_X1 _16437_ ( .A(_00633_ ), .B1(_00612_ ), .B2(_03090_ ), .C1(_00629_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16438_ ( .A(_03515_ ), .ZN(_00634_ ) );
OAI221_X1 _16439_ ( .A(_00634_ ), .B1(_00612_ ), .B2(_03091_ ), .C1(_03302_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
INV_X1 _16440_ ( .A(_03519_ ), .ZN(_00635_ ) );
OAI221_X1 _16441_ ( .A(_00635_ ), .B1(_00612_ ), .B2(_03092_ ), .C1(_03302_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
OAI21_X1 _16442_ ( .A(\IF_ID_inst [26] ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_00636_ ) );
OAI221_X1 _16443_ ( .A(_00636_ ), .B1(_03093_ ), .B2(_03557_ ), .C1(_03302_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
OAI21_X1 _16444_ ( .A(\IF_ID_inst [25] ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_00637_ ) );
OAI221_X1 _16445_ ( .A(_00637_ ), .B1(_03094_ ), .B2(_03557_ ), .C1(_03302_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16446_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03091_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16447_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03092_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16448_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03093_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16449_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03094_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16450_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03096_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16451_ ( .A(_00626_ ), .B(_00627_ ), .C1(_03097_ ), .C2(_00628_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16452_ ( .A(_00625_ ), .B(_00621_ ), .C1(_03098_ ), .C2(_00613_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OR2_X1 _16453_ ( .A1(_03087_ ), .A2(_03170_ ), .ZN(_00638_ ) );
OAI221_X1 _16454_ ( .A(_00638_ ), .B1(_03113_ ), .B2(_00612_ ), .C1(_00619_ ), .C2(_03096_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OR2_X1 _16455_ ( .A1(_03087_ ), .A2(_03181_ ), .ZN(_00639_ ) );
OAI221_X1 _16456_ ( .A(_00639_ ), .B1(_03114_ ), .B2(_00612_ ), .C1(_00619_ ), .C2(_03097_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16457_ ( .A(\IF_ID_inst [9] ), .B1(_03264_ ), .B2(_03265_ ), .ZN(_00640_ ) );
OAI221_X1 _16458_ ( .A(_00640_ ), .B1(_03182_ ), .B2(_03087_ ), .C1(_00619_ ), .C2(_03098_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16459_ ( .A1(_03153_ ), .A2(_03117_ ), .ZN(_00641_ ) );
OAI221_X1 _16460_ ( .A(_00641_ ), .B1(_03121_ ), .B2(_03087_ ), .C1(_00618_ ), .C2(_03089_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AND3_X1 _16461_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00642_ ) );
CLKBUF_X2 _16462_ ( .A(_06041_ ), .Z(_00643_ ) );
AND3_X1 _16463_ ( .A1(_00643_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00644_ ) );
BUF_X4 _16464_ ( .A(_06039_ ), .Z(_00645_ ) );
BUF_X4 _16465_ ( .A(_00645_ ), .Z(_00646_ ) );
AOI211_X1 _16466_ ( .A(_00642_ ), .B(_00644_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_00646_ ), .ZN(_00647_ ) );
NAND2_X1 _16467_ ( .A1(_00608_ ), .A2(\IF_ID_pc [2] ), .ZN(_00648_ ) );
BUF_X4 _16468_ ( .A(_00648_ ), .Z(_00649_ ) );
BUF_X4 _16469_ ( .A(_00649_ ), .Z(_00650_ ) );
NAND2_X1 _16470_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00651_ ) );
BUF_X4 _16471_ ( .A(_00651_ ), .Z(_00652_ ) );
BUF_X4 _16472_ ( .A(_00652_ ), .Z(_00653_ ) );
BUF_X4 _16473_ ( .A(_06046_ ), .Z(_00654_ ) );
BUF_X4 _16474_ ( .A(_00654_ ), .Z(_00655_ ) );
NAND3_X1 _16475_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00656_ ) );
NAND4_X1 _16476_ ( .A1(_00647_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00656_ ), .ZN(_00657_ ) );
NOR2_X1 _16477_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00658_ ) );
BUF_X2 _16478_ ( .A(_00658_ ), .Z(_00659_ ) );
BUF_X4 _16479_ ( .A(_00659_ ), .Z(_00660_ ) );
BUF_X4 _16480_ ( .A(_06041_ ), .Z(_00661_ ) );
BUF_X4 _16481_ ( .A(_00661_ ), .Z(_00662_ ) );
NAND3_X1 _16482_ ( .A1(_00662_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00663_ ) );
NAND3_X1 _16483_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00664_ ) );
AND2_X1 _16484_ ( .A1(_00663_ ), .A2(_00664_ ), .ZN(_00665_ ) );
NAND2_X1 _16485_ ( .A1(_00648_ ), .A2(_00651_ ), .ZN(_00666_ ) );
BUF_X4 _16486_ ( .A(_00666_ ), .Z(_00667_ ) );
BUF_X4 _16487_ ( .A(_00667_ ), .Z(_00668_ ) );
BUF_X4 _16488_ ( .A(_06047_ ), .Z(_00669_ ) );
NAND3_X1 _16489_ ( .A1(_00669_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00670_ ) );
BUF_X4 _16490_ ( .A(_06043_ ), .Z(_00671_ ) );
BUF_X4 _16491_ ( .A(_06045_ ), .Z(_00672_ ) );
BUF_X4 _16492_ ( .A(_00672_ ), .Z(_00673_ ) );
NAND3_X1 _16493_ ( .A1(_00671_ ), .A2(_00673_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00674_ ) );
NAND4_X1 _16494_ ( .A1(_00665_ ), .A2(_00668_ ), .A3(_00670_ ), .A4(_00674_ ), .ZN(_00675_ ) );
NAND3_X1 _16495_ ( .A1(_00657_ ), .A2(_00660_ ), .A3(_00675_ ), .ZN(_00676_ ) );
NAND2_X1 _16496_ ( .A1(_03816_ ), .A2(_03825_ ), .ZN(_00677_ ) );
XOR2_X1 _16497_ ( .A(\IF_ID_pc [2] ), .B(\myifu.tmp_offset [2] ), .Z(_00678_ ) );
NAND2_X1 _16498_ ( .A1(_03542_ ), .A2(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .ZN(_00679_ ) );
NOR2_X1 _16499_ ( .A1(_00678_ ), .A2(_00679_ ), .ZN(_00680_ ) );
INV_X1 _16500_ ( .A(_00680_ ), .ZN(_00681_ ) );
NOR2_X1 _16501_ ( .A1(_00677_ ), .A2(_00681_ ), .ZN(_00682_ ) );
BUF_X4 _16502_ ( .A(_00682_ ), .Z(_00683_ ) );
OAI21_X1 _16503_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03539_ ), .ZN(_00684_ ) );
BUF_X4 _16504_ ( .A(_00677_ ), .Z(_00685_ ) );
BUF_X4 _16505_ ( .A(_00685_ ), .Z(_00686_ ) );
BUF_X4 _16506_ ( .A(_00681_ ), .Z(_00687_ ) );
BUF_X4 _16507_ ( .A(_00687_ ), .Z(_00688_ ) );
NOR3_X1 _16508_ ( .A1(\myifu.data_in [8] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_00689_ ) );
OAI21_X1 _16509_ ( .A(_00676_ ), .B1(_00684_ ), .B2(_00689_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16510_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00690_ ) );
AND3_X1 _16511_ ( .A1(_00643_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00691_ ) );
AOI211_X1 _16512_ ( .A(_00690_ ), .B(_00691_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00646_ ), .ZN(_00692_ ) );
NAND3_X1 _16513_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00693_ ) );
NAND4_X1 _16514_ ( .A1(_00692_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00693_ ), .ZN(_00694_ ) );
BUF_X4 _16515_ ( .A(_00659_ ), .Z(_00695_ ) );
NAND3_X1 _16516_ ( .A1(_00662_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00696_ ) );
NAND3_X1 _16517_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00697_ ) );
AND2_X1 _16518_ ( .A1(_00696_ ), .A2(_00697_ ), .ZN(_00698_ ) );
NAND3_X1 _16519_ ( .A1(_00669_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00699_ ) );
NAND3_X1 _16520_ ( .A1(_00671_ ), .A2(_00673_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00700_ ) );
NAND4_X1 _16521_ ( .A1(_00698_ ), .A2(_00668_ ), .A3(_00699_ ), .A4(_00700_ ), .ZN(_00701_ ) );
NAND3_X1 _16522_ ( .A1(_00694_ ), .A2(_00695_ ), .A3(_00701_ ), .ZN(_00702_ ) );
AOI211_X1 _16523_ ( .A(_00687_ ), .B(_00685_ ), .C1(\io_master_arburst [0] ), .C2(_00507_ ), .ZN(_00703_ ) );
BUF_X4 _16524_ ( .A(_00682_ ), .Z(_00704_ ) );
OAI21_X1 _16525_ ( .A(\myifu.state [2] ), .B1(_00704_ ), .B2(_03269_ ), .ZN(_00705_ ) );
OAI21_X1 _16526_ ( .A(_00702_ ), .B1(_00703_ ), .B2(_00705_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
AND3_X1 _16527_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00706_ ) );
CLKBUF_X2 _16528_ ( .A(_06041_ ), .Z(_00707_ ) );
AND3_X1 _16529_ ( .A1(_00707_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00708_ ) );
AOI211_X1 _16530_ ( .A(_00706_ ), .B(_00708_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_00646_ ), .ZN(_00709_ ) );
NAND3_X1 _16531_ ( .A1(_00655_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00710_ ) );
NAND4_X1 _16532_ ( .A1(_00709_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00710_ ), .ZN(_00711_ ) );
NAND3_X1 _16533_ ( .A1(_00662_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00712_ ) );
NAND3_X1 _16534_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00713_ ) );
AND2_X1 _16535_ ( .A1(_00712_ ), .A2(_00713_ ), .ZN(_00714_ ) );
NAND3_X1 _16536_ ( .A1(_00669_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00715_ ) );
NAND3_X1 _16537_ ( .A1(_00671_ ), .A2(_00673_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00716_ ) );
NAND4_X1 _16538_ ( .A1(_00714_ ), .A2(_00668_ ), .A3(_00715_ ), .A4(_00716_ ), .ZN(_00717_ ) );
NAND3_X1 _16539_ ( .A1(_00711_ ), .A2(_00695_ ), .A3(_00717_ ), .ZN(_00718_ ) );
OAI21_X1 _16540_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03510_ ), .ZN(_00719_ ) );
NOR3_X1 _16541_ ( .A1(\myifu.data_in [30] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_00720_ ) );
OAI21_X1 _16542_ ( .A(_00718_ ), .B1(_00719_ ), .B2(_00720_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
INV_X1 _16543_ ( .A(\myifu.state [2] ), .ZN(_00721_ ) );
BUF_X4 _16544_ ( .A(_00721_ ), .Z(_00722_ ) );
NOR3_X1 _16545_ ( .A1(_00685_ ), .A2(\myifu.data_in [21] ), .A3(_00687_ ), .ZN(_00723_ ) );
INV_X1 _16546_ ( .A(_00682_ ), .ZN(_00724_ ) );
BUF_X4 _16547_ ( .A(_00724_ ), .Z(_00725_ ) );
AOI211_X1 _16548_ ( .A(_00722_ ), .B(_00723_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00725_ ), .ZN(_00726_ ) );
AND3_X1 _16549_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00727_ ) );
AND3_X1 _16550_ ( .A1(_06042_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00728_ ) );
AOI211_X1 _16551_ ( .A(_00727_ ), .B(_00728_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_00645_ ), .ZN(_00729_ ) );
NAND3_X1 _16552_ ( .A1(_00654_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00730_ ) );
NAND4_X1 _16553_ ( .A1(_00729_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_00730_ ), .ZN(_00731_ ) );
NAND3_X1 _16554_ ( .A1(_00661_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00732_ ) );
NAND3_X1 _16555_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00733_ ) );
AND2_X1 _16556_ ( .A1(_00732_ ), .A2(_00733_ ), .ZN(_00734_ ) );
NAND3_X1 _16557_ ( .A1(_06047_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00735_ ) );
NAND3_X1 _16558_ ( .A1(_06043_ ), .A2(_06046_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00736_ ) );
NAND4_X1 _16559_ ( .A1(_00734_ ), .A2(_00667_ ), .A3(_00735_ ), .A4(_00736_ ), .ZN(_00737_ ) );
AND3_X1 _16560_ ( .A1(_00731_ ), .A2(_00659_ ), .A3(_00737_ ), .ZN(_00738_ ) );
OR2_X1 _16561_ ( .A1(_00726_ ), .A2(_00738_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
AOI21_X1 _16562_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00739_ ) );
OAI21_X1 _16563_ ( .A(_00704_ ), .B1(_06090_ ), .B2(_00517_ ), .ZN(_00740_ ) );
NAND2_X1 _16564_ ( .A1(_00739_ ), .A2(_00740_ ), .ZN(_00741_ ) );
AND3_X1 _16565_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00742_ ) );
AND3_X1 _16566_ ( .A1(_06043_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00743_ ) );
AOI211_X1 _16567_ ( .A(_00742_ ), .B(_00743_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_06040_ ), .ZN(_00744_ ) );
BUF_X2 _16568_ ( .A(_00648_ ), .Z(_00745_ ) );
BUF_X4 _16569_ ( .A(_00652_ ), .Z(_00746_ ) );
NAND3_X1 _16570_ ( .A1(_06048_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00747_ ) );
NAND4_X1 _16571_ ( .A1(_00744_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_00747_ ), .ZN(_00748_ ) );
BUF_X4 _16572_ ( .A(_00661_ ), .Z(_00749_ ) );
NAND3_X1 _16573_ ( .A1(_00749_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00750_ ) );
NAND3_X1 _16574_ ( .A1(fanout_net_11 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00751_ ) );
AND2_X1 _16575_ ( .A1(_00750_ ), .A2(_00751_ ), .ZN(_00752_ ) );
BUF_X2 _16576_ ( .A(_00666_ ), .Z(_00753_ ) );
BUF_X4 _16577_ ( .A(_06046_ ), .Z(_00754_ ) );
BUF_X4 _16578_ ( .A(_00754_ ), .Z(_00755_ ) );
NAND3_X1 _16579_ ( .A1(_00755_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00756_ ) );
BUF_X4 _16580_ ( .A(_06047_ ), .Z(_00757_ ) );
NAND3_X1 _16581_ ( .A1(_06044_ ), .A2(_00757_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00758_ ) );
NAND4_X1 _16582_ ( .A1(_00752_ ), .A2(_00753_ ), .A3(_00756_ ), .A4(_00758_ ), .ZN(_00759_ ) );
NAND3_X1 _16583_ ( .A1(_00748_ ), .A2(_00660_ ), .A3(_00759_ ), .ZN(_00760_ ) );
NAND2_X1 _16584_ ( .A1(_00741_ ), .A2(_00760_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
BUF_X4 _16585_ ( .A(_00721_ ), .Z(_00761_ ) );
NOR3_X1 _16586_ ( .A1(\myifu.data_in [19] ), .A2(_00685_ ), .A3(_00687_ ), .ZN(_00762_ ) );
BUF_X4 _16587_ ( .A(_00724_ ), .Z(_00763_ ) );
AOI211_X1 _16588_ ( .A(_00761_ ), .B(_00762_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_00764_ ) );
AND3_X1 _16589_ ( .A1(fanout_net_12 ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00765_ ) );
AND3_X1 _16590_ ( .A1(_06042_ ), .A2(fanout_net_7 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00766_ ) );
AOI211_X1 _16591_ ( .A(_00765_ ), .B(_00766_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_00645_ ), .ZN(_00767_ ) );
NAND3_X1 _16592_ ( .A1(_00654_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00768_ ) );
NAND4_X1 _16593_ ( .A1(_00767_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_00768_ ), .ZN(_00769_ ) );
NAND3_X1 _16594_ ( .A1(_00661_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00770_ ) );
NAND3_X1 _16595_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00771_ ) );
AND2_X1 _16596_ ( .A1(_00770_ ), .A2(_00771_ ), .ZN(_00772_ ) );
NAND3_X1 _16597_ ( .A1(_06047_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00773_ ) );
NAND3_X1 _16598_ ( .A1(_06043_ ), .A2(_06046_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00774_ ) );
NAND4_X1 _16599_ ( .A1(_00772_ ), .A2(_00667_ ), .A3(_00773_ ), .A4(_00774_ ), .ZN(_00775_ ) );
AND3_X1 _16600_ ( .A1(_00769_ ), .A2(_00659_ ), .A3(_00775_ ), .ZN(_00776_ ) );
OR2_X1 _16601_ ( .A1(_00764_ ), .A2(_00776_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
NOR3_X1 _16602_ ( .A1(\myifu.data_in [18] ), .A2(_00685_ ), .A3(_00687_ ), .ZN(_00777_ ) );
AOI211_X1 _16603_ ( .A(_00761_ ), .B(_00777_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_00778_ ) );
NAND3_X1 _16604_ ( .A1(_00661_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00779_ ) );
NAND3_X1 _16605_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00780_ ) );
AND2_X1 _16606_ ( .A1(_00779_ ), .A2(_00780_ ), .ZN(_00781_ ) );
BUF_X4 _16607_ ( .A(_00666_ ), .Z(_00782_ ) );
NAND3_X1 _16608_ ( .A1(_00754_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00783_ ) );
BUF_X4 _16609_ ( .A(_06042_ ), .Z(_00784_ ) );
NAND3_X1 _16610_ ( .A1(_00784_ ), .A2(_06047_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00785_ ) );
NAND4_X1 _16611_ ( .A1(_00781_ ), .A2(_00782_ ), .A3(_00783_ ), .A4(_00785_ ), .ZN(_00786_ ) );
AND3_X1 _16612_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00787_ ) );
AND3_X1 _16613_ ( .A1(_06041_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00788_ ) );
AOI211_X1 _16614_ ( .A(_00787_ ), .B(_00788_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_06039_ ), .ZN(_00789_ ) );
NAND3_X1 _16615_ ( .A1(_00672_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00790_ ) );
NAND4_X1 _16616_ ( .A1(_00789_ ), .A2(_00648_ ), .A3(_00651_ ), .A4(_00790_ ), .ZN(_00791_ ) );
AND3_X1 _16617_ ( .A1(_00786_ ), .A2(_00659_ ), .A3(_00791_ ), .ZN(_00792_ ) );
OR2_X1 _16618_ ( .A1(_00778_ ), .A2(_00792_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
NOR3_X1 _16619_ ( .A1(_00685_ ), .A2(\myifu.data_in [17] ), .A3(_00687_ ), .ZN(_00793_ ) );
AOI211_X1 _16620_ ( .A(_00761_ ), .B(_00793_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_00794_ ) );
AND3_X1 _16621_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00795_ ) );
AND3_X1 _16622_ ( .A1(_06042_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00796_ ) );
AOI211_X1 _16623_ ( .A(_00795_ ), .B(_00796_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_00645_ ), .ZN(_00797_ ) );
NAND3_X1 _16624_ ( .A1(_00654_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00798_ ) );
NAND4_X1 _16625_ ( .A1(_00797_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_00798_ ), .ZN(_00799_ ) );
NAND3_X1 _16626_ ( .A1(_00661_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00800_ ) );
NAND3_X1 _16627_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00801_ ) );
AND2_X1 _16628_ ( .A1(_00800_ ), .A2(_00801_ ), .ZN(_00802_ ) );
NAND3_X1 _16629_ ( .A1(_00672_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00803_ ) );
NAND3_X1 _16630_ ( .A1(_06043_ ), .A2(_06046_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00804_ ) );
NAND4_X1 _16631_ ( .A1(_00802_ ), .A2(_00667_ ), .A3(_00803_ ), .A4(_00804_ ), .ZN(_00805_ ) );
AND3_X1 _16632_ ( .A1(_00799_ ), .A2(_00659_ ), .A3(_00805_ ), .ZN(_00806_ ) );
OR2_X1 _16633_ ( .A1(_00794_ ), .A2(_00806_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NOR3_X1 _16634_ ( .A1(_00685_ ), .A2(\myifu.data_in [16] ), .A3(_00687_ ), .ZN(_00807_ ) );
AOI211_X1 _16635_ ( .A(_00761_ ), .B(_00807_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_00808_ ) );
AND3_X1 _16636_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00809_ ) );
AND3_X1 _16637_ ( .A1(_06042_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00810_ ) );
AOI211_X1 _16638_ ( .A(_00809_ ), .B(_00810_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_00645_ ), .ZN(_00811_ ) );
NAND3_X1 _16639_ ( .A1(_00654_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00812_ ) );
NAND4_X1 _16640_ ( .A1(_00811_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_00812_ ), .ZN(_00813_ ) );
NAND3_X1 _16641_ ( .A1(_00661_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00814_ ) );
NAND3_X1 _16642_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00815_ ) );
AND2_X1 _16643_ ( .A1(_00814_ ), .A2(_00815_ ), .ZN(_00816_ ) );
NAND3_X1 _16644_ ( .A1(_00672_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00817_ ) );
NAND3_X1 _16645_ ( .A1(_06043_ ), .A2(_06046_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00818_ ) );
NAND4_X1 _16646_ ( .A1(_00816_ ), .A2(_00667_ ), .A3(_00817_ ), .A4(_00818_ ), .ZN(_00819_ ) );
AND3_X1 _16647_ ( .A1(_00813_ ), .A2(_00659_ ), .A3(_00819_ ), .ZN(_00820_ ) );
OR2_X1 _16648_ ( .A1(_00808_ ), .A2(_00820_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
AOI21_X1 _16649_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00821_ ) );
OAI21_X1 _16650_ ( .A(_00704_ ), .B1(_06090_ ), .B2(_00534_ ), .ZN(_00822_ ) );
NAND2_X1 _16651_ ( .A1(_00821_ ), .A2(_00822_ ), .ZN(_00823_ ) );
AND3_X1 _16652_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00824_ ) );
AND3_X1 _16653_ ( .A1(_00643_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00825_ ) );
AOI211_X1 _16654_ ( .A(_00824_ ), .B(_00825_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_06040_ ), .ZN(_00826_ ) );
NAND3_X1 _16655_ ( .A1(_06048_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00827_ ) );
NAND4_X1 _16656_ ( .A1(_00826_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_00827_ ), .ZN(_00828_ ) );
NAND3_X1 _16657_ ( .A1(_00749_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00829_ ) );
NAND3_X1 _16658_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00830_ ) );
AND2_X1 _16659_ ( .A1(_00829_ ), .A2(_00830_ ), .ZN(_00831_ ) );
NAND3_X1 _16660_ ( .A1(_00755_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00832_ ) );
NAND3_X1 _16661_ ( .A1(_06044_ ), .A2(_00757_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00833_ ) );
NAND4_X1 _16662_ ( .A1(_00831_ ), .A2(_00753_ ), .A3(_00832_ ), .A4(_00833_ ), .ZN(_00834_ ) );
NAND3_X1 _16663_ ( .A1(_00828_ ), .A2(_00660_ ), .A3(_00834_ ), .ZN(_00835_ ) );
NAND2_X1 _16664_ ( .A1(_00823_ ), .A2(_00835_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
AOI21_X1 _16665_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00836_ ) );
OAI21_X1 _16666_ ( .A(_00704_ ), .B1(_06082_ ), .B2(_00537_ ), .ZN(_00837_ ) );
NAND2_X1 _16667_ ( .A1(_00836_ ), .A2(_00837_ ), .ZN(_00838_ ) );
AND3_X1 _16668_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00839_ ) );
AND3_X1 _16669_ ( .A1(_00643_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00840_ ) );
AOI211_X1 _16670_ ( .A(_00839_ ), .B(_00840_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_06040_ ), .ZN(_00841_ ) );
NAND3_X1 _16671_ ( .A1(_06048_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00842_ ) );
NAND4_X1 _16672_ ( .A1(_00841_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_00842_ ), .ZN(_00843_ ) );
NAND3_X1 _16673_ ( .A1(_00749_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00844_ ) );
NAND3_X1 _16674_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00845_ ) );
AND2_X1 _16675_ ( .A1(_00844_ ), .A2(_00845_ ), .ZN(_00846_ ) );
NAND3_X1 _16676_ ( .A1(_00755_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00847_ ) );
NAND3_X1 _16677_ ( .A1(_06044_ ), .A2(_00757_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00848_ ) );
NAND4_X1 _16678_ ( .A1(_00846_ ), .A2(_00753_ ), .A3(_00847_ ), .A4(_00848_ ), .ZN(_00849_ ) );
NAND3_X1 _16679_ ( .A1(_00843_ ), .A2(_00660_ ), .A3(_00849_ ), .ZN(_00850_ ) );
NAND2_X1 _16680_ ( .A1(_00838_ ), .A2(_00850_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
NOR3_X1 _16681_ ( .A1(\myifu.data_in [13] ), .A2(_00685_ ), .A3(_00687_ ), .ZN(_00851_ ) );
AOI211_X1 _16682_ ( .A(_00761_ ), .B(_00851_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_00852_ ) );
AND3_X1 _16683_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00853_ ) );
AND3_X1 _16684_ ( .A1(_06042_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00854_ ) );
AOI211_X1 _16685_ ( .A(_00853_ ), .B(_00854_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_06039_ ), .ZN(_00855_ ) );
NAND3_X1 _16686_ ( .A1(_00654_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00856_ ) );
NAND4_X1 _16687_ ( .A1(_00855_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_00856_ ), .ZN(_00857_ ) );
NAND3_X1 _16688_ ( .A1(_06042_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00858_ ) );
NAND3_X1 _16689_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00859_ ) );
AND2_X1 _16690_ ( .A1(_00858_ ), .A2(_00859_ ), .ZN(_00860_ ) );
NAND3_X1 _16691_ ( .A1(_00672_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_00861_ ) );
NAND3_X1 _16692_ ( .A1(_06043_ ), .A2(_06046_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_00862_ ) );
NAND4_X1 _16693_ ( .A1(_00860_ ), .A2(_00667_ ), .A3(_00861_ ), .A4(_00862_ ), .ZN(_00863_ ) );
AND3_X1 _16694_ ( .A1(_00857_ ), .A2(_00659_ ), .A3(_00863_ ), .ZN(_00864_ ) );
OR2_X1 _16695_ ( .A1(_00852_ ), .A2(_00864_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
AOI21_X1 _16696_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00865_ ) );
OAI21_X1 _16697_ ( .A(_00704_ ), .B1(_06082_ ), .B2(_00544_ ), .ZN(_00866_ ) );
NAND2_X1 _16698_ ( .A1(_00865_ ), .A2(_00866_ ), .ZN(_00867_ ) );
AND3_X1 _16699_ ( .A1(fanout_net_12 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_00868_ ) );
AND3_X1 _16700_ ( .A1(_00643_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_00869_ ) );
AOI211_X1 _16701_ ( .A(_00868_ ), .B(_00869_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_06040_ ), .ZN(_00870_ ) );
NAND3_X1 _16702_ ( .A1(_06048_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_00871_ ) );
NAND4_X1 _16703_ ( .A1(_00870_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_00871_ ), .ZN(_00872_ ) );
NAND3_X1 _16704_ ( .A1(_00749_ ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_00873_ ) );
NAND3_X1 _16705_ ( .A1(fanout_net_13 ), .A2(fanout_net_8 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_00874_ ) );
AND2_X1 _16706_ ( .A1(_00873_ ), .A2(_00874_ ), .ZN(_00875_ ) );
NAND3_X1 _16707_ ( .A1(_00755_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_00876_ ) );
NAND3_X1 _16708_ ( .A1(_06044_ ), .A2(_00757_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_00877_ ) );
NAND4_X1 _16709_ ( .A1(_00875_ ), .A2(_00668_ ), .A3(_00876_ ), .A4(_00877_ ), .ZN(_00878_ ) );
NAND3_X1 _16710_ ( .A1(_00872_ ), .A2(_00660_ ), .A3(_00878_ ), .ZN(_00879_ ) );
NAND2_X1 _16711_ ( .A1(_00867_ ), .A2(_00879_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
AND3_X1 _16712_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_00880_ ) );
AND3_X1 _16713_ ( .A1(_00707_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_00881_ ) );
AOI211_X1 _16714_ ( .A(_00880_ ), .B(_00881_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_00646_ ), .ZN(_00882_ ) );
NAND3_X1 _16715_ ( .A1(_00655_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_00883_ ) );
NAND4_X1 _16716_ ( .A1(_00882_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00883_ ), .ZN(_00884_ ) );
NAND3_X1 _16717_ ( .A1(_00662_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_00885_ ) );
NAND3_X1 _16718_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_00886_ ) );
AND2_X1 _16719_ ( .A1(_00885_ ), .A2(_00886_ ), .ZN(_00887_ ) );
NAND3_X1 _16720_ ( .A1(_00669_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_00888_ ) );
NAND3_X1 _16721_ ( .A1(_00671_ ), .A2(_00673_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_00889_ ) );
NAND4_X1 _16722_ ( .A1(_00887_ ), .A2(_00668_ ), .A3(_00888_ ), .A4(_00889_ ), .ZN(_00890_ ) );
NAND3_X1 _16723_ ( .A1(_00884_ ), .A2(_00695_ ), .A3(_00890_ ), .ZN(_00891_ ) );
OAI21_X1 _16724_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03506_ ), .ZN(_00892_ ) );
NOR3_X1 _16725_ ( .A1(_00686_ ), .A2(\myifu.data_in [29] ), .A3(_00688_ ), .ZN(_00893_ ) );
OAI21_X1 _16726_ ( .A(_00891_ ), .B1(_00892_ ), .B2(_00893_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16727_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_00894_ ) );
AND3_X1 _16728_ ( .A1(_00707_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_00895_ ) );
AOI211_X1 _16729_ ( .A(_00894_ ), .B(_00895_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_00646_ ), .ZN(_00896_ ) );
NAND3_X1 _16730_ ( .A1(_00655_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_00897_ ) );
NAND4_X1 _16731_ ( .A1(_00896_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00897_ ), .ZN(_00898_ ) );
NAND3_X1 _16732_ ( .A1(_00662_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_00899_ ) );
NAND3_X1 _16733_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_00900_ ) );
AND2_X1 _16734_ ( .A1(_00899_ ), .A2(_00900_ ), .ZN(_00901_ ) );
NAND3_X1 _16735_ ( .A1(_00669_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_00902_ ) );
NAND3_X1 _16736_ ( .A1(_00671_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_00903_ ) );
NAND4_X1 _16737_ ( .A1(_00901_ ), .A2(_00782_ ), .A3(_00902_ ), .A4(_00903_ ), .ZN(_00904_ ) );
NAND3_X1 _16738_ ( .A1(_00898_ ), .A2(_00695_ ), .A3(_00904_ ), .ZN(_00905_ ) );
OAI21_X1 _16739_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03555_ ), .ZN(_00906_ ) );
NOR3_X1 _16740_ ( .A1(\myifu.data_in [11] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_00907_ ) );
OAI21_X1 _16741_ ( .A(_00905_ ), .B1(_00906_ ), .B2(_00907_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
AND3_X1 _16742_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_00908_ ) );
AND3_X1 _16743_ ( .A1(_00707_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_00909_ ) );
AOI211_X1 _16744_ ( .A(_00908_ ), .B(_00909_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_00646_ ), .ZN(_00910_ ) );
NAND3_X1 _16745_ ( .A1(_00655_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_00911_ ) );
NAND4_X1 _16746_ ( .A1(_00910_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00911_ ), .ZN(_00912_ ) );
NAND3_X1 _16747_ ( .A1(_00662_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_00913_ ) );
NAND3_X1 _16748_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_00914_ ) );
AND2_X1 _16749_ ( .A1(_00913_ ), .A2(_00914_ ), .ZN(_00915_ ) );
NAND3_X1 _16750_ ( .A1(_00669_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_00916_ ) );
NAND3_X1 _16751_ ( .A1(_00671_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_00917_ ) );
NAND4_X1 _16752_ ( .A1(_00915_ ), .A2(_00782_ ), .A3(_00916_ ), .A4(_00917_ ), .ZN(_00918_ ) );
NAND3_X1 _16753_ ( .A1(_00912_ ), .A2(_00695_ ), .A3(_00918_ ), .ZN(_00919_ ) );
OAI21_X1 _16754_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03548_ ), .ZN(_00920_ ) );
NOR3_X1 _16755_ ( .A1(\myifu.data_in [10] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_00921_ ) );
OAI21_X1 _16756_ ( .A(_00919_ ), .B1(_00920_ ), .B2(_00921_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
AND3_X1 _16757_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_00922_ ) );
AND3_X1 _16758_ ( .A1(_00707_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_00923_ ) );
AOI211_X1 _16759_ ( .A(_00922_ ), .B(_00923_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_00646_ ), .ZN(_00924_ ) );
NAND3_X1 _16760_ ( .A1(_00655_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_00925_ ) );
NAND4_X1 _16761_ ( .A1(_00924_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00925_ ), .ZN(_00926_ ) );
NAND3_X1 _16762_ ( .A1(_00784_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_00927_ ) );
NAND3_X1 _16763_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_00928_ ) );
AND2_X1 _16764_ ( .A1(_00927_ ), .A2(_00928_ ), .ZN(_00929_ ) );
NAND3_X1 _16765_ ( .A1(_00673_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_00930_ ) );
NAND3_X1 _16766_ ( .A1(_00671_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_00931_ ) );
NAND4_X1 _16767_ ( .A1(_00929_ ), .A2(_00782_ ), .A3(_00930_ ), .A4(_00931_ ), .ZN(_00932_ ) );
NAND3_X1 _16768_ ( .A1(_00926_ ), .A2(_00695_ ), .A3(_00932_ ), .ZN(_00933_ ) );
OAI21_X1 _16769_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03535_ ), .ZN(_00934_ ) );
NOR3_X1 _16770_ ( .A1(\myifu.data_in [9] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_00935_ ) );
OAI21_X1 _16771_ ( .A(_00933_ ), .B1(_00934_ ), .B2(_00935_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
NOR3_X1 _16772_ ( .A1(\myifu.data_in [7] ), .A2(_00677_ ), .A3(_00687_ ), .ZN(_00936_ ) );
AOI211_X1 _16773_ ( .A(_00761_ ), .B(_00936_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_00763_ ), .ZN(_00937_ ) );
AND3_X1 _16774_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_00938_ ) );
AND3_X1 _16775_ ( .A1(_06041_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_00939_ ) );
AOI211_X1 _16776_ ( .A(_00938_ ), .B(_00939_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_06039_ ), .ZN(_00940_ ) );
NAND3_X1 _16777_ ( .A1(_00654_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_00941_ ) );
NAND4_X1 _16778_ ( .A1(_00940_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_00941_ ), .ZN(_00942_ ) );
NAND3_X1 _16779_ ( .A1(_06042_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_00943_ ) );
NAND3_X1 _16780_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_00944_ ) );
AND2_X1 _16781_ ( .A1(_00943_ ), .A2(_00944_ ), .ZN(_00945_ ) );
NAND3_X1 _16782_ ( .A1(_00672_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_00946_ ) );
NAND3_X1 _16783_ ( .A1(_06043_ ), .A2(_06046_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_00947_ ) );
NAND4_X1 _16784_ ( .A1(_00945_ ), .A2(_00667_ ), .A3(_00946_ ), .A4(_00947_ ), .ZN(_00948_ ) );
AND3_X1 _16785_ ( .A1(_00942_ ), .A2(_00659_ ), .A3(_00948_ ), .ZN(_00949_ ) );
OR2_X1 _16786_ ( .A1(_00937_ ), .A2(_00949_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AND3_X1 _16787_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_00950_ ) );
AND3_X1 _16788_ ( .A1(_00707_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_00951_ ) );
AOI211_X1 _16789_ ( .A(_00950_ ), .B(_00951_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00645_ ), .ZN(_00952_ ) );
NAND3_X1 _16790_ ( .A1(_00757_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_00953_ ) );
NAND4_X1 _16791_ ( .A1(_00952_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_00953_ ), .ZN(_00954_ ) );
NAND3_X1 _16792_ ( .A1(_00784_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_00955_ ) );
NAND3_X1 _16793_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_00956_ ) );
AND2_X1 _16794_ ( .A1(_00955_ ), .A2(_00956_ ), .ZN(_00957_ ) );
NAND3_X1 _16795_ ( .A1(_00673_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_00958_ ) );
NAND3_X1 _16796_ ( .A1(_00749_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_00959_ ) );
NAND4_X1 _16797_ ( .A1(_00957_ ), .A2(_00782_ ), .A3(_00958_ ), .A4(_00959_ ), .ZN(_00960_ ) );
NAND3_X1 _16798_ ( .A1(_00954_ ), .A2(_00695_ ), .A3(_00960_ ), .ZN(_00961_ ) );
OAI21_X1 _16799_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03158_ ), .ZN(_00962_ ) );
NOR3_X1 _16800_ ( .A1(\myifu.data_in [6] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_00963_ ) );
OAI21_X1 _16801_ ( .A(_00961_ ), .B1(_00962_ ), .B2(_00963_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
AOI21_X1 _16802_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00964_ ) );
OAI21_X1 _16803_ ( .A(_00704_ ), .B1(_06082_ ), .B2(_00569_ ), .ZN(_00965_ ) );
NAND2_X1 _16804_ ( .A1(_00964_ ), .A2(_00965_ ), .ZN(_00966_ ) );
AND3_X1 _16805_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_00967_ ) );
AND3_X1 _16806_ ( .A1(_00643_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_00968_ ) );
AOI211_X1 _16807_ ( .A(_00967_ ), .B(_00968_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_06040_ ), .ZN(_00969_ ) );
NAND3_X1 _16808_ ( .A1(_06048_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_00970_ ) );
NAND4_X1 _16809_ ( .A1(_00969_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_00970_ ), .ZN(_00971_ ) );
NAND3_X1 _16810_ ( .A1(_00749_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_00972_ ) );
NAND3_X1 _16811_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_00973_ ) );
AND2_X1 _16812_ ( .A1(_00972_ ), .A2(_00973_ ), .ZN(_00974_ ) );
NAND3_X1 _16813_ ( .A1(_00755_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_00975_ ) );
NAND3_X1 _16814_ ( .A1(_06044_ ), .A2(_00757_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_00976_ ) );
NAND4_X1 _16815_ ( .A1(_00974_ ), .A2(_00668_ ), .A3(_00975_ ), .A4(_00976_ ), .ZN(_00977_ ) );
NAND3_X1 _16816_ ( .A1(_00971_ ), .A2(_00660_ ), .A3(_00977_ ), .ZN(_00978_ ) );
NAND2_X1 _16817_ ( .A1(_00966_ ), .A2(_00978_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
AOI21_X1 _16818_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00979_ ) );
OAI21_X1 _16819_ ( .A(_00704_ ), .B1(_06082_ ), .B2(_00572_ ), .ZN(_00980_ ) );
NAND2_X1 _16820_ ( .A1(_00979_ ), .A2(_00980_ ), .ZN(_00981_ ) );
AND3_X1 _16821_ ( .A1(fanout_net_14 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_00982_ ) );
AND3_X1 _16822_ ( .A1(_00643_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_00983_ ) );
AOI211_X1 _16823_ ( .A(_00982_ ), .B(_00983_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_06040_ ), .ZN(_00984_ ) );
NAND3_X1 _16824_ ( .A1(_00755_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_00985_ ) );
NAND4_X1 _16825_ ( .A1(_00984_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_00985_ ), .ZN(_00986_ ) );
NAND3_X1 _16826_ ( .A1(_00662_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_00987_ ) );
NAND3_X1 _16827_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_00988_ ) );
AND2_X1 _16828_ ( .A1(_00987_ ), .A2(_00988_ ), .ZN(_00989_ ) );
NAND3_X1 _16829_ ( .A1(_00755_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_00990_ ) );
NAND3_X1 _16830_ ( .A1(_06044_ ), .A2(_00669_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_00991_ ) );
NAND4_X1 _16831_ ( .A1(_00989_ ), .A2(_00668_ ), .A3(_00990_ ), .A4(_00991_ ), .ZN(_00992_ ) );
NAND3_X1 _16832_ ( .A1(_00986_ ), .A2(_00660_ ), .A3(_00992_ ), .ZN(_00993_ ) );
NAND2_X1 _16833_ ( .A1(_00981_ ), .A2(_00993_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _16834_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00994_ ) );
OAI21_X1 _16835_ ( .A(_00704_ ), .B1(_06082_ ), .B2(_00575_ ), .ZN(_00995_ ) );
NAND2_X1 _16836_ ( .A1(_00994_ ), .A2(_00995_ ), .ZN(_00996_ ) );
AND3_X1 _16837_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_00997_ ) );
AND3_X1 _16838_ ( .A1(_00643_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_00998_ ) );
AOI211_X1 _16839_ ( .A(_00997_ ), .B(_00998_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00646_ ), .ZN(_00999_ ) );
NAND3_X1 _16840_ ( .A1(_00755_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_01000_ ) );
NAND4_X1 _16841_ ( .A1(_00999_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_01000_ ), .ZN(_01001_ ) );
NAND3_X1 _16842_ ( .A1(_00662_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_01002_ ) );
NAND3_X1 _16843_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_01003_ ) );
AND2_X1 _16844_ ( .A1(_01002_ ), .A2(_01003_ ), .ZN(_01004_ ) );
NAND3_X1 _16845_ ( .A1(_00655_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_01005_ ) );
NAND3_X1 _16846_ ( .A1(_00671_ ), .A2(_00669_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_01006_ ) );
NAND4_X1 _16847_ ( .A1(_01004_ ), .A2(_00668_ ), .A3(_01005_ ), .A4(_01006_ ), .ZN(_01007_ ) );
NAND3_X1 _16848_ ( .A1(_01001_ ), .A2(_00660_ ), .A3(_01007_ ), .ZN(_01008_ ) );
NAND2_X1 _16849_ ( .A1(_00996_ ), .A2(_01008_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
AOI21_X1 _16850_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01009_ ) );
OAI21_X1 _16851_ ( .A(_00704_ ), .B1(_06082_ ), .B2(_00578_ ), .ZN(_01010_ ) );
NAND2_X1 _16852_ ( .A1(_01009_ ), .A2(_01010_ ), .ZN(_01011_ ) );
AND3_X1 _16853_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_01012_ ) );
AND3_X1 _16854_ ( .A1(_00643_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_01013_ ) );
AOI211_X1 _16855_ ( .A(_01012_ ), .B(_01013_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_00646_ ), .ZN(_01014_ ) );
NAND3_X1 _16856_ ( .A1(_00755_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_01015_ ) );
NAND4_X1 _16857_ ( .A1(_01014_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_01015_ ), .ZN(_01016_ ) );
NAND3_X1 _16858_ ( .A1(_00662_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_01017_ ) );
NAND3_X1 _16859_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_01018_ ) );
AND2_X1 _16860_ ( .A1(_01017_ ), .A2(_01018_ ), .ZN(_01019_ ) );
NAND3_X1 _16861_ ( .A1(_00655_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_01020_ ) );
NAND3_X1 _16862_ ( .A1(_00671_ ), .A2(_00669_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_01021_ ) );
NAND4_X1 _16863_ ( .A1(_01019_ ), .A2(_00668_ ), .A3(_01020_ ), .A4(_01021_ ), .ZN(_01022_ ) );
NAND3_X1 _16864_ ( .A1(_01016_ ), .A2(_00660_ ), .A3(_01022_ ), .ZN(_01023_ ) );
NAND2_X1 _16865_ ( .A1(_01011_ ), .A2(_01023_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
AOI21_X1 _16866_ ( .A(_00722_ ), .B1(_00725_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01024_ ) );
OAI21_X1 _16867_ ( .A(_00682_ ), .B1(_06082_ ), .B2(_00584_ ), .ZN(_01025_ ) );
NAND2_X1 _16868_ ( .A1(_01024_ ), .A2(_01025_ ), .ZN(_01026_ ) );
AND3_X1 _16869_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01027_ ) );
AND3_X1 _16870_ ( .A1(_00643_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01028_ ) );
AOI211_X1 _16871_ ( .A(_01027_ ), .B(_01028_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_00646_ ), .ZN(_01029_ ) );
NAND3_X1 _16872_ ( .A1(_00755_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01030_ ) );
NAND4_X1 _16873_ ( .A1(_01029_ ), .A2(_00745_ ), .A3(_00746_ ), .A4(_01030_ ), .ZN(_01031_ ) );
NAND3_X1 _16874_ ( .A1(_00662_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01032_ ) );
NAND3_X1 _16875_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01033_ ) );
AND2_X1 _16876_ ( .A1(_01032_ ), .A2(_01033_ ), .ZN(_01034_ ) );
NAND3_X1 _16877_ ( .A1(_00655_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01035_ ) );
NAND3_X1 _16878_ ( .A1(_00671_ ), .A2(_00669_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01036_ ) );
NAND4_X1 _16879_ ( .A1(_01034_ ), .A2(_00668_ ), .A3(_01035_ ), .A4(_01036_ ), .ZN(_01037_ ) );
NAND3_X1 _16880_ ( .A1(_01031_ ), .A2(_00660_ ), .A3(_01037_ ), .ZN(_01038_ ) );
NAND2_X1 _16881_ ( .A1(_01026_ ), .A2(_01038_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
AND3_X1 _16882_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01039_ ) );
AND3_X1 _16883_ ( .A1(_00707_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01040_ ) );
AOI211_X1 _16884_ ( .A(_01039_ ), .B(_01040_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00645_ ), .ZN(_01041_ ) );
NAND3_X1 _16885_ ( .A1(_00757_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01042_ ) );
NAND4_X1 _16886_ ( .A1(_01041_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_01042_ ), .ZN(_01043_ ) );
NAND3_X1 _16887_ ( .A1(_00784_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01044_ ) );
NAND3_X1 _16888_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01045_ ) );
AND2_X1 _16889_ ( .A1(_01044_ ), .A2(_01045_ ), .ZN(_01046_ ) );
NAND3_X1 _16890_ ( .A1(_00673_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01047_ ) );
NAND3_X1 _16891_ ( .A1(_00749_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01048_ ) );
NAND4_X1 _16892_ ( .A1(_01046_ ), .A2(_00782_ ), .A3(_01047_ ), .A4(_01048_ ), .ZN(_01049_ ) );
NAND3_X1 _16893_ ( .A1(_01043_ ), .A2(_00695_ ), .A3(_01049_ ), .ZN(_01050_ ) );
OAI21_X1 _16894_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03516_ ), .ZN(_01051_ ) );
NOR3_X1 _16895_ ( .A1(\myifu.data_in [28] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_01052_ ) );
OAI21_X1 _16896_ ( .A(_01050_ ), .B1(_01051_ ), .B2(_01052_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
NOR3_X1 _16897_ ( .A1(\myifu.data_in [0] ), .A2(_00677_ ), .A3(_00681_ ), .ZN(_01053_ ) );
AOI211_X1 _16898_ ( .A(_00761_ ), .B(_01053_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_01054_ ) );
NAND3_X1 _16899_ ( .A1(_00661_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01055_ ) );
NAND3_X1 _16900_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01056_ ) );
AND2_X1 _16901_ ( .A1(_01055_ ), .A2(_01056_ ), .ZN(_01057_ ) );
NAND3_X1 _16902_ ( .A1(_00654_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01058_ ) );
NAND3_X1 _16903_ ( .A1(_00784_ ), .A2(_06047_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01059_ ) );
NAND4_X1 _16904_ ( .A1(_01057_ ), .A2(_00782_ ), .A3(_01058_ ), .A4(_01059_ ), .ZN(_01060_ ) );
AND3_X1 _16905_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01061_ ) );
AND3_X1 _16906_ ( .A1(_06041_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01062_ ) );
AOI211_X1 _16907_ ( .A(_01061_ ), .B(_01062_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_06039_ ), .ZN(_01063_ ) );
NAND3_X1 _16908_ ( .A1(_00672_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01064_ ) );
NAND4_X1 _16909_ ( .A1(_01063_ ), .A2(_00648_ ), .A3(_00651_ ), .A4(_01064_ ), .ZN(_01065_ ) );
AND3_X1 _16910_ ( .A1(_01060_ ), .A2(_00658_ ), .A3(_01065_ ), .ZN(_01066_ ) );
OR2_X1 _16911_ ( .A1(_01054_ ), .A2(_01066_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
AND3_X1 _16912_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01067_ ) );
AND3_X1 _16913_ ( .A1(_00707_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01068_ ) );
AOI211_X1 _16914_ ( .A(_01067_ ), .B(_01068_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00645_ ), .ZN(_01069_ ) );
NAND3_X1 _16915_ ( .A1(_00757_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01070_ ) );
NAND4_X1 _16916_ ( .A1(_01069_ ), .A2(_00650_ ), .A3(_00653_ ), .A4(_01070_ ), .ZN(_01071_ ) );
NAND3_X1 _16917_ ( .A1(_00784_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01072_ ) );
NAND3_X1 _16918_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01073_ ) );
AND2_X1 _16919_ ( .A1(_01072_ ), .A2(_01073_ ), .ZN(_01074_ ) );
NAND3_X1 _16920_ ( .A1(_00673_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01075_ ) );
NAND3_X1 _16921_ ( .A1(_00749_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01076_ ) );
NAND4_X1 _16922_ ( .A1(_01074_ ), .A2(_00782_ ), .A3(_01075_ ), .A4(_01076_ ), .ZN(_01077_ ) );
NAND3_X1 _16923_ ( .A1(_01071_ ), .A2(_00695_ ), .A3(_01077_ ), .ZN(_01078_ ) );
OAI21_X1 _16924_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03520_ ), .ZN(_01079_ ) );
NOR3_X1 _16925_ ( .A1(\myifu.data_in [27] ), .A2(_00686_ ), .A3(_00688_ ), .ZN(_01080_ ) );
OAI21_X1 _16926_ ( .A(_01078_ ), .B1(_01079_ ), .B2(_01080_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
AND3_X1 _16927_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01081_ ) );
AND3_X1 _16928_ ( .A1(_00707_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01082_ ) );
AOI211_X1 _16929_ ( .A(_01081_ ), .B(_01082_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_00645_ ), .ZN(_01083_ ) );
NAND3_X1 _16930_ ( .A1(_00757_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01084_ ) );
NAND4_X1 _16931_ ( .A1(_01083_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_01084_ ), .ZN(_01085_ ) );
NAND3_X1 _16932_ ( .A1(_00784_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01086_ ) );
NAND3_X1 _16933_ ( .A1(\IF_ID_pc [4] ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01087_ ) );
AND2_X1 _16934_ ( .A1(_01086_ ), .A2(_01087_ ), .ZN(_01088_ ) );
NAND3_X1 _16935_ ( .A1(_00673_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01089_ ) );
NAND3_X1 _16936_ ( .A1(_00749_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01090_ ) );
NAND4_X1 _16937_ ( .A1(_01088_ ), .A2(_00782_ ), .A3(_01089_ ), .A4(_01090_ ), .ZN(_01091_ ) );
NAND3_X1 _16938_ ( .A1(_01085_ ), .A2(_00695_ ), .A3(_01091_ ), .ZN(_01092_ ) );
OAI21_X1 _16939_ ( .A(\myifu.state [2] ), .B1(_00683_ ), .B2(_03530_ ), .ZN(_01093_ ) );
NOR3_X1 _16940_ ( .A1(_00686_ ), .A2(\myifu.data_in [26] ), .A3(_00688_ ), .ZN(_01094_ ) );
OAI21_X1 _16941_ ( .A(_01092_ ), .B1(_01093_ ), .B2(_01094_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
AND3_X1 _16942_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01095_ ) );
AND3_X1 _16943_ ( .A1(_00707_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01096_ ) );
AOI211_X1 _16944_ ( .A(_01095_ ), .B(_01096_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00645_ ), .ZN(_01097_ ) );
NAND3_X1 _16945_ ( .A1(_00757_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01098_ ) );
NAND4_X1 _16946_ ( .A1(_01097_ ), .A2(_00649_ ), .A3(_00652_ ), .A4(_01098_ ), .ZN(_01099_ ) );
NAND3_X1 _16947_ ( .A1(_00784_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01100_ ) );
NAND3_X1 _16948_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01101_ ) );
AND2_X1 _16949_ ( .A1(_01100_ ), .A2(_01101_ ), .ZN(_01102_ ) );
NAND3_X1 _16950_ ( .A1(_00673_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01103_ ) );
NAND3_X1 _16951_ ( .A1(_00749_ ), .A2(_00754_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01104_ ) );
NAND4_X1 _16952_ ( .A1(_01102_ ), .A2(_00782_ ), .A3(_01103_ ), .A4(_01104_ ), .ZN(_01105_ ) );
NAND3_X1 _16953_ ( .A1(_01099_ ), .A2(_00659_ ), .A3(_01105_ ), .ZN(_01106_ ) );
OAI21_X1 _16954_ ( .A(\myifu.state [2] ), .B1(_00704_ ), .B2(_03524_ ), .ZN(_01107_ ) );
NOR3_X1 _16955_ ( .A1(\myifu.data_in [25] ), .A2(_00685_ ), .A3(_00687_ ), .ZN(_01108_ ) );
OAI21_X1 _16956_ ( .A(_01106_ ), .B1(_01107_ ), .B2(_01108_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
NOR3_X1 _16957_ ( .A1(_00685_ ), .A2(\myifu.data_in [24] ), .A3(_00681_ ), .ZN(_01109_ ) );
AOI211_X1 _16958_ ( .A(_00761_ ), .B(_01109_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_01110_ ) );
AND3_X1 _16959_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01111_ ) );
AND3_X1 _16960_ ( .A1(_06041_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01112_ ) );
AOI211_X1 _16961_ ( .A(_01111_ ), .B(_01112_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_06039_ ), .ZN(_01113_ ) );
NAND3_X1 _16962_ ( .A1(_06047_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01114_ ) );
NAND4_X1 _16963_ ( .A1(_01113_ ), .A2(_00649_ ), .A3(_00651_ ), .A4(_01114_ ), .ZN(_01115_ ) );
NAND3_X1 _16964_ ( .A1(_06042_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01116_ ) );
NAND3_X1 _16965_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01117_ ) );
AND2_X1 _16966_ ( .A1(_01116_ ), .A2(_01117_ ), .ZN(_01118_ ) );
NAND3_X1 _16967_ ( .A1(_00672_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01119_ ) );
NAND3_X1 _16968_ ( .A1(_06043_ ), .A2(_06046_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01120_ ) );
NAND4_X1 _16969_ ( .A1(_01118_ ), .A2(_00667_ ), .A3(_01119_ ), .A4(_01120_ ), .ZN(_01121_ ) );
AND3_X1 _16970_ ( .A1(_01115_ ), .A2(_00658_ ), .A3(_01121_ ), .ZN(_01122_ ) );
OR2_X1 _16971_ ( .A1(_01110_ ), .A2(_01122_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
NOR3_X1 _16972_ ( .A1(\myifu.data_in [23] ), .A2(_00677_ ), .A3(_00681_ ), .ZN(_01123_ ) );
AOI211_X1 _16973_ ( .A(_00761_ ), .B(_01123_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .C2(_00763_ ), .ZN(_01124_ ) );
NAND3_X1 _16974_ ( .A1(_00661_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01125_ ) );
NAND3_X1 _16975_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01126_ ) );
AND2_X1 _16976_ ( .A1(_01125_ ), .A2(_01126_ ), .ZN(_01127_ ) );
NAND3_X1 _16977_ ( .A1(_00654_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01128_ ) );
NAND3_X1 _16978_ ( .A1(_00784_ ), .A2(_06047_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01129_ ) );
NAND4_X1 _16979_ ( .A1(_01127_ ), .A2(_00667_ ), .A3(_01128_ ), .A4(_01129_ ), .ZN(_01130_ ) );
AND3_X1 _16980_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01131_ ) );
AND3_X1 _16981_ ( .A1(_06041_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01132_ ) );
AOI211_X1 _16982_ ( .A(_01131_ ), .B(_01132_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_06039_ ), .ZN(_01133_ ) );
NAND3_X1 _16983_ ( .A1(_00672_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01134_ ) );
NAND4_X1 _16984_ ( .A1(_01133_ ), .A2(_00648_ ), .A3(_00651_ ), .A4(_01134_ ), .ZN(_01135_ ) );
AND3_X1 _16985_ ( .A1(_01130_ ), .A2(_00658_ ), .A3(_01135_ ), .ZN(_01136_ ) );
OR2_X1 _16986_ ( .A1(_01124_ ), .A2(_01136_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
NOR3_X1 _16987_ ( .A1(\myifu.data_in [22] ), .A2(_00677_ ), .A3(_00681_ ), .ZN(_01137_ ) );
AOI211_X1 _16988_ ( .A(_00761_ ), .B(_01137_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .C2(_00763_ ), .ZN(_01138_ ) );
NAND3_X1 _16989_ ( .A1(_00661_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01139_ ) );
NAND3_X1 _16990_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01140_ ) );
AND2_X1 _16991_ ( .A1(_01139_ ), .A2(_01140_ ), .ZN(_01141_ ) );
NAND3_X1 _16992_ ( .A1(_00654_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01142_ ) );
NAND3_X1 _16993_ ( .A1(_00784_ ), .A2(_06047_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01143_ ) );
NAND4_X1 _16994_ ( .A1(_01141_ ), .A2(_00667_ ), .A3(_01142_ ), .A4(_01143_ ), .ZN(_01144_ ) );
AND3_X1 _16995_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01145_ ) );
AND3_X1 _16996_ ( .A1(_06041_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01146_ ) );
AOI211_X1 _16997_ ( .A(_01145_ ), .B(_01146_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_06039_ ), .ZN(_01147_ ) );
NAND3_X1 _16998_ ( .A1(_00672_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01148_ ) );
NAND4_X1 _16999_ ( .A1(_01147_ ), .A2(_00648_ ), .A3(_00651_ ), .A4(_01148_ ), .ZN(_01149_ ) );
AND3_X1 _17000_ ( .A1(_01144_ ), .A2(_00658_ ), .A3(_01149_ ), .ZN(_01150_ ) );
OR2_X1 _17001_ ( .A1(_01138_ ), .A2(_01150_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI211_X1 _17002_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_03228_ ), .C1(_03643_ ), .C2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17003_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01151_ ) );
AND4_X1 _17004_ ( .A1(_01151_ ), .A2(_01883_ ), .A3(\myifu.state [0] ), .A4(_01960_ ), .ZN(_01152_ ) );
AND3_X1 _17005_ ( .A1(_03816_ ), .A2(\myifu.state [2] ), .A3(_03825_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
AOI211_X1 _17006_ ( .A(_00501_ ), .B(_01152_ ), .C1(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .C2(_03822_ ), .ZN(_01153_ ) );
NOR2_X1 _17007_ ( .A1(_01153_ ), .A2(reset ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _17008_ ( .A1(_06027_ ), .A2(_01982_ ), .ZN(_01154_ ) );
INV_X1 _17009_ ( .A(_01154_ ), .ZN(_01155_ ) );
AND3_X1 _17010_ ( .A1(_01155_ ), .A2(_01151_ ), .A3(_01962_ ), .ZN(_01156_ ) );
AND2_X1 _17011_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01157_ ) );
OR4_X1 _17012_ ( .A1(reset ), .A2(_01156_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A4(_01157_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _17013_ ( .A1(_03826_ ), .A2(_01631_ ), .A3(\myifu.state [2] ), .ZN(_01158_ ) );
NAND2_X1 _17014_ ( .A1(_01154_ ), .A2(_02083_ ), .ZN(_01159_ ) );
NAND2_X1 _17015_ ( .A1(_01158_ ), .A2(_01159_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
INV_X1 _17016_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01160_ ) );
NOR3_X1 _17017_ ( .A1(_01160_ ), .A2(_00609_ ), .A3(_00753_ ), .ZN(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ) );
NOR3_X1 _17018_ ( .A1(_01160_ ), .A2(_00610_ ), .A3(_00753_ ), .ZN(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ) );
AND4_X1 _17019_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00753_ ), .ZN(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ) );
AND4_X1 _17020_ ( .A1(\IF_ID_pc [4] ), .A2(_06038_ ), .A3(_06048_ ), .A4(_00753_ ), .ZN(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ) );
NOR3_X1 _17021_ ( .A1(_01160_ ), .A2(_00607_ ), .A3(_00753_ ), .ZN(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ) );
AND4_X1 _17022_ ( .A1(_06044_ ), .A2(_06038_ ), .A3(\IF_ID_pc [3] ), .A4(_00753_ ), .ZN(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _17023_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06040_ ), .A3(_00753_ ), .ZN(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ) );
AND4_X1 _17024_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06040_ ), .A3(_00745_ ), .A4(_00746_ ), .ZN(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ) );
AND3_X1 _17025_ ( .A1(_02071_ ), .A2(_06040_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ) );
AND3_X1 _17026_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06044_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ) );
AND3_X1 _17027_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_06048_ ), .ZN(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ) );
AND3_X1 _17028_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ) );
NAND3_X1 _17029_ ( .A1(_01883_ ), .A2(_01960_ ), .A3(\myifu.state [0] ), .ZN(_01161_ ) );
AND2_X1 _17030_ ( .A1(_00503_ ), .A2(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01162_ ) );
NOR4_X1 _17031_ ( .A1(_01162_ ), .A2(_03229_ ), .A3(_00501_ ), .A4(_01157_ ), .ZN(_01163_ ) );
NAND2_X1 _17032_ ( .A1(_01161_ ), .A2(_01163_ ), .ZN(_01164_ ) );
AOI221_X4 _17033_ ( .A(_01164_ ), .B1(_01155_ ), .B2(\myifu.state [0] ), .C1(_01963_ ), .C2(_03826_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17034_ ( .A1(_03634_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03230_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
AOI211_X1 _17035_ ( .A(_00488_ ), .B(_00490_ ), .C1(_03087_ ), .C2(_03157_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
OR4_X1 _17036_ ( .A1(reset ), .A2(_01162_ ), .A3(_00501_ ), .A4(_01157_ ), .ZN(_01165_ ) );
AOI211_X1 _17037_ ( .A(_03229_ ), .B(_01165_ ), .C1(_01961_ ), .C2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
INV_X2 _17038_ ( .A(\mylsu.state [3] ), .ZN(_01166_ ) );
MUX2_X1 _17039_ ( .A(_01166_ ), .B(_01998_ ), .S(\mylsu.state [0] ), .Z(_01167_ ) );
AOI21_X1 _17040_ ( .A(_01167_ ), .B1(_06143_ ), .B2(\mylsu.state [3] ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ) );
AOI211_X1 _17041_ ( .A(_03890_ ), .B(_01167_ ), .C1(_06143_ ), .C2(\mylsu.state [3] ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
AND2_X1 _17042_ ( .A1(_03884_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
AND2_X1 _17043_ ( .A1(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .A2(_02041_ ), .ZN(_01168_ ) );
AND3_X1 _17044_ ( .A1(_02043_ ), .A2(_02056_ ), .A3(_01168_ ), .ZN(_01169_ ) );
INV_X1 _17045_ ( .A(_01169_ ), .ZN(_01170_ ) );
AOI22_X1 _17046_ ( .A1(_06122_ ), .A2(_06123_ ), .B1(_03812_ ), .B2(_06141_ ), .ZN(_01171_ ) );
AOI21_X1 _17047_ ( .A(_03813_ ), .B1(_06122_ ), .B2(_06123_ ), .ZN(_01172_ ) );
NOR2_X1 _17048_ ( .A1(_01171_ ), .A2(_01172_ ), .ZN(_01173_ ) );
AND3_X1 _17049_ ( .A1(_03825_ ), .A2(_01173_ ), .A3(\io_master_arid [1] ), .ZN(_01174_ ) );
OAI22_X1 _17050_ ( .A1(_06034_ ), .A2(_01170_ ), .B1(_01174_ ), .B2(_06068_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND2_X1 _17051_ ( .A1(_06124_ ), .A2(_03884_ ), .ZN(_01175_ ) );
INV_X1 _17052_ ( .A(io_master_wready ), .ZN(_01176_ ) );
NAND2_X1 _17053_ ( .A1(_06024_ ), .A2(_01176_ ), .ZN(_01177_ ) );
AND4_X1 _17054_ ( .A1(_01999_ ), .A2(_02068_ ), .A3(_01175_ ), .A4(_01177_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
INV_X1 _17055_ ( .A(_02067_ ), .ZN(_01178_ ) );
AND2_X1 _17056_ ( .A1(io_master_awready ), .A2(io_master_wready ), .ZN(_01179_ ) );
NOR2_X1 _17057_ ( .A1(_03841_ ), .A2(_01179_ ), .ZN(_01180_ ) );
AND4_X1 _17058_ ( .A1(io_master_awready ), .A2(_06126_ ), .A3(_03885_ ), .A4(_01180_ ), .ZN(_01181_ ) );
NAND3_X1 _17059_ ( .A1(_06066_ ), .A2(_01178_ ), .A3(_01181_ ), .ZN(_01182_ ) );
NAND3_X1 _17060_ ( .A1(_03885_ ), .A2(\mylsu.state [2] ), .A3(_01176_ ), .ZN(_01183_ ) );
NAND2_X1 _17061_ ( .A1(_01182_ ), .A2(_01183_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
NOR2_X1 _17062_ ( .A1(_03841_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01184_ ) );
AND4_X1 _17063_ ( .A1(\mylsu.state [0] ), .A2(_01175_ ), .A3(_01179_ ), .A4(_01184_ ), .ZN(_01185_ ) );
NAND3_X1 _17064_ ( .A1(_06066_ ), .A2(_01178_ ), .A3(_01185_ ), .ZN(_01186_ ) );
NAND3_X1 _17065_ ( .A1(_03885_ ), .A2(\mylsu.state [4] ), .A3(io_master_awready ), .ZN(_01187_ ) );
AND3_X1 _17066_ ( .A1(_03883_ ), .A2(io_master_wready ), .A3(_03067_ ), .ZN(_01188_ ) );
NAND2_X1 _17067_ ( .A1(_01188_ ), .A2(\mylsu.state [2] ), .ZN(_01189_ ) );
NAND3_X1 _17068_ ( .A1(_06138_ ), .A2(\mylsu.state [1] ), .A3(_03885_ ), .ZN(_01190_ ) );
NAND4_X1 _17069_ ( .A1(_01186_ ), .A2(_01187_ ), .A3(_01189_ ), .A4(_01190_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
NAND4_X1 _17070_ ( .A1(_03825_ ), .A2(_01173_ ), .A3(\io_master_arid [1] ), .A4(_00282_ ), .ZN(_01191_ ) );
OAI21_X1 _17071_ ( .A(_01169_ ), .B1(_06027_ ), .B2(_06032_ ), .ZN(_01192_ ) );
AND4_X1 _17072_ ( .A1(_02041_ ), .A2(_02040_ ), .A3(_02056_ ), .A4(_06036_ ), .ZN(_01193_ ) );
NAND2_X1 _17073_ ( .A1(_01193_ ), .A2(\mylsu.state [0] ), .ZN(_01194_ ) );
AND4_X1 _17074_ ( .A1(_02054_ ), .A2(_02053_ ), .A3(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .A4(_02041_ ), .ZN(_01195_ ) );
INV_X1 _17075_ ( .A(\mylsu.state [0] ), .ZN(_01196_ ) );
NOR4_X1 _17076_ ( .A1(_06037_ ), .A2(_01196_ ), .A3(_03831_ ), .A4(_01177_ ), .ZN(_01197_ ) );
NAND3_X1 _17077_ ( .A1(_01197_ ), .A2(_06066_ ), .A3(_01178_ ), .ZN(_01198_ ) );
AND3_X1 _17078_ ( .A1(_01178_ ), .A2(_06124_ ), .A3(_02040_ ), .ZN(_01199_ ) );
NAND4_X1 _17079_ ( .A1(_01199_ ), .A2(\mylsu.state [0] ), .A3(_01175_ ), .A4(_01184_ ), .ZN(_01200_ ) );
NAND3_X1 _17080_ ( .A1(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .A2(_03831_ ), .A3(_03845_ ), .ZN(_01201_ ) );
NAND3_X1 _17081_ ( .A1(_06135_ ), .A2(\mylsu.state [1] ), .A3(_06137_ ), .ZN(_01202_ ) );
NAND3_X1 _17082_ ( .A1(_03884_ ), .A2(_03841_ ), .A3(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_01203_ ) );
AND4_X1 _17083_ ( .A1(_03884_ ), .A2(_01201_ ), .A3(_01202_ ), .A4(_01203_ ), .ZN(_01204_ ) );
NAND4_X1 _17084_ ( .A1(_02067_ ), .A2(\mylsu.state [0] ), .A3(_01175_ ), .A4(_01184_ ), .ZN(_01205_ ) );
NAND4_X1 _17085_ ( .A1(_01198_ ), .A2(_01200_ ), .A3(_01204_ ), .A4(_01205_ ), .ZN(_01206_ ) );
AOI211_X1 _17086_ ( .A(_01195_ ), .B(_01206_ ), .C1(\mylsu.state [0] ), .C2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01207_ ) );
NAND4_X1 _17087_ ( .A1(_01191_ ), .A2(_01192_ ), .A3(_01194_ ), .A4(_01207_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND3_X1 _17088_ ( .A1(_03885_ ), .A2(\mylsu.state [4] ), .A3(_06024_ ), .ZN(_01208_ ) );
NOR2_X1 _17089_ ( .A1(_06025_ ), .A2(_01196_ ), .ZN(_01209_ ) );
NAND3_X1 _17090_ ( .A1(_01209_ ), .A2(_01184_ ), .A3(_01188_ ), .ZN(_01210_ ) );
OAI21_X1 _17091_ ( .A(_01208_ ), .B1(_02093_ ), .B2(_01210_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
MUX2_X1 _17092_ ( .A(\LS_WB_wdata_csreg [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_03835_ ), .Z(_01211_ ) );
INV_X1 _17093_ ( .A(_03842_ ), .ZN(_01212_ ) );
OR2_X1 _17094_ ( .A1(_03832_ ), .A2(_01212_ ), .ZN(_01213_ ) );
BUF_X4 _17095_ ( .A(_01213_ ), .Z(_01214_ ) );
BUF_X4 _17096_ ( .A(_01214_ ), .Z(_01215_ ) );
MUX2_X1 _17097_ ( .A(_01211_ ), .B(\EX_LS_pc [21] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
OAI22_X1 _17098_ ( .A1(_03835_ ), .A2(_02089_ ), .B1(_02025_ ), .B2(_06163_ ), .ZN(_01216_ ) );
MUX2_X1 _17099_ ( .A(_01216_ ), .B(\EX_LS_pc [20] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _17100_ ( .A(\LS_WB_wdata_csreg [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_03835_ ), .Z(_01217_ ) );
MUX2_X1 _17101_ ( .A(_01217_ ), .B(\EX_LS_pc [19] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
NAND2_X1 _17102_ ( .A1(\EX_LS_flag [2] ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_01218_ ) );
OAI21_X1 _17103_ ( .A(_01218_ ), .B1(_03835_ ), .B2(_02090_ ), .ZN(_01219_ ) );
MUX2_X1 _17104_ ( .A(_01219_ ), .B(\EX_LS_pc [18] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
AOI21_X1 _17105_ ( .A(\EX_LS_pc [17] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01220_ ) );
MUX2_X1 _17106_ ( .A(\LS_WB_wdata_csreg [17] ), .B(\EX_LS_result_csreg_mem [17] ), .S(_02128_ ), .Z(_01221_ ) );
NOR3_X1 _17107_ ( .A1(_03832_ ), .A2(_01212_ ), .A3(_01221_ ), .ZN(_01222_ ) );
NOR2_X1 _17108_ ( .A1(_01220_ ), .A2(_01222_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
BUF_X4 _17109_ ( .A(_02129_ ), .Z(_01223_ ) );
AOI221_X4 _17110_ ( .A(_01214_ ), .B1(\LS_WB_wdata_csreg [16] ), .B2(_01223_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [16] ), .ZN(_01224_ ) );
BUF_X4 _17111_ ( .A(_03833_ ), .Z(_01225_ ) );
BUF_X4 _17112_ ( .A(_03843_ ), .Z(_01226_ ) );
AOI21_X1 _17113_ ( .A(\EX_LS_pc [16] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01227_ ) );
NOR2_X1 _17114_ ( .A1(_01224_ ), .A2(_01227_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _17115_ ( .A(\LS_WB_wdata_csreg [15] ), .B(\EX_LS_result_csreg_mem [15] ), .S(_03835_ ), .Z(_01228_ ) );
MUX2_X1 _17116_ ( .A(_01228_ ), .B(\EX_LS_pc [15] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _17117_ ( .A(\LS_WB_wdata_csreg [14] ), .B(\EX_LS_result_csreg_mem [14] ), .S(_03835_ ), .Z(_01229_ ) );
MUX2_X1 _17118_ ( .A(_01229_ ), .B(\EX_LS_pc [14] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _17119_ ( .A(\LS_WB_wdata_csreg [13] ), .B(\EX_LS_result_csreg_mem [13] ), .S(_03835_ ), .Z(_01230_ ) );
MUX2_X1 _17120_ ( .A(_01230_ ), .B(\EX_LS_pc [13] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
AOI21_X1 _17121_ ( .A(\EX_LS_pc [12] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01231_ ) );
BUF_X4 _17122_ ( .A(_02129_ ), .Z(_01232_ ) );
OAI21_X1 _17123_ ( .A(_03843_ ), .B1(_01232_ ), .B2(_06164_ ), .ZN(_01233_ ) );
AOI221_X4 _17124_ ( .A(_01233_ ), .B1(\LS_WB_wdata_csreg [12] ), .B2(_01232_ ), .C1(_02093_ ), .C2(_06124_ ), .ZN(_01234_ ) );
NOR2_X1 _17125_ ( .A1(_01231_ ), .A2(_01234_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _17126_ ( .A(\EX_LS_pc [30] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01235_ ) );
OAI21_X1 _17127_ ( .A(_03843_ ), .B1(_01232_ ), .B2(_07414_ ), .ZN(_01236_ ) );
AOI221_X4 _17128_ ( .A(_01236_ ), .B1(\LS_WB_wdata_csreg [30] ), .B2(_01232_ ), .C1(_02093_ ), .C2(_06124_ ), .ZN(_01237_ ) );
NOR2_X1 _17129_ ( .A1(_01235_ ), .A2(_01237_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
AOI221_X4 _17130_ ( .A(_01214_ ), .B1(\LS_WB_wdata_csreg [11] ), .B2(_01223_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [11] ), .ZN(_01238_ ) );
AOI21_X1 _17131_ ( .A(\EX_LS_pc [11] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01239_ ) );
NOR2_X1 _17132_ ( .A1(_01238_ ), .A2(_01239_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _17133_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_02128_ ), .Z(_01240_ ) );
MUX2_X1 _17134_ ( .A(_01240_ ), .B(\EX_LS_pc [10] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
AOI221_X4 _17135_ ( .A(_01214_ ), .B1(\LS_WB_wdata_csreg [9] ), .B2(_01223_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [9] ), .ZN(_01241_ ) );
AOI21_X1 _17136_ ( .A(\EX_LS_pc [9] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01242_ ) );
NOR2_X1 _17137_ ( .A1(_01241_ ), .A2(_01242_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
AOI221_X4 _17138_ ( .A(_01214_ ), .B1(\LS_WB_wdata_csreg [8] ), .B2(_01223_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [8] ), .ZN(_01243_ ) );
AOI21_X1 _17139_ ( .A(\EX_LS_pc [8] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01244_ ) );
NOR2_X1 _17140_ ( .A1(_01243_ ), .A2(_01244_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
AOI21_X1 _17141_ ( .A(\EX_LS_pc [7] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01245_ ) );
OAI21_X1 _17142_ ( .A(_03843_ ), .B1(_01232_ ), .B2(_06157_ ), .ZN(_01246_ ) );
AOI221_X4 _17143_ ( .A(_01246_ ), .B1(\LS_WB_wdata_csreg [7] ), .B2(_01232_ ), .C1(_02093_ ), .C2(_06124_ ), .ZN(_01247_ ) );
NOR2_X1 _17144_ ( .A1(_01245_ ), .A2(_01247_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
AOI21_X1 _17145_ ( .A(\EX_LS_pc [6] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01248_ ) );
OAI21_X1 _17146_ ( .A(_03843_ ), .B1(_02129_ ), .B2(_05720_ ), .ZN(_01249_ ) );
AOI221_X4 _17147_ ( .A(_01249_ ), .B1(\LS_WB_wdata_csreg [6] ), .B2(_01232_ ), .C1(_02093_ ), .C2(_06124_ ), .ZN(_01250_ ) );
NOR2_X1 _17148_ ( .A1(_01248_ ), .A2(_01250_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
OAI22_X1 _17149_ ( .A1(_03835_ ), .A2(_02086_ ), .B1(_02025_ ), .B2(_06147_ ), .ZN(_01251_ ) );
MUX2_X1 _17150_ ( .A(_01251_ ), .B(\EX_LS_pc [5] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _17151_ ( .A(\LS_WB_wdata_csreg [4] ), .B(\EX_LS_result_csreg_mem [4] ), .S(_02128_ ), .Z(_01252_ ) );
MUX2_X1 _17152_ ( .A(_01252_ ), .B(\EX_LS_pc [4] ), .S(_01215_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
AOI221_X4 _17153_ ( .A(_01214_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [3] ), .C1(\LS_WB_wdata_csreg [3] ), .C2(_01223_ ), .ZN(_01253_ ) );
AOI21_X1 _17154_ ( .A(\EX_LS_pc [3] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01254_ ) );
NOR2_X1 _17155_ ( .A1(_01253_ ), .A2(_01254_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
AOI21_X1 _17156_ ( .A(\EX_LS_pc [2] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01255_ ) );
OAI21_X1 _17157_ ( .A(_03843_ ), .B1(_02129_ ), .B2(_06148_ ), .ZN(_01256_ ) );
AOI221_X4 _17158_ ( .A(_01256_ ), .B1(\LS_WB_wdata_csreg [2] ), .B2(_01232_ ), .C1(_02093_ ), .C2(_06124_ ), .ZN(_01257_ ) );
NOR2_X1 _17159_ ( .A1(_01255_ ), .A2(_01257_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _17160_ ( .A(\LS_WB_wdata_csreg [29] ), .B(\EX_LS_result_csreg_mem [29] ), .S(_02128_ ), .Z(_01258_ ) );
MUX2_X1 _17161_ ( .A(_01258_ ), .B(\EX_LS_pc [29] ), .S(_01214_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
AOI221_X4 _17162_ ( .A(_01214_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [1] ), .C1(\LS_WB_wdata_csreg [1] ), .C2(_01223_ ), .ZN(_01259_ ) );
AOI21_X1 _17163_ ( .A(\EX_LS_pc [1] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01260_ ) );
NOR2_X1 _17164_ ( .A1(_01259_ ), .A2(_01260_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI221_X4 _17165_ ( .A(_01214_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [0] ), .C1(\LS_WB_wdata_csreg [0] ), .C2(_01223_ ), .ZN(_01261_ ) );
AOI21_X1 _17166_ ( .A(\EX_LS_pc [0] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01262_ ) );
NOR2_X1 _17167_ ( .A1(_01261_ ), .A2(_01262_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
AOI21_X1 _17168_ ( .A(\EX_LS_pc [28] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01263_ ) );
OAI21_X1 _17169_ ( .A(_03843_ ), .B1(_02129_ ), .B2(_05623_ ), .ZN(_01264_ ) );
AOI221_X4 _17170_ ( .A(_01264_ ), .B1(\LS_WB_wdata_csreg [28] ), .B2(_01232_ ), .C1(_02093_ ), .C2(_06124_ ), .ZN(_01265_ ) );
NOR2_X1 _17171_ ( .A1(_01263_ ), .A2(_01265_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _17172_ ( .A(\EX_LS_pc [27] ), .B1(_03834_ ), .B2(_03844_ ), .ZN(_01266_ ) );
OAI21_X1 _17173_ ( .A(_03842_ ), .B1(_02129_ ), .B2(_05852_ ), .ZN(_01267_ ) );
AOI221_X4 _17174_ ( .A(_01267_ ), .B1(\LS_WB_wdata_csreg [27] ), .B2(_01232_ ), .C1(_02093_ ), .C2(_06124_ ), .ZN(_01268_ ) );
NOR2_X1 _17175_ ( .A1(_01266_ ), .A2(_01268_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI221_X4 _17176_ ( .A(_01214_ ), .B1(\LS_WB_wdata_csreg [26] ), .B2(_01223_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [26] ), .ZN(_01269_ ) );
AOI21_X1 _17177_ ( .A(\EX_LS_pc [26] ), .B1(_03833_ ), .B2(_01226_ ), .ZN(_01270_ ) );
NOR2_X1 _17178_ ( .A1(_01269_ ), .A2(_01270_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI21_X1 _17179_ ( .A(\EX_LS_pc [25] ), .B1(_01225_ ), .B2(_03844_ ), .ZN(_01271_ ) );
MUX2_X1 _17180_ ( .A(\LS_WB_wdata_csreg [25] ), .B(\EX_LS_result_csreg_mem [25] ), .S(_02128_ ), .Z(_01272_ ) );
NOR3_X1 _17181_ ( .A1(_03832_ ), .A2(_01212_ ), .A3(_01272_ ), .ZN(_01273_ ) );
NOR2_X1 _17182_ ( .A1(_01271_ ), .A2(_01273_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI221_X4 _17183_ ( .A(_01213_ ), .B1(\LS_WB_wdata_csreg [24] ), .B2(_01223_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [24] ), .ZN(_01274_ ) );
AOI21_X1 _17184_ ( .A(\EX_LS_pc [24] ), .B1(_03833_ ), .B2(_03843_ ), .ZN(_01275_ ) );
NOR2_X1 _17185_ ( .A1(_01274_ ), .A2(_01275_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _17186_ ( .A(\EX_LS_pc [23] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01276_ ) );
MUX2_X1 _17187_ ( .A(\LS_WB_wdata_csreg [23] ), .B(\EX_LS_result_csreg_mem [23] ), .S(_02128_ ), .Z(_01277_ ) );
NOR3_X1 _17188_ ( .A1(_03832_ ), .A2(_01212_ ), .A3(_01277_ ), .ZN(_01278_ ) );
NOR2_X1 _17189_ ( .A1(_01276_ ), .A2(_01278_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
AOI221_X4 _17190_ ( .A(_01213_ ), .B1(\LS_WB_wdata_csreg [22] ), .B2(_01223_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [22] ), .ZN(_01279_ ) );
AOI21_X1 _17191_ ( .A(\EX_LS_pc [22] ), .B1(_03833_ ), .B2(_03843_ ), .ZN(_01280_ ) );
NOR2_X1 _17192_ ( .A1(_01279_ ), .A2(_01280_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
AOI21_X1 _17193_ ( .A(\EX_LS_pc [31] ), .B1(_01225_ ), .B2(_01226_ ), .ZN(_01281_ ) );
MUX2_X1 _17194_ ( .A(\LS_WB_wdata_csreg [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_02128_ ), .Z(_01282_ ) );
NOR3_X1 _17195_ ( .A1(_03832_ ), .A2(_01212_ ), .A3(_01282_ ), .ZN(_01283_ ) );
NOR2_X1 _17196_ ( .A1(_01281_ ), .A2(_01283_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17197_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01284_ ) );
INV_X1 _17198_ ( .A(_01284_ ), .ZN(_01285_ ) );
OR3_X1 _17199_ ( .A1(_00534_ ), .A2(_06029_ ), .A3(_01285_ ), .ZN(_01286_ ) );
NAND3_X1 _17200_ ( .A1(_00507_ ), .A2(_06028_ ), .A3(_01285_ ), .ZN(_01287_ ) );
AND2_X1 _17201_ ( .A1(_01286_ ), .A2(_01287_ ), .ZN(_01288_ ) );
AND2_X1 _17202_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01289_ ) );
BUF_X4 _17203_ ( .A(_01289_ ), .Z(_01290_ ) );
INV_X1 _17204_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01291_ ) );
AND2_X2 _17205_ ( .A1(_01290_ ), .A2(_01291_ ), .ZN(_01292_ ) );
AND2_X1 _17206_ ( .A1(_01288_ ), .A2(_01292_ ), .ZN(_01293_ ) );
AND2_X1 _17207_ ( .A1(_01291_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01294_ ) );
INV_X1 _17208_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_01295_ ) );
AND2_X2 _17209_ ( .A1(_01294_ ), .A2(_01295_ ), .ZN(_01296_ ) );
NAND2_X1 _17210_ ( .A1(_01295_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01297_ ) );
NOR2_X1 _17211_ ( .A1(_01297_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01298_ ) );
OR2_X2 _17212_ ( .A1(_01296_ ), .A2(_01298_ ), .ZN(_01299_ ) );
NOR2_X2 _17213_ ( .A1(_01293_ ), .A2(_01299_ ), .ZN(_01300_ ) );
AND2_X1 _17214_ ( .A1(_01289_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01301_ ) );
BUF_X2 _17215_ ( .A(_01301_ ), .Z(_01302_ ) );
NOR4_X1 _17216_ ( .A1(_00513_ ), .A2(_00514_ ), .A3(_06031_ ), .A4(_01302_ ), .ZN(_01303_ ) );
BUF_X4 _17217_ ( .A(_01292_ ), .Z(_01304_ ) );
OAI21_X1 _17218_ ( .A(_01300_ ), .B1(_01303_ ), .B2(_01304_ ), .ZN(_01305_ ) );
INV_X1 _17219_ ( .A(_01296_ ), .ZN(_01306_ ) );
BUF_X4 _17220_ ( .A(_01306_ ), .Z(_01307_ ) );
NOR2_X1 _17221_ ( .A1(_00534_ ), .A2(_06030_ ), .ZN(_01308_ ) );
NOR2_X1 _17222_ ( .A1(_06077_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01309_ ) );
NOR2_X1 _17223_ ( .A1(_00602_ ), .A2(_06030_ ), .ZN(_01310_ ) );
NOR2_X1 _17224_ ( .A1(_06074_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01311_ ) );
AOI22_X1 _17225_ ( .A1(_01308_ ), .A2(_01309_ ), .B1(_01310_ ), .B2(_01311_ ), .ZN(_01312_ ) );
AND3_X1 _17226_ ( .A1(_00561_ ), .A2(_00563_ ), .A3(_06028_ ), .ZN(_01313_ ) );
NAND2_X1 _17227_ ( .A1(_01313_ ), .A2(_01284_ ), .ZN(_01314_ ) );
NAND4_X1 _17228_ ( .A1(_00507_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_06028_ ), .ZN(_01315_ ) );
AND3_X1 _17229_ ( .A1(_01312_ ), .A2(_01314_ ), .A3(_01315_ ), .ZN(_01316_ ) );
BUF_X4 _17230_ ( .A(_01316_ ), .Z(_01317_ ) );
OAI21_X1 _17231_ ( .A(_01305_ ), .B1(_01307_ ), .B2(_01317_ ), .ZN(_01318_ ) );
MUX2_X1 _17232_ ( .A(\EX_LS_result_reg [21] ), .B(_01318_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
INV_X1 _17233_ ( .A(_01302_ ), .ZN(_01319_ ) );
AND2_X2 _17234_ ( .A1(_01300_ ), .A2(_01319_ ), .ZN(_01320_ ) );
NOR2_X2 _17235_ ( .A1(_00517_ ), .A2(_06029_ ), .ZN(_01321_ ) );
OAI21_X1 _17236_ ( .A(_01320_ ), .B1(_01290_ ), .B2(_01321_ ), .ZN(_01322_ ) );
OAI21_X1 _17237_ ( .A(_01322_ ), .B1(_01307_ ), .B2(_01317_ ), .ZN(_01323_ ) );
MUX2_X1 _17238_ ( .A(\EX_LS_result_reg [20] ), .B(_01323_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
AND4_X1 _17239_ ( .A1(\io_master_arid [1] ), .A2(_00519_ ), .A3(_00522_ ), .A4(_01319_ ), .ZN(_01324_ ) );
OAI21_X1 _17240_ ( .A(_01300_ ), .B1(_01304_ ), .B2(_01324_ ), .ZN(_01325_ ) );
NOR2_X1 _17241_ ( .A1(_01316_ ), .A2(_01306_ ), .ZN(_01326_ ) );
NOR2_X2 _17242_ ( .A1(_01326_ ), .A2(_01166_ ), .ZN(_01327_ ) );
BUF_X4 _17243_ ( .A(_01166_ ), .Z(_01328_ ) );
AOI22_X1 _17244_ ( .A1(_01325_ ), .A2(_01327_ ), .B1(_01328_ ), .B2(_04652_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
AND4_X1 _17245_ ( .A1(\io_master_arid [1] ), .A2(_00523_ ), .A3(_00525_ ), .A4(_01319_ ), .ZN(_01329_ ) );
OAI21_X1 _17246_ ( .A(_01300_ ), .B1(_01304_ ), .B2(_01329_ ), .ZN(_01330_ ) );
OAI21_X1 _17247_ ( .A(_01330_ ), .B1(_01307_ ), .B2(_01317_ ), .ZN(_01331_ ) );
MUX2_X1 _17248_ ( .A(\EX_LS_result_reg [18] ), .B(_01331_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NOR4_X1 _17249_ ( .A1(_00527_ ), .A2(_00528_ ), .A3(_06032_ ), .A4(_01302_ ), .ZN(_01332_ ) );
OAI21_X1 _17250_ ( .A(_01300_ ), .B1(_01304_ ), .B2(_01332_ ), .ZN(_01333_ ) );
AOI22_X1 _17251_ ( .A1(_01333_ ), .A2(_01327_ ), .B1(_01328_ ), .B2(_04724_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NOR4_X1 _17252_ ( .A1(_00530_ ), .A2(_00531_ ), .A3(_06031_ ), .A4(_01302_ ), .ZN(_01334_ ) );
OAI21_X1 _17253_ ( .A(_01300_ ), .B1(_01304_ ), .B2(_01334_ ), .ZN(_01335_ ) );
OAI21_X1 _17254_ ( .A(_01335_ ), .B1(_01307_ ), .B2(_01317_ ), .ZN(_01336_ ) );
MUX2_X1 _17255_ ( .A(\EX_LS_result_reg [16] ), .B(_01336_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
INV_X1 _17256_ ( .A(_01290_ ), .ZN(_01337_ ) );
AOI21_X1 _17257_ ( .A(_01337_ ), .B1(_01286_ ), .B2(_01287_ ), .ZN(_01338_ ) );
NOR3_X1 _17258_ ( .A1(_01296_ ), .A2(_01290_ ), .A3(_01298_ ), .ZN(_01339_ ) );
AOI21_X1 _17259_ ( .A(_01338_ ), .B1(_01308_ ), .B2(_01339_ ), .ZN(_01340_ ) );
AOI22_X1 _17260_ ( .A1(_01327_ ), .A2(_01340_ ), .B1(_01328_ ), .B2(_04232_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
NOR2_X1 _17261_ ( .A1(_01337_ ), .A2(_01284_ ), .ZN(_01341_ ) );
INV_X1 _17262_ ( .A(_01341_ ), .ZN(_01342_ ) );
NOR3_X1 _17263_ ( .A1(_00511_ ), .A2(_06031_ ), .A3(_01342_ ), .ZN(_01343_ ) );
NOR2_X1 _17264_ ( .A1(_00537_ ), .A2(_06029_ ), .ZN(_01344_ ) );
AOI21_X1 _17265_ ( .A(_01343_ ), .B1(_01344_ ), .B2(_01342_ ), .ZN(_01345_ ) );
OAI22_X1 _17266_ ( .A1(_01317_ ), .A2(_01307_ ), .B1(_01299_ ), .B2(_01345_ ), .ZN(_01346_ ) );
MUX2_X1 _17267_ ( .A(\EX_LS_result_reg [14] ), .B(_01346_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
NAND2_X1 _17268_ ( .A1(\io_master_arid [1] ), .A2(_01342_ ), .ZN(_01347_ ) );
NOR2_X1 _17269_ ( .A1(_01347_ ), .A2(_01299_ ), .ZN(_01348_ ) );
AND3_X1 _17270_ ( .A1(_00538_ ), .A2(_00541_ ), .A3(_01348_ ), .ZN(_01349_ ) );
AND2_X1 _17271_ ( .A1(_00546_ ), .A2(_00547_ ), .ZN(_01350_ ) );
NOR2_X1 _17272_ ( .A1(_01350_ ), .A2(_06032_ ), .ZN(_01351_ ) );
AOI21_X1 _17273_ ( .A(_01349_ ), .B1(_01351_ ), .B2(_01341_ ), .ZN(_01352_ ) );
AOI22_X1 _17274_ ( .A1(_01327_ ), .A2(_01352_ ), .B1(_01328_ ), .B2(_04285_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
OR3_X1 _17275_ ( .A1(_00581_ ), .A2(_06031_ ), .A3(_01342_ ), .ZN(_01353_ ) );
OR4_X1 _17276_ ( .A1(_06031_ ), .A2(_00544_ ), .A3(_01299_ ), .A4(_01341_ ), .ZN(_01354_ ) );
OAI211_X1 _17277_ ( .A(_01353_ ), .B(_01354_ ), .C1(_01317_ ), .C2(_01307_ ), .ZN(_01355_ ) );
MUX2_X1 _17278_ ( .A(\EX_LS_result_reg [12] ), .B(_01355_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
NOR2_X1 _17279_ ( .A1(_00511_ ), .A2(_06029_ ), .ZN(_01356_ ) );
OAI21_X1 _17280_ ( .A(_01320_ ), .B1(_01290_ ), .B2(_01356_ ), .ZN(_01357_ ) );
OAI21_X1 _17281_ ( .A(_01357_ ), .B1(_01307_ ), .B2(_01317_ ), .ZN(_01358_ ) );
MUX2_X1 _17282_ ( .A(\EX_LS_result_reg [30] ), .B(_01358_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _17283_ ( .A1(_00548_ ), .A2(_00550_ ), .A3(_01348_ ), .ZN(_01359_ ) );
NAND2_X1 _17284_ ( .A1(_00588_ ), .A2(_00590_ ), .ZN(_01360_ ) );
OR2_X1 _17285_ ( .A1(_01360_ ), .A2(_06031_ ), .ZN(_01361_ ) );
OAI221_X1 _17286_ ( .A(_01359_ ), .B1(_01342_ ), .B2(_01361_ ), .C1(_01316_ ), .C2(_01306_ ), .ZN(_01362_ ) );
MUX2_X1 _17287_ ( .A(\EX_LS_result_reg [11] ), .B(_01362_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
AND2_X1 _17288_ ( .A1(_00592_ ), .A2(_00593_ ), .ZN(_01363_ ) );
OR3_X1 _17289_ ( .A1(_01363_ ), .A2(_06031_ ), .A3(_01342_ ), .ZN(_01364_ ) );
NAND3_X1 _17290_ ( .A1(_00551_ ), .A2(_00553_ ), .A3(_01348_ ), .ZN(_01365_ ) );
OAI211_X1 _17291_ ( .A(_01364_ ), .B(_01365_ ), .C1(_01317_ ), .C2(_01306_ ), .ZN(_01366_ ) );
MUX2_X1 _17292_ ( .A(\EX_LS_result_reg [10] ), .B(_01366_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17293_ ( .A1(_00555_ ), .A2(_00557_ ), .A3(_01348_ ), .ZN(_01367_ ) );
NAND2_X1 _17294_ ( .A1(_00594_ ), .A2(_00596_ ), .ZN(_01368_ ) );
NOR2_X1 _17295_ ( .A1(_01368_ ), .A2(_06032_ ), .ZN(_01369_ ) );
AOI21_X1 _17296_ ( .A(_01367_ ), .B1(_01369_ ), .B2(_01341_ ), .ZN(_01370_ ) );
AOI22_X1 _17297_ ( .A1(_01327_ ), .A2(_01370_ ), .B1(_01328_ ), .B2(_04101_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17298_ ( .A1(_00558_ ), .A2(_00560_ ), .A3(_01348_ ), .ZN(_01371_ ) );
AND2_X1 _17299_ ( .A1(_00598_ ), .A2(_00599_ ), .ZN(_01372_ ) );
NOR2_X1 _17300_ ( .A1(_01372_ ), .A2(_06032_ ), .ZN(_01373_ ) );
AOI21_X1 _17301_ ( .A(_01371_ ), .B1(_01373_ ), .B2(_01341_ ), .ZN(_01374_ ) );
AOI22_X1 _17302_ ( .A1(_01327_ ), .A2(_01374_ ), .B1(_01328_ ), .B2(_04146_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
AND4_X1 _17303_ ( .A1(_01299_ ), .A2(_01312_ ), .A3(_01314_ ), .A4(_01315_ ), .ZN(_01375_ ) );
NOR3_X1 _17304_ ( .A1(_00602_ ), .A2(_06031_ ), .A3(_01342_ ), .ZN(_01376_ ) );
AOI211_X1 _17305_ ( .A(_01299_ ), .B(_01376_ ), .C1(_01313_ ), .C2(_01342_ ), .ZN(_01377_ ) );
OR3_X1 _17306_ ( .A1(_01375_ ), .A2(_01166_ ), .A3(_01377_ ), .ZN(_01378_ ) );
OAI21_X1 _17307_ ( .A(_01378_ ), .B1(\mylsu.state [3] ), .B2(_04923_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
NOR2_X2 _17308_ ( .A1(_00566_ ), .A2(_06029_ ), .ZN(_01379_ ) );
NOR2_X2 _17309_ ( .A1(_00605_ ), .A2(_06029_ ), .ZN(_01380_ ) );
MUX2_X1 _17310_ ( .A(_01356_ ), .B(_01380_ ), .S(_01311_ ), .Z(_01381_ ) );
INV_X1 _17311_ ( .A(_01309_ ), .ZN(_01382_ ) );
MUX2_X2 _17312_ ( .A(_01344_ ), .B(_01381_ ), .S(_01382_ ), .Z(_01383_ ) );
MUX2_X1 _17313_ ( .A(_01379_ ), .B(_01383_ ), .S(_01285_ ), .Z(_01384_ ) );
MUX2_X1 _17314_ ( .A(_01379_ ), .B(_01380_ ), .S(_01285_ ), .Z(_01385_ ) );
MUX2_X1 _17315_ ( .A(_01379_ ), .B(_01385_ ), .S(_01301_ ), .Z(_01386_ ) );
MUX2_X1 _17316_ ( .A(_01386_ ), .B(_01385_ ), .S(_01292_ ), .Z(_01387_ ) );
MUX2_X1 _17317_ ( .A(_01387_ ), .B(_01384_ ), .S(_01298_ ), .Z(_01388_ ) );
MUX2_X1 _17318_ ( .A(_01384_ ), .B(_01388_ ), .S(_01306_ ), .Z(_01389_ ) );
MUX2_X1 _17319_ ( .A(\EX_LS_result_reg [6] ), .B(_01389_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _17320_ ( .A1(_01166_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01390_ ) );
NOR2_X1 _17321_ ( .A1(_01339_ ), .A2(_01284_ ), .ZN(_01391_ ) );
INV_X1 _17322_ ( .A(_01391_ ), .ZN(_01392_ ) );
AOI211_X1 _17323_ ( .A(_01166_ ), .B(_06032_ ), .C1(_00569_ ), .C2(_01392_ ), .ZN(_01393_ ) );
AND2_X1 _17324_ ( .A1(_01299_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01394_ ) );
NOR2_X1 _17325_ ( .A1(_01392_ ), .A2(_01394_ ), .ZN(_01395_ ) );
OAI21_X1 _17326_ ( .A(_01395_ ), .B1(_00513_ ), .B2(_00514_ ), .ZN(_01396_ ) );
NAND2_X1 _17327_ ( .A1(_01393_ ), .A2(_01396_ ), .ZN(_01397_ ) );
NAND3_X1 _17328_ ( .A1(_00538_ ), .A2(_00541_ ), .A3(_06074_ ), .ZN(_01398_ ) );
NAND3_X1 _17329_ ( .A1(_06122_ ), .A2(_06123_ ), .A3(_00545_ ), .ZN(_01399_ ) );
OAI211_X1 _17330_ ( .A(\mylsu.araddr_tmp [1] ), .B(_01399_ ), .C1(_00554_ ), .C2(\io_master_rdata [29] ), .ZN(_01400_ ) );
AND3_X1 _17331_ ( .A1(_01398_ ), .A2(_01394_ ), .A3(_01400_ ), .ZN(_01401_ ) );
OAI21_X1 _17332_ ( .A(_01390_ ), .B1(_01397_ ), .B2(_01401_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
OR3_X1 _17333_ ( .A1(_00572_ ), .A2(_06030_ ), .A3(_01285_ ), .ZN(_01402_ ) );
NOR3_X1 _17334_ ( .A1(_00544_ ), .A2(_06030_ ), .A3(_01382_ ), .ZN(_01403_ ) );
NOR2_X1 _17335_ ( .A1(_00581_ ), .A2(_06029_ ), .ZN(_01404_ ) );
MUX2_X1 _17336_ ( .A(_01404_ ), .B(_01321_ ), .S(_01311_ ), .Z(_01405_ ) );
AOI21_X1 _17337_ ( .A(_01403_ ), .B1(_01405_ ), .B2(_01382_ ), .ZN(_01406_ ) );
OAI21_X1 _17338_ ( .A(_01402_ ), .B1(_01406_ ), .B2(_01284_ ), .ZN(_01407_ ) );
NOR2_X2 _17339_ ( .A1(_00572_ ), .A2(_06029_ ), .ZN(_01408_ ) );
MUX2_X2 _17340_ ( .A(_01408_ ), .B(_01321_ ), .S(_01285_ ), .Z(_01409_ ) );
MUX2_X1 _17341_ ( .A(_01408_ ), .B(_01409_ ), .S(_01301_ ), .Z(_01410_ ) );
MUX2_X1 _17342_ ( .A(_01410_ ), .B(_01409_ ), .S(_01292_ ), .Z(_01411_ ) );
MUX2_X1 _17343_ ( .A(_01411_ ), .B(_01407_ ), .S(_01298_ ), .Z(_01412_ ) );
MUX2_X1 _17344_ ( .A(_01407_ ), .B(_01412_ ), .S(_01306_ ), .Z(_01413_ ) );
MUX2_X1 _17345_ ( .A(\EX_LS_result_reg [4] ), .B(_01413_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
NOR3_X1 _17346_ ( .A1(_01360_ ), .A2(_06030_ ), .A3(_01311_ ), .ZN(_01414_ ) );
AND4_X1 _17347_ ( .A1(_06028_ ), .A2(_00519_ ), .A3(_00522_ ), .A4(_01311_ ), .ZN(_01415_ ) );
OAI21_X1 _17348_ ( .A(_01382_ ), .B1(_01414_ ), .B2(_01415_ ), .ZN(_01416_ ) );
NAND4_X1 _17349_ ( .A1(_00548_ ), .A2(_00550_ ), .A3(\io_master_arid [1] ), .A4(_01309_ ), .ZN(_01417_ ) );
AOI21_X1 _17350_ ( .A(_01284_ ), .B1(_01416_ ), .B2(_01417_ ), .ZN(_01418_ ) );
NOR3_X1 _17351_ ( .A1(_00575_ ), .A2(_06030_ ), .A3(_01285_ ), .ZN(_01419_ ) );
OAI21_X1 _17352_ ( .A(_01296_ ), .B1(_01418_ ), .B2(_01419_ ), .ZN(_01420_ ) );
AND4_X1 _17353_ ( .A1(_06028_ ), .A2(_00519_ ), .A3(_00522_ ), .A4(_01285_ ), .ZN(_01421_ ) );
OR2_X1 _17354_ ( .A1(_01419_ ), .A2(_01421_ ), .ZN(_01422_ ) );
AND2_X1 _17355_ ( .A1(_01422_ ), .A2(_01292_ ), .ZN(_01423_ ) );
OAI21_X1 _17356_ ( .A(_01302_ ), .B1(_01419_ ), .B2(_01421_ ), .ZN(_01424_ ) );
OR3_X1 _17357_ ( .A1(_00575_ ), .A2(_06030_ ), .A3(_01302_ ), .ZN(_01425_ ) );
AOI21_X1 _17358_ ( .A(_01304_ ), .B1(_01424_ ), .B2(_01425_ ), .ZN(_01426_ ) );
OAI22_X1 _17359_ ( .A1(_01423_ ), .A2(_01426_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01297_ ), .ZN(_01427_ ) );
OAI21_X1 _17360_ ( .A(_01298_ ), .B1(_01418_ ), .B2(_01419_ ), .ZN(_01428_ ) );
AND2_X1 _17361_ ( .A1(_01427_ ), .A2(_01428_ ), .ZN(_01429_ ) );
OAI21_X1 _17362_ ( .A(_01420_ ), .B1(_01429_ ), .B2(_01296_ ), .ZN(_01430_ ) );
MUX2_X1 _17363_ ( .A(\EX_LS_result_reg [3] ), .B(_01430_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
AOI211_X1 _17364_ ( .A(_06030_ ), .B(_01311_ ), .C1(_00592_ ), .C2(_00593_ ), .ZN(_01431_ ) );
AND4_X1 _17365_ ( .A1(_06028_ ), .A2(_00523_ ), .A3(_00525_ ), .A4(_01311_ ), .ZN(_01432_ ) );
OAI21_X1 _17366_ ( .A(_01382_ ), .B1(_01431_ ), .B2(_01432_ ), .ZN(_01433_ ) );
NAND4_X1 _17367_ ( .A1(_00551_ ), .A2(_00553_ ), .A3(_06028_ ), .A4(_01309_ ), .ZN(_01434_ ) );
AOI21_X1 _17368_ ( .A(_01284_ ), .B1(_01433_ ), .B2(_01434_ ), .ZN(_01435_ ) );
NOR3_X1 _17369_ ( .A1(_00578_ ), .A2(_06029_ ), .A3(_01285_ ), .ZN(_01436_ ) );
OAI21_X1 _17370_ ( .A(_01296_ ), .B1(_01435_ ), .B2(_01436_ ), .ZN(_01437_ ) );
AND4_X1 _17371_ ( .A1(_06028_ ), .A2(_00523_ ), .A3(_00525_ ), .A4(_01285_ ), .ZN(_01438_ ) );
OR2_X1 _17372_ ( .A1(_01436_ ), .A2(_01438_ ), .ZN(_01439_ ) );
AND2_X1 _17373_ ( .A1(_01439_ ), .A2(_01292_ ), .ZN(_01440_ ) );
OAI21_X1 _17374_ ( .A(_01302_ ), .B1(_01436_ ), .B2(_01438_ ), .ZN(_01441_ ) );
OR3_X1 _17375_ ( .A1(_00578_ ), .A2(_06030_ ), .A3(_01302_ ), .ZN(_01442_ ) );
AOI21_X1 _17376_ ( .A(_01304_ ), .B1(_01441_ ), .B2(_01442_ ), .ZN(_01443_ ) );
OAI22_X1 _17377_ ( .A1(_01440_ ), .A2(_01443_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01297_ ), .ZN(_01444_ ) );
OAI21_X1 _17378_ ( .A(_01298_ ), .B1(_01435_ ), .B2(_01436_ ), .ZN(_01445_ ) );
AND2_X1 _17379_ ( .A1(_01444_ ), .A2(_01445_ ), .ZN(_01446_ ) );
OAI21_X1 _17380_ ( .A(_01437_ ), .B1(_01446_ ), .B2(_01296_ ), .ZN(_01447_ ) );
MUX2_X1 _17381_ ( .A(\EX_LS_result_reg [2] ), .B(_01447_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
OAI21_X1 _17382_ ( .A(_01320_ ), .B1(_01290_ ), .B2(_01351_ ), .ZN(_01448_ ) );
OAI21_X1 _17383_ ( .A(_01448_ ), .B1(_01307_ ), .B2(_01317_ ), .ZN(_01449_ ) );
MUX2_X1 _17384_ ( .A(\EX_LS_result_reg [29] ), .B(_01449_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
NAND2_X1 _17385_ ( .A1(_00584_ ), .A2(_01392_ ), .ZN(_01450_ ) );
AND2_X1 _17386_ ( .A1(\io_master_arid [1] ), .A2(\mylsu.state [3] ), .ZN(_01451_ ) );
OAI21_X1 _17387_ ( .A(_01395_ ), .B1(_00527_ ), .B2(_00528_ ), .ZN(_01452_ ) );
NAND3_X1 _17388_ ( .A1(_01450_ ), .A2(_01451_ ), .A3(_01452_ ), .ZN(_01453_ ) );
NAND3_X1 _17389_ ( .A1(_00594_ ), .A2(_00596_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01454_ ) );
NAND3_X1 _17390_ ( .A1(_00555_ ), .A2(_00557_ ), .A3(_06074_ ), .ZN(_01455_ ) );
AND3_X1 _17391_ ( .A1(_01454_ ), .A2(_01455_ ), .A3(_01394_ ), .ZN(_01456_ ) );
OAI22_X1 _17392_ ( .A1(_01453_ ), .A2(_01456_ ), .B1(\mylsu.state [3] ), .B2(_04340_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
NAND2_X1 _17393_ ( .A1(_01166_ ), .A2(\EX_LS_result_reg [0] ), .ZN(_01457_ ) );
OR2_X1 _17394_ ( .A1(_01372_ ), .A2(_06074_ ), .ZN(_01458_ ) );
NAND3_X1 _17395_ ( .A1(_00558_ ), .A2(_00560_ ), .A3(_06074_ ), .ZN(_01459_ ) );
AND3_X1 _17396_ ( .A1(_01458_ ), .A2(_01394_ ), .A3(_01459_ ), .ZN(_01460_ ) );
NAND2_X1 _17397_ ( .A1(_00587_ ), .A2(_01392_ ), .ZN(_01461_ ) );
OAI21_X1 _17398_ ( .A(_01395_ ), .B1(_00530_ ), .B2(_00531_ ), .ZN(_01462_ ) );
NAND3_X1 _17399_ ( .A1(_01461_ ), .A2(_01451_ ), .A3(_01462_ ), .ZN(_01463_ ) );
OAI21_X1 _17400_ ( .A(_01457_ ), .B1(_01460_ ), .B2(_01463_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
NOR3_X1 _17401_ ( .A1(_00581_ ), .A2(_06032_ ), .A3(_01302_ ), .ZN(_01464_ ) );
OAI21_X1 _17402_ ( .A(_01300_ ), .B1(_01304_ ), .B2(_01464_ ), .ZN(_01465_ ) );
OAI21_X1 _17403_ ( .A(_01465_ ), .B1(_01307_ ), .B2(_01317_ ), .ZN(_01466_ ) );
MUX2_X1 _17404_ ( .A(\EX_LS_result_reg [28] ), .B(_01466_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
OR4_X1 _17405_ ( .A1(_01302_ ), .A2(_01293_ ), .A3(_01299_ ), .A4(_01361_ ), .ZN(_01467_ ) );
NOR4_X1 _17406_ ( .A1(_01288_ ), .A2(\mylsu.typ_tmp [0] ), .A3(_01337_ ), .A4(_01299_ ), .ZN(_01468_ ) );
NOR3_X1 _17407_ ( .A1(_01326_ ), .A2(_01468_ ), .A3(_01166_ ), .ZN(_01469_ ) );
AOI22_X1 _17408_ ( .A1(_01467_ ), .A2(_01469_ ), .B1(_01328_ ), .B2(_04593_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
AOI211_X1 _17409_ ( .A(_06032_ ), .B(_01290_ ), .C1(_00592_ ), .C2(_00593_ ), .ZN(_01470_ ) );
OAI21_X1 _17410_ ( .A(_01300_ ), .B1(_01304_ ), .B2(_01470_ ), .ZN(_01471_ ) );
AOI22_X1 _17411_ ( .A1(_01471_ ), .A2(_01327_ ), .B1(_01328_ ), .B2(_04569_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
OAI21_X1 _17412_ ( .A(_01320_ ), .B1(_01290_ ), .B2(_01369_ ), .ZN(_01472_ ) );
AOI22_X1 _17413_ ( .A1(_01472_ ), .A2(_01327_ ), .B1(_01328_ ), .B2(_04643_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
NAND3_X1 _17414_ ( .A1(_01300_ ), .A2(_01319_ ), .A3(_01373_ ), .ZN(_01473_ ) );
AOI22_X1 _17415_ ( .A1(_01469_ ), .A2(_01473_ ), .B1(_01328_ ), .B2(_04619_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
OAI21_X1 _17416_ ( .A(_01320_ ), .B1(_01290_ ), .B2(_01310_ ), .ZN(_01474_ ) );
AOI22_X1 _17417_ ( .A1(_01474_ ), .A2(_01327_ ), .B1(_01166_ ), .B2(_04794_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
OAI21_X1 _17418_ ( .A(_01320_ ), .B1(_01290_ ), .B2(_01380_ ), .ZN(_01475_ ) );
AOI22_X1 _17419_ ( .A1(_01475_ ), .A2(_01327_ ), .B1(_01166_ ), .B2(_04750_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17420_ ( .A1(_00507_ ), .A2(\io_master_arid [1] ), .A3(_01337_ ), .ZN(_01476_ ) );
OAI21_X1 _17421_ ( .A(_01300_ ), .B1(_01304_ ), .B2(_01476_ ), .ZN(_01477_ ) );
OAI21_X1 _17422_ ( .A(_01477_ ), .B1(_01307_ ), .B2(_01316_ ), .ZN(_01478_ ) );
MUX2_X1 _17423_ ( .A(\EX_LS_result_reg [31] ), .B(_01478_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17424_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(\LS_WB_waddr_reg [1] ), .ZN(_01479_ ) );
INV_X1 _17425_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01480_ ) );
INV_X1 _17426_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01481_ ) );
NAND3_X1 _17427_ ( .A1(_01479_ ), .A2(_01480_ ), .A3(_01481_ ), .ZN(_01482_ ) );
AND2_X1 _17428_ ( .A1(_01558_ ), .A2(LS_WB_wen_reg ), .ZN(_01483_ ) );
NAND2_X1 _17429_ ( .A1(_01482_ ), .A2(_01483_ ), .ZN(_01484_ ) );
BUF_X4 _17430_ ( .A(_01484_ ), .Z(_01485_ ) );
INV_X1 _17431_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01486_ ) );
AOI21_X1 _17432_ ( .A(_01485_ ), .B1(_01486_ ), .B2(_01481_ ), .ZN(_01487_ ) );
NOR2_X1 _17433_ ( .A1(_01484_ ), .A2(_01480_ ), .ZN(_01488_ ) );
INV_X1 _17434_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01489_ ) );
NOR4_X1 _17435_ ( .A1(_01487_ ), .A2(_01488_ ), .A3(_01489_ ), .A4(_01485_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _17436_ ( .A1(_01485_ ), .A2(_01489_ ), .ZN(_01490_ ) );
NOR2_X1 _17437_ ( .A1(_01485_ ), .A2(_01481_ ), .ZN(_01491_ ) );
AND4_X1 _17438_ ( .A1(_01480_ ), .A2(_01490_ ), .A3(_01491_ ), .A4(_01486_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _17439_ ( .A1(_01489_ ), .A2(_01488_ ), .A3(_01491_ ), .A4(_01486_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR2_X1 _17440_ ( .A1(_01484_ ), .A2(_01486_ ), .ZN(_01492_ ) );
AND4_X1 _17441_ ( .A1(_01489_ ), .A2(_01488_ ), .A3(_01492_ ), .A4(_01481_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
CLKBUF_X1 _17442_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
AOI21_X1 _17443_ ( .A(_01485_ ), .B1(_01480_ ), .B2(_01489_ ), .ZN(_01493_ ) );
NOR4_X1 _17444_ ( .A1(_01493_ ), .A2(_01492_ ), .A3(_01481_ ), .A4(_01485_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17445_ ( .A1(_01493_ ), .A2(_01491_ ), .A3(_01486_ ), .A4(_01485_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17446_ ( .A1(_01480_ ), .A2(_01490_ ), .A3(_01492_ ), .A4(_01481_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17447_ ( .A1(_01480_ ), .A2(_01490_ ), .A3(_01492_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _17448_ ( .A1(_01487_ ), .A2(_01490_ ), .A3(_01480_ ), .A4(_01485_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
NOR4_X1 _17449_ ( .A1(_01487_ ), .A2(_01480_ ), .A3(_01489_ ), .A4(_01485_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17450_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01488_ ), .A3(_01491_ ), .A4(_01486_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17451_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01488_ ), .A3(_01492_ ), .A4(_01481_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17452_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01488_ ), .A3(_01491_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17453_ ( .A1(_01489_ ), .A2(_01488_ ), .A3(_01492_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17454_ ( .A1(_01493_ ), .A2(_01486_ ), .A3(_01481_ ), .A4(_01485_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17455_ ( .A1(_01964_ ), .A2(_01631_ ), .A3(_01971_ ), .ZN(_01494_ ) );
NAND2_X1 _17456_ ( .A1(_01494_ ), .A2(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17457_ ( .A(reset ), .B(_01964_ ), .C1(_01965_ ), .C2(_06085_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17458_ ( .A(_01482_ ), .Z(_01495_ ) );
CLKBUF_X2 _17459_ ( .A(_01483_ ), .Z(_01496_ ) );
AND3_X1 _17460_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17461_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17462_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17463_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17464_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17465_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17466_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17467_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17468_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17469_ ( .A1(_01495_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01496_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17470_ ( .A(_01482_ ), .Z(_01497_ ) );
CLKBUF_X2 _17471_ ( .A(_01483_ ), .Z(_01498_ ) );
AND3_X1 _17472_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17473_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17474_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17475_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17476_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17477_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17478_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17479_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17480_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17481_ ( .A1(_01497_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01498_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17482_ ( .A(_01482_ ), .Z(_01499_ ) );
CLKBUF_X2 _17483_ ( .A(_01483_ ), .Z(_01500_ ) );
AND3_X1 _17484_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17485_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17486_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17487_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17488_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17489_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17490_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17491_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17492_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17493_ ( .A1(_01499_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01500_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17494_ ( .A1(_01482_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01483_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17495_ ( .A1(_01482_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01483_ ), .ZN(\myreg.Reg[3]_$_DFFE_PP__Q_D ) );
AND3_X1 _17496_ ( .A1(_01631_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17497_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01501_ ) );
AND2_X1 _17498_ ( .A1(_01501_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01502_ ) );
INV_X1 _17499_ ( .A(_01502_ ), .ZN(_01503_ ) );
NOR2_X1 _17500_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01504_ ) );
OAI211_X1 _17501_ ( .A(_01558_ ), .B(\mysc.state [0] ), .C1(_01503_ ), .C2(_01504_ ), .ZN(_01505_ ) );
INV_X1 _17502_ ( .A(_01505_ ), .ZN(_01506_ ) );
OR3_X1 _17503_ ( .A1(_01506_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17504_ ( .A1(_01503_ ), .A2(reset ), .A3(_01504_ ), .ZN(_01507_ ) );
NAND2_X1 _17505_ ( .A1(_01507_ ), .A2(\mysc.state [0] ), .ZN(_01508_ ) );
OR3_X1 _17506_ ( .A1(_03871_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01509_ ) );
NAND2_X1 _17507_ ( .A1(_01508_ ), .A2(_01509_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17508_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07984_ ) );
CLKGATE_X1 _17509_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_07985_ ) );
CLKGATE_X1 _17510_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07986_ ) );
CLKGATE_X1 _17511_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07987_ ) );
CLKGATE_X1 _17512_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07988_ ) );
CLKGATE_X1 _17513_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07989_ ) );
CLKGATE_X1 _17514_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_07990_ ) );
CLKGATE_X1 _17515_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_07991_ ) );
CLKGATE_X1 _17516_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_07992_ ) );
CLKGATE_X1 _17517_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_07993_ ) );
CLKGATE_X1 _17518_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_07994_ ) );
CLKGATE_X1 _17519_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07995_ ) );
CLKGATE_X1 _17520_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07996_ ) );
CLKGATE_X1 _17521_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07997_ ) );
CLKGATE_X1 _17522_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_07998_ ) );
CLKGATE_X1 _17523_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07999_ ) );
CLKGATE_X1 _17524_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_08000_ ) );
CLKGATE_X1 _17525_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08001_ ) );
CLKGATE_X1 _17526_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_08002_ ) );
CLKGATE_X1 _17527_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ), .GCK(_08003_ ) );
CLKGATE_X1 _17528_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .GCK(_08004_ ) );
CLKGATE_X1 _17529_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08005_ ) );
CLKGATE_X1 _17530_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_2_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_08006_ ) );
CLKGATE_X1 _17531_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_08007_ ) );
CLKGATE_X1 _17532_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_08008_ ) );
CLKGATE_X1 _17533_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_08009_ ) );
CLKGATE_X1 _17534_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_08010_ ) );
CLKGATE_X1 _17535_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_08011_ ) );
CLKGATE_X1 _17536_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_08012_ ) );
CLKGATE_X1 _17537_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_08013_ ) );
CLKGATE_X1 _17538_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_08014_ ) );
CLKGATE_X1 _17539_ ( .CK(clock ), .E(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ), .GCK(_08015_ ) );
CLKGATE_X1 _17540_ ( .CK(clock ), .E(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ), .GCK(_08016_ ) );
CLKGATE_X1 _17541_ ( .CK(clock ), .E(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ), .GCK(_08017_ ) );
CLKGATE_X1 _17542_ ( .CK(clock ), .E(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ), .GCK(_08018_ ) );
CLKGATE_X1 _17543_ ( .CK(clock ), .E(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ), .GCK(_08019_ ) );
CLKGATE_X1 _17544_ ( .CK(clock ), .E(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ), .GCK(_08020_ ) );
CLKGATE_X1 _17545_ ( .CK(clock ), .E(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ), .GCK(_08021_ ) );
CLKGATE_X1 _17546_ ( .CK(clock ), .E(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ), .GCK(_08022_ ) );
CLKGATE_X1 _17547_ ( .CK(clock ), .E(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ), .GCK(_08023_ ) );
CLKGATE_X1 _17548_ ( .CK(clock ), .E(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ), .GCK(_08024_ ) );
CLKGATE_X1 _17549_ ( .CK(clock ), .E(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ), .GCK(_08025_ ) );
CLKGATE_X1 _17550_ ( .CK(clock ), .E(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ), .GCK(_08026_ ) );
CLKGATE_X1 _17551_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08027_ ) );
CLKGATE_X1 _17552_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08028_ ) );
CLKGATE_X1 _17553_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_08029_ ) );
CLKGATE_X1 _17554_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08030_ ) );
CLKGATE_X1 _17555_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08031_ ) );
CLKGATE_X1 _17556_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08032_ ) );
CLKGATE_X1 _17557_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08033_ ) );
CLKGATE_X1 _17558_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08034_ ) );
CLKGATE_X1 _17559_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_08035_ ) );
CLKGATE_X1 _17560_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08036_ ) );
CLKGATE_X1 _17561_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08037_ ) );
CLKGATE_X1 _17562_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08038_ ) );
CLKGATE_X1 _17563_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08039_ ) );
CLKGATE_X1 _17564_ ( .CK(clock ), .E(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08040_ ) );
CLKGATE_X1 _17565_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_08041_ ) );
CLKGATE_X1 _17566_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ), .GCK(_08042_ ) );
CLKGATE_X1 _17567_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08043_ ) );
CLKGATE_X1 _17568_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08044_ ) );
CLKGATE_X1 _17569_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFFE_PP0P__Q_E ), .GCK(_08045_ ) );
CLKGATE_X1 _17570_ ( .CK(clock ), .E(\mycsreg.CSReg[3]_$_DFFE_PP__Q_E ), .GCK(_08046_ ) );
CLKGATE_X1 _17571_ ( .CK(clock ), .E(\mycsreg.CSReg[2]_$_DFFE_PP__Q_E ), .GCK(_08047_ ) );
CLKGATE_X1 _17572_ ( .CK(clock ), .E(\mycsreg.CSReg[1]_$_DFFE_PP__Q_E ), .GCK(_08048_ ) );
CLKGATE_X1 _17573_ ( .CK(clock ), .E(\mycsreg.CSReg[0]_$_DFFE_PP__Q_E ), .GCK(_08049_ ) );
LOGIC1_X1 _17574_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17575_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08280_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08281_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08282_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08283_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08284_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08285_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08286_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08287_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08288_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08289_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08290_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08291_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08292_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08293_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08294_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08295_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08296_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08297_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08298_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08299_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08300_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08301_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08302_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08303_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08304_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08305_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08306_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08307_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08308_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08309_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08310_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08049_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08311_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08048_ ), .Q(\mtvec [31] ), .QN(_08312_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08048_ ), .Q(\mtvec [30] ), .QN(_08313_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08048_ ), .Q(\mtvec [21] ), .QN(_08314_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08048_ ), .Q(\mtvec [20] ), .QN(_08315_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08048_ ), .Q(\mtvec [19] ), .QN(_08316_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08048_ ), .Q(\mtvec [18] ), .QN(_08317_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08048_ ), .Q(\mtvec [17] ), .QN(_08318_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08048_ ), .Q(\mtvec [16] ), .QN(_08319_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08048_ ), .Q(\mtvec [15] ), .QN(_08320_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08048_ ), .Q(\mtvec [14] ), .QN(_08321_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08048_ ), .Q(\mtvec [13] ), .QN(_08322_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08048_ ), .Q(\mtvec [12] ), .QN(_08323_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08048_ ), .Q(\mtvec [29] ), .QN(_08324_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08048_ ), .Q(\mtvec [11] ), .QN(_08325_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08048_ ), .Q(\mtvec [10] ), .QN(_08326_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08048_ ), .Q(\mtvec [9] ), .QN(_08327_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08048_ ), .Q(\mtvec [8] ), .QN(_08328_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08048_ ), .Q(\mtvec [7] ), .QN(_08329_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08048_ ), .Q(\mtvec [6] ), .QN(_08330_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08048_ ), .Q(\mtvec [5] ), .QN(_08331_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08048_ ), .Q(\mtvec [4] ), .QN(_08332_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08048_ ), .Q(\mtvec [3] ), .QN(_08333_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08048_ ), .Q(\mtvec [2] ), .QN(_08334_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08048_ ), .Q(\mtvec [28] ), .QN(_08335_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08048_ ), .Q(\mtvec [1] ), .QN(_08336_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08048_ ), .Q(\mtvec [0] ), .QN(_08337_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08048_ ), .Q(\mtvec [27] ), .QN(_08338_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08048_ ), .Q(\mtvec [26] ), .QN(_08339_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08048_ ), .Q(\mtvec [25] ), .QN(_08340_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08048_ ), .Q(\mtvec [24] ), .QN(_08341_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08048_ ), .Q(\mtvec [23] ), .QN(_08342_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08048_ ), .Q(\mtvec [22] ), .QN(_08343_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_08047_ ), .Q(\mepc [31] ), .QN(_08344_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_08047_ ), .Q(\mepc [30] ), .QN(_08345_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_08047_ ), .Q(\mepc [21] ), .QN(_08346_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_08047_ ), .Q(\mepc [20] ), .QN(_08347_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_08047_ ), .Q(\mepc [19] ), .QN(_08348_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_08047_ ), .Q(\mepc [18] ), .QN(_08349_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_08047_ ), .Q(\mepc [17] ), .QN(_08350_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_08047_ ), .Q(\mepc [16] ), .QN(_08351_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_08047_ ), .Q(\mepc [15] ), .QN(_08352_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_08047_ ), .Q(\mepc [14] ), .QN(_08353_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_08047_ ), .Q(\mepc [13] ), .QN(_08354_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_08047_ ), .Q(\mepc [12] ), .QN(_08355_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_08047_ ), .Q(\mepc [29] ), .QN(_08356_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_08047_ ), .Q(\mepc [11] ), .QN(_08357_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_08047_ ), .Q(\mepc [10] ), .QN(_08358_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_08047_ ), .Q(\mepc [9] ), .QN(_08359_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_08047_ ), .Q(\mepc [8] ), .QN(_08360_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_08047_ ), .Q(\mepc [7] ), .QN(_08361_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_08047_ ), .Q(\mepc [6] ), .QN(_08362_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_08047_ ), .Q(\mepc [5] ), .QN(_08363_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_08047_ ), .Q(\mepc [4] ), .QN(_08364_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_08047_ ), .Q(\mepc [3] ), .QN(_08365_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_08047_ ), .Q(\mepc [2] ), .QN(_08366_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_08047_ ), .Q(\mepc [28] ), .QN(_08367_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_08047_ ), .Q(\mepc [1] ), .QN(_08368_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_08047_ ), .Q(\mepc [0] ), .QN(_08369_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_08047_ ), .Q(\mepc [27] ), .QN(_08370_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_08047_ ), .Q(\mepc [26] ), .QN(_08371_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_08047_ ), .Q(\mepc [25] ), .QN(_08372_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_08047_ ), .Q(\mepc [24] ), .QN(_08373_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_08047_ ), .Q(\mepc [23] ), .QN(_08374_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_08047_ ), .Q(\mepc [22] ), .QN(_08375_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08376_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08377_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08378_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08279_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08278_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08277_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08276_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08275_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08274_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08273_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08272_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08271_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08270_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08269_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08268_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08267_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08266_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08265_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08264_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08263_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08262_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08261_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08260_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08259_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08258_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00086_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08257_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00087_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08256_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00088_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08255_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00089_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08254_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00090_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08253_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00091_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08252_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00092_ ), .CK(_08046_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08251_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFFE_PP0P__Q ( .D(\mylsu.wen_reg_$_ANDNOT__A_Y_$_NAND__A_B ), .CK(_08045_ ), .Q(excp_written ), .QN(_08379_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08380_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08381_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08382_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08383_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08384_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08385_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08386_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08387_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08388_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08389_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08390_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08391_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08392_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08393_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08394_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08395_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08396_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08397_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08398_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08399_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08400_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08401_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08402_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08403_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08404_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08405_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08406_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08407_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08408_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08409_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08410_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08044_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08250_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00093_ ), .CK(_08043_ ), .Q(\myec.state [1] ), .QN(_08249_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00094_ ), .CK(_08043_ ), .Q(\myec.state [0] ), .QN(_08411_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PN0__Q ( .D(_00095_ ), .CK(clock ), .Q(check_quest ), .QN(_08412_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08248_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08413_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08414_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08415_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08416_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08417_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08418_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08419_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08420_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08421_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08422_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08247_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00096_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08246_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00097_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08245_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00098_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08244_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00099_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08243_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00100_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08242_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00101_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08241_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00102_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08240_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00103_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08239_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00104_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08238_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00105_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08237_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00106_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08236_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00107_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08235_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00108_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08234_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00109_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08233_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00110_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08232_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00111_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08231_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00112_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08230_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00113_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08229_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00114_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08228_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00115_ ), .CK(_08042_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08227_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q ( .D(_00116_ ), .CK(_08041_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08226_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_1 ( .D(_00117_ ), .CK(_08041_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08225_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_2 ( .D(_00118_ ), .CK(_08041_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08224_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_3 ( .D(_00119_ ), .CK(_08041_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08223_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_4 ( .D(_00120_ ), .CK(_08041_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08222_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q ( .D(_00121_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [30] ), .QN(_08221_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_1 ( .D(_00122_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [29] ), .QN(_08220_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_10 ( .D(_00123_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [20] ), .QN(_08219_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_11 ( .D(_00124_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [19] ), .QN(_08218_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_12 ( .D(_00125_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [18] ), .QN(_08217_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_13 ( .D(_00126_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [17] ), .QN(_08216_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_14 ( .D(_00127_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [16] ), .QN(_08215_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_15 ( .D(_00128_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [15] ), .QN(_08214_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_16 ( .D(_00129_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [14] ), .QN(_08213_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_17 ( .D(_00130_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [13] ), .QN(_08212_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_18 ( .D(_00131_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [12] ), .QN(_08211_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_19 ( .D(_00132_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [11] ), .QN(_08210_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_2 ( .D(_00133_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [28] ), .QN(_08209_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_20 ( .D(_00134_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [10] ), .QN(_08208_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_21 ( .D(_00135_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [9] ), .QN(_08207_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_22 ( .D(_00136_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [8] ), .QN(_08206_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_23 ( .D(_00137_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [7] ), .QN(_08205_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_24 ( .D(_00138_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [6] ), .QN(_08204_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_25 ( .D(_00139_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [5] ), .QN(_08203_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_26 ( .D(_00140_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [4] ), .QN(_08202_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_27 ( .D(_00141_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [3] ), .QN(_08201_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_28 ( .D(_00142_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [2] ), .QN(_08200_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_29 ( .D(_00143_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [1] ), .QN(_08199_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_3 ( .D(_00144_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [27] ), .QN(_08198_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_30 ( .D(_00145_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [0] ), .QN(_08197_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_4 ( .D(_00146_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [26] ), .QN(_08196_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_5 ( .D(_00147_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [25] ), .QN(_08195_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_6 ( .D(_00148_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [24] ), .QN(_08194_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_7 ( .D(_00149_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [23] ), .QN(_08193_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_8 ( .D(_00150_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [22] ), .QN(_08192_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_9 ( .D(_00151_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [21] ), .QN(_08191_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN1P__Q ( .D(_00152_ ), .CK(_08040_ ), .Q(\myexu.pc_jump [31] ), .QN(_08190_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q ( .D(_00153_ ), .CK(_08041_ ), .Q(\EX_LS_pc [31] ), .QN(_08189_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_1 ( .D(_00154_ ), .CK(_08041_ ), .Q(\EX_LS_pc [30] ), .QN(_08188_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_10 ( .D(_00155_ ), .CK(_08041_ ), .Q(\EX_LS_pc [21] ), .QN(_08187_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_11 ( .D(_00156_ ), .CK(_08041_ ), .Q(\EX_LS_pc [20] ), .QN(_08186_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_12 ( .D(_00157_ ), .CK(_08041_ ), .Q(\EX_LS_pc [19] ), .QN(_08185_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_13 ( .D(_00158_ ), .CK(_08041_ ), .Q(\EX_LS_pc [18] ), .QN(_08184_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_14 ( .D(_00159_ ), .CK(_08041_ ), .Q(\EX_LS_pc [17] ), .QN(_08183_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_15 ( .D(_00160_ ), .CK(_08041_ ), .Q(\EX_LS_pc [16] ), .QN(_08182_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_16 ( .D(_00161_ ), .CK(_08041_ ), .Q(\EX_LS_pc [15] ), .QN(_08181_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_17 ( .D(_00162_ ), .CK(_08041_ ), .Q(\EX_LS_pc [14] ), .QN(_08180_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_18 ( .D(_00163_ ), .CK(_08041_ ), .Q(\EX_LS_pc [13] ), .QN(_08179_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_19 ( .D(_00164_ ), .CK(_08041_ ), .Q(\EX_LS_pc [12] ), .QN(_08178_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_2 ( .D(_00165_ ), .CK(_08041_ ), .Q(\EX_LS_pc [29] ), .QN(_08177_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_20 ( .D(_00166_ ), .CK(_08041_ ), .Q(\EX_LS_pc [11] ), .QN(_08176_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_21 ( .D(_00167_ ), .CK(_08041_ ), .Q(\EX_LS_pc [10] ), .QN(_08175_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_22 ( .D(_00168_ ), .CK(_08041_ ), .Q(\EX_LS_pc [9] ), .QN(_08174_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_23 ( .D(_00169_ ), .CK(_08041_ ), .Q(\EX_LS_pc [8] ), .QN(_08173_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_24 ( .D(_00170_ ), .CK(_08041_ ), .Q(\EX_LS_pc [7] ), .QN(_08172_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_25 ( .D(_00171_ ), .CK(_08041_ ), .Q(\EX_LS_pc [6] ), .QN(_08171_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_26 ( .D(_00172_ ), .CK(_08041_ ), .Q(\EX_LS_pc [5] ), .QN(_08170_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_27 ( .D(_00173_ ), .CK(_08041_ ), .Q(\EX_LS_pc [4] ), .QN(_08169_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_28 ( .D(_00174_ ), .CK(_08041_ ), .Q(\EX_LS_pc [3] ), .QN(_08168_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_29 ( .D(_00175_ ), .CK(_08041_ ), .Q(\EX_LS_pc [2] ), .QN(_08167_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_3 ( .D(_00176_ ), .CK(_08041_ ), .Q(\EX_LS_pc [28] ), .QN(_08166_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_30 ( .D(_00177_ ), .CK(_08041_ ), .Q(\EX_LS_pc [1] ), .QN(_08165_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_31 ( .D(_00178_ ), .CK(_08041_ ), .Q(\EX_LS_pc [0] ), .QN(_08164_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_4 ( .D(_00179_ ), .CK(_08041_ ), .Q(\EX_LS_pc [27] ), .QN(_08163_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_5 ( .D(_00180_ ), .CK(_08041_ ), .Q(\EX_LS_pc [26] ), .QN(_08162_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_6 ( .D(_00181_ ), .CK(_08041_ ), .Q(\EX_LS_pc [25] ), .QN(_08161_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_7 ( .D(_00182_ ), .CK(_08041_ ), .Q(\EX_LS_pc [24] ), .QN(_08160_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_8 ( .D(_00183_ ), .CK(_08041_ ), .Q(\EX_LS_pc [23] ), .QN(_08159_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_9 ( .D(_00184_ ), .CK(_08041_ ), .Q(\EX_LS_pc [22] ), .QN(_08423_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08424_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08425_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08426_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08427_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08428_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08429_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08430_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08431_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08432_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08433_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08434_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08435_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08436_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08437_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08438_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08439_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08440_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08441_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08442_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08443_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08444_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08445_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08446_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08447_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08448_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08449_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08450_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08451_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08452_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08453_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08454_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08042_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08455_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08042_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PN0__Q ( .D(_00186_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q ( .D(_00185_ ), .CK(_08041_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_1 ( .D(_00187_ ), .CK(_08041_ ), .Q(\EX_LS_flag [1] ), .QN(_08158_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_2 ( .D(_00188_ ), .CK(_08041_ ), .Q(\EX_LS_flag [0] ), .QN(_08157_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_3 ( .D(_00189_ ), .CK(_08041_ ), .Q(\EX_LS_typ [4] ), .QN(_08156_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_4 ( .D(_00190_ ), .CK(_08041_ ), .Q(\EX_LS_typ [3] ), .QN(_08155_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_5 ( .D(_00191_ ), .CK(_08041_ ), .Q(\EX_LS_typ [2] ), .QN(_08154_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_6 ( .D(_00192_ ), .CK(_08041_ ), .Q(\EX_LS_typ [1] ), .QN(_08153_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_7 ( .D(_00193_ ), .CK(_08041_ ), .Q(\EX_LS_typ [0] ), .QN(_08152_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00194_ ), .CK(_08039_ ), .Q(\ID_EX_csr [11] ), .QN(_08151_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00195_ ), .CK(_08039_ ), .Q(\ID_EX_csr [10] ), .QN(_08150_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00196_ ), .CK(_08039_ ), .Q(\ID_EX_csr [1] ), .QN(_08149_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00197_ ), .CK(_08039_ ), .Q(\ID_EX_csr [0] ), .QN(_08148_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00198_ ), .CK(_08039_ ), .Q(\ID_EX_csr [9] ), .QN(_08147_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00199_ ), .CK(_08039_ ), .Q(\ID_EX_csr [8] ), .QN(_08146_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00200_ ), .CK(_08039_ ), .Q(\ID_EX_csr [7] ), .QN(_08145_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00201_ ), .CK(_08039_ ), .Q(\ID_EX_csr [6] ), .QN(_08144_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00202_ ), .CK(_08039_ ), .Q(\ID_EX_csr [5] ), .QN(_08143_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00203_ ), .CK(_08039_ ), .Q(\ID_EX_csr [4] ), .QN(_08142_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00204_ ), .CK(_08039_ ), .Q(\ID_EX_csr [3] ), .QN(_08141_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00205_ ), .CK(_08039_ ), .Q(\ID_EX_csr [2] ), .QN(_08140_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00206_ ), .CK(_08038_ ), .Q(exception_quest_IDU ), .QN(_08139_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00207_ ), .CK(_08037_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08036_ ), .Q(\ID_EX_imm [31] ), .QN(_08456_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08036_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08036_ ), .Q(\ID_EX_imm [21] ), .QN(_08457_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08036_ ), .Q(\ID_EX_imm [20] ), .QN(_08458_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08036_ ), .Q(\ID_EX_imm [19] ), .QN(_08459_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08036_ ), .Q(\ID_EX_imm [18] ), .QN(_08460_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08036_ ), .Q(\ID_EX_imm [17] ), .QN(_08461_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08036_ ), .Q(\ID_EX_imm [16] ), .QN(_08462_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08036_ ), .Q(\ID_EX_imm [15] ), .QN(_08463_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08036_ ), .Q(\ID_EX_imm [14] ), .QN(_08464_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08036_ ), .Q(\ID_EX_imm [13] ), .QN(_08465_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08036_ ), .Q(\ID_EX_imm [12] ), .QN(_08466_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08036_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08036_ ), .Q(\ID_EX_imm [11] ), .QN(_08467_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08036_ ), .Q(\ID_EX_imm [10] ), .QN(_08468_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08036_ ), .Q(\ID_EX_imm [9] ), .QN(_08469_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08036_ ), .Q(\ID_EX_imm [8] ), .QN(_08470_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08036_ ), .Q(\ID_EX_imm [7] ), .QN(_08471_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08036_ ), .Q(\ID_EX_imm [6] ), .QN(_08472_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08036_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08036_ ), .Q(\ID_EX_imm [4] ), .QN(_08473_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08036_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08036_ ), .Q(\ID_EX_imm [2] ), .QN(_08474_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08036_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08036_ ), .Q(\ID_EX_imm [1] ), .QN(_08475_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08036_ ), .Q(\ID_EX_imm [0] ), .QN(_08476_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08036_ ), .Q(\ID_EX_imm [27] ), .QN(_08477_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08036_ ), .Q(\ID_EX_imm [26] ), .QN(_08478_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08036_ ), .Q(\ID_EX_imm [25] ), .QN(_08479_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08036_ ), .Q(\ID_EX_imm [24] ), .QN(_08480_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08036_ ), .Q(\ID_EX_imm [23] ), .QN(_08481_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08036_ ), .Q(\ID_EX_imm [22] ), .QN(_08482_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08035_ ), .Q(\ID_EX_pc [31] ), .QN(_08483_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08035_ ), .Q(\ID_EX_pc [30] ), .QN(_08484_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08035_ ), .Q(\ID_EX_pc [21] ), .QN(_08485_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08035_ ), .Q(\ID_EX_pc [20] ), .QN(_08486_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08035_ ), .Q(\ID_EX_pc [19] ), .QN(_08487_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08035_ ), .Q(\ID_EX_pc [18] ), .QN(_08488_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08035_ ), .Q(\ID_EX_pc [17] ), .QN(_08489_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08035_ ), .Q(\ID_EX_pc [16] ), .QN(_08490_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08035_ ), .Q(\ID_EX_pc [15] ), .QN(_08491_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08035_ ), .Q(\ID_EX_pc [14] ), .QN(_08492_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08035_ ), .Q(\ID_EX_pc [13] ), .QN(_08493_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08035_ ), .Q(\ID_EX_pc [12] ), .QN(_08494_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08035_ ), .Q(\ID_EX_pc [29] ), .QN(_08495_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08035_ ), .Q(\ID_EX_pc [11] ), .QN(_08496_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08035_ ), .Q(\ID_EX_pc [10] ), .QN(_08497_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08035_ ), .Q(\ID_EX_pc [9] ), .QN(_08498_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08035_ ), .Q(\ID_EX_pc [8] ), .QN(_08499_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08035_ ), .Q(\ID_EX_pc [7] ), .QN(_08500_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08035_ ), .Q(\ID_EX_pc [6] ), .QN(_08501_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08035_ ), .Q(\ID_EX_pc [5] ), .QN(_08502_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08035_ ), .Q(\ID_EX_pc [4] ), .QN(_08503_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08035_ ), .Q(\ID_EX_pc [3] ), .QN(_08504_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08035_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08035_ ), .Q(\ID_EX_pc [28] ), .QN(_08505_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08035_ ), .Q(\ID_EX_pc [1] ), .QN(_08506_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08035_ ), .Q(\ID_EX_pc [0] ), .QN(_08507_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08035_ ), .Q(\ID_EX_pc [27] ), .QN(_08508_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08035_ ), .Q(\ID_EX_pc [26] ), .QN(_08509_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08035_ ), .Q(\ID_EX_pc [25] ), .QN(_08510_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08035_ ), .Q(\ID_EX_pc [24] ), .QN(_08511_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08035_ ), .Q(\ID_EX_pc [23] ), .QN(_08512_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08035_ ), .Q(\ID_EX_pc [22] ), .QN(_08138_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00208_ ), .CK(_08034_ ), .Q(\ID_EX_rd [4] ), .QN(_08137_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00209_ ), .CK(_08034_ ), .Q(\ID_EX_rd [3] ), .QN(_08136_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00210_ ), .CK(_08034_ ), .Q(\ID_EX_rd [2] ), .QN(_08135_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00211_ ), .CK(_08034_ ), .Q(\ID_EX_rd [1] ), .QN(_08134_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00212_ ), .CK(_08034_ ), .Q(\ID_EX_rd [0] ), .QN(_08133_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00213_ ), .CK(_08033_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08132_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00214_ ), .CK(_08033_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08131_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00216_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08129_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00215_ ), .CK(_08033_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08130_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00218_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08127_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00217_ ), .CK(_08033_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08128_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00220_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08125_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00219_ ), .CK(_08033_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08126_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00222_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08123_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00221_ ), .CK(_08032_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08124_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00223_ ), .CK(_08032_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08122_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00225_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08120_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00224_ ), .CK(_08032_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08121_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00227_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08118_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00226_ ), .CK(_08032_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08119_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00229_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08116_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00228_ ), .CK(_08032_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08117_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00231_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08114_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00230_ ), .CK(_08031_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08115_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00232_ ), .CK(_08030_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08113_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08514_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00233_ ), .CK(_08029_ ), .Q(\ID_EX_typ [7] ), .QN(_08513_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00234_ ), .CK(_08029_ ), .Q(\ID_EX_typ [6] ), .QN(_08112_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00235_ ), .CK(_08029_ ), .Q(\ID_EX_typ [5] ), .QN(_08111_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00236_ ), .CK(_08029_ ), .Q(\ID_EX_typ [4] ), .QN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00237_ ), .CK(_08029_ ), .Q(\ID_EX_typ [3] ), .QN(_08110_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00238_ ), .CK(_08029_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00239_ ), .CK(_08029_ ), .Q(\ID_EX_typ [1] ), .QN(_08109_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00240_ ), .CK(_08029_ ), .Q(\ID_EX_typ [0] ), .QN(_08515_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08028_ ), .Q(check_assert ), .QN(_08516_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08027_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08027_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08027_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08027_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08027_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08027_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08027_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08027_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08027_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08027_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08027_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08027_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08027_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08027_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08027_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08027_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08027_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08027_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08027_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08027_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08027_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08027_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08027_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08027_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08027_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08027_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08027_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08027_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08027_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08027_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08027_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08027_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08517_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08518_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08519_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08520_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08521_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08522_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08523_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08524_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08525_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08526_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08527_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08528_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08529_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08530_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08531_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08532_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08533_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08534_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08535_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08536_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08537_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08538_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08539_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08540_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08541_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08542_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08543_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08544_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08545_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08546_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08547_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08026_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08548_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08549_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08550_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08551_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08552_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08553_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08554_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08555_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08556_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08557_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08558_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08559_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08560_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08561_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08562_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08563_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08564_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08565_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08566_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08567_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08025_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08024_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08023_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08022_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08021_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08020_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08019_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08018_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08017_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08016_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08855_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08856_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08857_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08858_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08859_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08860_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08861_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08862_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08863_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08864_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08865_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08866_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08867_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08868_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08869_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08870_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08871_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08872_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08873_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08874_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08875_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08876_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08877_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08878_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08879_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08015_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08108_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00241_ ), .CK(_08014_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08107_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00242_ ), .CK(_08013_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08106_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00243_ ), .CK(_08012_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08880_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_08011_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08105_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00244_ ), .CK(_08010_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00245_ ), .CK(_08009_ ), .Q(\IF_ID_pc [30] ), .QN(_08104_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00246_ ), .CK(_08009_ ), .Q(\IF_ID_pc [21] ), .QN(_08103_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00247_ ), .CK(_08009_ ), .Q(\IF_ID_pc [20] ), .QN(_08102_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00248_ ), .CK(_08009_ ), .Q(\IF_ID_pc [19] ), .QN(_08101_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00249_ ), .CK(_08009_ ), .Q(\IF_ID_pc [18] ), .QN(_08100_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00250_ ), .CK(_08009_ ), .Q(\IF_ID_pc [17] ), .QN(_08099_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00251_ ), .CK(_08009_ ), .Q(\IF_ID_pc [16] ), .QN(_08098_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00252_ ), .CK(_08009_ ), .Q(\IF_ID_pc [15] ), .QN(_08097_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00253_ ), .CK(_08009_ ), .Q(\IF_ID_pc [14] ), .QN(_08096_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00254_ ), .CK(_08009_ ), .Q(\IF_ID_pc [13] ), .QN(_08095_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00255_ ), .CK(_08009_ ), .Q(\IF_ID_pc [12] ), .QN(_08094_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00256_ ), .CK(_08009_ ), .Q(\IF_ID_pc [29] ), .QN(_08093_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00257_ ), .CK(_08009_ ), .Q(\IF_ID_pc [11] ), .QN(_08092_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00258_ ), .CK(_08009_ ), .Q(\IF_ID_pc [10] ), .QN(_08091_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00259_ ), .CK(_08009_ ), .Q(\IF_ID_pc [9] ), .QN(_08090_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00260_ ), .CK(_08009_ ), .Q(\IF_ID_pc [8] ), .QN(_08089_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00261_ ), .CK(_08009_ ), .Q(\IF_ID_pc [7] ), .QN(_08088_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00262_ ), .CK(_08009_ ), .Q(\IF_ID_pc [6] ), .QN(_08087_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00263_ ), .CK(_08009_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00264_ ), .CK(_08009_ ), .Q(\IF_ID_pc [4] ), .QN(_08086_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00266_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08085_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00265_ ), .CK(_08009_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00268_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08083_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00267_ ), .CK(_08009_ ), .Q(\IF_ID_pc [2] ), .QN(_08084_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00269_ ), .CK(_08009_ ), .Q(\IF_ID_pc [28] ), .QN(_08082_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00270_ ), .CK(_08009_ ), .Q(\IF_ID_pc [1] ), .QN(_08081_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00271_ ), .CK(_08009_ ), .Q(\IF_ID_pc [27] ), .QN(_08080_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00272_ ), .CK(_08009_ ), .Q(\IF_ID_pc [26] ), .QN(_08079_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00273_ ), .CK(_08009_ ), .Q(\IF_ID_pc [25] ), .QN(_08078_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00274_ ), .CK(_08009_ ), .Q(\IF_ID_pc [24] ), .QN(_08077_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00275_ ), .CK(_08009_ ), .Q(\IF_ID_pc [23] ), .QN(_08076_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00276_ ), .CK(_08009_ ), .Q(\IF_ID_pc [22] ), .QN(_08075_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00277_ ), .CK(_08009_ ), .Q(\IF_ID_pc [31] ), .QN(_08074_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08882_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08073_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00278_ ), .CK(_08008_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08881_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00280_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00279_ ), .CK(_08007_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08072_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08883_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08884_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08885_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08886_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08887_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08888_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08889_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08890_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08891_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08892_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08893_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08894_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08895_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08896_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08897_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08898_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08899_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08900_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08901_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08902_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08903_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08904_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08905_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08906_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08907_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08908_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08909_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08910_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08911_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08912_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08913_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08006_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08914_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08915_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08916_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08917_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08918_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08919_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08920_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08921_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08922_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08923_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08924_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08925_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08926_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08927_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08928_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08929_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08930_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08931_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08932_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08933_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08934_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08935_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08936_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08937_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08938_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08939_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08940_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08941_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08942_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08943_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08944_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08945_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08005_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08071_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PN0P__Q ( .D(_00281_ ), .CK(_08004_ ), .Q(LS_WB_pc ), .QN(_08070_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PN0P__Q ( .D(_00282_ ), .CK(_08003_ ), .Q(\mylsu.previous_load_done ), .QN(_08946_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08947_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08948_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08949_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_08006_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_08006_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08950_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_08006_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08069_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00283_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08068_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00284_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08067_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00285_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08066_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00286_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08065_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00287_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08064_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00288_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08063_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00289_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08062_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00290_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08061_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00291_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08060_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00292_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08059_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00293_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08058_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00294_ ), .CK(_08006_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08951_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_08006_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08952_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_08006_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08953_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_08006_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08954_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_08006_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08955_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08956_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08957_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08958_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08959_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08960_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08961_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08962_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08963_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08964_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08965_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08966_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08967_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08968_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08969_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08970_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08971_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08972_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08973_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08974_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08975_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08976_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08977_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08978_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08979_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08980_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08981_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08982_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08983_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08984_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08985_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08986_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_08006_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08987_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08988_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_08989_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_08990_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_08991_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_08992_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_08993_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_08994_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_08995_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_08996_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_08997_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_08998_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_08999_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_09000_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_09001_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_09002_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_09003_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_09004_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_09005_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_09006_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_09007_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_09008_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_09009_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_09010_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_09011_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_09012_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_09013_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_09014_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_09015_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_09016_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_09017_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_09018_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_08002_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08057_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q ( .D(_00295_ ), .CK(_08001_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_08056_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_1 ( .D(_00296_ ), .CK(_08001_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08055_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_2 ( .D(_00297_ ), .CK(_08001_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08054_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_3 ( .D(_00298_ ), .CK(_08001_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08053_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_4 ( .D(_00299_ ), .CK(_08001_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08052_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_5 ( .D(_00300_ ), .CK(_08001_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08051_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PN0P__Q ( .D(_00301_ ), .CK(_08001_ ), .Q(LS_WB_wen_reg ), .QN(_09019_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_09020_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_09021_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_08000_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07999_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07998_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07997_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07996_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07995_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07994_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07993_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07992_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07991_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07990_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07989_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07988_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07987_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07986_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_1_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_10_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_11_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_12_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_13_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_14_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_15_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_16_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_17_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_18_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_19_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_2_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_20_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_21_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_22_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_23_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_24_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_25_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_26_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_27_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_28_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_29_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_3_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_30_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_31_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_4_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_5_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_6_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_7_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_8_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[3]_$_DFFE_PP__Q_9_D ), .CK(_07985_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00302_ ), .CK(_07984_ ), .Q(loaduse_clear ), .QN(_09022_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_09023_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_09024_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08050_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\ID_EX_typ [2] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_41 ) );

endmodule
