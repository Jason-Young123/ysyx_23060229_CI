//Generate the verilog at 2025-09-29T16:33:38 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire _09036_ ;
wire _09037_ ;
wire _09038_ ;
wire _09039_ ;
wire _09040_ ;
wire _09041_ ;
wire _09042_ ;
wire _09043_ ;
wire _09044_ ;
wire _09045_ ;
wire _09046_ ;
wire _09047_ ;
wire _09048_ ;
wire _09049_ ;
wire _09050_ ;
wire _09051_ ;
wire _09052_ ;
wire _09053_ ;
wire _09054_ ;
wire _09055_ ;
wire _09056_ ;
wire _09057_ ;
wire _09058_ ;
wire _09059_ ;
wire _09060_ ;
wire _09061_ ;
wire _09062_ ;
wire _09063_ ;
wire _09064_ ;
wire _09065_ ;
wire _09066_ ;
wire _09067_ ;
wire _09068_ ;
wire _09069_ ;
wire _09070_ ;
wire _09071_ ;
wire _09072_ ;
wire _09073_ ;
wire _09074_ ;
wire _09075_ ;
wire _09076_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.excp_written_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_NOR__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_B_$_MUX__Y_A_$_NOR__B_Y ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[5]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire fanout_net_45 ;
wire fanout_net_46 ;
wire fanout_net_47 ;
wire fanout_net_48 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

INV_X1 _09077_ ( .A(\LS_WB_wdata_csreg [31] ), .ZN(_01633_ ) );
NOR2_X1 _09078_ ( .A1(_01633_ ), .A2(fanout_net_1 ), .ZN(_00000_ ) );
INV_X2 _09079_ ( .A(fanout_net_1 ), .ZN(_01634_ ) );
BUF_X4 _09080_ ( .A(_01634_ ), .Z(_01635_ ) );
AND3_X4 _09081_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01636_ ) );
AND3_X4 _09082_ ( .A1(_01636_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01637_ ) );
AND3_X4 _09083_ ( .A1(_01637_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01638_ ) );
AND3_X4 _09084_ ( .A1(_01638_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01639_ ) );
AND3_X4 _09085_ ( .A1(_01639_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01640_ ) );
AND3_X4 _09086_ ( .A1(_01640_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01641_ ) );
AND3_X4 _09087_ ( .A1(_01641_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01642_ ) );
AND3_X4 _09088_ ( .A1(_01642_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01643_ ) );
AND3_X4 _09089_ ( .A1(_01643_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01644_ ) );
AND3_X4 _09090_ ( .A1(_01644_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01645_ ) );
AND3_X4 _09091_ ( .A1(_01645_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01646_ ) );
AND3_X4 _09092_ ( .A1(_01646_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01647_ ) );
AND3_X4 _09093_ ( .A1(_01647_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01648_ ) );
AND2_X4 _09094_ ( .A1(_01648_ ), .A2(\myclint.mtime [27] ), .ZN(_01649_ ) );
AND2_X1 _09095_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01650_ ) );
AND2_X1 _09096_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01651_ ) );
AND4_X2 _09097_ ( .A1(\myclint.mtime [33] ), .A2(_01649_ ), .A3(_01650_ ), .A4(_01651_ ), .ZN(_01652_ ) );
AND3_X4 _09098_ ( .A1(_01652_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01653_ ) );
AND3_X4 _09099_ ( .A1(_01653_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [35] ), .ZN(_01654_ ) );
AND2_X2 _09100_ ( .A1(_01654_ ), .A2(\myclint.mtime [37] ), .ZN(_01655_ ) );
AND2_X1 _09101_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [39] ), .ZN(_01656_ ) );
AND2_X1 _09102_ ( .A1(_01655_ ), .A2(_01656_ ), .ZN(_01657_ ) );
AND2_X1 _09103_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_01658_ ) );
AND2_X2 _09104_ ( .A1(_01657_ ), .A2(_01658_ ), .ZN(_01659_ ) );
AND2_X2 _09105_ ( .A1(\myclint.mtime [42] ), .A2(\myclint.mtime [43] ), .ZN(_01660_ ) );
AND2_X2 _09106_ ( .A1(_01659_ ), .A2(_01660_ ), .ZN(_01661_ ) );
AND2_X1 _09107_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01662_ ) );
AND3_X1 _09108_ ( .A1(_01662_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01663_ ) );
NAND2_X1 _09109_ ( .A1(_01661_ ), .A2(_01663_ ), .ZN(_01664_ ) );
AND2_X1 _09110_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01665_ ) );
INV_X1 _09111_ ( .A(_01665_ ), .ZN(_01666_ ) );
NOR2_X1 _09112_ ( .A1(_01664_ ), .A2(_01666_ ), .ZN(_01667_ ) );
AND2_X1 _09113_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01668_ ) );
AND2_X1 _09114_ ( .A1(_01667_ ), .A2(_01668_ ), .ZN(_01669_ ) );
AND2_X1 _09115_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01670_ ) );
AND2_X2 _09116_ ( .A1(_01669_ ), .A2(_01670_ ), .ZN(_01671_ ) );
AND2_X1 _09117_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01672_ ) );
NAND2_X2 _09118_ ( .A1(_01671_ ), .A2(_01672_ ), .ZN(_01673_ ) );
AND2_X1 _09119_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01674_ ) );
INV_X1 _09120_ ( .A(_01674_ ), .ZN(_01675_ ) );
NOR2_X2 _09121_ ( .A1(_01673_ ), .A2(_01675_ ), .ZN(_01676_ ) );
AND2_X1 _09122_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01677_ ) );
AND2_X1 _09123_ ( .A1(_01676_ ), .A2(_01677_ ), .ZN(_01678_ ) );
NAND3_X1 _09124_ ( .A1(_01678_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01679_ ) );
NOR2_X1 _09125_ ( .A1(_01679_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01680_ ) );
OAI21_X1 _09126_ ( .A(_01635_ ), .B1(_01680_ ), .B2(\myclint.mtime [63] ), .ZN(_01681_ ) );
AND3_X4 _09127_ ( .A1(_01648_ ), .A2(\myclint.mtime [28] ), .A3(\myclint.mtime [27] ), .ZN(_01682_ ) );
AND2_X4 _09128_ ( .A1(_01682_ ), .A2(\myclint.mtime [29] ), .ZN(_01683_ ) );
AND2_X1 _09129_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01684_ ) );
AND3_X4 _09130_ ( .A1(_01683_ ), .A2(_01684_ ), .A3(_01650_ ), .ZN(_01685_ ) );
AND3_X4 _09131_ ( .A1(_01685_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01686_ ) );
AND2_X4 _09132_ ( .A1(_01686_ ), .A2(\myclint.mtime [36] ), .ZN(_01687_ ) );
AND2_X4 _09133_ ( .A1(_01687_ ), .A2(\myclint.mtime [37] ), .ZN(_01688_ ) );
AND2_X1 _09134_ ( .A1(_01688_ ), .A2(_01656_ ), .ZN(_01689_ ) );
AND2_X2 _09135_ ( .A1(_01689_ ), .A2(_01658_ ), .ZN(_01690_ ) );
AND2_X2 _09136_ ( .A1(_01690_ ), .A2(_01660_ ), .ZN(_01691_ ) );
AND2_X2 _09137_ ( .A1(_01691_ ), .A2(_01663_ ), .ZN(_01692_ ) );
AND2_X2 _09138_ ( .A1(_01692_ ), .A2(_01665_ ), .ZN(_01693_ ) );
AND2_X1 _09139_ ( .A1(_01693_ ), .A2(_01668_ ), .ZN(_01694_ ) );
AND2_X2 _09140_ ( .A1(_01694_ ), .A2(_01670_ ), .ZN(_01695_ ) );
AND2_X2 _09141_ ( .A1(_01695_ ), .A2(_01672_ ), .ZN(_01696_ ) );
AND2_X2 _09142_ ( .A1(_01696_ ), .A2(_01674_ ), .ZN(_01697_ ) );
AND2_X2 _09143_ ( .A1(_01697_ ), .A2(_01677_ ), .ZN(_01698_ ) );
NAND3_X1 _09144_ ( .A1(_01698_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01699_ ) );
NOR2_X1 _09145_ ( .A1(_01699_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01700_ ) );
AOI21_X1 _09146_ ( .A(_01681_ ), .B1(_01700_ ), .B2(\myclint.mtime [63] ), .ZN(_00001_ ) );
AND2_X1 _09147_ ( .A1(_01638_ ), .A2(\myclint.mtime [7] ), .ZN(_01701_ ) );
AND4_X1 _09148_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01702_ ) );
AND2_X1 _09149_ ( .A1(\myclint.mtime [10] ), .A2(\myclint.mtime [11] ), .ZN(_01703_ ) );
AND4_X1 _09150_ ( .A1(\myclint.mtime [8] ), .A2(_01702_ ), .A3(\myclint.mtime [9] ), .A4(_01703_ ), .ZN(_01704_ ) );
AND2_X1 _09151_ ( .A1(_01701_ ), .A2(_01704_ ), .ZN(_01705_ ) );
AND2_X1 _09152_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_01706_ ) );
AND3_X1 _09153_ ( .A1(_01706_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01707_ ) );
AND4_X1 _09154_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01708_ ) );
AND2_X1 _09155_ ( .A1(_01707_ ), .A2(_01708_ ), .ZN(_01709_ ) );
AND2_X1 _09156_ ( .A1(\myclint.mtime [26] ), .A2(\myclint.mtime [27] ), .ZN(_01710_ ) );
AND3_X1 _09157_ ( .A1(_01710_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_01711_ ) );
AND4_X1 _09158_ ( .A1(_01650_ ), .A2(_01709_ ), .A3(_01651_ ), .A4(_01711_ ), .ZN(_01712_ ) );
AND2_X2 _09159_ ( .A1(_01705_ ), .A2(_01712_ ), .ZN(_01713_ ) );
AND3_X1 _09160_ ( .A1(_01684_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01714_ ) );
AND2_X1 _09161_ ( .A1(_01660_ ), .A2(_01658_ ), .ZN(_01715_ ) );
AND4_X1 _09162_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01716_ ) );
AND4_X1 _09163_ ( .A1(_01663_ ), .A2(_01714_ ), .A3(_01715_ ), .A4(_01716_ ), .ZN(_01717_ ) );
AND2_X1 _09164_ ( .A1(_01713_ ), .A2(_01717_ ), .ZN(_01718_ ) );
AND4_X1 _09165_ ( .A1(_01672_ ), .A2(_01670_ ), .A3(_01668_ ), .A4(_01665_ ), .ZN(_01719_ ) );
AND2_X1 _09166_ ( .A1(_01718_ ), .A2(_01719_ ), .ZN(_01720_ ) );
AND4_X1 _09167_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01721_ ) );
AND2_X1 _09168_ ( .A1(_01720_ ), .A2(_01721_ ), .ZN(_01722_ ) );
AND3_X1 _09169_ ( .A1(_01722_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01723_ ) );
XNOR2_X1 _09170_ ( .A(_01723_ ), .B(\myclint.mtime [62] ), .ZN(_01724_ ) );
NOR2_X1 _09171_ ( .A1(_01724_ ), .A2(fanout_net_1 ), .ZN(_00002_ ) );
INV_X1 _09172_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01725_ ) );
AND3_X1 _09173_ ( .A1(_01667_ ), .A2(_01725_ ), .A3(_01668_ ), .ZN(_01726_ ) );
OAI21_X1 _09174_ ( .A(_01635_ ), .B1(_01726_ ), .B2(\myclint.mtime [53] ), .ZN(_01727_ ) );
AND3_X1 _09175_ ( .A1(_01693_ ), .A2(_01725_ ), .A3(_01668_ ), .ZN(_01728_ ) );
AOI21_X1 _09176_ ( .A(_01727_ ), .B1(_01728_ ), .B2(\myclint.mtime [53] ), .ZN(_00003_ ) );
AND2_X1 _09177_ ( .A1(_01668_ ), .A2(_01665_ ), .ZN(_01729_ ) );
AND2_X1 _09178_ ( .A1(_01718_ ), .A2(_01729_ ), .ZN(_01730_ ) );
XNOR2_X1 _09179_ ( .A(_01730_ ), .B(\myclint.mtime [52] ), .ZN(_01731_ ) );
NOR2_X1 _09180_ ( .A1(_01731_ ), .A2(fanout_net_1 ), .ZN(_00004_ ) );
NOR3_X1 _09181_ ( .A1(_01664_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01666_ ), .ZN(_01732_ ) );
OAI21_X1 _09182_ ( .A(_01635_ ), .B1(_01732_ ), .B2(\myclint.mtime [51] ), .ZN(_01733_ ) );
INV_X1 _09183_ ( .A(_01692_ ), .ZN(_01734_ ) );
NOR3_X1 _09184_ ( .A1(_01734_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01666_ ), .ZN(_01735_ ) );
AOI21_X1 _09185_ ( .A(_01733_ ), .B1(_01735_ ), .B2(\myclint.mtime [51] ), .ZN(_00005_ ) );
INV_X1 _09186_ ( .A(_01713_ ), .ZN(_01736_ ) );
INV_X1 _09187_ ( .A(_01717_ ), .ZN(_01737_ ) );
OR4_X1 _09188_ ( .A1(\myclint.mtime [50] ), .A2(_01736_ ), .A3(_01666_ ), .A4(_01737_ ), .ZN(_01738_ ) );
AND3_X1 _09189_ ( .A1(_01713_ ), .A2(_01665_ ), .A3(_01717_ ), .ZN(_01739_ ) );
INV_X1 _09190_ ( .A(_01739_ ), .ZN(_01740_ ) );
NAND2_X1 _09191_ ( .A1(_01740_ ), .A2(\myclint.mtime [50] ), .ZN(_01741_ ) );
AOI21_X1 _09192_ ( .A(fanout_net_1 ), .B1(_01738_ ), .B2(_01741_ ), .ZN(_00006_ ) );
INV_X1 _09193_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01742_ ) );
AND4_X1 _09194_ ( .A1(\myclint.mtime [49] ), .A2(_01691_ ), .A3(_01742_ ), .A4(_01663_ ), .ZN(_01743_ ) );
BUF_X4 _09195_ ( .A(_01634_ ), .Z(_01744_ ) );
AND3_X1 _09196_ ( .A1(_01661_ ), .A2(_01742_ ), .A3(_01663_ ), .ZN(_01745_ ) );
OAI21_X1 _09197_ ( .A(_01744_ ), .B1(_01745_ ), .B2(\myclint.mtime [49] ), .ZN(_01746_ ) );
NOR2_X1 _09198_ ( .A1(_01743_ ), .A2(_01746_ ), .ZN(_00007_ ) );
INV_X1 _09199_ ( .A(_01705_ ), .ZN(_01747_ ) );
INV_X1 _09200_ ( .A(_01712_ ), .ZN(_01748_ ) );
OR4_X1 _09201_ ( .A1(\myclint.mtime [48] ), .A2(_01747_ ), .A3(_01748_ ), .A4(_01737_ ), .ZN(_01749_ ) );
OAI21_X1 _09202_ ( .A(\myclint.mtime [48] ), .B1(_01736_ ), .B2(_01737_ ), .ZN(_01750_ ) );
AOI21_X1 _09203_ ( .A(fanout_net_1 ), .B1(_01749_ ), .B2(_01750_ ), .ZN(_00008_ ) );
NAND3_X1 _09204_ ( .A1(_01659_ ), .A2(_01662_ ), .A3(_01660_ ), .ZN(_01751_ ) );
NOR2_X1 _09205_ ( .A1(_01751_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01752_ ) );
OAI21_X1 _09206_ ( .A(_01635_ ), .B1(_01752_ ), .B2(\myclint.mtime [47] ), .ZN(_01753_ ) );
NAND3_X1 _09207_ ( .A1(_01690_ ), .A2(\myclint.mtime [44] ), .A3(_01660_ ), .ZN(_01754_ ) );
INV_X1 _09208_ ( .A(\myclint.mtime [45] ), .ZN(_01755_ ) );
NOR3_X1 _09209_ ( .A1(_01754_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01755_ ), .ZN(_01756_ ) );
AOI21_X1 _09210_ ( .A(_01753_ ), .B1(_01756_ ), .B2(\myclint.mtime [47] ), .ZN(_00009_ ) );
AND2_X1 _09211_ ( .A1(_01714_ ), .A2(_01716_ ), .ZN(_01757_ ) );
AND2_X1 _09212_ ( .A1(_01713_ ), .A2(_01757_ ), .ZN(_01758_ ) );
AND3_X1 _09213_ ( .A1(_01758_ ), .A2(_01662_ ), .A3(_01715_ ), .ZN(_01759_ ) );
XNOR2_X1 _09214_ ( .A(_01759_ ), .B(\myclint.mtime [46] ), .ZN(_01760_ ) );
NOR2_X1 _09215_ ( .A1(_01760_ ), .A2(fanout_net_1 ), .ZN(_00010_ ) );
INV_X1 _09216_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01761_ ) );
NAND3_X1 _09217_ ( .A1(_01659_ ), .A2(_01761_ ), .A3(_01660_ ), .ZN(_01762_ ) );
AOI21_X1 _09218_ ( .A(fanout_net_1 ), .B1(_01762_ ), .B2(_01755_ ), .ZN(_01763_ ) );
NAND4_X1 _09219_ ( .A1(_01690_ ), .A2(\myclint.mtime [45] ), .A3(_01761_ ), .A4(_01660_ ), .ZN(_01764_ ) );
AND2_X1 _09220_ ( .A1(_01763_ ), .A2(_01764_ ), .ZN(_00011_ ) );
AND2_X1 _09221_ ( .A1(_01758_ ), .A2(_01715_ ), .ZN(_01765_ ) );
XNOR2_X1 _09222_ ( .A(_01765_ ), .B(\myclint.mtime [44] ), .ZN(_01766_ ) );
NOR2_X1 _09223_ ( .A1(_01766_ ), .A2(fanout_net_1 ), .ZN(_00012_ ) );
INV_X1 _09224_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01767_ ) );
AND3_X1 _09225_ ( .A1(_01676_ ), .A2(_01767_ ), .A3(_01677_ ), .ZN(_01768_ ) );
OAI21_X1 _09226_ ( .A(_01635_ ), .B1(_01768_ ), .B2(\myclint.mtime [61] ), .ZN(_01769_ ) );
AND3_X1 _09227_ ( .A1(_01697_ ), .A2(_01767_ ), .A3(_01677_ ), .ZN(_01770_ ) );
AOI21_X1 _09228_ ( .A(_01769_ ), .B1(_01770_ ), .B2(\myclint.mtime [61] ), .ZN(_00013_ ) );
NAND3_X1 _09229_ ( .A1(_01713_ ), .A2(_01658_ ), .A3(_01757_ ), .ZN(_01771_ ) );
OR3_X1 _09230_ ( .A1(_01771_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [43] ), .ZN(_01772_ ) );
OAI21_X1 _09231_ ( .A(\myclint.mtime [43] ), .B1(_01771_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01773_ ) );
AOI21_X1 _09232_ ( .A(fanout_net_1 ), .B1(_01772_ ), .B2(_01773_ ), .ZN(_00014_ ) );
OR2_X1 _09233_ ( .A1(_01771_ ), .A2(\myclint.mtime [42] ), .ZN(_01774_ ) );
NAND2_X1 _09234_ ( .A1(_01771_ ), .A2(\myclint.mtime [42] ), .ZN(_01775_ ) );
AOI21_X1 _09235_ ( .A(fanout_net_1 ), .B1(_01774_ ), .B2(_01775_ ), .ZN(_00015_ ) );
INV_X1 _09236_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01776_ ) );
AND4_X1 _09237_ ( .A1(\myclint.mtime [41] ), .A2(_01688_ ), .A3(_01776_ ), .A4(_01656_ ), .ZN(_01777_ ) );
AND3_X1 _09238_ ( .A1(_01655_ ), .A2(_01776_ ), .A3(_01656_ ), .ZN(_01778_ ) );
OAI21_X1 _09239_ ( .A(_01744_ ), .B1(_01778_ ), .B2(\myclint.mtime [41] ), .ZN(_01779_ ) );
NOR2_X1 _09240_ ( .A1(_01777_ ), .A2(_01779_ ), .ZN(_00016_ ) );
XNOR2_X1 _09241_ ( .A(_01758_ ), .B(\myclint.mtime [40] ), .ZN(_01780_ ) );
NOR2_X1 _09242_ ( .A1(_01780_ ), .A2(fanout_net_1 ), .ZN(_00017_ ) );
INV_X1 _09243_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01781_ ) );
AND4_X1 _09244_ ( .A1(_01781_ ), .A2(_01687_ ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01782_ ) );
AND3_X1 _09245_ ( .A1(_01654_ ), .A2(_01781_ ), .A3(\myclint.mtime [37] ), .ZN(_01783_ ) );
OAI21_X1 _09246_ ( .A(_01744_ ), .B1(_01783_ ), .B2(\myclint.mtime [39] ), .ZN(_01784_ ) );
NOR2_X1 _09247_ ( .A1(_01782_ ), .A2(_01784_ ), .ZN(_00018_ ) );
AND2_X1 _09248_ ( .A1(_01713_ ), .A2(_01714_ ), .ZN(_01785_ ) );
AND3_X1 _09249_ ( .A1(_01785_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .ZN(_01786_ ) );
XNOR2_X1 _09250_ ( .A(_01786_ ), .B(\myclint.mtime [38] ), .ZN(_01787_ ) );
NOR2_X1 _09251_ ( .A1(_01787_ ), .A2(fanout_net_1 ), .ZN(_00019_ ) );
NAND3_X1 _09252_ ( .A1(_01652_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01788_ ) );
INV_X1 _09253_ ( .A(\myclint.mtime [35] ), .ZN(_01789_ ) );
NOR3_X1 _09254_ ( .A1(_01788_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01789_ ), .ZN(_01790_ ) );
OAI21_X1 _09255_ ( .A(_01635_ ), .B1(_01790_ ), .B2(\myclint.mtime [37] ), .ZN(_01791_ ) );
NAND2_X1 _09256_ ( .A1(_01685_ ), .A2(\myclint.mtime [34] ), .ZN(_01792_ ) );
NOR3_X1 _09257_ ( .A1(_01792_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01789_ ), .ZN(_01793_ ) );
AOI21_X1 _09258_ ( .A(_01791_ ), .B1(\myclint.mtime [37] ), .B2(_01793_ ), .ZN(_00020_ ) );
BUF_X2 _09259_ ( .A(_01634_ ), .Z(_01794_ ) );
NOR2_X1 _09260_ ( .A1(_01788_ ), .A2(_01789_ ), .ZN(_01795_ ) );
OAI21_X1 _09261_ ( .A(_01794_ ), .B1(_01795_ ), .B2(\myclint.mtime [36] ), .ZN(_01796_ ) );
NOR2_X1 _09262_ ( .A1(_01796_ ), .A2(_01654_ ), .ZN(_00021_ ) );
NAND3_X1 _09263_ ( .A1(_01705_ ), .A2(_01684_ ), .A3(_01712_ ), .ZN(_01797_ ) );
NOR2_X1 _09264_ ( .A1(_01797_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01798_ ) );
XNOR2_X1 _09265_ ( .A(_01798_ ), .B(\myclint.mtime [35] ), .ZN(_01799_ ) );
NOR2_X1 _09266_ ( .A1(_01799_ ), .A2(fanout_net_1 ), .ZN(_00022_ ) );
BUF_X4 _09267_ ( .A(_01634_ ), .Z(_01800_ ) );
OAI21_X1 _09268_ ( .A(_01800_ ), .B1(_01685_ ), .B2(\myclint.mtime [34] ), .ZN(_01801_ ) );
NOR2_X1 _09269_ ( .A1(_01801_ ), .A2(_01653_ ), .ZN(_00023_ ) );
XNOR2_X1 _09270_ ( .A(_01722_ ), .B(\myclint.mtime [60] ), .ZN(_01802_ ) );
NOR2_X1 _09271_ ( .A1(_01802_ ), .A2(fanout_net_1 ), .ZN(_00024_ ) );
AND2_X1 _09272_ ( .A1(_01649_ ), .A2(_01651_ ), .ZN(_01803_ ) );
INV_X1 _09273_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01804_ ) );
AND3_X1 _09274_ ( .A1(_01803_ ), .A2(_01804_ ), .A3(_01650_ ), .ZN(_01805_ ) );
OAI21_X1 _09275_ ( .A(_01800_ ), .B1(_01805_ ), .B2(\myclint.mtime [33] ), .ZN(_01806_ ) );
AND4_X1 _09276_ ( .A1(_01804_ ), .A2(_01683_ ), .A3(\myclint.mtime [33] ), .A4(_01650_ ), .ZN(_01807_ ) );
NOR2_X1 _09277_ ( .A1(_01806_ ), .A2(_01807_ ), .ZN(_00025_ ) );
XNOR2_X1 _09278_ ( .A(_01713_ ), .B(\myclint.mtime [32] ), .ZN(_01808_ ) );
NOR2_X1 _09279_ ( .A1(_01808_ ), .A2(fanout_net_1 ), .ZN(_00026_ ) );
AND2_X1 _09280_ ( .A1(_01705_ ), .A2(_01709_ ), .ZN(_01809_ ) );
NAND3_X1 _09281_ ( .A1(_01809_ ), .A2(_01651_ ), .A3(_01711_ ), .ZN(_01810_ ) );
NOR2_X1 _09282_ ( .A1(_01810_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01811_ ) );
XNOR2_X1 _09283_ ( .A(_01811_ ), .B(\myclint.mtime [31] ), .ZN(_01812_ ) );
NOR2_X1 _09284_ ( .A1(_01812_ ), .A2(fanout_net_1 ), .ZN(_00027_ ) );
OR2_X1 _09285_ ( .A1(_01810_ ), .A2(\myclint.mtime [30] ), .ZN(_01813_ ) );
NAND2_X1 _09286_ ( .A1(_01810_ ), .A2(\myclint.mtime [30] ), .ZN(_01814_ ) );
AOI21_X1 _09287_ ( .A(fanout_net_1 ), .B1(_01813_ ), .B2(_01814_ ), .ZN(_00028_ ) );
INV_X1 _09288_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01815_ ) );
AND3_X1 _09289_ ( .A1(_01648_ ), .A2(_01815_ ), .A3(\myclint.mtime [27] ), .ZN(_01816_ ) );
AND2_X1 _09290_ ( .A1(_01816_ ), .A2(\myclint.mtime [29] ), .ZN(_01817_ ) );
OAI21_X1 _09291_ ( .A(_01744_ ), .B1(_01816_ ), .B2(\myclint.mtime [29] ), .ZN(_01818_ ) );
NOR2_X1 _09292_ ( .A1(_01817_ ), .A2(_01818_ ), .ZN(_00029_ ) );
NAND2_X1 _09293_ ( .A1(_01809_ ), .A2(_01711_ ), .ZN(_01819_ ) );
XNOR2_X1 _09294_ ( .A(_01819_ ), .B(\myclint.mtime [28] ), .ZN(_01820_ ) );
AND2_X1 _09295_ ( .A1(_01820_ ), .A2(_01794_ ), .ZN(_00030_ ) );
NAND3_X1 _09296_ ( .A1(_01809_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_01821_ ) );
OR3_X1 _09297_ ( .A1(_01821_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01822_ ) );
OAI21_X1 _09298_ ( .A(\myclint.mtime [27] ), .B1(_01821_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01823_ ) );
AOI21_X1 _09299_ ( .A(fanout_net_1 ), .B1(_01822_ ), .B2(_01823_ ), .ZN(_00031_ ) );
AND2_X1 _09300_ ( .A1(_01647_ ), .A2(\myclint.mtime [25] ), .ZN(_01824_ ) );
OAI21_X1 _09301_ ( .A(_01800_ ), .B1(_01824_ ), .B2(\myclint.mtime [26] ), .ZN(_01825_ ) );
NOR2_X1 _09302_ ( .A1(_01825_ ), .A2(_01648_ ), .ZN(_00032_ ) );
INV_X1 _09303_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01826_ ) );
AND3_X1 _09304_ ( .A1(_01646_ ), .A2(_01826_ ), .A3(\myclint.mtime [23] ), .ZN(_01827_ ) );
AND2_X1 _09305_ ( .A1(_01827_ ), .A2(\myclint.mtime [25] ), .ZN(_01828_ ) );
OAI21_X1 _09306_ ( .A(_01744_ ), .B1(_01827_ ), .B2(\myclint.mtime [25] ), .ZN(_01829_ ) );
NOR2_X1 _09307_ ( .A1(_01828_ ), .A2(_01829_ ), .ZN(_00033_ ) );
AND2_X1 _09308_ ( .A1(_01646_ ), .A2(\myclint.mtime [23] ), .ZN(_01830_ ) );
OAI21_X1 _09309_ ( .A(_01800_ ), .B1(_01830_ ), .B2(\myclint.mtime [24] ), .ZN(_01831_ ) );
NOR2_X1 _09310_ ( .A1(_01831_ ), .A2(_01647_ ), .ZN(_00034_ ) );
NOR3_X1 _09311_ ( .A1(_01673_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01675_ ), .ZN(_01832_ ) );
OAI21_X1 _09312_ ( .A(_01635_ ), .B1(_01832_ ), .B2(\myclint.mtime [59] ), .ZN(_01833_ ) );
INV_X1 _09313_ ( .A(_01696_ ), .ZN(_01834_ ) );
NOR3_X1 _09314_ ( .A1(_01834_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01675_ ), .ZN(_01835_ ) );
AOI21_X1 _09315_ ( .A(_01833_ ), .B1(_01835_ ), .B2(\myclint.mtime [59] ), .ZN(_00035_ ) );
AND2_X1 _09316_ ( .A1(_01705_ ), .A2(_01707_ ), .ZN(_01836_ ) );
NAND3_X1 _09317_ ( .A1(_01836_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01837_ ) );
OR3_X1 _09318_ ( .A1(_01837_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01838_ ) );
OAI21_X1 _09319_ ( .A(\myclint.mtime [23] ), .B1(_01837_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01839_ ) );
AOI21_X1 _09320_ ( .A(fanout_net_1 ), .B1(_01838_ ), .B2(_01839_ ), .ZN(_00036_ ) );
AND2_X1 _09321_ ( .A1(_01645_ ), .A2(\myclint.mtime [21] ), .ZN(_01840_ ) );
OAI21_X1 _09322_ ( .A(_01800_ ), .B1(_01840_ ), .B2(\myclint.mtime [22] ), .ZN(_01841_ ) );
NOR2_X1 _09323_ ( .A1(_01841_ ), .A2(_01646_ ), .ZN(_00037_ ) );
INV_X1 _09324_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01842_ ) );
AND3_X1 _09325_ ( .A1(_01644_ ), .A2(_01842_ ), .A3(\myclint.mtime [19] ), .ZN(_01843_ ) );
AND2_X1 _09326_ ( .A1(_01843_ ), .A2(\myclint.mtime [21] ), .ZN(_01844_ ) );
OAI21_X1 _09327_ ( .A(_01744_ ), .B1(_01843_ ), .B2(\myclint.mtime [21] ), .ZN(_01845_ ) );
NOR2_X1 _09328_ ( .A1(_01844_ ), .A2(_01845_ ), .ZN(_00038_ ) );
AND2_X1 _09329_ ( .A1(_01644_ ), .A2(\myclint.mtime [19] ), .ZN(_01846_ ) );
OAI21_X1 _09330_ ( .A(_01800_ ), .B1(_01846_ ), .B2(\myclint.mtime [20] ), .ZN(_01847_ ) );
NOR2_X1 _09331_ ( .A1(_01847_ ), .A2(_01645_ ), .ZN(_00039_ ) );
NAND3_X1 _09332_ ( .A1(_01705_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_01848_ ) );
OR3_X1 _09333_ ( .A1(_01848_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01849_ ) );
OAI21_X1 _09334_ ( .A(\myclint.mtime [19] ), .B1(_01848_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01850_ ) );
AOI21_X1 _09335_ ( .A(fanout_net_1 ), .B1(_01849_ ), .B2(_01850_ ), .ZN(_00040_ ) );
AND2_X1 _09336_ ( .A1(_01643_ ), .A2(\myclint.mtime [17] ), .ZN(_01851_ ) );
OAI21_X1 _09337_ ( .A(_01800_ ), .B1(_01851_ ), .B2(\myclint.mtime [18] ), .ZN(_01852_ ) );
NOR2_X1 _09338_ ( .A1(_01852_ ), .A2(_01644_ ), .ZN(_00041_ ) );
INV_X1 _09339_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01853_ ) );
AND3_X1 _09340_ ( .A1(_01642_ ), .A2(_01853_ ), .A3(\myclint.mtime [15] ), .ZN(_01854_ ) );
AND2_X1 _09341_ ( .A1(_01854_ ), .A2(\myclint.mtime [17] ), .ZN(_01855_ ) );
OAI21_X1 _09342_ ( .A(_01635_ ), .B1(_01854_ ), .B2(\myclint.mtime [17] ), .ZN(_01856_ ) );
NOR2_X1 _09343_ ( .A1(_01855_ ), .A2(_01856_ ), .ZN(_00042_ ) );
AND2_X1 _09344_ ( .A1(_01642_ ), .A2(\myclint.mtime [15] ), .ZN(_01857_ ) );
OAI21_X1 _09345_ ( .A(_01800_ ), .B1(_01857_ ), .B2(\myclint.mtime [16] ), .ZN(_01858_ ) );
NOR2_X1 _09346_ ( .A1(_01858_ ), .A2(_01643_ ), .ZN(_00043_ ) );
AND3_X1 _09347_ ( .A1(_01703_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01859_ ) );
AND2_X1 _09348_ ( .A1(_01701_ ), .A2(_01859_ ), .ZN(_01860_ ) );
NAND3_X1 _09349_ ( .A1(_01860_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01861_ ) );
OR3_X1 _09350_ ( .A1(_01861_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01862_ ) );
OAI21_X1 _09351_ ( .A(\myclint.mtime [15] ), .B1(_01861_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01863_ ) );
AOI21_X1 _09352_ ( .A(fanout_net_1 ), .B1(_01862_ ), .B2(_01863_ ), .ZN(_00044_ ) );
AND2_X1 _09353_ ( .A1(_01641_ ), .A2(\myclint.mtime [13] ), .ZN(_01864_ ) );
OAI21_X1 _09354_ ( .A(_01800_ ), .B1(_01864_ ), .B2(\myclint.mtime [14] ), .ZN(_01865_ ) );
NOR2_X1 _09355_ ( .A1(_01865_ ), .A2(_01642_ ), .ZN(_00045_ ) );
NAND3_X1 _09356_ ( .A1(_01718_ ), .A2(_01674_ ), .A3(_01719_ ), .ZN(_01866_ ) );
OR2_X1 _09357_ ( .A1(_01866_ ), .A2(\myclint.mtime [58] ), .ZN(_01867_ ) );
NAND2_X1 _09358_ ( .A1(_01866_ ), .A2(\myclint.mtime [58] ), .ZN(_01868_ ) );
AOI21_X1 _09359_ ( .A(fanout_net_1 ), .B1(_01867_ ), .B2(_01868_ ), .ZN(_00046_ ) );
INV_X1 _09360_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01869_ ) );
AND3_X1 _09361_ ( .A1(_01640_ ), .A2(_01869_ ), .A3(\myclint.mtime [11] ), .ZN(_01870_ ) );
AND2_X1 _09362_ ( .A1(_01870_ ), .A2(\myclint.mtime [13] ), .ZN(_01871_ ) );
OAI21_X1 _09363_ ( .A(_01635_ ), .B1(_01870_ ), .B2(\myclint.mtime [13] ), .ZN(_01872_ ) );
NOR2_X1 _09364_ ( .A1(_01871_ ), .A2(_01872_ ), .ZN(_00047_ ) );
AND2_X1 _09365_ ( .A1(_01640_ ), .A2(\myclint.mtime [11] ), .ZN(_01873_ ) );
OAI21_X1 _09366_ ( .A(_01800_ ), .B1(_01873_ ), .B2(\myclint.mtime [12] ), .ZN(_01874_ ) );
NOR2_X1 _09367_ ( .A1(_01874_ ), .A2(_01641_ ), .ZN(_00048_ ) );
NAND3_X1 _09368_ ( .A1(_01701_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_01875_ ) );
OR3_X1 _09369_ ( .A1(_01875_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_01876_ ) );
OAI21_X1 _09370_ ( .A(\myclint.mtime [11] ), .B1(_01875_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01877_ ) );
AOI21_X1 _09371_ ( .A(fanout_net_1 ), .B1(_01876_ ), .B2(_01877_ ), .ZN(_00049_ ) );
AND2_X1 _09372_ ( .A1(_01639_ ), .A2(\myclint.mtime [9] ), .ZN(_01878_ ) );
OAI21_X1 _09373_ ( .A(_01744_ ), .B1(_01878_ ), .B2(\myclint.mtime [10] ), .ZN(_01879_ ) );
NOR2_X1 _09374_ ( .A1(_01879_ ), .A2(_01640_ ), .ZN(_00050_ ) );
INV_X1 _09375_ ( .A(_01701_ ), .ZN(_01880_ ) );
OR3_X1 _09376_ ( .A1(_01880_ ), .A2(\myclint.mtime [9] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01881_ ) );
OAI21_X1 _09377_ ( .A(\myclint.mtime [9] ), .B1(_01880_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01882_ ) );
AOI21_X1 _09378_ ( .A(fanout_net_1 ), .B1(_01881_ ), .B2(_01882_ ), .ZN(_00051_ ) );
OAI21_X1 _09379_ ( .A(_01744_ ), .B1(_01701_ ), .B2(\myclint.mtime [8] ), .ZN(_01883_ ) );
NOR2_X1 _09380_ ( .A1(_01883_ ), .A2(_01639_ ), .ZN(_00052_ ) );
AND2_X1 _09381_ ( .A1(_01637_ ), .A2(\myclint.mtime [5] ), .ZN(_01884_ ) );
INV_X1 _09382_ ( .A(_01884_ ), .ZN(_01885_ ) );
OR3_X1 _09383_ ( .A1(_01885_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [7] ), .ZN(_01886_ ) );
OAI21_X1 _09384_ ( .A(\myclint.mtime [7] ), .B1(_01885_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01887_ ) );
AOI21_X1 _09385_ ( .A(fanout_net_1 ), .B1(_01886_ ), .B2(_01887_ ), .ZN(_00053_ ) );
OAI21_X1 _09386_ ( .A(_01744_ ), .B1(_01884_ ), .B2(\myclint.mtime [6] ), .ZN(_01888_ ) );
NOR2_X1 _09387_ ( .A1(_01888_ ), .A2(_01638_ ), .ZN(_00054_ ) );
AND2_X1 _09388_ ( .A1(_01636_ ), .A2(\myclint.mtime [3] ), .ZN(_01889_ ) );
INV_X1 _09389_ ( .A(_01889_ ), .ZN(_01890_ ) );
OR3_X1 _09390_ ( .A1(_01890_ ), .A2(\myclint.mtime [5] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01891_ ) );
OAI21_X1 _09391_ ( .A(\myclint.mtime [5] ), .B1(_01890_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01892_ ) );
AOI21_X1 _09392_ ( .A(fanout_net_1 ), .B1(_01891_ ), .B2(_01892_ ), .ZN(_00055_ ) );
OAI21_X1 _09393_ ( .A(_01744_ ), .B1(_01889_ ), .B2(\myclint.mtime [4] ), .ZN(_01893_ ) );
NOR2_X1 _09394_ ( .A1(_01893_ ), .A2(_01637_ ), .ZN(_00056_ ) );
INV_X1 _09395_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01894_ ) );
AND3_X1 _09396_ ( .A1(_01671_ ), .A2(_01894_ ), .A3(_01672_ ), .ZN(_01895_ ) );
OAI21_X1 _09397_ ( .A(_01635_ ), .B1(_01895_ ), .B2(\myclint.mtime [57] ), .ZN(_01896_ ) );
AND3_X1 _09398_ ( .A1(_01695_ ), .A2(_01894_ ), .A3(_01672_ ), .ZN(_01897_ ) );
AOI21_X1 _09399_ ( .A(_01896_ ), .B1(_01897_ ), .B2(\myclint.mtime [57] ), .ZN(_00057_ ) );
AND2_X1 _09400_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01898_ ) );
INV_X1 _09401_ ( .A(_01898_ ), .ZN(_01899_ ) );
OR3_X1 _09402_ ( .A1(_01899_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01900_ ) );
OAI21_X1 _09403_ ( .A(\myclint.mtime [3] ), .B1(_01899_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01901_ ) );
AOI21_X1 _09404_ ( .A(fanout_net_1 ), .B1(_01900_ ), .B2(_01901_ ), .ZN(_00058_ ) );
AOI21_X1 _09405_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01902_ ) );
NOR3_X1 _09406_ ( .A1(_01636_ ), .A2(_01902_ ), .A3(fanout_net_1 ), .ZN(_00059_ ) );
NOR2_X1 _09407_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01903_ ) );
NOR3_X1 _09408_ ( .A1(_01898_ ), .A2(_01903_ ), .A3(fanout_net_1 ), .ZN(_00060_ ) );
AND2_X1 _09409_ ( .A1(_01794_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_00061_ ) );
XNOR2_X1 _09410_ ( .A(_01720_ ), .B(\myclint.mtime [56] ), .ZN(_01904_ ) );
NOR2_X1 _09411_ ( .A1(_01904_ ), .A2(fanout_net_2 ), .ZN(_00062_ ) );
NAND3_X1 _09412_ ( .A1(_01718_ ), .A2(_01670_ ), .A3(_01729_ ), .ZN(_01905_ ) );
OR3_X1 _09413_ ( .A1(_01905_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01906_ ) );
OAI21_X1 _09414_ ( .A(\myclint.mtime [55] ), .B1(_01905_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01907_ ) );
AOI21_X1 _09415_ ( .A(fanout_net_2 ), .B1(_01906_ ), .B2(_01907_ ), .ZN(_00063_ ) );
OR2_X1 _09416_ ( .A1(_01905_ ), .A2(\myclint.mtime [54] ), .ZN(_01908_ ) );
NAND2_X1 _09417_ ( .A1(_01905_ ), .A2(\myclint.mtime [54] ), .ZN(_01909_ ) );
AOI21_X1 _09418_ ( .A(fanout_net_2 ), .B1(_01908_ ), .B2(_01909_ ), .ZN(_00064_ ) );
INV_X1 _09419_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01910_ ) );
MUX2_X1 _09420_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(fanout_net_47 ), .Z(_01911_ ) );
INV_X32 _09421_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01912_ ) );
BUF_X2 _09422_ ( .A(_01912_ ), .Z(_01913_ ) );
AND2_X1 _09423_ ( .A1(_01911_ ), .A2(_01913_ ), .ZN(_01914_ ) );
MUX2_X1 _09424_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(fanout_net_47 ), .Z(_01915_ ) );
AOI21_X1 _09425_ ( .A(_01914_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01915_ ), .ZN(_01916_ ) );
NOR2_X1 _09426_ ( .A1(_01916_ ), .A2(\IF_ID_pc [20] ), .ZN(_01917_ ) );
MUX2_X1 _09427_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(fanout_net_47 ), .Z(_01918_ ) );
AND2_X1 _09428_ ( .A1(_01918_ ), .A2(_01913_ ), .ZN(_01919_ ) );
MUX2_X1 _09429_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(fanout_net_47 ), .Z(_01920_ ) );
AOI21_X1 _09430_ ( .A(_01919_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01920_ ), .ZN(_01921_ ) );
AOI21_X1 _09431_ ( .A(_01917_ ), .B1(\IF_ID_pc [18] ), .B2(_01921_ ), .ZN(_01922_ ) );
MUX2_X1 _09432_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(fanout_net_47 ), .Z(_01923_ ) );
OR2_X1 _09433_ ( .A1(_01923_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01924_ ) );
MUX2_X1 _09434_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(fanout_net_47 ), .Z(_01925_ ) );
OAI21_X1 _09435_ ( .A(_01924_ ), .B1(_01913_ ), .B2(_01925_ ), .ZN(_01926_ ) );
INV_X1 _09436_ ( .A(\IF_ID_pc [27] ), .ZN(_01927_ ) );
MUX2_X1 _09437_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(fanout_net_47 ), .Z(_01928_ ) );
MUX2_X1 _09438_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(fanout_net_47 ), .Z(_01929_ ) );
MUX2_X1 _09439_ ( .A(_01928_ ), .B(_01929_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01930_ ) );
OAI221_X1 _09440_ ( .A(_01922_ ), .B1(\IF_ID_pc [29] ), .B2(_01926_ ), .C1(_01927_ ), .C2(_01930_ ), .ZN(_01931_ ) );
INV_X1 _09441_ ( .A(\IF_ID_pc [24] ), .ZN(_01932_ ) );
MUX2_X1 _09442_ ( .A(\myifu.myicache.tag[2][19] ), .B(\myifu.myicache.tag[3][19] ), .S(fanout_net_47 ), .Z(_01933_ ) );
BUF_X8 _09443_ ( .A(_01912_ ), .Z(_01934_ ) );
OR2_X2 _09444_ ( .A1(_01933_ ), .A2(_01934_ ), .ZN(_01935_ ) );
MUX2_X1 _09445_ ( .A(\myifu.myicache.tag[0][19] ), .B(\myifu.myicache.tag[1][19] ), .S(fanout_net_47 ), .Z(_01936_ ) );
OR2_X4 _09446_ ( .A1(_01936_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01937_ ) );
AOI21_X1 _09447_ ( .A(_01932_ ), .B1(_01935_ ), .B2(_01937_ ), .ZN(_01938_ ) );
INV_X1 _09448_ ( .A(\IF_ID_pc [23] ), .ZN(_01939_ ) );
MUX2_X1 _09449_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(fanout_net_47 ), .Z(_01940_ ) );
MUX2_X1 _09450_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(fanout_net_47 ), .Z(_01941_ ) );
MUX2_X1 _09451_ ( .A(_01940_ ), .B(_01941_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01942_ ) );
AOI21_X1 _09452_ ( .A(_01938_ ), .B1(_01939_ ), .B2(_01942_ ), .ZN(_01943_ ) );
INV_X1 _09453_ ( .A(\IF_ID_pc [16] ), .ZN(_01944_ ) );
MUX2_X1 _09454_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_47 ), .Z(_01945_ ) );
MUX2_X1 _09455_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_47 ), .Z(_01946_ ) );
MUX2_X1 _09456_ ( .A(_01945_ ), .B(_01946_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01947_ ) );
OAI221_X1 _09457_ ( .A(_01943_ ), .B1(\IF_ID_pc [18] ), .B2(_01921_ ), .C1(_01944_ ), .C2(_01947_ ), .ZN(_01948_ ) );
NAND2_X1 _09458_ ( .A1(_01930_ ), .A2(_01927_ ), .ZN(_01949_ ) );
INV_X32 _09459_ ( .A(fanout_net_47 ), .ZN(_01950_ ) );
BUF_X32 _09460_ ( .A(_01950_ ), .Z(_01951_ ) );
OR2_X4 _09461_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[1][3] ), .ZN(_01952_ ) );
OAI211_X1 _09462_ ( .A(_01952_ ), .B(_01913_ ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[0][3] ), .ZN(_01953_ ) );
OR2_X1 _09463_ ( .A1(fanout_net_47 ), .A2(\myifu.myicache.tag[2][3] ), .ZN(_01954_ ) );
BUF_X8 _09464_ ( .A(_01950_ ), .Z(_01955_ ) );
OAI211_X1 _09465_ ( .A(_01954_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01955_ ), .C2(\myifu.myicache.tag[3][3] ), .ZN(_01956_ ) );
NAND3_X1 _09466_ ( .A1(_01953_ ), .A2(\IF_ID_pc [8] ), .A3(_01956_ ), .ZN(_01957_ ) );
OR2_X1 _09467_ ( .A1(fanout_net_47 ), .A2(\myifu.myicache.tag[0][2] ), .ZN(_01958_ ) );
OAI211_X1 _09468_ ( .A(_01958_ ), .B(_01913_ ), .C1(_01955_ ), .C2(\myifu.myicache.tag[1][2] ), .ZN(_01959_ ) );
OR2_X1 _09469_ ( .A1(fanout_net_47 ), .A2(\myifu.myicache.tag[2][2] ), .ZN(_01960_ ) );
OAI211_X1 _09470_ ( .A(_01960_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01955_ ), .C2(\myifu.myicache.tag[3][2] ), .ZN(_01961_ ) );
INV_X1 _09471_ ( .A(\IF_ID_pc [7] ), .ZN(_01962_ ) );
AND3_X1 _09472_ ( .A1(_01959_ ), .A2(_01961_ ), .A3(_01962_ ), .ZN(_01963_ ) );
AOI21_X1 _09473_ ( .A(_01962_ ), .B1(_01959_ ), .B2(_01961_ ), .ZN(_01964_ ) );
OAI211_X1 _09474_ ( .A(_01949_ ), .B(_01957_ ), .C1(_01963_ ), .C2(_01964_ ), .ZN(_01965_ ) );
INV_X1 _09475_ ( .A(\IF_ID_pc [30] ), .ZN(_01966_ ) );
MUX2_X1 _09476_ ( .A(\myifu.myicache.tag[2][25] ), .B(\myifu.myicache.tag[3][25] ), .S(fanout_net_47 ), .Z(_01967_ ) );
OR2_X1 _09477_ ( .A1(_01967_ ), .A2(_01934_ ), .ZN(_01968_ ) );
MUX2_X1 _09478_ ( .A(\myifu.myicache.tag[0][25] ), .B(\myifu.myicache.tag[1][25] ), .S(fanout_net_47 ), .Z(_01969_ ) );
OR2_X1 _09479_ ( .A1(_01969_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01970_ ) );
AOI21_X1 _09480_ ( .A(_01966_ ), .B1(_01968_ ), .B2(_01970_ ), .ZN(_01971_ ) );
AND3_X1 _09481_ ( .A1(_01968_ ), .A2(_01970_ ), .A3(_01966_ ), .ZN(_01972_ ) );
AND3_X4 _09482_ ( .A1(_01935_ ), .A2(_01937_ ), .A3(_01932_ ), .ZN(_01973_ ) );
AOI21_X1 _09483_ ( .A(\IF_ID_pc [8] ), .B1(_01953_ ), .B2(_01956_ ), .ZN(_01974_ ) );
OR4_X4 _09484_ ( .A1(_01971_ ), .A2(_01972_ ), .A3(_01973_ ), .A4(_01974_ ), .ZN(_01975_ ) );
NOR4_X4 _09485_ ( .A1(_01931_ ), .A2(_01948_ ), .A3(_01965_ ), .A4(_01975_ ), .ZN(_01976_ ) );
OR2_X1 _09486_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[1][17] ), .ZN(_01977_ ) );
OAI211_X1 _09487_ ( .A(_01977_ ), .B(_01934_ ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[0][17] ), .ZN(_01978_ ) );
OR2_X1 _09488_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[3][17] ), .ZN(_01979_ ) );
OAI211_X1 _09489_ ( .A(_01979_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[2][17] ), .ZN(_01980_ ) );
NAND2_X1 _09490_ ( .A1(_01978_ ), .A2(_01980_ ), .ZN(_01981_ ) );
XOR2_X1 _09491_ ( .A(_01981_ ), .B(\IF_ID_pc [22] ), .Z(_01982_ ) );
OR2_X1 _09492_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[1][21] ), .ZN(_01983_ ) );
OAI211_X1 _09493_ ( .A(_01983_ ), .B(_01934_ ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[0][21] ), .ZN(_01984_ ) );
OR2_X1 _09494_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[3][21] ), .ZN(_01985_ ) );
OAI211_X1 _09495_ ( .A(_01985_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[2][21] ), .ZN(_01986_ ) );
INV_X1 _09496_ ( .A(\IF_ID_pc [26] ), .ZN(_01987_ ) );
AND3_X1 _09497_ ( .A1(_01984_ ), .A2(_01986_ ), .A3(_01987_ ), .ZN(_01988_ ) );
AOI21_X1 _09498_ ( .A(_01987_ ), .B1(_01984_ ), .B2(_01986_ ), .ZN(_01989_ ) );
OR2_X1 _09499_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[1][0] ), .ZN(_01990_ ) );
OAI211_X1 _09500_ ( .A(_01990_ ), .B(_01934_ ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[0][0] ), .ZN(_01991_ ) );
OR2_X1 _09501_ ( .A1(fanout_net_47 ), .A2(\myifu.myicache.tag[2][0] ), .ZN(_01992_ ) );
OAI211_X1 _09502_ ( .A(_01992_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01951_ ), .C2(\myifu.myicache.tag[3][0] ), .ZN(_01993_ ) );
AND3_X1 _09503_ ( .A1(_01991_ ), .A2(_01993_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01994_ ) );
AOI21_X1 _09504_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_01991_ ), .B2(_01993_ ), .ZN(_01995_ ) );
OAI22_X1 _09505_ ( .A1(_01988_ ), .A2(_01989_ ), .B1(_01994_ ), .B2(_01995_ ), .ZN(_01996_ ) );
OR2_X1 _09506_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[1][4] ), .ZN(_01997_ ) );
OAI211_X1 _09507_ ( .A(_01997_ ), .B(_01913_ ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[0][4] ), .ZN(_01998_ ) );
OR2_X1 _09508_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[3][4] ), .ZN(_01999_ ) );
OAI211_X1 _09509_ ( .A(_01999_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[2][4] ), .ZN(_02000_ ) );
AND3_X1 _09510_ ( .A1(_01998_ ), .A2(_02000_ ), .A3(\IF_ID_pc [9] ), .ZN(_02001_ ) );
AOI21_X1 _09511_ ( .A(\IF_ID_pc [9] ), .B1(_01998_ ), .B2(_02000_ ), .ZN(_02002_ ) );
OR4_X1 _09512_ ( .A1(_01982_ ), .A2(_01996_ ), .A3(_02001_ ), .A4(_02002_ ), .ZN(_02003_ ) );
OR2_X1 _09513_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_02004_ ) );
OAI211_X1 _09514_ ( .A(_02004_ ), .B(_01913_ ), .C1(fanout_net_47 ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_02005_ ) );
OR2_X1 _09515_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[3][12] ), .ZN(_02006_ ) );
OAI211_X1 _09516_ ( .A(_02006_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][12] ), .ZN(_02007_ ) );
NAND2_X1 _09517_ ( .A1(_02005_ ), .A2(_02007_ ), .ZN(_02008_ ) );
XNOR2_X1 _09518_ ( .A(_02008_ ), .B(\IF_ID_pc [17] ), .ZN(_02009_ ) );
MUX2_X1 _09519_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02010_ ) );
MUX2_X1 _09520_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02011_ ) );
MUX2_X1 _09521_ ( .A(_02010_ ), .B(_02011_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02012_ ) );
MUX2_X1 _09522_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02013_ ) );
MUX2_X1 _09523_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02014_ ) );
MUX2_X1 _09524_ ( .A(_02013_ ), .B(_02014_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02015_ ) );
INV_X1 _09525_ ( .A(\IF_ID_pc [14] ), .ZN(_02016_ ) );
NAND2_X1 _09526_ ( .A1(_02015_ ), .A2(_02016_ ), .ZN(_02017_ ) );
AND3_X1 _09527_ ( .A1(_02009_ ), .A2(_02012_ ), .A3(_02017_ ), .ZN(_02018_ ) );
MUX2_X1 _09528_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02019_ ) );
MUX2_X1 _09529_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02020_ ) );
MUX2_X1 _09530_ ( .A(_02019_ ), .B(_02020_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02021_ ) );
XNOR2_X1 _09531_ ( .A(_02021_ ), .B(\IF_ID_pc [10] ), .ZN(_02022_ ) );
INV_X1 _09532_ ( .A(\IF_ID_pc [12] ), .ZN(_02023_ ) );
MUX2_X1 _09533_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02024_ ) );
MUX2_X1 _09534_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02025_ ) );
MUX2_X1 _09535_ ( .A(_02024_ ), .B(_02025_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02026_ ) );
AOI22_X1 _09536_ ( .A1(_01916_ ), .A2(\IF_ID_pc [20] ), .B1(_02023_ ), .B2(_02026_ ), .ZN(_02027_ ) );
NAND3_X1 _09537_ ( .A1(_02018_ ), .A2(_02022_ ), .A3(_02027_ ), .ZN(_02028_ ) );
OR2_X1 _09538_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[1][1] ), .ZN(_02029_ ) );
OAI211_X1 _09539_ ( .A(_02029_ ), .B(_01934_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][1] ), .ZN(_02030_ ) );
OR2_X1 _09540_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][1] ), .ZN(_02031_ ) );
OAI211_X1 _09541_ ( .A(_02031_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01955_ ), .C2(\myifu.myicache.tag[3][1] ), .ZN(_02032_ ) );
INV_X1 _09542_ ( .A(\IF_ID_pc [6] ), .ZN(_02033_ ) );
AND3_X1 _09543_ ( .A1(_02030_ ), .A2(_02032_ ), .A3(_02033_ ), .ZN(_02034_ ) );
AOI21_X1 _09544_ ( .A(_02033_ ), .B1(_02030_ ), .B2(_02032_ ), .ZN(_02035_ ) );
OR2_X1 _09545_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[3][8] ), .ZN(_02036_ ) );
OAI211_X1 _09546_ ( .A(_02036_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][8] ), .ZN(_02037_ ) );
INV_X1 _09547_ ( .A(\IF_ID_pc [13] ), .ZN(_02038_ ) );
OR2_X1 _09548_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][8] ), .ZN(_02039_ ) );
OAI211_X1 _09549_ ( .A(_02039_ ), .B(_01934_ ), .C1(_01955_ ), .C2(\myifu.myicache.tag[1][8] ), .ZN(_02040_ ) );
AND3_X1 _09550_ ( .A1(_02037_ ), .A2(_02038_ ), .A3(_02040_ ), .ZN(_02041_ ) );
AOI21_X1 _09551_ ( .A(_02038_ ), .B1(_02037_ ), .B2(_02040_ ), .ZN(_02042_ ) );
OAI22_X1 _09552_ ( .A1(_02034_ ), .A2(_02035_ ), .B1(_02041_ ), .B2(_02042_ ), .ZN(_02043_ ) );
OR2_X1 _09553_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][10] ), .ZN(_02044_ ) );
OAI211_X1 _09554_ ( .A(_02044_ ), .B(_01934_ ), .C1(_01955_ ), .C2(\myifu.myicache.tag[1][10] ), .ZN(_02045_ ) );
OR2_X1 _09555_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][10] ), .ZN(_02046_ ) );
OAI211_X1 _09556_ ( .A(_02046_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01955_ ), .C2(\myifu.myicache.tag[3][10] ), .ZN(_02047_ ) );
NAND2_X1 _09557_ ( .A1(_02045_ ), .A2(_02047_ ), .ZN(_02048_ ) );
INV_X1 _09558_ ( .A(\IF_ID_pc [15] ), .ZN(_02049_ ) );
XNOR2_X1 _09559_ ( .A(_02048_ ), .B(_02049_ ), .ZN(_02050_ ) );
OR2_X1 _09560_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[1][26] ), .ZN(_02051_ ) );
OAI211_X1 _09561_ ( .A(_02051_ ), .B(_01913_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][26] ), .ZN(_02052_ ) );
OR2_X1 _09562_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[3][26] ), .ZN(_02053_ ) );
OAI211_X1 _09563_ ( .A(_02053_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][26] ), .ZN(_02054_ ) );
AOI21_X1 _09564_ ( .A(\IF_ID_pc [31] ), .B1(_02052_ ), .B2(_02054_ ), .ZN(_02055_ ) );
AND3_X1 _09565_ ( .A1(_02052_ ), .A2(_02054_ ), .A3(\IF_ID_pc [31] ), .ZN(_02056_ ) );
OR4_X1 _09566_ ( .A1(_02043_ ), .A2(_02050_ ), .A3(_02055_ ), .A4(_02056_ ), .ZN(_02057_ ) );
NOR3_X1 _09567_ ( .A1(_02003_ ), .A2(_02028_ ), .A3(_02057_ ), .ZN(_02058_ ) );
MUX2_X1 _09568_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02059_ ) );
MUX2_X1 _09569_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02060_ ) );
MUX2_X2 _09570_ ( .A(_02059_ ), .B(_02060_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02061_ ) );
INV_X1 _09571_ ( .A(\IF_ID_pc [21] ), .ZN(_02062_ ) );
NOR2_X1 _09572_ ( .A1(_02061_ ), .A2(_02062_ ), .ZN(_02063_ ) );
OR2_X1 _09573_ ( .A1(_01950_ ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_02064_ ) );
OAI211_X1 _09574_ ( .A(_02064_ ), .B(_01934_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_02065_ ) );
OR2_X1 _09575_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][6] ), .ZN(_02066_ ) );
OAI211_X1 _09576_ ( .A(_02066_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01955_ ), .C2(\myifu.myicache.tag[3][6] ), .ZN(_02067_ ) );
AOI21_X1 _09577_ ( .A(\IF_ID_pc [11] ), .B1(_02065_ ), .B2(_02067_ ), .ZN(_02068_ ) );
NOR2_X1 _09578_ ( .A1(_02063_ ), .A2(_02068_ ), .ZN(_02069_ ) );
MUX2_X1 _09579_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02070_ ) );
AND2_X1 _09580_ ( .A1(_02070_ ), .A2(_01913_ ), .ZN(_02071_ ) );
MUX2_X1 _09581_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02072_ ) );
AOI21_X1 _09582_ ( .A(_02071_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_02072_ ), .ZN(_02073_ ) );
OAI221_X1 _09583_ ( .A(_02069_ ), .B1(_01939_ ), .B2(_01942_ ), .C1(\IF_ID_pc [25] ), .C2(_02073_ ), .ZN(_02074_ ) );
AOI22_X1 _09584_ ( .A1(_02073_ ), .A2(\IF_ID_pc [25] ), .B1(_01944_ ), .B2(_01947_ ), .ZN(_02075_ ) );
NAND2_X1 _09585_ ( .A1(_01926_ ), .A2(\IF_ID_pc [29] ), .ZN(_02076_ ) );
OAI211_X1 _09586_ ( .A(_02075_ ), .B(_02076_ ), .C1(_02016_ ), .C2(_02015_ ), .ZN(_02077_ ) );
NOR2_X1 _09587_ ( .A1(_02026_ ), .A2(_02023_ ), .ZN(_02078_ ) );
OR2_X1 _09588_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][14] ), .ZN(_02079_ ) );
OAI211_X1 _09589_ ( .A(_02079_ ), .B(_01934_ ), .C1(_01955_ ), .C2(\myifu.myicache.tag[1][14] ), .ZN(_02080_ ) );
OR2_X1 _09590_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][14] ), .ZN(_02081_ ) );
OAI211_X1 _09591_ ( .A(_02081_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01955_ ), .C2(\myifu.myicache.tag[3][14] ), .ZN(_02082_ ) );
AND3_X1 _09592_ ( .A1(_02080_ ), .A2(_02082_ ), .A3(\IF_ID_pc [19] ), .ZN(_02083_ ) );
AND3_X1 _09593_ ( .A1(_02065_ ), .A2(_02067_ ), .A3(\IF_ID_pc [11] ), .ZN(_02084_ ) );
AOI21_X1 _09594_ ( .A(\IF_ID_pc [19] ), .B1(_02080_ ), .B2(_02082_ ), .ZN(_02085_ ) );
OR4_X1 _09595_ ( .A1(_02078_ ), .A2(_02083_ ), .A3(_02084_ ), .A4(_02085_ ), .ZN(_02086_ ) );
AND2_X2 _09596_ ( .A1(_02061_ ), .A2(_02062_ ), .ZN(_02087_ ) );
OR2_X1 _09597_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[1][23] ), .ZN(_02088_ ) );
OAI211_X1 _09598_ ( .A(_02088_ ), .B(_01913_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][23] ), .ZN(_02089_ ) );
OR2_X1 _09599_ ( .A1(_01951_ ), .A2(\myifu.myicache.tag[3][23] ), .ZN(_02090_ ) );
OAI211_X1 _09600_ ( .A(_02090_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][23] ), .ZN(_02091_ ) );
AOI21_X1 _09601_ ( .A(\IF_ID_pc [28] ), .B1(_02089_ ), .B2(_02091_ ), .ZN(_02092_ ) );
AND3_X1 _09602_ ( .A1(_02089_ ), .A2(_02091_ ), .A3(\IF_ID_pc [28] ), .ZN(_02093_ ) );
OR3_X1 _09603_ ( .A1(_02087_ ), .A2(_02092_ ), .A3(_02093_ ), .ZN(_02094_ ) );
NOR4_X1 _09604_ ( .A1(_02074_ ), .A2(_02077_ ), .A3(_02086_ ), .A4(_02094_ ), .ZN(_02095_ ) );
NAND3_X2 _09605_ ( .A1(_01976_ ), .A2(_02058_ ), .A3(_02095_ ), .ZN(_02096_ ) );
AND2_X4 _09606_ ( .A1(_02096_ ), .A2(\myifu.state [0] ), .ZN(_02097_ ) );
INV_X2 _09607_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_02098_ ) );
NOR2_X4 _09608_ ( .A1(_02097_ ), .A2(_02098_ ), .ZN(_02099_ ) );
NOR2_X1 _09609_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_02100_ ) );
NOR2_X4 _09610_ ( .A1(_02099_ ), .A2(_02100_ ), .ZN(_02101_ ) );
CLKBUF_X2 _09611_ ( .A(_02101_ ), .Z(_02102_ ) );
CLKBUF_X2 _09612_ ( .A(_02102_ ), .Z(_02103_ ) );
CLKBUF_X2 _09613_ ( .A(_02103_ ), .Z(_02104_ ) );
INV_X32 _09614_ ( .A(\EX_LS_flag [2] ), .ZN(_02105_ ) );
NAND4_X1 _09615_ ( .A1(_02105_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(\mylsu.state [0] ), .ZN(_02106_ ) );
INV_X1 _09616_ ( .A(EXU_valid_LSU ), .ZN(_02107_ ) );
NOR2_X1 _09617_ ( .A1(_02106_ ), .A2(_02107_ ), .ZN(_02108_ ) );
BUF_X4 _09618_ ( .A(_02108_ ), .Z(_02109_ ) );
BUF_X4 _09619_ ( .A(_02109_ ), .Z(_02110_ ) );
AND2_X1 _09620_ ( .A1(fanout_net_7 ), .A2(\EX_LS_typ [1] ), .ZN(_02111_ ) );
NOR2_X1 _09621_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02112_ ) );
NAND3_X1 _09622_ ( .A1(_02111_ ), .A2(_02112_ ), .A3(\EX_LS_typ [0] ), .ZN(_02113_ ) );
NOR2_X1 _09623_ ( .A1(fanout_net_7 ), .A2(\EX_LS_dest_csreg_mem [1] ), .ZN(_02114_ ) );
INV_X1 _09624_ ( .A(\EX_LS_typ [2] ), .ZN(_02115_ ) );
NOR4_X1 _09625_ ( .A1(_02114_ ), .A2(_02115_ ), .A3(\EX_LS_typ [1] ), .A4(\EX_LS_typ [3] ), .ZN(_02116_ ) );
AOI21_X1 _09626_ ( .A(_02116_ ), .B1(_02112_ ), .B2(_02111_ ), .ZN(_02117_ ) );
OAI21_X1 _09627_ ( .A(_02113_ ), .B1(_02117_ ), .B2(\EX_LS_typ [0] ), .ZN(_02118_ ) );
AND2_X4 _09628_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02119_ ) );
AND2_X4 _09629_ ( .A1(_02119_ ), .A2(_02105_ ), .ZN(_02120_ ) );
INV_X1 _09630_ ( .A(\EX_LS_typ [4] ), .ZN(_02121_ ) );
AND2_X1 _09631_ ( .A1(_02120_ ), .A2(_02121_ ), .ZN(_02122_ ) );
AND2_X1 _09632_ ( .A1(_02118_ ), .A2(_02122_ ), .ZN(_02123_ ) );
OR2_X1 _09633_ ( .A1(\EX_LS_dest_csreg_mem [26] ), .A2(\EX_LS_dest_csreg_mem [24] ), .ZN(_02124_ ) );
NOR3_X1 _09634_ ( .A1(_02124_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\EX_LS_dest_csreg_mem [25] ), .ZN(_02125_ ) );
NOR4_X1 _09635_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\EX_LS_dest_csreg_mem [29] ), .A4(\EX_LS_dest_csreg_mem [28] ), .ZN(_02126_ ) );
AND2_X1 _09636_ ( .A1(_02125_ ), .A2(_02126_ ), .ZN(_02127_ ) );
AND2_X1 _09637_ ( .A1(_02127_ ), .A2(_02120_ ), .ZN(_02128_ ) );
NOR2_X1 _09638_ ( .A1(_02123_ ), .A2(_02128_ ), .ZN(_02129_ ) );
INV_X32 _09639_ ( .A(\EX_LS_flag [1] ), .ZN(_02130_ ) );
NOR2_X4 _09640_ ( .A1(_02130_ ), .A2(\EX_LS_flag [0] ), .ZN(_02131_ ) );
AND2_X2 _09641_ ( .A1(_02131_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02132_ ) );
AND2_X1 _09642_ ( .A1(_02127_ ), .A2(_02132_ ), .ZN(_02133_ ) );
NAND3_X1 _09643_ ( .A1(_02105_ ), .A2(_02121_ ), .A3(\EX_LS_typ [0] ), .ZN(_02134_ ) );
NOR3_X1 _09644_ ( .A1(_02134_ ), .A2(_02130_ ), .A3(\EX_LS_flag [0] ), .ZN(_02135_ ) );
INV_X1 _09645_ ( .A(_02135_ ), .ZN(_02136_ ) );
INV_X1 _09646_ ( .A(_02114_ ), .ZN(_02137_ ) );
AND3_X1 _09647_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02138_ ) );
AOI22_X1 _09648_ ( .A1(_02137_ ), .A2(_02138_ ), .B1(_02111_ ), .B2(_02112_ ), .ZN(_02139_ ) );
NOR2_X1 _09649_ ( .A1(_02136_ ), .A2(_02139_ ), .ZN(_02140_ ) );
NOR2_X1 _09650_ ( .A1(_02133_ ), .A2(_02140_ ), .ZN(_02141_ ) );
AND2_X1 _09651_ ( .A1(_02129_ ), .A2(_02141_ ), .ZN(_02142_ ) );
AOI211_X1 _09652_ ( .A(_01910_ ), .B(_02104_ ), .C1(_02110_ ), .C2(_02142_ ), .ZN(_02143_ ) );
NOR2_X1 _09653_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02144_ ) );
AND3_X1 _09654_ ( .A1(_02096_ ), .A2(\myifu.state [0] ), .A3(_02144_ ), .ZN(_02145_ ) );
NOR4_X1 _09655_ ( .A1(_02099_ ), .A2(_02098_ ), .A3(_02100_ ), .A4(_02145_ ), .ZN(_02146_ ) );
NOR2_X1 _09656_ ( .A1(_02143_ ), .A2(_02146_ ), .ZN(_02147_ ) );
NOR2_X1 _09657_ ( .A1(_02108_ ), .A2(_01910_ ), .ZN(_02148_ ) );
NOR2_X4 _09658_ ( .A1(_02101_ ), .A2(_02148_ ), .ZN(_02149_ ) );
BUF_X8 _09659_ ( .A(_02149_ ), .Z(_02150_ ) );
CLKBUF_X2 _09660_ ( .A(_02106_ ), .Z(_02151_ ) );
CLKBUF_X2 _09661_ ( .A(_02107_ ), .Z(_02152_ ) );
OR3_X1 _09662_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(_02152_ ), .ZN(_02153_ ) );
OAI211_X1 _09663_ ( .A(_02150_ ), .B(_02153_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_02110_ ), .ZN(_02154_ ) );
INV_X4 _09664_ ( .A(_02101_ ), .ZN(_02155_ ) );
BUF_X4 _09665_ ( .A(_02155_ ), .Z(_02156_ ) );
OAI21_X1 _09666_ ( .A(_02154_ ), .B1(_01944_ ), .B2(_02156_ ), .ZN(\io_master_araddr [16] ) );
OR3_X1 _09667_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(_02107_ ), .ZN(_02157_ ) );
OAI211_X1 _09668_ ( .A(_02149_ ), .B(_02157_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_02108_ ), .ZN(_02158_ ) );
OAI21_X1 _09669_ ( .A(_02158_ ), .B1(_01939_ ), .B2(_02155_ ), .ZN(\io_master_araddr [23] ) );
OR3_X1 _09670_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(_02107_ ), .ZN(_02159_ ) );
OAI211_X1 _09671_ ( .A(_02149_ ), .B(_02159_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_02108_ ), .ZN(_02160_ ) );
INV_X1 _09672_ ( .A(\IF_ID_pc [29] ), .ZN(_02161_ ) );
OAI21_X1 _09673_ ( .A(_02160_ ), .B1(_02161_ ), .B2(_02155_ ), .ZN(\io_master_araddr [29] ) );
OR3_X1 _09674_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(_02152_ ), .ZN(_02162_ ) );
OAI211_X1 _09675_ ( .A(_02150_ ), .B(_02162_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_02109_ ), .ZN(_02163_ ) );
OAI21_X1 _09676_ ( .A(_02163_ ), .B1(_01987_ ), .B2(_02155_ ), .ZN(\io_master_araddr [26] ) );
OR4_X1 _09677_ ( .A1(\io_master_araddr [16] ), .A2(\io_master_araddr [23] ), .A3(\io_master_araddr [29] ), .A4(\io_master_araddr [26] ), .ZN(_02164_ ) );
OR3_X1 _09678_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(_02107_ ), .ZN(_02165_ ) );
OAI211_X1 _09679_ ( .A(_02149_ ), .B(_02165_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_02108_ ), .ZN(_02166_ ) );
OAI221_X1 _09680_ ( .A(\IF_ID_pc [22] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_02167_ ) );
AND2_X1 _09681_ ( .A1(_02166_ ), .A2(_02167_ ), .ZN(_02168_ ) );
OR3_X1 _09682_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [25] ), .A3(_02152_ ), .ZN(_02169_ ) );
OAI211_X2 _09683_ ( .A(_02150_ ), .B(_02169_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_02110_ ), .ZN(_02170_ ) );
INV_X1 _09684_ ( .A(\IF_ID_pc [25] ), .ZN(_02171_ ) );
OAI21_X2 _09685_ ( .A(_02170_ ), .B1(_02171_ ), .B2(_02156_ ), .ZN(\io_master_araddr [25] ) );
NAND2_X1 _09686_ ( .A1(_02168_ ), .A2(\io_master_araddr [25] ), .ZN(_02172_ ) );
OR3_X1 _09687_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(_02152_ ), .ZN(_02173_ ) );
OAI211_X1 _09688_ ( .A(_02149_ ), .B(_02173_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_02109_ ), .ZN(_02174_ ) );
OAI21_X1 _09689_ ( .A(_02174_ ), .B1(_01966_ ), .B2(_02155_ ), .ZN(\io_master_araddr [30] ) );
OR3_X1 _09690_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(_02152_ ), .ZN(_02175_ ) );
OAI211_X1 _09691_ ( .A(_02150_ ), .B(_02175_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_02109_ ), .ZN(_02176_ ) );
OAI221_X1 _09692_ ( .A(\IF_ID_pc [24] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_02177_ ) );
AND2_X1 _09693_ ( .A1(_02176_ ), .A2(_02177_ ), .ZN(_02178_ ) );
INV_X1 _09694_ ( .A(_02178_ ), .ZN(\io_master_araddr [24] ) );
NOR4_X2 _09695_ ( .A1(_02164_ ), .A2(_02172_ ), .A3(\io_master_araddr [30] ), .A4(\io_master_araddr [24] ), .ZN(_02179_ ) );
OR3_X1 _09696_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(_02152_ ), .ZN(_02180_ ) );
OAI211_X1 _09697_ ( .A(_02149_ ), .B(_02180_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_02109_ ), .ZN(_02181_ ) );
INV_X1 _09698_ ( .A(\IF_ID_pc [28] ), .ZN(_02182_ ) );
OAI21_X1 _09699_ ( .A(_02181_ ), .B1(_02182_ ), .B2(_02155_ ), .ZN(\io_master_araddr [28] ) );
OR3_X1 _09700_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(_02152_ ), .ZN(_02183_ ) );
OAI211_X1 _09701_ ( .A(_02150_ ), .B(_02183_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_02109_ ), .ZN(_02184_ ) );
INV_X1 _09702_ ( .A(\IF_ID_pc [18] ), .ZN(_02185_ ) );
OAI21_X1 _09703_ ( .A(_02184_ ), .B1(_02185_ ), .B2(_02156_ ), .ZN(\io_master_araddr [18] ) );
CLKBUF_X2 _09704_ ( .A(_02152_ ), .Z(_02186_ ) );
OR3_X1 _09705_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(_02186_ ), .ZN(_02187_ ) );
OAI211_X1 _09706_ ( .A(_02150_ ), .B(_02187_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_02110_ ), .ZN(_02188_ ) );
OAI21_X1 _09707_ ( .A(_02188_ ), .B1(_01927_ ), .B2(_02156_ ), .ZN(\io_master_araddr [27] ) );
OR3_X1 _09708_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(_02152_ ), .ZN(_02189_ ) );
OAI211_X1 _09709_ ( .A(_02149_ ), .B(_02189_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_02109_ ), .ZN(_02190_ ) );
OAI21_X1 _09710_ ( .A(_02190_ ), .B1(_02062_ ), .B2(_02155_ ), .ZN(\io_master_araddr [21] ) );
NOR4_X1 _09711_ ( .A1(\io_master_araddr [28] ), .A2(\io_master_araddr [18] ), .A3(\io_master_araddr [27] ), .A4(\io_master_araddr [21] ), .ZN(_02191_ ) );
OR3_X1 _09712_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(_02186_ ), .ZN(_02192_ ) );
OAI211_X1 _09713_ ( .A(_02150_ ), .B(_02192_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_02110_ ), .ZN(_02193_ ) );
INV_X1 _09714_ ( .A(\IF_ID_pc [19] ), .ZN(_02194_ ) );
OAI21_X1 _09715_ ( .A(_02193_ ), .B1(_02194_ ), .B2(_02156_ ), .ZN(\io_master_araddr [19] ) );
OR3_X1 _09716_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(_02107_ ), .ZN(_02195_ ) );
OAI211_X1 _09717_ ( .A(_02149_ ), .B(_02195_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_02109_ ), .ZN(_02196_ ) );
INV_X1 _09718_ ( .A(\IF_ID_pc [20] ), .ZN(_02197_ ) );
OAI21_X1 _09719_ ( .A(_02196_ ), .B1(_02197_ ), .B2(_02155_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09720_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(_02152_ ), .ZN(_02198_ ) );
OAI211_X1 _09721_ ( .A(_02150_ ), .B(_02198_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_02109_ ), .ZN(_02199_ ) );
INV_X1 _09722_ ( .A(\IF_ID_pc [17] ), .ZN(_02200_ ) );
OAI21_X1 _09723_ ( .A(_02199_ ), .B1(_02200_ ), .B2(_02156_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09724_ ( .A1(_02106_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(_02107_ ), .ZN(_02201_ ) );
OAI211_X1 _09725_ ( .A(_02149_ ), .B(_02201_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_02109_ ), .ZN(_02202_ ) );
OAI221_X1 _09726_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_02203_ ) );
NAND2_X1 _09727_ ( .A1(_02202_ ), .A2(_02203_ ), .ZN(\io_master_araddr [31] ) );
NOR4_X1 _09728_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [17] ), .A4(\io_master_araddr [31] ), .ZN(_02204_ ) );
AND2_X1 _09729_ ( .A1(_02191_ ), .A2(_02204_ ), .ZN(_02205_ ) );
AND3_X1 _09730_ ( .A1(_02179_ ), .A2(\myclint.rvalid ), .A3(_02205_ ), .ZN(_02206_ ) );
AND2_X1 _09731_ ( .A1(_02179_ ), .A2(_02205_ ), .ZN(_02207_ ) );
INV_X1 _09732_ ( .A(_02207_ ), .ZN(_02208_ ) );
AOI21_X1 _09733_ ( .A(_02104_ ), .B1(_02110_ ), .B2(_02142_ ), .ZN(_02209_ ) );
AOI211_X1 _09734_ ( .A(_02100_ ), .B(_02099_ ), .C1(\myifu.state [0] ), .C2(_02144_ ), .ZN(_02210_ ) );
OR3_X1 _09735_ ( .A1(_02208_ ), .A2(_02209_ ), .A3(_02210_ ), .ZN(_02211_ ) );
INV_X1 _09736_ ( .A(\myclint.rvalid ), .ZN(_02212_ ) );
AOI221_X4 _09737_ ( .A(fanout_net_2 ), .B1(_02147_ ), .B2(_02206_ ), .C1(_02211_ ), .C2(_02212_ ), .ZN(_00065_ ) );
INV_X1 _09738_ ( .A(\LS_WB_wdata_csreg [30] ), .ZN(_02213_ ) );
NOR2_X1 _09739_ ( .A1(_02213_ ), .A2(fanout_net_2 ), .ZN(_00066_ ) );
INV_X1 _09740_ ( .A(\LS_WB_wdata_csreg [21] ), .ZN(_02214_ ) );
NOR2_X1 _09741_ ( .A1(_02214_ ), .A2(fanout_net_2 ), .ZN(_00067_ ) );
INV_X1 _09742_ ( .A(\LS_WB_wdata_csreg [20] ), .ZN(_02215_ ) );
NOR2_X1 _09743_ ( .A1(_02215_ ), .A2(fanout_net_2 ), .ZN(_00068_ ) );
INV_X1 _09744_ ( .A(\LS_WB_wdata_csreg [19] ), .ZN(_02216_ ) );
NOR2_X1 _09745_ ( .A1(_02216_ ), .A2(fanout_net_2 ), .ZN(_00069_ ) );
INV_X1 _09746_ ( .A(\LS_WB_wdata_csreg [18] ), .ZN(_02217_ ) );
NOR2_X1 _09747_ ( .A1(_02217_ ), .A2(fanout_net_2 ), .ZN(_00070_ ) );
INV_X1 _09748_ ( .A(\LS_WB_wdata_csreg [17] ), .ZN(_02218_ ) );
NOR2_X1 _09749_ ( .A1(_02218_ ), .A2(fanout_net_2 ), .ZN(_00071_ ) );
INV_X1 _09750_ ( .A(\LS_WB_wdata_csreg [16] ), .ZN(_02219_ ) );
NOR2_X1 _09751_ ( .A1(_02219_ ), .A2(fanout_net_2 ), .ZN(_00072_ ) );
INV_X1 _09752_ ( .A(\LS_WB_wdata_csreg [15] ), .ZN(_02220_ ) );
NOR2_X1 _09753_ ( .A1(_02220_ ), .A2(fanout_net_2 ), .ZN(_00073_ ) );
INV_X1 _09754_ ( .A(\LS_WB_wdata_csreg [14] ), .ZN(_02221_ ) );
NOR2_X1 _09755_ ( .A1(_02221_ ), .A2(fanout_net_2 ), .ZN(_00074_ ) );
INV_X1 _09756_ ( .A(\LS_WB_wdata_csreg [13] ), .ZN(_02222_ ) );
NOR2_X1 _09757_ ( .A1(_02222_ ), .A2(fanout_net_2 ), .ZN(_00075_ ) );
INV_X1 _09758_ ( .A(\LS_WB_wdata_csreg [12] ), .ZN(_02223_ ) );
NOR2_X1 _09759_ ( .A1(_02223_ ), .A2(fanout_net_2 ), .ZN(_00076_ ) );
INV_X1 _09760_ ( .A(\LS_WB_wdata_csreg [29] ), .ZN(_02224_ ) );
NOR2_X1 _09761_ ( .A1(_02224_ ), .A2(fanout_net_2 ), .ZN(_00077_ ) );
INV_X1 _09762_ ( .A(\LS_WB_wdata_csreg [11] ), .ZN(_02225_ ) );
NOR2_X1 _09763_ ( .A1(_02225_ ), .A2(fanout_net_2 ), .ZN(_00078_ ) );
INV_X1 _09764_ ( .A(\LS_WB_wdata_csreg [10] ), .ZN(_02226_ ) );
NOR2_X1 _09765_ ( .A1(_02226_ ), .A2(fanout_net_2 ), .ZN(_00079_ ) );
INV_X1 _09766_ ( .A(\LS_WB_wdata_csreg [9] ), .ZN(_02227_ ) );
NOR2_X1 _09767_ ( .A1(_02227_ ), .A2(fanout_net_2 ), .ZN(_00080_ ) );
INV_X1 _09768_ ( .A(\LS_WB_wdata_csreg [8] ), .ZN(_02228_ ) );
NOR2_X1 _09769_ ( .A1(_02228_ ), .A2(fanout_net_2 ), .ZN(_00081_ ) );
INV_X1 _09770_ ( .A(\LS_WB_wdata_csreg [7] ), .ZN(_02229_ ) );
NOR2_X1 _09771_ ( .A1(_02229_ ), .A2(fanout_net_2 ), .ZN(_00082_ ) );
INV_X1 _09772_ ( .A(\LS_WB_wdata_csreg [6] ), .ZN(_02230_ ) );
NOR2_X1 _09773_ ( .A1(_02230_ ), .A2(fanout_net_2 ), .ZN(_00083_ ) );
INV_X1 _09774_ ( .A(\LS_WB_wdata_csreg [5] ), .ZN(_02231_ ) );
NOR2_X1 _09775_ ( .A1(_02231_ ), .A2(fanout_net_2 ), .ZN(_00084_ ) );
INV_X1 _09776_ ( .A(\LS_WB_wdata_csreg [4] ), .ZN(_02232_ ) );
NOR2_X1 _09777_ ( .A1(_02232_ ), .A2(fanout_net_2 ), .ZN(_00085_ ) );
INV_X1 _09778_ ( .A(\LS_WB_wdata_csreg [3] ), .ZN(_02233_ ) );
NOR2_X1 _09779_ ( .A1(_02233_ ), .A2(fanout_net_2 ), .ZN(_00086_ ) );
INV_X1 _09780_ ( .A(\LS_WB_wdata_csreg [2] ), .ZN(_02234_ ) );
NOR2_X1 _09781_ ( .A1(_02234_ ), .A2(fanout_net_2 ), .ZN(_00087_ ) );
INV_X1 _09782_ ( .A(\LS_WB_wdata_csreg [28] ), .ZN(_02235_ ) );
NOR2_X1 _09783_ ( .A1(_02235_ ), .A2(fanout_net_2 ), .ZN(_00088_ ) );
INV_X1 _09784_ ( .A(\LS_WB_wdata_csreg [1] ), .ZN(_02236_ ) );
NOR2_X1 _09785_ ( .A1(_02236_ ), .A2(fanout_net_2 ), .ZN(_00089_ ) );
INV_X1 _09786_ ( .A(\LS_WB_wdata_csreg [0] ), .ZN(_02237_ ) );
NOR2_X1 _09787_ ( .A1(_02237_ ), .A2(fanout_net_2 ), .ZN(_00090_ ) );
INV_X1 _09788_ ( .A(\LS_WB_wdata_csreg [27] ), .ZN(_02238_ ) );
NOR2_X1 _09789_ ( .A1(_02238_ ), .A2(fanout_net_3 ), .ZN(_00091_ ) );
INV_X1 _09790_ ( .A(\LS_WB_wdata_csreg [26] ), .ZN(_02239_ ) );
NOR2_X1 _09791_ ( .A1(_02239_ ), .A2(fanout_net_3 ), .ZN(_00092_ ) );
INV_X1 _09792_ ( .A(\LS_WB_wdata_csreg [25] ), .ZN(_02240_ ) );
NOR2_X1 _09793_ ( .A1(_02240_ ), .A2(fanout_net_3 ), .ZN(_00093_ ) );
INV_X1 _09794_ ( .A(\LS_WB_wdata_csreg [24] ), .ZN(_02241_ ) );
NOR2_X1 _09795_ ( .A1(_02241_ ), .A2(fanout_net_3 ), .ZN(_00094_ ) );
INV_X1 _09796_ ( .A(\LS_WB_wdata_csreg [23] ), .ZN(_02242_ ) );
NOR2_X1 _09797_ ( .A1(_02242_ ), .A2(fanout_net_3 ), .ZN(_00095_ ) );
INV_X1 _09798_ ( .A(\LS_WB_wdata_csreg [22] ), .ZN(_02243_ ) );
NOR2_X1 _09799_ ( .A1(_02243_ ), .A2(fanout_net_3 ), .ZN(_00096_ ) );
NOR3_X1 _09800_ ( .A1(_01633_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00097_ ) );
NOR3_X1 _09801_ ( .A1(_02213_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00098_ ) );
NOR3_X1 _09802_ ( .A1(_02214_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00099_ ) );
NOR3_X1 _09803_ ( .A1(_02215_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00100_ ) );
NOR3_X1 _09804_ ( .A1(_02216_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00101_ ) );
NOR3_X1 _09805_ ( .A1(_02217_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00102_ ) );
NOR3_X1 _09806_ ( .A1(_02218_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00103_ ) );
NOR3_X1 _09807_ ( .A1(_02219_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00104_ ) );
NOR3_X1 _09808_ ( .A1(_02220_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00105_ ) );
NOR3_X1 _09809_ ( .A1(_02221_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00106_ ) );
NOR3_X1 _09810_ ( .A1(_02222_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00107_ ) );
NOR3_X1 _09811_ ( .A1(_02223_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00108_ ) );
NOR3_X1 _09812_ ( .A1(_02224_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00109_ ) );
NOR3_X1 _09813_ ( .A1(_02225_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00110_ ) );
NOR3_X1 _09814_ ( .A1(_02226_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00111_ ) );
NOR3_X1 _09815_ ( .A1(_02227_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00112_ ) );
NOR3_X1 _09816_ ( .A1(_02228_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00113_ ) );
NOR3_X1 _09817_ ( .A1(_02229_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00114_ ) );
NOR3_X1 _09818_ ( .A1(_02230_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00115_ ) );
NOR3_X1 _09819_ ( .A1(_02231_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00116_ ) );
NOR3_X1 _09820_ ( .A1(_02232_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00117_ ) );
INV_X1 _09821_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02244_ ) );
NOR2_X1 _09822_ ( .A1(_02244_ ), .A2(\LS_WB_wen_csreg [3] ), .ZN(_02245_ ) );
AOI211_X1 _09823_ ( .A(fanout_net_3 ), .B(_02245_ ), .C1(_02233_ ), .C2(_02244_ ), .ZN(_00118_ ) );
NOR2_X1 _09824_ ( .A1(_02244_ ), .A2(\LS_WB_wen_csreg [2] ), .ZN(_02246_ ) );
AOI211_X1 _09825_ ( .A(fanout_net_3 ), .B(_02246_ ), .C1(_02234_ ), .C2(_02244_ ), .ZN(_00119_ ) );
NOR3_X1 _09826_ ( .A1(_02235_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00120_ ) );
NOR2_X1 _09827_ ( .A1(_02244_ ), .A2(\LS_WB_wen_csreg [1] ), .ZN(_02247_ ) );
AOI211_X1 _09828_ ( .A(fanout_net_4 ), .B(_02247_ ), .C1(_02236_ ), .C2(_02244_ ), .ZN(_00121_ ) );
NOR2_X1 _09829_ ( .A1(_02244_ ), .A2(\LS_WB_wen_csreg [0] ), .ZN(_02248_ ) );
AOI211_X1 _09830_ ( .A(fanout_net_4 ), .B(_02248_ ), .C1(_02237_ ), .C2(_02244_ ), .ZN(_00122_ ) );
NOR3_X1 _09831_ ( .A1(_02238_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00123_ ) );
NOR3_X1 _09832_ ( .A1(_02239_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00124_ ) );
NOR3_X1 _09833_ ( .A1(_02240_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00125_ ) );
NOR3_X1 _09834_ ( .A1(_02241_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00126_ ) );
NOR3_X1 _09835_ ( .A1(_02242_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00127_ ) );
NOR3_X1 _09836_ ( .A1(_02243_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00128_ ) );
AND3_X1 _09837_ ( .A1(_01794_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00129_ ) );
NOR2_X1 _09838_ ( .A1(\myec.state [1] ), .A2(\myec.state [0] ), .ZN(_02249_ ) );
OR2_X1 _09839_ ( .A1(\myexu.pc_jump [25] ), .A2(\myexu.pc_jump [24] ), .ZN(_02250_ ) );
OR3_X1 _09840_ ( .A1(_02250_ ), .A2(\myexu.pc_jump [27] ), .A3(\myexu.pc_jump [26] ), .ZN(_02251_ ) );
OR4_X1 _09841_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02252_ ) );
NOR2_X1 _09842_ ( .A1(_02251_ ), .A2(_02252_ ), .ZN(_02253_ ) );
INV_X1 _09843_ ( .A(_02253_ ), .ZN(_02254_ ) );
NOR2_X1 _09844_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02255_ ) );
AOI21_X1 _09845_ ( .A(exception_quest_IDU ), .B1(_02254_ ), .B2(_02255_ ), .ZN(_02256_ ) );
OAI211_X1 _09846_ ( .A(_01634_ ), .B(_02249_ ), .C1(_02256_ ), .C2(exception_quest_IDU ), .ZN(_02257_ ) );
INV_X2 _09847_ ( .A(_02141_ ), .ZN(_02258_ ) );
NOR4_X1 _09848_ ( .A1(_02257_ ), .A2(_02258_ ), .A3(_02128_ ), .A4(_02123_ ), .ZN(_00130_ ) );
INV_X1 _09849_ ( .A(_02249_ ), .ZN(_02259_ ) );
AOI211_X1 _09850_ ( .A(fanout_net_4 ), .B(_02259_ ), .C1(_02142_ ), .C2(exception_quest_IDU ), .ZN(_00131_ ) );
INV_X1 _09851_ ( .A(IDU_valid_EXU ), .ZN(_02260_ ) );
NOR2_X1 _09852_ ( .A1(_02260_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _09853_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_02261_ ) );
INV_X1 _09854_ ( .A(\ID_EX_typ [5] ), .ZN(_02262_ ) );
NOR2_X1 _09855_ ( .A1(_02262_ ), .A2(\ID_EX_typ [6] ), .ZN(_02263_ ) );
AND3_X1 _09856_ ( .A1(_02263_ ), .A2(\ID_EX_typ [7] ), .A3(fanout_net_8 ), .ZN(_02264_ ) );
INV_X1 _09857_ ( .A(check_quest ), .ZN(_02265_ ) );
NOR2_X1 _09858_ ( .A1(_02265_ ), .A2(check_assert ), .ZN(_02266_ ) );
INV_X1 _09859_ ( .A(\ID_EX_typ [6] ), .ZN(_02267_ ) );
NAND3_X1 _09860_ ( .A1(_02267_ ), .A2(_02262_ ), .A3(\ID_EX_typ [7] ), .ZN(_02268_ ) );
MUX2_X1 _09861_ ( .A(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .B(_02266_ ), .S(_02268_ ), .Z(_02269_ ) );
INV_X1 _09862_ ( .A(\ID_EX_typ [7] ), .ZN(_02270_ ) );
NOR2_X1 _09863_ ( .A1(_02270_ ), .A2(\ID_EX_typ [6] ), .ZN(_02271_ ) );
AND2_X2 _09864_ ( .A1(_02271_ ), .A2(\ID_EX_typ [5] ), .ZN(_02272_ ) );
INV_X1 _09865_ ( .A(_02272_ ), .ZN(_02273_ ) );
BUF_X4 _09866_ ( .A(_02273_ ), .Z(_02274_ ) );
BUF_X4 _09867_ ( .A(_02274_ ), .Z(_02275_ ) );
AOI211_X1 _09868_ ( .A(_02261_ ), .B(_02264_ ), .C1(_02269_ ), .C2(_02275_ ), .ZN(_02276_ ) );
NOR2_X1 _09869_ ( .A1(fanout_net_4 ), .A2(fanout_net_20 ), .ZN(_02277_ ) );
BUF_X2 _09870_ ( .A(_02277_ ), .Z(_02278_ ) );
CLKBUF_X2 _09871_ ( .A(_02278_ ), .Z(_02279_ ) );
OAI21_X1 _09872_ ( .A(_02279_ ), .B1(\myexu.state_$_ANDNOT__B_Y ), .B2(_02266_ ), .ZN(_02280_ ) );
NOR2_X1 _09873_ ( .A1(_02276_ ), .A2(_02280_ ), .ZN(_00132_ ) );
INV_X32 _09874_ ( .A(fanout_net_21 ), .ZN(_02281_ ) );
BUF_X4 _09875_ ( .A(_02281_ ), .Z(_02282_ ) );
BUF_X4 _09876_ ( .A(_02282_ ), .Z(_02283_ ) );
BUF_X8 _09877_ ( .A(_02283_ ), .Z(_02284_ ) );
BUF_X2 _09878_ ( .A(_02284_ ), .Z(_02285_ ) );
BUF_X4 _09879_ ( .A(_02285_ ), .Z(_02286_ ) );
BUF_X4 _09880_ ( .A(_02286_ ), .Z(_02287_ ) );
NOR2_X1 _09881_ ( .A1(_02287_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02288_ ) );
OAI21_X1 _09882_ ( .A(fanout_net_29 ), .B1(fanout_net_21 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02289_ ) );
NOR2_X1 _09883_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02290_ ) );
INV_X2 _09884_ ( .A(fanout_net_29 ), .ZN(_02291_ ) );
BUF_X4 _09885_ ( .A(_02291_ ), .Z(_02292_ ) );
BUF_X4 _09886_ ( .A(_02292_ ), .Z(_02293_ ) );
BUF_X4 _09887_ ( .A(_02293_ ), .Z(_02294_ ) );
BUF_X4 _09888_ ( .A(_02294_ ), .Z(_02295_ ) );
BUF_X4 _09889_ ( .A(_02295_ ), .Z(_02296_ ) );
BUF_X4 _09890_ ( .A(_02296_ ), .Z(_02297_ ) );
BUF_X2 _09891_ ( .A(_02284_ ), .Z(_02298_ ) );
BUF_X8 _09892_ ( .A(_02298_ ), .Z(_02299_ ) );
BUF_X4 _09893_ ( .A(_02299_ ), .Z(_02300_ ) );
BUF_X4 _09894_ ( .A(_02300_ ), .Z(_02301_ ) );
OAI21_X1 _09895_ ( .A(_02297_ ), .B1(_02301_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02302_ ) );
OAI221_X1 _09896_ ( .A(fanout_net_32 ), .B1(_02288_ ), .B2(_02289_ ), .C1(_02290_ ), .C2(_02302_ ), .ZN(_02303_ ) );
MUX2_X1 _09897_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02304_ ) );
MUX2_X1 _09898_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02305_ ) );
MUX2_X1 _09899_ ( .A(_02304_ ), .B(_02305_ ), .S(_02297_ ), .Z(_02306_ ) );
OAI211_X1 _09900_ ( .A(fanout_net_34 ), .B(_02303_ ), .C1(_02306_ ), .C2(fanout_net_32 ), .ZN(_02307_ ) );
MUX2_X1 _09901_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02308_ ) );
AND2_X1 _09902_ ( .A1(_02308_ ), .A2(_02297_ ), .ZN(_02309_ ) );
MUX2_X1 _09903_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02310_ ) );
AOI211_X1 _09904_ ( .A(fanout_net_32 ), .B(_02309_ ), .C1(fanout_net_29 ), .C2(_02310_ ), .ZN(_02311_ ) );
INV_X1 _09905_ ( .A(fanout_net_34 ), .ZN(_02312_ ) );
BUF_X4 _09906_ ( .A(_02312_ ), .Z(_02313_ ) );
BUF_X4 _09907_ ( .A(_02313_ ), .Z(_02314_ ) );
BUF_X4 _09908_ ( .A(_02314_ ), .Z(_02315_ ) );
MUX2_X1 _09909_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02316_ ) );
MUX2_X1 _09910_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02317_ ) );
MUX2_X1 _09911_ ( .A(_02316_ ), .B(_02317_ ), .S(fanout_net_29 ), .Z(_02318_ ) );
INV_X2 _09912_ ( .A(fanout_net_32 ), .ZN(_02319_ ) );
BUF_X4 _09913_ ( .A(_02319_ ), .Z(_02320_ ) );
BUF_X4 _09914_ ( .A(_02320_ ), .Z(_02321_ ) );
BUF_X4 _09915_ ( .A(_02321_ ), .Z(_02322_ ) );
BUF_X4 _09916_ ( .A(_02322_ ), .Z(_02323_ ) );
BUF_X4 _09917_ ( .A(_02323_ ), .Z(_02324_ ) );
OAI21_X1 _09918_ ( .A(_02315_ ), .B1(_02318_ ), .B2(_02324_ ), .ZN(_02325_ ) );
AND3_X1 _09919_ ( .A1(_02130_ ), .A2(\EX_LS_flag [0] ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02326_ ) );
INV_X1 _09920_ ( .A(\EX_LS_flag [0] ), .ZN(_02327_ ) );
NOR2_X1 _09921_ ( .A1(_02327_ ), .A2(\EX_LS_flag [1] ), .ZN(_02328_ ) );
AOI211_X2 _09922_ ( .A(_02326_ ), .B(_02120_ ), .C1(\EX_LS_flag [2] ), .C2(_02328_ ), .ZN(_02329_ ) );
AND2_X4 _09923_ ( .A1(_02131_ ), .A2(\EX_LS_flag [2] ), .ZN(_02330_ ) );
BUF_X16 _09924_ ( .A(_02330_ ), .Z(_02331_ ) );
INV_X8 _09925_ ( .A(_02331_ ), .ZN(_02332_ ) );
NAND2_X4 _09926_ ( .A1(_02329_ ), .A2(_02332_ ), .ZN(_02333_ ) );
XNOR2_X1 _09927_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02334_ ) );
OR4_X4 _09928_ ( .A1(\EX_LS_dest_reg [3] ), .A2(\EX_LS_dest_reg [2] ), .A3(\EX_LS_dest_reg [1] ), .A4(\EX_LS_dest_reg [0] ), .ZN(_02335_ ) );
OR2_X4 _09929_ ( .A1(_02335_ ), .A2(\EX_LS_dest_reg [4] ), .ZN(_02336_ ) );
INV_X1 _09930_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02337_ ) );
NAND2_X1 _09931_ ( .A1(_02337_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02338_ ) );
NAND4_X4 _09932_ ( .A1(_02333_ ), .A2(_02334_ ), .A3(_02336_ ), .A4(_02338_ ), .ZN(_02339_ ) );
BUF_X8 _09933_ ( .A(_02339_ ), .Z(_02340_ ) );
BUF_X8 _09934_ ( .A(_02340_ ), .Z(_02341_ ) );
BUF_X4 _09935_ ( .A(_02341_ ), .Z(_02342_ ) );
BUF_X2 _09936_ ( .A(_02342_ ), .Z(_02343_ ) );
XNOR2_X1 _09937_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .ZN(_02344_ ) );
XNOR2_X1 _09938_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .ZN(_02345_ ) );
INV_X1 _09939_ ( .A(\EX_LS_dest_reg [3] ), .ZN(_02346_ ) );
INV_X2 _09940_ ( .A(\ID_EX_rs1 [1] ), .ZN(_02347_ ) );
AOI22_X1 _09941_ ( .A1(\ID_EX_rs1 [3] ), .A2(_02346_ ), .B1(_02347_ ), .B2(\EX_LS_dest_reg [1] ), .ZN(_02348_ ) );
INV_X2 _09942_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .ZN(_02349_ ) );
INV_X1 _09943_ ( .A(\ID_EX_rs1 [3] ), .ZN(_02350_ ) );
AOI21_X1 _09944_ ( .A(_02349_ ), .B1(_02350_ ), .B2(\EX_LS_dest_reg [3] ), .ZN(_02351_ ) );
NAND4_X4 _09945_ ( .A1(_02344_ ), .A2(_02345_ ), .A3(_02348_ ), .A4(_02351_ ), .ZN(_02352_ ) );
BUF_X2 _09946_ ( .A(_02352_ ), .Z(_02353_ ) );
BUF_X2 _09947_ ( .A(_02353_ ), .Z(_02354_ ) );
BUF_X2 _09948_ ( .A(_02354_ ), .Z(_02355_ ) );
OAI221_X1 _09949_ ( .A(_02307_ ), .B1(_02311_ ), .B2(_02325_ ), .C1(_02343_ ), .C2(_02355_ ), .ZN(_02356_ ) );
OR3_X1 _09950_ ( .A1(_02343_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02357_ ) );
AND2_X2 _09951_ ( .A1(_02356_ ), .A2(_02357_ ), .ZN(_02358_ ) );
INV_X1 _09952_ ( .A(\ID_EX_imm [30] ), .ZN(_02359_ ) );
XNOR2_X1 _09953_ ( .A(_02358_ ), .B(_02359_ ), .ZN(_02360_ ) );
INV_X1 _09954_ ( .A(_02360_ ), .ZN(_02361_ ) );
OR3_X1 _09955_ ( .A1(_02342_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02354_ ), .ZN(_02362_ ) );
OR2_X1 _09956_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02363_ ) );
BUF_X4 _09957_ ( .A(_02295_ ), .Z(_02364_ ) );
OAI211_X1 _09958_ ( .A(_02363_ ), .B(_02364_ ), .C1(_02287_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02365_ ) );
OR2_X1 _09959_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02366_ ) );
OAI211_X1 _09960_ ( .A(_02366_ ), .B(fanout_net_29 ), .C1(_02300_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02367_ ) );
NAND3_X1 _09961_ ( .A1(_02365_ ), .A2(_02367_ ), .A3(fanout_net_32 ), .ZN(_02368_ ) );
MUX2_X1 _09962_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02369_ ) );
MUX2_X1 _09963_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02370_ ) );
MUX2_X1 _09964_ ( .A(_02369_ ), .B(_02370_ ), .S(_02296_ ), .Z(_02371_ ) );
OAI211_X1 _09965_ ( .A(_02315_ ), .B(_02368_ ), .C1(_02371_ ), .C2(fanout_net_32 ), .ZN(_02372_ ) );
NOR2_X1 _09966_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02373_ ) );
OAI21_X1 _09967_ ( .A(_02296_ ), .B1(_02286_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02374_ ) );
INV_X1 _09968_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02375_ ) );
INV_X1 _09969_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02376_ ) );
MUX2_X1 _09970_ ( .A(_02375_ ), .B(_02376_ ), .S(fanout_net_21 ), .Z(_02377_ ) );
BUF_X4 _09971_ ( .A(_02295_ ), .Z(_02378_ ) );
OAI221_X1 _09972_ ( .A(_02323_ ), .B1(_02373_ ), .B2(_02374_ ), .C1(_02377_ ), .C2(_02378_ ), .ZN(_02379_ ) );
MUX2_X1 _09973_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02380_ ) );
MUX2_X1 _09974_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02381_ ) );
MUX2_X1 _09975_ ( .A(_02380_ ), .B(_02381_ ), .S(fanout_net_29 ), .Z(_02382_ ) );
BUF_X4 _09976_ ( .A(_02323_ ), .Z(_02383_ ) );
OAI211_X1 _09977_ ( .A(fanout_net_34 ), .B(_02379_ ), .C1(_02382_ ), .C2(_02383_ ), .ZN(_02384_ ) );
BUF_X8 _09978_ ( .A(_02342_ ), .Z(_02385_ ) );
BUF_X2 _09979_ ( .A(_02354_ ), .Z(_02386_ ) );
OAI211_X1 _09980_ ( .A(_02372_ ), .B(_02384_ ), .C1(_02385_ ), .C2(_02386_ ), .ZN(_02387_ ) );
NAND2_X1 _09981_ ( .A1(_02362_ ), .A2(_02387_ ), .ZN(_02388_ ) );
XNOR2_X1 _09982_ ( .A(_02388_ ), .B(\ID_EX_imm [28] ), .ZN(_02389_ ) );
OR3_X1 _09983_ ( .A1(_02342_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02354_ ), .ZN(_02390_ ) );
OR2_X1 _09984_ ( .A1(_02285_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02391_ ) );
OAI211_X1 _09985_ ( .A(_02391_ ), .B(_02296_ ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02392_ ) );
OR2_X1 _09986_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02393_ ) );
OAI211_X1 _09987_ ( .A(_02393_ ), .B(fanout_net_29 ), .C1(_02286_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02394_ ) );
NAND3_X1 _09988_ ( .A1(_02392_ ), .A2(_02323_ ), .A3(_02394_ ), .ZN(_02395_ ) );
MUX2_X1 _09989_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02396_ ) );
MUX2_X1 _09990_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02397_ ) );
MUX2_X1 _09991_ ( .A(_02396_ ), .B(_02397_ ), .S(_02295_ ), .Z(_02398_ ) );
OAI211_X1 _09992_ ( .A(_02314_ ), .B(_02395_ ), .C1(_02398_ ), .C2(_02383_ ), .ZN(_02399_ ) );
OR2_X1 _09993_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02400_ ) );
OAI211_X1 _09994_ ( .A(_02400_ ), .B(fanout_net_29 ), .C1(_02286_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02401_ ) );
OR2_X1 _09995_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02402_ ) );
OAI211_X1 _09996_ ( .A(_02402_ ), .B(_02296_ ), .C1(_02286_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02403_ ) );
NAND3_X1 _09997_ ( .A1(_02401_ ), .A2(_02403_ ), .A3(fanout_net_32 ), .ZN(_02404_ ) );
MUX2_X1 _09998_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02405_ ) );
MUX2_X1 _09999_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02406_ ) );
MUX2_X1 _10000_ ( .A(_02405_ ), .B(_02406_ ), .S(fanout_net_29 ), .Z(_02407_ ) );
OAI211_X1 _10001_ ( .A(fanout_net_34 ), .B(_02404_ ), .C1(_02407_ ), .C2(fanout_net_32 ), .ZN(_02408_ ) );
OAI211_X1 _10002_ ( .A(_02399_ ), .B(_02408_ ), .C1(_02385_ ), .C2(_02386_ ), .ZN(_02409_ ) );
NAND2_X1 _10003_ ( .A1(_02390_ ), .A2(_02409_ ), .ZN(_02410_ ) );
BUF_X4 _10004_ ( .A(_02410_ ), .Z(_02411_ ) );
INV_X1 _10005_ ( .A(\ID_EX_imm [22] ), .ZN(_02412_ ) );
XNOR2_X1 _10006_ ( .A(_02411_ ), .B(_02412_ ), .ZN(_02413_ ) );
BUF_X2 _10007_ ( .A(_02352_ ), .Z(_02414_ ) );
BUF_X8 _10008_ ( .A(_02414_ ), .Z(_02415_ ) );
OR3_X4 _10009_ ( .A1(_02342_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02415_ ), .ZN(_02416_ ) );
OR2_X1 _10010_ ( .A1(_02298_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02417_ ) );
OAI211_X1 _10011_ ( .A(_02417_ ), .B(fanout_net_29 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02418_ ) );
OR2_X1 _10012_ ( .A1(fanout_net_21 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02419_ ) );
OAI211_X1 _10013_ ( .A(_02419_ ), .B(_02295_ ), .C1(_02299_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02420_ ) );
NAND3_X1 _10014_ ( .A1(_02418_ ), .A2(_02323_ ), .A3(_02420_ ), .ZN(_02421_ ) );
MUX2_X1 _10015_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02422_ ) );
MUX2_X1 _10016_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02423_ ) );
MUX2_X1 _10017_ ( .A(_02422_ ), .B(_02423_ ), .S(_02295_ ), .Z(_02424_ ) );
OAI211_X1 _10018_ ( .A(_02314_ ), .B(_02421_ ), .C1(_02424_ ), .C2(_02323_ ), .ZN(_02425_ ) );
OR2_X1 _10019_ ( .A1(_02298_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02426_ ) );
OAI211_X1 _10020_ ( .A(_02426_ ), .B(fanout_net_29 ), .C1(fanout_net_21 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02427_ ) );
OR2_X1 _10021_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02428_ ) );
OAI211_X1 _10022_ ( .A(_02428_ ), .B(_02295_ ), .C1(_02299_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02429_ ) );
NAND3_X1 _10023_ ( .A1(_02427_ ), .A2(fanout_net_32 ), .A3(_02429_ ), .ZN(_02430_ ) );
MUX2_X1 _10024_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02431_ ) );
MUX2_X1 _10025_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02432_ ) );
MUX2_X1 _10026_ ( .A(_02431_ ), .B(_02432_ ), .S(fanout_net_29 ), .Z(_02433_ ) );
OAI211_X1 _10027_ ( .A(fanout_net_34 ), .B(_02430_ ), .C1(_02433_ ), .C2(fanout_net_32 ), .ZN(_02434_ ) );
OAI211_X1 _10028_ ( .A(_02425_ ), .B(_02434_ ), .C1(_02342_ ), .C2(_02354_ ), .ZN(_02435_ ) );
INV_X1 _10029_ ( .A(\ID_EX_imm [23] ), .ZN(_02436_ ) );
NAND3_X1 _10030_ ( .A1(_02416_ ), .A2(_02435_ ), .A3(_02436_ ), .ZN(_02437_ ) );
NAND2_X2 _10031_ ( .A1(_02416_ ), .A2(_02435_ ), .ZN(_02438_ ) );
NAND2_X1 _10032_ ( .A1(_02438_ ), .A2(\ID_EX_imm [23] ), .ZN(_02439_ ) );
AND3_X1 _10033_ ( .A1(_02413_ ), .A2(_02437_ ), .A3(_02439_ ), .ZN(_02440_ ) );
OR3_X1 _10034_ ( .A1(_02342_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02354_ ), .ZN(_02441_ ) );
INV_X1 _10035_ ( .A(\ID_EX_imm [21] ), .ZN(_02442_ ) );
OR2_X1 _10036_ ( .A1(_02285_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02443_ ) );
OAI211_X1 _10037_ ( .A(_02443_ ), .B(fanout_net_29 ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02444_ ) );
OR2_X1 _10038_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02445_ ) );
OAI211_X1 _10039_ ( .A(_02445_ ), .B(_02296_ ), .C1(_02286_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02446_ ) );
NAND3_X1 _10040_ ( .A1(_02444_ ), .A2(_02323_ ), .A3(_02446_ ), .ZN(_02447_ ) );
MUX2_X1 _10041_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02448_ ) );
MUX2_X1 _10042_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02449_ ) );
MUX2_X1 _10043_ ( .A(_02448_ ), .B(_02449_ ), .S(_02295_ ), .Z(_02450_ ) );
OAI211_X1 _10044_ ( .A(_02314_ ), .B(_02447_ ), .C1(_02450_ ), .C2(_02383_ ), .ZN(_02451_ ) );
OR2_X1 _10045_ ( .A1(_02285_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02452_ ) );
OAI211_X1 _10046_ ( .A(_02452_ ), .B(_02296_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02453_ ) );
OR2_X1 _10047_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02454_ ) );
OAI211_X1 _10048_ ( .A(_02454_ ), .B(fanout_net_29 ), .C1(_02286_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02455_ ) );
NAND3_X1 _10049_ ( .A1(_02453_ ), .A2(fanout_net_32 ), .A3(_02455_ ), .ZN(_02456_ ) );
MUX2_X1 _10050_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02457_ ) );
MUX2_X1 _10051_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02458_ ) );
MUX2_X1 _10052_ ( .A(_02457_ ), .B(_02458_ ), .S(fanout_net_29 ), .Z(_02459_ ) );
OAI211_X1 _10053_ ( .A(fanout_net_34 ), .B(_02456_ ), .C1(_02459_ ), .C2(fanout_net_32 ), .ZN(_02460_ ) );
OAI211_X1 _10054_ ( .A(_02451_ ), .B(_02460_ ), .C1(_02342_ ), .C2(_02354_ ), .ZN(_02461_ ) );
AND3_X1 _10055_ ( .A1(_02441_ ), .A2(_02442_ ), .A3(_02461_ ), .ZN(_02462_ ) );
AOI21_X1 _10056_ ( .A(_02442_ ), .B1(_02441_ ), .B2(_02461_ ), .ZN(_02463_ ) );
NOR2_X1 _10057_ ( .A1(_02462_ ), .A2(_02463_ ), .ZN(_02464_ ) );
OR3_X1 _10058_ ( .A1(_02385_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02386_ ), .ZN(_02465_ ) );
OR2_X1 _10059_ ( .A1(_02286_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02466_ ) );
OAI211_X1 _10060_ ( .A(_02466_ ), .B(_02378_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02467_ ) );
OR2_X1 _10061_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02468_ ) );
OAI211_X1 _10062_ ( .A(_02468_ ), .B(fanout_net_29 ), .C1(_02287_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02469_ ) );
NAND3_X1 _10063_ ( .A1(_02467_ ), .A2(fanout_net_32 ), .A3(_02469_ ), .ZN(_02470_ ) );
MUX2_X1 _10064_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02471_ ) );
MUX2_X1 _10065_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02472_ ) );
MUX2_X1 _10066_ ( .A(_02471_ ), .B(_02472_ ), .S(_02364_ ), .Z(_02473_ ) );
OAI211_X1 _10067_ ( .A(_02315_ ), .B(_02470_ ), .C1(_02473_ ), .C2(fanout_net_32 ), .ZN(_02474_ ) );
NOR2_X1 _10068_ ( .A1(_02300_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02475_ ) );
OAI21_X1 _10069_ ( .A(fanout_net_29 ), .B1(fanout_net_22 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02476_ ) );
NOR2_X1 _10070_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02477_ ) );
OAI21_X1 _10071_ ( .A(_02364_ ), .B1(_02300_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02478_ ) );
OAI221_X1 _10072_ ( .A(_02383_ ), .B1(_02475_ ), .B2(_02476_ ), .C1(_02477_ ), .C2(_02478_ ), .ZN(_02479_ ) );
MUX2_X1 _10073_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02480_ ) );
MUX2_X1 _10074_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02481_ ) );
MUX2_X1 _10075_ ( .A(_02480_ ), .B(_02481_ ), .S(fanout_net_29 ), .Z(_02482_ ) );
OAI211_X1 _10076_ ( .A(fanout_net_34 ), .B(_02479_ ), .C1(_02482_ ), .C2(_02324_ ), .ZN(_02483_ ) );
OAI211_X1 _10077_ ( .A(_02474_ ), .B(_02483_ ), .C1(_02385_ ), .C2(_02386_ ), .ZN(_02484_ ) );
NAND2_X2 _10078_ ( .A1(_02465_ ), .A2(_02484_ ), .ZN(_02485_ ) );
XOR2_X1 _10079_ ( .A(_02485_ ), .B(\ID_EX_imm [20] ), .Z(_02486_ ) );
NAND3_X1 _10080_ ( .A1(_02440_ ), .A2(_02464_ ), .A3(_02486_ ), .ZN(_02487_ ) );
OR3_X1 _10081_ ( .A1(_02341_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02415_ ), .ZN(_02488_ ) );
OR2_X1 _10082_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02489_ ) );
BUF_X4 _10083_ ( .A(_02293_ ), .Z(_02490_ ) );
BUF_X4 _10084_ ( .A(_02490_ ), .Z(_02491_ ) );
OAI211_X1 _10085_ ( .A(_02489_ ), .B(_02491_ ), .C1(_02285_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02492_ ) );
OR2_X1 _10086_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02493_ ) );
OAI211_X1 _10087_ ( .A(_02493_ ), .B(fanout_net_29 ), .C1(_02285_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02494_ ) );
NAND3_X1 _10088_ ( .A1(_02492_ ), .A2(_02494_ ), .A3(_02322_ ), .ZN(_02495_ ) );
MUX2_X1 _10089_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02496_ ) );
MUX2_X1 _10090_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02497_ ) );
MUX2_X1 _10091_ ( .A(_02496_ ), .B(_02497_ ), .S(_02491_ ), .Z(_02498_ ) );
OAI211_X1 _10092_ ( .A(_02314_ ), .B(_02495_ ), .C1(_02498_ ), .C2(_02322_ ), .ZN(_02499_ ) );
OR2_X1 _10093_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02500_ ) );
OAI211_X1 _10094_ ( .A(_02500_ ), .B(fanout_net_29 ), .C1(_02285_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02501_ ) );
OR2_X1 _10095_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02502_ ) );
OAI211_X1 _10096_ ( .A(_02502_ ), .B(_02491_ ), .C1(_02285_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02503_ ) );
NAND3_X1 _10097_ ( .A1(_02501_ ), .A2(_02503_ ), .A3(fanout_net_32 ), .ZN(_02504_ ) );
MUX2_X1 _10098_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02505_ ) );
MUX2_X1 _10099_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02506_ ) );
MUX2_X1 _10100_ ( .A(_02505_ ), .B(_02506_ ), .S(fanout_net_29 ), .Z(_02507_ ) );
OAI211_X1 _10101_ ( .A(fanout_net_34 ), .B(_02504_ ), .C1(_02507_ ), .C2(fanout_net_32 ), .ZN(_02508_ ) );
OAI211_X1 _10102_ ( .A(_02499_ ), .B(_02508_ ), .C1(_02341_ ), .C2(_02354_ ), .ZN(_02509_ ) );
NAND2_X2 _10103_ ( .A1(_02488_ ), .A2(_02509_ ), .ZN(_02510_ ) );
INV_X1 _10104_ ( .A(\ID_EX_imm [18] ), .ZN(_02511_ ) );
XNOR2_X1 _10105_ ( .A(_02510_ ), .B(_02511_ ), .ZN(_02512_ ) );
OR3_X1 _10106_ ( .A1(_02341_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02415_ ), .ZN(_02513_ ) );
OR2_X1 _10107_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02514_ ) );
OAI211_X1 _10108_ ( .A(_02514_ ), .B(_02491_ ), .C1(_02298_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02515_ ) );
OR2_X1 _10109_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02516_ ) );
OAI211_X1 _10110_ ( .A(_02516_ ), .B(fanout_net_29 ), .C1(_02298_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02517_ ) );
NAND3_X1 _10111_ ( .A1(_02515_ ), .A2(_02517_ ), .A3(_02322_ ), .ZN(_02518_ ) );
MUX2_X1 _10112_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02519_ ) );
MUX2_X1 _10113_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02520_ ) );
MUX2_X1 _10114_ ( .A(_02519_ ), .B(_02520_ ), .S(_02491_ ), .Z(_02521_ ) );
OAI211_X1 _10115_ ( .A(_02314_ ), .B(_02518_ ), .C1(_02521_ ), .C2(_02322_ ), .ZN(_02522_ ) );
OR2_X1 _10116_ ( .A1(_02284_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02523_ ) );
OAI211_X1 _10117_ ( .A(_02523_ ), .B(_02491_ ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02524_ ) );
OR2_X1 _10118_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02525_ ) );
OAI211_X1 _10119_ ( .A(_02525_ ), .B(fanout_net_29 ), .C1(_02298_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02526_ ) );
NAND3_X1 _10120_ ( .A1(_02524_ ), .A2(fanout_net_32 ), .A3(_02526_ ), .ZN(_02527_ ) );
MUX2_X1 _10121_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02528_ ) );
MUX2_X1 _10122_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02529_ ) );
MUX2_X1 _10123_ ( .A(_02528_ ), .B(_02529_ ), .S(fanout_net_29 ), .Z(_02530_ ) );
OAI211_X1 _10124_ ( .A(fanout_net_34 ), .B(_02527_ ), .C1(_02530_ ), .C2(fanout_net_32 ), .ZN(_02531_ ) );
OAI211_X1 _10125_ ( .A(_02522_ ), .B(_02531_ ), .C1(_02341_ ), .C2(_02415_ ), .ZN(_02532_ ) );
NAND2_X2 _10126_ ( .A1(_02513_ ), .A2(_02532_ ), .ZN(_02533_ ) );
INV_X1 _10127_ ( .A(\ID_EX_imm [19] ), .ZN(_02534_ ) );
XNOR2_X1 _10128_ ( .A(_02533_ ), .B(_02534_ ), .ZN(_02535_ ) );
AND2_X1 _10129_ ( .A1(_02512_ ), .A2(_02535_ ), .ZN(_02536_ ) );
OR3_X1 _10130_ ( .A1(_02385_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02386_ ), .ZN(_02537_ ) );
OR2_X1 _10131_ ( .A1(_02299_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02538_ ) );
OAI211_X1 _10132_ ( .A(_02538_ ), .B(fanout_net_29 ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02539_ ) );
OR2_X1 _10133_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02540_ ) );
OAI211_X1 _10134_ ( .A(_02540_ ), .B(_02364_ ), .C1(_02287_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02541_ ) );
NAND3_X1 _10135_ ( .A1(_02539_ ), .A2(_02383_ ), .A3(_02541_ ), .ZN(_02542_ ) );
MUX2_X1 _10136_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02543_ ) );
MUX2_X1 _10137_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02544_ ) );
MUX2_X1 _10138_ ( .A(_02543_ ), .B(_02544_ ), .S(_02364_ ), .Z(_02545_ ) );
OAI211_X1 _10139_ ( .A(_02315_ ), .B(_02542_ ), .C1(_02545_ ), .C2(_02324_ ), .ZN(_02546_ ) );
OR2_X1 _10140_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02547_ ) );
OAI211_X1 _10141_ ( .A(_02547_ ), .B(fanout_net_29 ), .C1(_02287_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02548_ ) );
OR2_X1 _10142_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02549_ ) );
OAI211_X1 _10143_ ( .A(_02549_ ), .B(_02364_ ), .C1(_02287_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02550_ ) );
NAND3_X1 _10144_ ( .A1(_02548_ ), .A2(_02550_ ), .A3(fanout_net_32 ), .ZN(_02551_ ) );
MUX2_X1 _10145_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02552_ ) );
MUX2_X1 _10146_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02553_ ) );
MUX2_X1 _10147_ ( .A(_02552_ ), .B(_02553_ ), .S(fanout_net_29 ), .Z(_02554_ ) );
OAI211_X1 _10148_ ( .A(fanout_net_34 ), .B(_02551_ ), .C1(_02554_ ), .C2(fanout_net_32 ), .ZN(_02555_ ) );
OAI211_X1 _10149_ ( .A(_02546_ ), .B(_02555_ ), .C1(_02385_ ), .C2(_02386_ ), .ZN(_02556_ ) );
NAND2_X2 _10150_ ( .A1(_02537_ ), .A2(_02556_ ), .ZN(_02557_ ) );
INV_X1 _10151_ ( .A(\ID_EX_imm [17] ), .ZN(_02558_ ) );
XNOR2_X2 _10152_ ( .A(_02557_ ), .B(_02558_ ), .ZN(_02559_ ) );
OR3_X1 _10153_ ( .A1(_02343_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02355_ ), .ZN(_02560_ ) );
OR2_X1 _10154_ ( .A1(_02300_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02561_ ) );
OAI211_X1 _10155_ ( .A(_02561_ ), .B(_02297_ ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02562_ ) );
OR2_X1 _10156_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02563_ ) );
OAI211_X1 _10157_ ( .A(_02563_ ), .B(fanout_net_29 ), .C1(_02301_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02564_ ) );
NAND3_X1 _10158_ ( .A1(_02562_ ), .A2(_02324_ ), .A3(_02564_ ), .ZN(_02565_ ) );
MUX2_X1 _10159_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02566_ ) );
MUX2_X1 _10160_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02567_ ) );
MUX2_X1 _10161_ ( .A(_02566_ ), .B(_02567_ ), .S(_02378_ ), .Z(_02568_ ) );
OAI211_X1 _10162_ ( .A(_02315_ ), .B(_02565_ ), .C1(_02568_ ), .C2(_02324_ ), .ZN(_02569_ ) );
OR2_X1 _10163_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02570_ ) );
OAI211_X1 _10164_ ( .A(_02570_ ), .B(fanout_net_29 ), .C1(_02301_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02571_ ) );
OR2_X1 _10165_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02572_ ) );
OAI211_X1 _10166_ ( .A(_02572_ ), .B(_02297_ ), .C1(_02301_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02573_ ) );
NAND3_X1 _10167_ ( .A1(_02571_ ), .A2(_02573_ ), .A3(fanout_net_32 ), .ZN(_02574_ ) );
MUX2_X1 _10168_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02575_ ) );
MUX2_X1 _10169_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02576_ ) );
MUX2_X1 _10170_ ( .A(_02575_ ), .B(_02576_ ), .S(fanout_net_29 ), .Z(_02577_ ) );
OAI211_X1 _10171_ ( .A(fanout_net_34 ), .B(_02574_ ), .C1(_02577_ ), .C2(fanout_net_32 ), .ZN(_02578_ ) );
OAI211_X1 _10172_ ( .A(_02569_ ), .B(_02578_ ), .C1(_02343_ ), .C2(_02355_ ), .ZN(_02579_ ) );
NAND2_X2 _10173_ ( .A1(_02560_ ), .A2(_02579_ ), .ZN(_02580_ ) );
INV_X1 _10174_ ( .A(\ID_EX_imm [16] ), .ZN(_02581_ ) );
XNOR2_X1 _10175_ ( .A(_02580_ ), .B(_02581_ ), .ZN(_02582_ ) );
NAND3_X1 _10176_ ( .A1(_02536_ ), .A2(_02559_ ), .A3(_02582_ ), .ZN(_02583_ ) );
OR3_X4 _10177_ ( .A1(_02340_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02414_ ), .ZN(_02584_ ) );
OR2_X1 _10178_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02585_ ) );
OAI211_X1 _10179_ ( .A(_02585_ ), .B(_02293_ ), .C1(_02284_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02586_ ) );
OR2_X1 _10180_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02587_ ) );
BUF_X4 _10181_ ( .A(_02283_ ), .Z(_02588_ ) );
OAI211_X1 _10182_ ( .A(_02587_ ), .B(fanout_net_30 ), .C1(_02588_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02589_ ) );
NAND3_X1 _10183_ ( .A1(_02586_ ), .A2(_02589_ ), .A3(_02320_ ), .ZN(_02590_ ) );
MUX2_X1 _10184_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02591_ ) );
MUX2_X1 _10185_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02592_ ) );
MUX2_X1 _10186_ ( .A(_02591_ ), .B(_02592_ ), .S(_02293_ ), .Z(_02593_ ) );
OAI211_X1 _10187_ ( .A(_02313_ ), .B(_02590_ ), .C1(_02593_ ), .C2(_02320_ ), .ZN(_02594_ ) );
OR2_X1 _10188_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02595_ ) );
OAI211_X1 _10189_ ( .A(_02595_ ), .B(fanout_net_30 ), .C1(_02588_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02596_ ) );
OR2_X1 _10190_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02597_ ) );
OAI211_X1 _10191_ ( .A(_02597_ ), .B(_02293_ ), .C1(_02588_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02598_ ) );
NAND3_X1 _10192_ ( .A1(_02596_ ), .A2(_02598_ ), .A3(fanout_net_32 ), .ZN(_02599_ ) );
MUX2_X1 _10193_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02600_ ) );
MUX2_X1 _10194_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02601_ ) );
MUX2_X1 _10195_ ( .A(_02600_ ), .B(_02601_ ), .S(fanout_net_30 ), .Z(_02602_ ) );
OAI211_X1 _10196_ ( .A(fanout_net_34 ), .B(_02599_ ), .C1(_02602_ ), .C2(fanout_net_32 ), .ZN(_02603_ ) );
OAI211_X1 _10197_ ( .A(_02594_ ), .B(_02603_ ), .C1(_02340_ ), .C2(_02414_ ), .ZN(_02604_ ) );
NAND2_X2 _10198_ ( .A1(_02584_ ), .A2(_02604_ ), .ZN(_02605_ ) );
BUF_X4 _10199_ ( .A(_02605_ ), .Z(_02606_ ) );
XOR2_X1 _10200_ ( .A(_02606_ ), .B(\ID_EX_imm [15] ), .Z(_02607_ ) );
OR3_X1 _10201_ ( .A1(_02341_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02415_ ), .ZN(_02608_ ) );
OR2_X1 _10202_ ( .A1(_02284_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02609_ ) );
OAI211_X1 _10203_ ( .A(_02609_ ), .B(_02491_ ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02610_ ) );
OR2_X1 _10204_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02611_ ) );
OAI211_X1 _10205_ ( .A(_02611_ ), .B(fanout_net_30 ), .C1(_02298_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02612_ ) );
NAND3_X1 _10206_ ( .A1(_02610_ ), .A2(fanout_net_32 ), .A3(_02612_ ), .ZN(_02613_ ) );
MUX2_X1 _10207_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02614_ ) );
MUX2_X1 _10208_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02615_ ) );
MUX2_X1 _10209_ ( .A(_02614_ ), .B(_02615_ ), .S(_02491_ ), .Z(_02616_ ) );
OAI211_X1 _10210_ ( .A(_02314_ ), .B(_02613_ ), .C1(_02616_ ), .C2(fanout_net_32 ), .ZN(_02617_ ) );
NOR2_X1 _10211_ ( .A1(_02298_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02618_ ) );
OAI21_X1 _10212_ ( .A(fanout_net_30 ), .B1(fanout_net_24 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02619_ ) );
NOR2_X1 _10213_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02620_ ) );
OAI21_X1 _10214_ ( .A(_02491_ ), .B1(_02298_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02621_ ) );
OAI221_X1 _10215_ ( .A(_02322_ ), .B1(_02618_ ), .B2(_02619_ ), .C1(_02620_ ), .C2(_02621_ ), .ZN(_02622_ ) );
MUX2_X1 _10216_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02623_ ) );
MUX2_X1 _10217_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02624_ ) );
MUX2_X1 _10218_ ( .A(_02623_ ), .B(_02624_ ), .S(fanout_net_30 ), .Z(_02625_ ) );
OAI211_X1 _10219_ ( .A(fanout_net_34 ), .B(_02622_ ), .C1(_02625_ ), .C2(_02322_ ), .ZN(_02626_ ) );
OAI211_X1 _10220_ ( .A(_02617_ ), .B(_02626_ ), .C1(_02341_ ), .C2(_02415_ ), .ZN(_02627_ ) );
NAND2_X1 _10221_ ( .A1(_02608_ ), .A2(_02627_ ), .ZN(_02628_ ) );
BUF_X2 _10222_ ( .A(_02628_ ), .Z(_02629_ ) );
XOR2_X1 _10223_ ( .A(_02629_ ), .B(\ID_EX_imm [14] ), .Z(_02630_ ) );
AND2_X1 _10224_ ( .A1(_02607_ ), .A2(_02630_ ), .ZN(_02631_ ) );
OR2_X1 _10225_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02632_ ) );
OAI211_X1 _10226_ ( .A(_02632_ ), .B(_02293_ ), .C1(_02284_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02633_ ) );
OR2_X1 _10227_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02634_ ) );
OAI211_X1 _10228_ ( .A(_02634_ ), .B(fanout_net_30 ), .C1(_02588_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02635_ ) );
NAND3_X1 _10229_ ( .A1(_02633_ ), .A2(_02635_ ), .A3(fanout_net_32 ), .ZN(_02636_ ) );
MUX2_X1 _10230_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02637_ ) );
MUX2_X1 _10231_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02638_ ) );
MUX2_X1 _10232_ ( .A(_02637_ ), .B(_02638_ ), .S(_02293_ ), .Z(_02639_ ) );
OAI211_X1 _10233_ ( .A(_02313_ ), .B(_02636_ ), .C1(_02639_ ), .C2(fanout_net_32 ), .ZN(_02640_ ) );
INV_X1 _10234_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02641_ ) );
AOI21_X1 _10235_ ( .A(fanout_net_30 ), .B1(_02641_ ), .B2(fanout_net_24 ), .ZN(_02642_ ) );
OR2_X1 _10236_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02643_ ) );
MUX2_X1 _10237_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02644_ ) );
AOI221_X4 _10238_ ( .A(fanout_net_32 ), .B1(_02642_ ), .B2(_02643_ ), .C1(_02644_ ), .C2(fanout_net_30 ), .ZN(_02645_ ) );
MUX2_X1 _10239_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02646_ ) );
MUX2_X1 _10240_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02647_ ) );
MUX2_X1 _10241_ ( .A(_02646_ ), .B(_02647_ ), .S(fanout_net_30 ), .Z(_02648_ ) );
OAI21_X1 _10242_ ( .A(fanout_net_34 ), .B1(_02648_ ), .B2(_02320_ ), .ZN(_02649_ ) );
OAI221_X1 _10243_ ( .A(_02640_ ), .B1(_02645_ ), .B2(_02649_ ), .C1(_02340_ ), .C2(_02353_ ), .ZN(_02650_ ) );
OR3_X1 _10244_ ( .A1(_02340_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02414_ ), .ZN(_02651_ ) );
NAND2_X4 _10245_ ( .A1(_02650_ ), .A2(_02651_ ), .ZN(_02652_ ) );
XNOR2_X1 _10246_ ( .A(_02652_ ), .B(\ID_EX_imm [5] ), .ZN(_02653_ ) );
BUF_X4 _10247_ ( .A(_02339_ ), .Z(_02654_ ) );
OR3_X1 _10248_ ( .A1(_02654_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02414_ ), .ZN(_02655_ ) );
CLKBUF_X2 _10249_ ( .A(_02282_ ), .Z(_02656_ ) );
OR2_X1 _10250_ ( .A1(_02656_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02657_ ) );
OAI211_X1 _10251_ ( .A(_02657_ ), .B(_02490_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02658_ ) );
OR2_X1 _10252_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02659_ ) );
OAI211_X1 _10253_ ( .A(_02659_ ), .B(fanout_net_30 ), .C1(_02284_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02660_ ) );
NAND3_X1 _10254_ ( .A1(_02658_ ), .A2(_02321_ ), .A3(_02660_ ), .ZN(_02661_ ) );
MUX2_X1 _10255_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02662_ ) );
MUX2_X1 _10256_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02663_ ) );
MUX2_X1 _10257_ ( .A(_02662_ ), .B(_02663_ ), .S(_02490_ ), .Z(_02664_ ) );
OAI211_X1 _10258_ ( .A(_02313_ ), .B(_02661_ ), .C1(_02664_ ), .C2(_02321_ ), .ZN(_02665_ ) );
OR2_X1 _10259_ ( .A1(_02656_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02666_ ) );
OAI211_X1 _10260_ ( .A(_02666_ ), .B(fanout_net_30 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02667_ ) );
OR2_X1 _10261_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02668_ ) );
OAI211_X1 _10262_ ( .A(_02668_ ), .B(_02490_ ), .C1(_02284_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02669_ ) );
NAND3_X1 _10263_ ( .A1(_02667_ ), .A2(fanout_net_32 ), .A3(_02669_ ), .ZN(_02670_ ) );
MUX2_X1 _10264_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02671_ ) );
MUX2_X1 _10265_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02672_ ) );
MUX2_X1 _10266_ ( .A(_02671_ ), .B(_02672_ ), .S(fanout_net_30 ), .Z(_02673_ ) );
OAI211_X1 _10267_ ( .A(fanout_net_34 ), .B(_02670_ ), .C1(_02673_ ), .C2(fanout_net_33 ), .ZN(_02674_ ) );
OAI211_X1 _10268_ ( .A(_02665_ ), .B(_02674_ ), .C1(_02654_ ), .C2(_02353_ ), .ZN(_02675_ ) );
NAND2_X2 _10269_ ( .A1(_02655_ ), .A2(_02675_ ), .ZN(_02676_ ) );
BUF_X4 _10270_ ( .A(_02676_ ), .Z(_02677_ ) );
AND2_X1 _10271_ ( .A1(_02677_ ), .A2(\ID_EX_imm [4] ), .ZN(_02678_ ) );
INV_X1 _10272_ ( .A(_02678_ ), .ZN(_02679_ ) );
NOR2_X1 _10273_ ( .A1(_02653_ ), .A2(_02679_ ), .ZN(_02680_ ) );
INV_X1 _10274_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02681_ ) );
AOI21_X1 _10275_ ( .A(_02680_ ), .B1(_02681_ ), .B2(_02652_ ), .ZN(_02682_ ) );
NOR2_X2 _10276_ ( .A1(_02340_ ), .A2(_02414_ ), .ZN(_02683_ ) );
NAND2_X2 _10277_ ( .A1(_02683_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02684_ ) );
OR2_X1 _10278_ ( .A1(_02283_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02685_ ) );
OAI211_X1 _10279_ ( .A(_02685_ ), .B(_02292_ ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02686_ ) );
OR2_X1 _10280_ ( .A1(fanout_net_24 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02687_ ) );
OAI211_X1 _10281_ ( .A(_02687_ ), .B(fanout_net_30 ), .C1(_02656_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02688_ ) );
NAND3_X1 _10282_ ( .A1(_02686_ ), .A2(_02319_ ), .A3(_02688_ ), .ZN(_02689_ ) );
MUX2_X1 _10283_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02690_ ) );
MUX2_X1 _10284_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02691_ ) );
MUX2_X1 _10285_ ( .A(_02690_ ), .B(_02691_ ), .S(_02292_ ), .Z(_02692_ ) );
OAI211_X1 _10286_ ( .A(_02313_ ), .B(_02689_ ), .C1(_02692_ ), .C2(_02320_ ), .ZN(_02693_ ) );
OR2_X1 _10287_ ( .A1(fanout_net_24 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02694_ ) );
OAI211_X1 _10288_ ( .A(_02694_ ), .B(fanout_net_30 ), .C1(_02656_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02695_ ) );
OR2_X1 _10289_ ( .A1(fanout_net_24 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02696_ ) );
OAI211_X1 _10290_ ( .A(_02696_ ), .B(_02292_ ), .C1(_02283_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02697_ ) );
NAND3_X1 _10291_ ( .A1(_02695_ ), .A2(_02697_ ), .A3(fanout_net_33 ), .ZN(_02698_ ) );
MUX2_X1 _10292_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02699_ ) );
MUX2_X1 _10293_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02700_ ) );
MUX2_X1 _10294_ ( .A(_02699_ ), .B(_02700_ ), .S(fanout_net_30 ), .Z(_02701_ ) );
OAI211_X1 _10295_ ( .A(fanout_net_34 ), .B(_02698_ ), .C1(_02701_ ), .C2(fanout_net_33 ), .ZN(_02702_ ) );
NAND2_X1 _10296_ ( .A1(_02693_ ), .A2(_02702_ ), .ZN(_02703_ ) );
OAI21_X1 _10297_ ( .A(_02703_ ), .B1(_02340_ ), .B2(_02414_ ), .ZN(_02704_ ) );
AND2_X2 _10298_ ( .A1(_02684_ ), .A2(_02704_ ), .ZN(_02705_ ) );
BUF_X8 _10299_ ( .A(_02705_ ), .Z(_02706_ ) );
XNOR2_X1 _10300_ ( .A(_02706_ ), .B(\ID_EX_imm [7] ), .ZN(_02707_ ) );
INV_X1 _10301_ ( .A(_02707_ ), .ZN(_02708_ ) );
OR3_X1 _10302_ ( .A1(_02341_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02415_ ), .ZN(_02709_ ) );
OR2_X1 _10303_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02710_ ) );
OAI211_X1 _10304_ ( .A(_02710_ ), .B(_02295_ ), .C1(_02299_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02711_ ) );
OR2_X1 _10305_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02712_ ) );
OAI211_X1 _10306_ ( .A(_02712_ ), .B(fanout_net_30 ), .C1(_02285_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02713_ ) );
NAND3_X1 _10307_ ( .A1(_02711_ ), .A2(_02713_ ), .A3(_02322_ ), .ZN(_02714_ ) );
MUX2_X1 _10308_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02715_ ) );
MUX2_X1 _10309_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02716_ ) );
MUX2_X1 _10310_ ( .A(_02715_ ), .B(_02716_ ), .S(_02491_ ), .Z(_02717_ ) );
OAI211_X1 _10311_ ( .A(_02314_ ), .B(_02714_ ), .C1(_02717_ ), .C2(_02323_ ), .ZN(_02718_ ) );
OR2_X1 _10312_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02719_ ) );
OAI211_X1 _10313_ ( .A(_02719_ ), .B(fanout_net_30 ), .C1(_02299_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02720_ ) );
OR2_X1 _10314_ ( .A1(fanout_net_25 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02721_ ) );
OAI211_X1 _10315_ ( .A(_02721_ ), .B(_02295_ ), .C1(_02285_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02722_ ) );
NAND3_X1 _10316_ ( .A1(_02720_ ), .A2(_02722_ ), .A3(fanout_net_33 ), .ZN(_02723_ ) );
MUX2_X1 _10317_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02724_ ) );
MUX2_X1 _10318_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02725_ ) );
MUX2_X1 _10319_ ( .A(_02724_ ), .B(_02725_ ), .S(fanout_net_30 ), .Z(_02726_ ) );
OAI211_X1 _10320_ ( .A(fanout_net_34 ), .B(_02723_ ), .C1(_02726_ ), .C2(fanout_net_33 ), .ZN(_02727_ ) );
OAI211_X1 _10321_ ( .A(_02718_ ), .B(_02727_ ), .C1(_02342_ ), .C2(_02354_ ), .ZN(_02728_ ) );
NAND2_X2 _10322_ ( .A1(_02709_ ), .A2(_02728_ ), .ZN(_02729_ ) );
INV_X1 _10323_ ( .A(\ID_EX_imm [6] ), .ZN(_02730_ ) );
XNOR2_X1 _10324_ ( .A(_02729_ ), .B(_02730_ ), .ZN(_02731_ ) );
NAND2_X1 _10325_ ( .A1(_02708_ ), .A2(_02731_ ), .ZN(_02732_ ) );
OR2_X1 _10326_ ( .A1(_02682_ ), .A2(_02732_ ), .ZN(_02733_ ) );
INV_X2 _10327_ ( .A(_02706_ ), .ZN(_02734_ ) );
OR2_X1 _10328_ ( .A1(_02734_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02735_ ) );
NAND2_X1 _10329_ ( .A1(_02729_ ), .A2(\ID_EX_imm [6] ), .ZN(_02736_ ) );
OR2_X1 _10330_ ( .A1(_02707_ ), .A2(_02736_ ), .ZN(_02737_ ) );
AND3_X1 _10331_ ( .A1(_02733_ ), .A2(_02735_ ), .A3(_02737_ ), .ZN(_02738_ ) );
OR3_X4 _10332_ ( .A1(_02339_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02352_ ), .ZN(_02739_ ) );
OR2_X1 _10333_ ( .A1(fanout_net_25 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02740_ ) );
OAI211_X1 _10334_ ( .A(_02740_ ), .B(_02291_ ), .C1(_02282_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02741_ ) );
OR2_X1 _10335_ ( .A1(fanout_net_25 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02742_ ) );
OAI211_X1 _10336_ ( .A(_02742_ ), .B(fanout_net_30 ), .C1(_02282_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02743_ ) );
NAND3_X1 _10337_ ( .A1(_02741_ ), .A2(_02743_ ), .A3(_02319_ ), .ZN(_02744_ ) );
MUX2_X1 _10338_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02745_ ) );
MUX2_X1 _10339_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02746_ ) );
MUX2_X1 _10340_ ( .A(_02745_ ), .B(_02746_ ), .S(_02291_ ), .Z(_02747_ ) );
OAI211_X1 _10341_ ( .A(fanout_net_34 ), .B(_02744_ ), .C1(_02747_ ), .C2(_02319_ ), .ZN(_02748_ ) );
NOR2_X1 _10342_ ( .A1(_02281_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02749_ ) );
OAI21_X1 _10343_ ( .A(fanout_net_30 ), .B1(fanout_net_25 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02750_ ) );
NOR2_X1 _10344_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(fanout_net_25 ), .ZN(_02751_ ) );
OAI21_X1 _10345_ ( .A(_02291_ ), .B1(_02281_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02752_ ) );
OAI221_X1 _10346_ ( .A(_02319_ ), .B1(_02749_ ), .B2(_02750_ ), .C1(_02751_ ), .C2(_02752_ ), .ZN(_02753_ ) );
MUX2_X1 _10347_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02754_ ) );
MUX2_X1 _10348_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02755_ ) );
MUX2_X1 _10349_ ( .A(_02754_ ), .B(_02755_ ), .S(_02291_ ), .Z(_02756_ ) );
OAI211_X1 _10350_ ( .A(_02312_ ), .B(_02753_ ), .C1(_02756_ ), .C2(_02319_ ), .ZN(_02757_ ) );
OAI211_X4 _10351_ ( .A(_02748_ ), .B(_02757_ ), .C1(_02339_ ), .C2(_02352_ ), .ZN(_02758_ ) );
AOI21_X1 _10352_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B1(_02739_ ), .B2(_02758_ ), .ZN(_02759_ ) );
NAND2_X4 _10353_ ( .A1(_02739_ ), .A2(_02758_ ), .ZN(_02760_ ) );
INV_X1 _10354_ ( .A(\ID_EX_imm [1] ), .ZN(_02761_ ) );
XNOR2_X1 _10355_ ( .A(_02760_ ), .B(_02761_ ), .ZN(_02762_ ) );
INV_X1 _10356_ ( .A(\ID_EX_imm [0] ), .ZN(_02763_ ) );
OR3_X2 _10357_ ( .A1(_02339_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_02352_ ), .ZN(_02764_ ) );
OR2_X1 _10358_ ( .A1(fanout_net_25 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02765_ ) );
OAI211_X1 _10359_ ( .A(_02765_ ), .B(_02291_ ), .C1(_02282_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02766_ ) );
OR2_X1 _10360_ ( .A1(fanout_net_25 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02767_ ) );
OAI211_X1 _10361_ ( .A(_02767_ ), .B(fanout_net_30 ), .C1(_02282_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02768_ ) );
NAND3_X1 _10362_ ( .A1(_02766_ ), .A2(_02768_ ), .A3(fanout_net_33 ), .ZN(_02769_ ) );
MUX2_X1 _10363_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02770_ ) );
MUX2_X1 _10364_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02771_ ) );
MUX2_X1 _10365_ ( .A(_02770_ ), .B(_02771_ ), .S(_02291_ ), .Z(_02772_ ) );
OAI211_X1 _10366_ ( .A(_02312_ ), .B(_02769_ ), .C1(_02772_ ), .C2(fanout_net_33 ), .ZN(_02773_ ) );
NOR2_X1 _10367_ ( .A1(_02282_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02774_ ) );
OAI21_X1 _10368_ ( .A(fanout_net_30 ), .B1(fanout_net_25 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02775_ ) );
NOR2_X1 _10369_ ( .A1(fanout_net_25 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02776_ ) );
OAI21_X1 _10370_ ( .A(_02291_ ), .B1(_02282_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02777_ ) );
OAI221_X1 _10371_ ( .A(_02319_ ), .B1(_02774_ ), .B2(_02775_ ), .C1(_02776_ ), .C2(_02777_ ), .ZN(_02778_ ) );
MUX2_X1 _10372_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02779_ ) );
MUX2_X1 _10373_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02780_ ) );
MUX2_X1 _10374_ ( .A(_02779_ ), .B(_02780_ ), .S(fanout_net_30 ), .Z(_02781_ ) );
OAI211_X1 _10375_ ( .A(fanout_net_34 ), .B(_02778_ ), .C1(_02781_ ), .C2(_02319_ ), .ZN(_02782_ ) );
OAI211_X1 _10376_ ( .A(_02773_ ), .B(_02782_ ), .C1(_02339_ ), .C2(_02352_ ), .ZN(_02783_ ) );
AOI21_X1 _10377_ ( .A(_02763_ ), .B1(_02764_ ), .B2(_02783_ ), .ZN(_02784_ ) );
AOI21_X1 _10378_ ( .A(_02759_ ), .B1(_02762_ ), .B2(_02784_ ), .ZN(_02785_ ) );
OR3_X1 _10379_ ( .A1(_02339_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02352_ ), .ZN(_02786_ ) );
OR2_X1 _10380_ ( .A1(fanout_net_25 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02787_ ) );
OAI211_X1 _10381_ ( .A(_02787_ ), .B(_02292_ ), .C1(_02283_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02788_ ) );
OR2_X1 _10382_ ( .A1(fanout_net_25 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02789_ ) );
OAI211_X1 _10383_ ( .A(_02789_ ), .B(fanout_net_30 ), .C1(_02283_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02790_ ) );
NAND3_X1 _10384_ ( .A1(_02788_ ), .A2(_02790_ ), .A3(_02319_ ), .ZN(_02791_ ) );
MUX2_X1 _10385_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02792_ ) );
MUX2_X1 _10386_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02793_ ) );
MUX2_X1 _10387_ ( .A(_02792_ ), .B(_02793_ ), .S(_02292_ ), .Z(_02794_ ) );
OAI211_X1 _10388_ ( .A(_02312_ ), .B(_02791_ ), .C1(_02794_ ), .C2(_02320_ ), .ZN(_02795_ ) );
OR2_X1 _10389_ ( .A1(_02282_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02796_ ) );
OAI211_X1 _10390_ ( .A(_02796_ ), .B(fanout_net_30 ), .C1(fanout_net_26 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02797_ ) );
OR2_X1 _10391_ ( .A1(fanout_net_26 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02798_ ) );
OAI211_X1 _10392_ ( .A(_02798_ ), .B(_02292_ ), .C1(_02283_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02799_ ) );
NAND3_X1 _10393_ ( .A1(_02797_ ), .A2(fanout_net_33 ), .A3(_02799_ ), .ZN(_02800_ ) );
MUX2_X1 _10394_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02801_ ) );
MUX2_X1 _10395_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02802_ ) );
MUX2_X1 _10396_ ( .A(_02801_ ), .B(_02802_ ), .S(fanout_net_30 ), .Z(_02803_ ) );
OAI211_X1 _10397_ ( .A(fanout_net_34 ), .B(_02800_ ), .C1(_02803_ ), .C2(fanout_net_33 ), .ZN(_02804_ ) );
OAI211_X1 _10398_ ( .A(_02795_ ), .B(_02804_ ), .C1(_02339_ ), .C2(_02352_ ), .ZN(_02805_ ) );
NAND2_X4 _10399_ ( .A1(_02786_ ), .A2(_02805_ ), .ZN(_02806_ ) );
XOR2_X1 _10400_ ( .A(_02806_ ), .B(\ID_EX_imm [2] ), .Z(_02807_ ) );
INV_X1 _10401_ ( .A(_02807_ ), .ZN(_02808_ ) );
OR3_X2 _10402_ ( .A1(_02340_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02414_ ), .ZN(_02809_ ) );
OR2_X1 _10403_ ( .A1(fanout_net_26 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02810_ ) );
OAI211_X1 _10404_ ( .A(_02810_ ), .B(_02293_ ), .C1(_02588_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02811_ ) );
OR2_X1 _10405_ ( .A1(fanout_net_26 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02812_ ) );
OAI211_X1 _10406_ ( .A(_02812_ ), .B(fanout_net_30 ), .C1(_02588_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02813_ ) );
NAND3_X1 _10407_ ( .A1(_02811_ ), .A2(_02813_ ), .A3(_02320_ ), .ZN(_02814_ ) );
MUX2_X1 _10408_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02815_ ) );
MUX2_X1 _10409_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02816_ ) );
MUX2_X1 _10410_ ( .A(_02815_ ), .B(_02816_ ), .S(_02293_ ), .Z(_02817_ ) );
OAI211_X1 _10411_ ( .A(_02313_ ), .B(_02814_ ), .C1(_02817_ ), .C2(_02320_ ), .ZN(_02818_ ) );
OR2_X1 _10412_ ( .A1(fanout_net_26 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02819_ ) );
OAI211_X1 _10413_ ( .A(_02819_ ), .B(fanout_net_30 ), .C1(_02588_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02820_ ) );
OR2_X1 _10414_ ( .A1(fanout_net_26 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02821_ ) );
OAI211_X1 _10415_ ( .A(_02821_ ), .B(_02293_ ), .C1(_02656_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02822_ ) );
NAND3_X1 _10416_ ( .A1(_02820_ ), .A2(_02822_ ), .A3(fanout_net_33 ), .ZN(_02823_ ) );
MUX2_X1 _10417_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02824_ ) );
MUX2_X1 _10418_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02825_ ) );
MUX2_X1 _10419_ ( .A(_02824_ ), .B(_02825_ ), .S(fanout_net_30 ), .Z(_02826_ ) );
OAI211_X1 _10420_ ( .A(fanout_net_34 ), .B(_02823_ ), .C1(_02826_ ), .C2(fanout_net_33 ), .ZN(_02827_ ) );
OAI211_X1 _10421_ ( .A(_02818_ ), .B(_02827_ ), .C1(_02340_ ), .C2(_02414_ ), .ZN(_02828_ ) );
NAND2_X4 _10422_ ( .A1(_02809_ ), .A2(_02828_ ), .ZN(_02829_ ) );
XNOR2_X1 _10423_ ( .A(_02829_ ), .B(\ID_EX_imm [3] ), .ZN(_02830_ ) );
NOR3_X2 _10424_ ( .A1(_02785_ ), .A2(_02808_ ), .A3(_02830_ ), .ZN(_02831_ ) );
NAND2_X1 _10425_ ( .A1(_02806_ ), .A2(\ID_EX_imm [2] ), .ZN(_02832_ ) );
INV_X4 _10426_ ( .A(_02829_ ), .ZN(_02833_ ) );
OAI22_X1 _10427_ ( .A1(_02830_ ), .A2(_02832_ ), .B1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B2(_02833_ ), .ZN(_02834_ ) );
OR2_X1 _10428_ ( .A1(_02831_ ), .A2(_02834_ ), .ZN(_02835_ ) );
INV_X1 _10429_ ( .A(_02653_ ), .ZN(_02836_ ) );
XOR2_X1 _10430_ ( .A(_02677_ ), .B(\ID_EX_imm [4] ), .Z(_02837_ ) );
AND2_X1 _10431_ ( .A1(_02836_ ), .A2(_02837_ ), .ZN(_02838_ ) );
NAND4_X1 _10432_ ( .A1(_02835_ ), .A2(_02708_ ), .A3(_02731_ ), .A4(_02838_ ), .ZN(_02839_ ) );
AND2_X2 _10433_ ( .A1(_02738_ ), .A2(_02839_ ), .ZN(_02840_ ) );
INV_X1 _10434_ ( .A(_02840_ ), .ZN(_02841_ ) );
OR3_X1 _10435_ ( .A1(_02654_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02353_ ), .ZN(_02842_ ) );
OR2_X1 _10436_ ( .A1(_02656_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02843_ ) );
OAI211_X1 _10437_ ( .A(_02843_ ), .B(_02490_ ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02844_ ) );
OR2_X1 _10438_ ( .A1(_02656_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02845_ ) );
OAI211_X1 _10439_ ( .A(_02845_ ), .B(fanout_net_31 ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02846_ ) );
NAND3_X1 _10440_ ( .A1(_02844_ ), .A2(_02846_ ), .A3(fanout_net_33 ), .ZN(_02847_ ) );
MUX2_X1 _10441_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02848_ ) );
MUX2_X1 _10442_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02849_ ) );
MUX2_X1 _10443_ ( .A(_02848_ ), .B(_02849_ ), .S(_02490_ ), .Z(_02850_ ) );
OAI211_X1 _10444_ ( .A(_02313_ ), .B(_02847_ ), .C1(_02850_ ), .C2(fanout_net_33 ), .ZN(_02851_ ) );
NOR2_X1 _10445_ ( .A1(_02284_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02852_ ) );
OAI21_X1 _10446_ ( .A(fanout_net_31 ), .B1(fanout_net_26 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02853_ ) );
NOR2_X1 _10447_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02854_ ) );
OAI21_X1 _10448_ ( .A(_02490_ ), .B1(_02284_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02855_ ) );
OAI221_X1 _10449_ ( .A(_02320_ ), .B1(_02852_ ), .B2(_02853_ ), .C1(_02854_ ), .C2(_02855_ ), .ZN(_02856_ ) );
MUX2_X1 _10450_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02857_ ) );
MUX2_X1 _10451_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02858_ ) );
MUX2_X1 _10452_ ( .A(_02857_ ), .B(_02858_ ), .S(fanout_net_31 ), .Z(_02859_ ) );
OAI211_X1 _10453_ ( .A(fanout_net_34 ), .B(_02856_ ), .C1(_02859_ ), .C2(_02321_ ), .ZN(_02860_ ) );
OAI211_X1 _10454_ ( .A(_02851_ ), .B(_02860_ ), .C1(_02654_ ), .C2(_02353_ ), .ZN(_02861_ ) );
NAND2_X1 _10455_ ( .A1(_02842_ ), .A2(_02861_ ), .ZN(_02862_ ) );
BUF_X4 _10456_ ( .A(_02862_ ), .Z(_02863_ ) );
INV_X1 _10457_ ( .A(\ID_EX_imm [12] ), .ZN(_02864_ ) );
XNOR2_X1 _10458_ ( .A(_02863_ ), .B(_02864_ ), .ZN(_02865_ ) );
OR3_X1 _10459_ ( .A1(_02654_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02353_ ), .ZN(_02866_ ) );
INV_X1 _10460_ ( .A(\ID_EX_imm [13] ), .ZN(_02867_ ) );
OR2_X1 _10461_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02868_ ) );
OAI211_X1 _10462_ ( .A(_02868_ ), .B(_02294_ ), .C1(_02298_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02869_ ) );
OR2_X1 _10463_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02870_ ) );
BUF_X4 _10464_ ( .A(_02588_ ), .Z(_02871_ ) );
OAI211_X1 _10465_ ( .A(_02870_ ), .B(fanout_net_31 ), .C1(_02871_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02872_ ) );
NAND3_X1 _10466_ ( .A1(_02869_ ), .A2(_02872_ ), .A3(_02321_ ), .ZN(_02873_ ) );
MUX2_X1 _10467_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02874_ ) );
MUX2_X1 _10468_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02875_ ) );
MUX2_X1 _10469_ ( .A(_02874_ ), .B(_02875_ ), .S(_02294_ ), .Z(_02876_ ) );
OAI211_X1 _10470_ ( .A(_02314_ ), .B(_02873_ ), .C1(_02876_ ), .C2(_02322_ ), .ZN(_02877_ ) );
OR2_X1 _10471_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02878_ ) );
OAI211_X1 _10472_ ( .A(_02878_ ), .B(fanout_net_31 ), .C1(_02871_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02879_ ) );
OR2_X1 _10473_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02880_ ) );
OAI211_X1 _10474_ ( .A(_02880_ ), .B(_02294_ ), .C1(_02871_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02881_ ) );
NAND3_X1 _10475_ ( .A1(_02879_ ), .A2(_02881_ ), .A3(fanout_net_33 ), .ZN(_02882_ ) );
MUX2_X1 _10476_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02883_ ) );
MUX2_X1 _10477_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02884_ ) );
MUX2_X1 _10478_ ( .A(_02883_ ), .B(_02884_ ), .S(fanout_net_31 ), .Z(_02885_ ) );
OAI211_X1 _10479_ ( .A(fanout_net_34 ), .B(_02882_ ), .C1(_02885_ ), .C2(fanout_net_33 ), .ZN(_02886_ ) );
OAI211_X1 _10480_ ( .A(_02877_ ), .B(_02886_ ), .C1(_02341_ ), .C2(_02415_ ), .ZN(_02887_ ) );
AND3_X1 _10481_ ( .A1(_02866_ ), .A2(_02867_ ), .A3(_02887_ ), .ZN(_02888_ ) );
AOI21_X1 _10482_ ( .A(_02867_ ), .B1(_02866_ ), .B2(_02887_ ), .ZN(_02889_ ) );
NOR2_X1 _10483_ ( .A1(_02888_ ), .A2(_02889_ ), .ZN(_02890_ ) );
AND2_X1 _10484_ ( .A1(_02865_ ), .A2(_02890_ ), .ZN(_02891_ ) );
OR3_X1 _10485_ ( .A1(_02654_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02353_ ), .ZN(_02892_ ) );
OR2_X1 _10486_ ( .A1(fanout_net_26 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02893_ ) );
OAI211_X1 _10487_ ( .A(_02893_ ), .B(_02294_ ), .C1(_02871_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02894_ ) );
OR2_X1 _10488_ ( .A1(fanout_net_26 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02895_ ) );
OAI211_X1 _10489_ ( .A(_02895_ ), .B(fanout_net_31 ), .C1(_02871_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02896_ ) );
NAND3_X1 _10490_ ( .A1(_02894_ ), .A2(_02896_ ), .A3(_02321_ ), .ZN(_02897_ ) );
MUX2_X1 _10491_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02898_ ) );
MUX2_X1 _10492_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02899_ ) );
MUX2_X1 _10493_ ( .A(_02898_ ), .B(_02899_ ), .S(_02490_ ), .Z(_02900_ ) );
OAI211_X1 _10494_ ( .A(_02313_ ), .B(_02897_ ), .C1(_02900_ ), .C2(_02321_ ), .ZN(_02901_ ) );
OR2_X1 _10495_ ( .A1(_02656_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02902_ ) );
OAI211_X1 _10496_ ( .A(_02902_ ), .B(_02294_ ), .C1(fanout_net_27 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02903_ ) );
OR2_X1 _10497_ ( .A1(fanout_net_27 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02904_ ) );
OAI211_X1 _10498_ ( .A(_02904_ ), .B(fanout_net_31 ), .C1(_02871_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02905_ ) );
NAND3_X1 _10499_ ( .A1(_02903_ ), .A2(fanout_net_33 ), .A3(_02905_ ), .ZN(_02906_ ) );
MUX2_X1 _10500_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02907_ ) );
MUX2_X1 _10501_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02908_ ) );
MUX2_X1 _10502_ ( .A(_02907_ ), .B(_02908_ ), .S(fanout_net_31 ), .Z(_02909_ ) );
OAI211_X1 _10503_ ( .A(fanout_net_34 ), .B(_02906_ ), .C1(_02909_ ), .C2(fanout_net_33 ), .ZN(_02910_ ) );
OAI211_X1 _10504_ ( .A(_02901_ ), .B(_02910_ ), .C1(_02654_ ), .C2(_02353_ ), .ZN(_02911_ ) );
NAND2_X2 _10505_ ( .A1(_02892_ ), .A2(_02911_ ), .ZN(_02912_ ) );
INV_X1 _10506_ ( .A(\ID_EX_imm [10] ), .ZN(_02913_ ) );
XNOR2_X1 _10507_ ( .A(_02912_ ), .B(_02913_ ), .ZN(_02914_ ) );
OR3_X2 _10508_ ( .A1(_02654_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_02353_ ), .ZN(_02915_ ) );
OR2_X1 _10509_ ( .A1(_02588_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02916_ ) );
OAI211_X1 _10510_ ( .A(_02916_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02917_ ) );
OR2_X1 _10511_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02918_ ) );
OAI211_X1 _10512_ ( .A(_02918_ ), .B(_02294_ ), .C1(_02871_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02919_ ) );
NAND3_X1 _10513_ ( .A1(_02917_ ), .A2(_02321_ ), .A3(_02919_ ), .ZN(_02920_ ) );
MUX2_X1 _10514_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02921_ ) );
MUX2_X1 _10515_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02922_ ) );
MUX2_X1 _10516_ ( .A(_02921_ ), .B(_02922_ ), .S(_02294_ ), .Z(_02923_ ) );
OAI211_X1 _10517_ ( .A(_02313_ ), .B(_02920_ ), .C1(_02923_ ), .C2(_02322_ ), .ZN(_02924_ ) );
OR2_X1 _10518_ ( .A1(_02588_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02925_ ) );
OAI211_X1 _10519_ ( .A(_02925_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02926_ ) );
OR2_X1 _10520_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02927_ ) );
OAI211_X1 _10521_ ( .A(_02927_ ), .B(_02294_ ), .C1(_02871_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02928_ ) );
NAND3_X1 _10522_ ( .A1(_02926_ ), .A2(fanout_net_33 ), .A3(_02928_ ), .ZN(_02929_ ) );
MUX2_X1 _10523_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02930_ ) );
MUX2_X1 _10524_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02931_ ) );
MUX2_X1 _10525_ ( .A(_02930_ ), .B(_02931_ ), .S(fanout_net_31 ), .Z(_02932_ ) );
OAI211_X1 _10526_ ( .A(fanout_net_34 ), .B(_02929_ ), .C1(_02932_ ), .C2(fanout_net_33 ), .ZN(_02933_ ) );
OAI211_X4 _10527_ ( .A(_02924_ ), .B(_02933_ ), .C1(_02341_ ), .C2(_02415_ ), .ZN(_02934_ ) );
NAND2_X2 _10528_ ( .A1(_02915_ ), .A2(_02934_ ), .ZN(_02935_ ) );
BUF_X4 _10529_ ( .A(_02935_ ), .Z(_02936_ ) );
INV_X1 _10530_ ( .A(\ID_EX_imm [11] ), .ZN(_02937_ ) );
XNOR2_X1 _10531_ ( .A(_02936_ ), .B(_02937_ ), .ZN(_02938_ ) );
AND2_X1 _10532_ ( .A1(_02914_ ), .A2(_02938_ ), .ZN(_02939_ ) );
OR3_X4 _10533_ ( .A1(_02654_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02353_ ), .ZN(_02940_ ) );
OR2_X1 _10534_ ( .A1(_02656_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02941_ ) );
OAI211_X1 _10535_ ( .A(_02941_ ), .B(_02294_ ), .C1(fanout_net_27 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02942_ ) );
OR2_X1 _10536_ ( .A1(_02656_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02943_ ) );
OAI211_X1 _10537_ ( .A(_02943_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02944_ ) );
NAND3_X1 _10538_ ( .A1(_02942_ ), .A2(_02944_ ), .A3(_02321_ ), .ZN(_02945_ ) );
MUX2_X1 _10539_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02946_ ) );
MUX2_X1 _10540_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02947_ ) );
MUX2_X1 _10541_ ( .A(_02946_ ), .B(_02947_ ), .S(_02490_ ), .Z(_02948_ ) );
OAI211_X1 _10542_ ( .A(_02313_ ), .B(_02945_ ), .C1(_02948_ ), .C2(_02321_ ), .ZN(_02949_ ) );
OR2_X1 _10543_ ( .A1(fanout_net_27 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02950_ ) );
OAI211_X1 _10544_ ( .A(_02950_ ), .B(fanout_net_31 ), .C1(_02871_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02951_ ) );
OR2_X1 _10545_ ( .A1(fanout_net_27 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02952_ ) );
OAI211_X1 _10546_ ( .A(_02952_ ), .B(_02490_ ), .C1(_02871_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02953_ ) );
NAND3_X1 _10547_ ( .A1(_02951_ ), .A2(_02953_ ), .A3(fanout_net_33 ), .ZN(_02954_ ) );
MUX2_X1 _10548_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02955_ ) );
MUX2_X1 _10549_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02956_ ) );
MUX2_X1 _10550_ ( .A(_02955_ ), .B(_02956_ ), .S(fanout_net_31 ), .Z(_02957_ ) );
OAI211_X1 _10551_ ( .A(fanout_net_34 ), .B(_02954_ ), .C1(_02957_ ), .C2(fanout_net_33 ), .ZN(_02958_ ) );
OAI211_X1 _10552_ ( .A(_02949_ ), .B(_02958_ ), .C1(_02654_ ), .C2(_02415_ ), .ZN(_02959_ ) );
NAND2_X2 _10553_ ( .A1(_02940_ ), .A2(_02959_ ), .ZN(_02960_ ) );
INV_X1 _10554_ ( .A(\ID_EX_imm [8] ), .ZN(_02961_ ) );
XNOR2_X1 _10555_ ( .A(_02960_ ), .B(_02961_ ), .ZN(_02962_ ) );
OR3_X1 _10556_ ( .A1(_02339_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02352_ ), .ZN(_02963_ ) );
OR2_X1 _10557_ ( .A1(fanout_net_27 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02964_ ) );
OAI211_X1 _10558_ ( .A(_02964_ ), .B(_02292_ ), .C1(_02283_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02965_ ) );
OR2_X1 _10559_ ( .A1(fanout_net_27 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02966_ ) );
OAI211_X1 _10560_ ( .A(_02966_ ), .B(fanout_net_31 ), .C1(_02283_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02967_ ) );
NAND3_X1 _10561_ ( .A1(_02965_ ), .A2(_02967_ ), .A3(_02319_ ), .ZN(_02968_ ) );
MUX2_X1 _10562_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02969_ ) );
MUX2_X1 _10563_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02970_ ) );
MUX2_X1 _10564_ ( .A(_02969_ ), .B(_02970_ ), .S(_02292_ ), .Z(_02971_ ) );
OAI211_X1 _10565_ ( .A(_02312_ ), .B(_02968_ ), .C1(_02971_ ), .C2(_02320_ ), .ZN(_02972_ ) );
OR2_X1 _10566_ ( .A1(_02282_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02973_ ) );
OAI211_X1 _10567_ ( .A(_02973_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02974_ ) );
OR2_X1 _10568_ ( .A1(fanout_net_27 ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02975_ ) );
OAI211_X1 _10569_ ( .A(_02975_ ), .B(_02292_ ), .C1(_02283_ ), .C2(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02976_ ) );
NAND3_X1 _10570_ ( .A1(_02974_ ), .A2(fanout_net_33 ), .A3(_02976_ ), .ZN(_02977_ ) );
MUX2_X1 _10571_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02978_ ) );
MUX2_X1 _10572_ ( .A(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02979_ ) );
MUX2_X1 _10573_ ( .A(_02978_ ), .B(_02979_ ), .S(fanout_net_31 ), .Z(_02980_ ) );
OAI211_X1 _10574_ ( .A(fanout_net_34 ), .B(_02977_ ), .C1(_02980_ ), .C2(fanout_net_33 ), .ZN(_02981_ ) );
OAI211_X2 _10575_ ( .A(_02972_ ), .B(_02981_ ), .C1(_02340_ ), .C2(_02414_ ), .ZN(_02982_ ) );
NAND2_X4 _10576_ ( .A1(_02963_ ), .A2(_02982_ ), .ZN(_02983_ ) );
INV_X1 _10577_ ( .A(\ID_EX_imm [9] ), .ZN(_02984_ ) );
XNOR2_X1 _10578_ ( .A(_02983_ ), .B(_02984_ ), .ZN(_02985_ ) );
AND2_X1 _10579_ ( .A1(_02962_ ), .A2(_02985_ ), .ZN(_02986_ ) );
AND2_X1 _10580_ ( .A1(_02939_ ), .A2(_02986_ ), .ZN(_02987_ ) );
AND4_X2 _10581_ ( .A1(_02631_ ), .A2(_02841_ ), .A3(_02891_ ), .A4(_02987_ ), .ZN(_02988_ ) );
INV_X1 _10582_ ( .A(_02988_ ), .ZN(_02989_ ) );
AND2_X1 _10583_ ( .A1(_02960_ ), .A2(\ID_EX_imm [8] ), .ZN(_02990_ ) );
AND2_X1 _10584_ ( .A1(_02985_ ), .A2(_02990_ ), .ZN(_02991_ ) );
AOI21_X1 _10585_ ( .A(_02991_ ), .B1(\ID_EX_imm [9] ), .B2(_02983_ ), .ZN(_02992_ ) );
INV_X1 _10586_ ( .A(_02992_ ), .ZN(_02993_ ) );
AND2_X1 _10587_ ( .A1(_02993_ ), .A2(_02939_ ), .ZN(_02994_ ) );
AOI21_X1 _10588_ ( .A(_02937_ ), .B1(_02915_ ), .B2(_02934_ ), .ZN(_02995_ ) );
AND2_X1 _10589_ ( .A1(_02912_ ), .A2(\ID_EX_imm [10] ), .ZN(_02996_ ) );
AND2_X1 _10590_ ( .A1(_02938_ ), .A2(_02996_ ), .ZN(_02997_ ) );
NOR3_X1 _10591_ ( .A1(_02994_ ), .A2(_02995_ ), .A3(_02997_ ), .ZN(_02998_ ) );
INV_X1 _10592_ ( .A(_02998_ ), .ZN(_02999_ ) );
AND3_X1 _10593_ ( .A1(_02891_ ), .A2(_02607_ ), .A3(_02630_ ), .ZN(_03000_ ) );
NAND2_X1 _10594_ ( .A1(_02999_ ), .A2(_03000_ ), .ZN(_03001_ ) );
OAI211_X1 _10595_ ( .A(\ID_EX_imm [14] ), .B(_02629_ ), .C1(_02606_ ), .C2(\ID_EX_imm [15] ), .ZN(_03002_ ) );
NAND2_X1 _10596_ ( .A1(_02863_ ), .A2(\ID_EX_imm [12] ), .ZN(_03003_ ) );
NOR3_X1 _10597_ ( .A1(_03003_ ), .A2(_02888_ ), .A3(_02889_ ), .ZN(_03004_ ) );
OR2_X1 _10598_ ( .A1(_03004_ ), .A2(_02889_ ), .ZN(_03005_ ) );
AOI22_X1 _10599_ ( .A1(_03005_ ), .A2(_02631_ ), .B1(\ID_EX_imm [15] ), .B2(_02606_ ), .ZN(_03006_ ) );
AND3_X1 _10600_ ( .A1(_03001_ ), .A2(_03002_ ), .A3(_03006_ ), .ZN(_03007_ ) );
AOI211_X1 _10601_ ( .A(_02487_ ), .B(_02583_ ), .C1(_02989_ ), .C2(_03007_ ), .ZN(_03008_ ) );
AND2_X1 _10602_ ( .A1(_02580_ ), .A2(\ID_EX_imm [16] ), .ZN(_03009_ ) );
AND2_X1 _10603_ ( .A1(_02559_ ), .A2(_03009_ ), .ZN(_03010_ ) );
AOI21_X1 _10604_ ( .A(_03010_ ), .B1(\ID_EX_imm [17] ), .B2(_02557_ ), .ZN(_03011_ ) );
INV_X1 _10605_ ( .A(_03011_ ), .ZN(_03012_ ) );
NAND2_X1 _10606_ ( .A1(_03012_ ), .A2(_02536_ ), .ZN(_03013_ ) );
AND2_X1 _10607_ ( .A1(_02510_ ), .A2(\ID_EX_imm [18] ), .ZN(_03014_ ) );
AND2_X1 _10608_ ( .A1(_02535_ ), .A2(_03014_ ), .ZN(_03015_ ) );
AOI21_X1 _10609_ ( .A(_03015_ ), .B1(\ID_EX_imm [19] ), .B2(_02533_ ), .ZN(_03016_ ) );
AND2_X2 _10610_ ( .A1(_03013_ ), .A2(_03016_ ), .ZN(_03017_ ) );
OR2_X1 _10611_ ( .A1(_03017_ ), .A2(_02487_ ), .ZN(_03018_ ) );
NAND2_X1 _10612_ ( .A1(_02485_ ), .A2(\ID_EX_imm [20] ), .ZN(_03019_ ) );
NOR3_X1 _10613_ ( .A1(_03019_ ), .A2(_02462_ ), .A3(_02463_ ), .ZN(_03020_ ) );
OR2_X1 _10614_ ( .A1(_03020_ ), .A2(_02463_ ), .ZN(_03021_ ) );
NAND2_X1 _10615_ ( .A1(_03021_ ), .A2(_02440_ ), .ZN(_03022_ ) );
NAND4_X1 _10616_ ( .A1(_02439_ ), .A2(\ID_EX_imm [22] ), .A3(_02437_ ), .A4(_02411_ ), .ZN(_03023_ ) );
NAND4_X1 _10617_ ( .A1(_03018_ ), .A2(_02439_ ), .A3(_03022_ ), .A4(_03023_ ), .ZN(_03024_ ) );
OR2_X1 _10618_ ( .A1(_03008_ ), .A2(_03024_ ), .ZN(_03025_ ) );
OR3_X1 _10619_ ( .A1(_02343_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02355_ ), .ZN(_03026_ ) );
OR2_X1 _10620_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03027_ ) );
OAI211_X1 _10621_ ( .A(_03027_ ), .B(_02297_ ), .C1(_02301_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03028_ ) );
OR2_X1 _10622_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03029_ ) );
OAI211_X1 _10623_ ( .A(_03029_ ), .B(fanout_net_31 ), .C1(_02301_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03030_ ) );
NAND3_X1 _10624_ ( .A1(_03028_ ), .A2(_03030_ ), .A3(fanout_net_33 ), .ZN(_03031_ ) );
MUX2_X1 _10625_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03032_ ) );
MUX2_X1 _10626_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03033_ ) );
MUX2_X1 _10627_ ( .A(_03032_ ), .B(_03033_ ), .S(_02378_ ), .Z(_03034_ ) );
OAI211_X1 _10628_ ( .A(_02315_ ), .B(_03031_ ), .C1(_03034_ ), .C2(fanout_net_33 ), .ZN(_03035_ ) );
NOR2_X1 _10629_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03036_ ) );
OAI21_X1 _10630_ ( .A(_02378_ ), .B1(_02287_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03037_ ) );
INV_X1 _10631_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03038_ ) );
INV_X1 _10632_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03039_ ) );
MUX2_X1 _10633_ ( .A(_03038_ ), .B(_03039_ ), .S(fanout_net_28 ), .Z(_03040_ ) );
OAI221_X1 _10634_ ( .A(_02383_ ), .B1(_03036_ ), .B2(_03037_ ), .C1(_03040_ ), .C2(_02297_ ), .ZN(_03041_ ) );
MUX2_X1 _10635_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03042_ ) );
MUX2_X1 _10636_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03043_ ) );
MUX2_X1 _10637_ ( .A(_03042_ ), .B(_03043_ ), .S(fanout_net_31 ), .Z(_03044_ ) );
OAI211_X1 _10638_ ( .A(fanout_net_34 ), .B(_03041_ ), .C1(_03044_ ), .C2(_02324_ ), .ZN(_03045_ ) );
OAI211_X1 _10639_ ( .A(_03035_ ), .B(_03045_ ), .C1(_02343_ ), .C2(_02355_ ), .ZN(_03046_ ) );
NAND2_X1 _10640_ ( .A1(_03026_ ), .A2(_03046_ ), .ZN(_03047_ ) );
INV_X1 _10641_ ( .A(\ID_EX_imm [24] ), .ZN(_03048_ ) );
XNOR2_X1 _10642_ ( .A(_03047_ ), .B(_03048_ ), .ZN(_03049_ ) );
AND2_X2 _10643_ ( .A1(_03025_ ), .A2(_03049_ ), .ZN(_03050_ ) );
AOI21_X1 _10644_ ( .A(_03048_ ), .B1(_03026_ ), .B2(_03046_ ), .ZN(_03051_ ) );
NOR2_X2 _10645_ ( .A1(_03050_ ), .A2(_03051_ ), .ZN(_03052_ ) );
OR3_X1 _10646_ ( .A1(_02343_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02355_ ), .ZN(_03053_ ) );
OR2_X1 _10647_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03054_ ) );
OAI211_X1 _10648_ ( .A(_03054_ ), .B(_02297_ ), .C1(_02301_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03055_ ) );
OR2_X1 _10649_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03056_ ) );
OAI211_X1 _10650_ ( .A(_03056_ ), .B(fanout_net_31 ), .C1(_02301_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03057_ ) );
NAND3_X1 _10651_ ( .A1(_03055_ ), .A2(_03057_ ), .A3(_02324_ ), .ZN(_03058_ ) );
MUX2_X1 _10652_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03059_ ) );
MUX2_X1 _10653_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03060_ ) );
MUX2_X1 _10654_ ( .A(_03059_ ), .B(_03060_ ), .S(_02378_ ), .Z(_03061_ ) );
OAI211_X1 _10655_ ( .A(_02315_ ), .B(_03058_ ), .C1(_03061_ ), .C2(_02324_ ), .ZN(_03062_ ) );
OR2_X1 _10656_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03063_ ) );
OAI211_X1 _10657_ ( .A(_03063_ ), .B(_02378_ ), .C1(_02287_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03064_ ) );
NOR2_X1 _10658_ ( .A1(_02301_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03065_ ) );
OAI21_X1 _10659_ ( .A(fanout_net_31 ), .B1(fanout_net_28 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03066_ ) );
OAI211_X1 _10660_ ( .A(_03064_ ), .B(fanout_net_33 ), .C1(_03065_ ), .C2(_03066_ ), .ZN(_03067_ ) );
MUX2_X1 _10661_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03068_ ) );
MUX2_X1 _10662_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03069_ ) );
MUX2_X1 _10663_ ( .A(_03068_ ), .B(_03069_ ), .S(fanout_net_31 ), .Z(_03070_ ) );
OAI211_X1 _10664_ ( .A(fanout_net_34 ), .B(_03067_ ), .C1(_03070_ ), .C2(fanout_net_33 ), .ZN(_03071_ ) );
OAI211_X1 _10665_ ( .A(_03062_ ), .B(_03071_ ), .C1(_02343_ ), .C2(_02355_ ), .ZN(_03072_ ) );
NAND2_X1 _10666_ ( .A1(_03053_ ), .A2(_03072_ ), .ZN(_03073_ ) );
NAND2_X1 _10667_ ( .A1(_03073_ ), .A2(\ID_EX_imm [25] ), .ZN(_03074_ ) );
NAND2_X2 _10668_ ( .A1(_03052_ ), .A2(_03074_ ), .ZN(_03075_ ) );
OR3_X1 _10669_ ( .A1(_02342_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02354_ ), .ZN(_03076_ ) );
INV_X1 _10670_ ( .A(\ID_EX_imm [27] ), .ZN(_03077_ ) );
OR2_X1 _10671_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03078_ ) );
OAI211_X1 _10672_ ( .A(_03078_ ), .B(_02364_ ), .C1(_02287_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03079_ ) );
OR2_X1 _10673_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03080_ ) );
OAI211_X1 _10674_ ( .A(_03080_ ), .B(fanout_net_31 ), .C1(_02300_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03081_ ) );
NAND3_X1 _10675_ ( .A1(_03079_ ), .A2(_03081_ ), .A3(_02383_ ), .ZN(_03082_ ) );
MUX2_X1 _10676_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03083_ ) );
MUX2_X1 _10677_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03084_ ) );
MUX2_X1 _10678_ ( .A(_03083_ ), .B(_03084_ ), .S(_02296_ ), .Z(_03085_ ) );
OAI211_X1 _10679_ ( .A(_02314_ ), .B(_03082_ ), .C1(_03085_ ), .C2(_02383_ ), .ZN(_03086_ ) );
OR2_X1 _10680_ ( .A1(_02299_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03087_ ) );
OAI211_X1 _10681_ ( .A(_03087_ ), .B(_02364_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03088_ ) );
OR2_X1 _10682_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03089_ ) );
OAI211_X1 _10683_ ( .A(_03089_ ), .B(fanout_net_31 ), .C1(_02300_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03090_ ) );
NAND3_X1 _10684_ ( .A1(_03088_ ), .A2(fanout_net_33 ), .A3(_03090_ ), .ZN(_03091_ ) );
MUX2_X1 _10685_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03092_ ) );
MUX2_X1 _10686_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03093_ ) );
MUX2_X1 _10687_ ( .A(_03092_ ), .B(_03093_ ), .S(fanout_net_31 ), .Z(_03094_ ) );
OAI211_X1 _10688_ ( .A(fanout_net_34 ), .B(_03091_ ), .C1(_03094_ ), .C2(fanout_net_33 ), .ZN(_03095_ ) );
OAI211_X1 _10689_ ( .A(_03086_ ), .B(_03095_ ), .C1(_02385_ ), .C2(_02386_ ), .ZN(_03096_ ) );
AND3_X1 _10690_ ( .A1(_03076_ ), .A2(_03077_ ), .A3(_03096_ ), .ZN(_03097_ ) );
AOI21_X1 _10691_ ( .A(_03077_ ), .B1(_03076_ ), .B2(_03096_ ), .ZN(_03098_ ) );
NOR2_X1 _10692_ ( .A1(_03097_ ), .A2(_03098_ ), .ZN(_03099_ ) );
OR3_X4 _10693_ ( .A1(_02385_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02386_ ), .ZN(_03100_ ) );
OR2_X1 _10694_ ( .A1(_02286_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03101_ ) );
OAI211_X1 _10695_ ( .A(_03101_ ), .B(_02378_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03102_ ) );
OR2_X1 _10696_ ( .A1(_02299_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03103_ ) );
OAI211_X1 _10697_ ( .A(_03103_ ), .B(fanout_net_31 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03104_ ) );
NAND3_X1 _10698_ ( .A1(_03102_ ), .A2(_03104_ ), .A3(fanout_net_33 ), .ZN(_03105_ ) );
MUX2_X1 _10699_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03106_ ) );
MUX2_X1 _10700_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_03107_ ) );
MUX2_X1 _10701_ ( .A(_03106_ ), .B(_03107_ ), .S(_02364_ ), .Z(_03108_ ) );
OAI211_X1 _10702_ ( .A(_02315_ ), .B(_03105_ ), .C1(_03108_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03109_ ) );
NOR2_X1 _10703_ ( .A1(_02300_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03110_ ) );
OAI21_X1 _10704_ ( .A(fanout_net_31 ), .B1(fanout_net_28 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03111_ ) );
NOR2_X1 _10705_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03112_ ) );
OAI21_X1 _10706_ ( .A(_02296_ ), .B1(_02300_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03113_ ) );
OAI221_X1 _10707_ ( .A(_02323_ ), .B1(_03110_ ), .B2(_03111_ ), .C1(_03112_ ), .C2(_03113_ ), .ZN(_03114_ ) );
MUX2_X1 _10708_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03115_ ) );
MUX2_X1 _10709_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03116_ ) );
MUX2_X1 _10710_ ( .A(_03115_ ), .B(_03116_ ), .S(fanout_net_31 ), .Z(_03117_ ) );
OAI211_X1 _10711_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03114_ ), .C1(_03117_ ), .C2(_02383_ ), .ZN(_03118_ ) );
OAI211_X1 _10712_ ( .A(_03109_ ), .B(_03118_ ), .C1(_02343_ ), .C2(_02355_ ), .ZN(_03119_ ) );
NAND2_X1 _10713_ ( .A1(_03100_ ), .A2(_03119_ ), .ZN(_03120_ ) );
INV_X1 _10714_ ( .A(\ID_EX_imm [26] ), .ZN(_03121_ ) );
XNOR2_X1 _10715_ ( .A(_03120_ ), .B(_03121_ ), .ZN(_03122_ ) );
INV_X1 _10716_ ( .A(\ID_EX_imm [25] ), .ZN(_03123_ ) );
NAND3_X1 _10717_ ( .A1(_03053_ ), .A2(_03123_ ), .A3(_03072_ ), .ZN(_03124_ ) );
NAND4_X1 _10718_ ( .A1(_03075_ ), .A2(_03099_ ), .A3(_03122_ ), .A4(_03124_ ), .ZN(_03125_ ) );
INV_X1 _10719_ ( .A(_03120_ ), .ZN(_03126_ ) );
NOR4_X1 _10720_ ( .A1(_03097_ ), .A2(_03126_ ), .A3(_03098_ ), .A4(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03127_ ) );
NOR2_X1 _10721_ ( .A1(_03127_ ), .A2(_03098_ ), .ZN(_03128_ ) );
AOI21_X2 _10722_ ( .A(_02389_ ), .B1(_03125_ ), .B2(_03128_ ), .ZN(_03129_ ) );
OR3_X1 _10723_ ( .A1(_02385_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02386_ ), .ZN(_03130_ ) );
OR2_X1 _10724_ ( .A1(_02299_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03131_ ) );
OAI211_X1 _10725_ ( .A(_03131_ ), .B(_02378_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03132_ ) );
OR2_X1 _10726_ ( .A1(_02299_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03133_ ) );
OAI211_X1 _10727_ ( .A(_03133_ ), .B(fanout_net_31 ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03134_ ) );
NAND3_X1 _10728_ ( .A1(_03132_ ), .A2(_03134_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03135_ ) );
MUX2_X1 _10729_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03136_ ) );
MUX2_X1 _10730_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03137_ ) );
MUX2_X1 _10731_ ( .A(_03136_ ), .B(_03137_ ), .S(_02364_ ), .Z(_03138_ ) );
OAI211_X1 _10732_ ( .A(_02315_ ), .B(_03135_ ), .C1(_03138_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03139_ ) );
NOR2_X1 _10733_ ( .A1(_02286_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03140_ ) );
OAI21_X1 _10734_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03141_ ) );
NOR2_X1 _10735_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03142_ ) );
OAI21_X1 _10736_ ( .A(_02296_ ), .B1(_02300_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03143_ ) );
OAI221_X1 _10737_ ( .A(_02323_ ), .B1(_03140_ ), .B2(_03141_ ), .C1(_03142_ ), .C2(_03143_ ), .ZN(_03144_ ) );
MUX2_X1 _10738_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03145_ ) );
MUX2_X1 _10739_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03146_ ) );
MUX2_X1 _10740_ ( .A(_03145_ ), .B(_03146_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03147_ ) );
OAI211_X1 _10741_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03144_ ), .C1(_03147_ ), .C2(_02383_ ), .ZN(_03148_ ) );
OAI211_X1 _10742_ ( .A(_03139_ ), .B(_03148_ ), .C1(_02385_ ), .C2(_02386_ ), .ZN(_03149_ ) );
NAND2_X1 _10743_ ( .A1(_03130_ ), .A2(_03149_ ), .ZN(_03150_ ) );
INV_X1 _10744_ ( .A(\ID_EX_imm [29] ), .ZN(_03151_ ) );
XNOR2_X1 _10745_ ( .A(_03150_ ), .B(_03151_ ), .ZN(_03152_ ) );
AND2_X2 _10746_ ( .A1(_03129_ ), .A2(_03152_ ), .ZN(_03153_ ) );
AOI21_X1 _10747_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02362_ ), .B2(_02387_ ), .ZN(_03154_ ) );
NAND2_X1 _10748_ ( .A1(_03152_ ), .A2(_03154_ ), .ZN(_03155_ ) );
INV_X1 _10749_ ( .A(_03150_ ), .ZN(_03156_ ) );
OAI21_X1 _10750_ ( .A(_03155_ ), .B1(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_03156_ ), .ZN(_03157_ ) );
OAI21_X1 _10751_ ( .A(_02361_ ), .B1(_03153_ ), .B2(_03157_ ), .ZN(_03158_ ) );
OR2_X1 _10752_ ( .A1(_02358_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03159_ ) );
AND2_X2 _10753_ ( .A1(_03158_ ), .A2(_03159_ ), .ZN(_03160_ ) );
NAND2_X1 _10754_ ( .A1(_02683_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_03161_ ) );
OR2_X1 _10755_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03162_ ) );
OAI211_X1 _10756_ ( .A(_03162_ ), .B(_02297_ ), .C1(_02301_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03163_ ) );
INV_X1 _10757_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03164_ ) );
NAND2_X1 _10758_ ( .A1(_03164_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .ZN(_03165_ ) );
OAI211_X1 _10759_ ( .A(_03165_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03166_ ) );
NAND3_X1 _10760_ ( .A1(_03163_ ), .A2(_03166_ ), .A3(_02324_ ), .ZN(_03167_ ) );
MUX2_X1 _10761_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03168_ ) );
MUX2_X1 _10762_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03169_ ) );
MUX2_X1 _10763_ ( .A(_03168_ ), .B(_03169_ ), .S(_02378_ ), .Z(_03170_ ) );
OAI211_X1 _10764_ ( .A(_02315_ ), .B(_03167_ ), .C1(_03170_ ), .C2(_02324_ ), .ZN(_03171_ ) );
OR2_X1 _10765_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03172_ ) );
OAI211_X1 _10766_ ( .A(_03172_ ), .B(_02297_ ), .C1(_02287_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03173_ ) );
INV_X1 _10767_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03174_ ) );
NAND2_X1 _10768_ ( .A1(_03174_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .ZN(_03175_ ) );
OAI211_X1 _10769_ ( .A(_03175_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03176_ ) );
NAND3_X1 _10770_ ( .A1(_03173_ ), .A2(_03176_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03177_ ) );
MUX2_X1 _10771_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03178_ ) );
MUX2_X1 _10772_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03179_ ) );
MUX2_X1 _10773_ ( .A(_03178_ ), .B(_03179_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03180_ ) );
OAI211_X1 _10774_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03177_ ), .C1(_03180_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03181_ ) );
NAND2_X1 _10775_ ( .A1(_03171_ ), .A2(_03181_ ), .ZN(_03182_ ) );
OAI21_X1 _10776_ ( .A(_03182_ ), .B1(_02343_ ), .B2(_02355_ ), .ZN(_03183_ ) );
AND2_X1 _10777_ ( .A1(_03161_ ), .A2(_03183_ ), .ZN(_03184_ ) );
BUF_X2 _10778_ ( .A(_03184_ ), .Z(_03185_ ) );
XNOR2_X1 _10779_ ( .A(_03185_ ), .B(\ID_EX_imm [31] ), .ZN(_03186_ ) );
XNOR2_X1 _10780_ ( .A(_03160_ ), .B(_03186_ ), .ZN(_03187_ ) );
AND2_X1 _10781_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_03188_ ) );
BUF_X4 _10782_ ( .A(_03188_ ), .Z(_03189_ ) );
BUF_X4 _10783_ ( .A(_03189_ ), .Z(_03190_ ) );
NOR2_X1 _10784_ ( .A1(_03187_ ), .A2(_03190_ ), .ZN(_00133_ ) );
OR3_X1 _10785_ ( .A1(_03153_ ), .A2(_03157_ ), .A3(_02361_ ), .ZN(_03191_ ) );
INV_X1 _10786_ ( .A(_03189_ ), .ZN(_03192_ ) );
CLKBUF_X2 _10787_ ( .A(_03192_ ), .Z(_03193_ ) );
AND3_X1 _10788_ ( .A1(_03191_ ), .A2(_03193_ ), .A3(_03158_ ), .ZN(_00134_ ) );
AOI21_X1 _10789_ ( .A(_02583_ ), .B1(_02989_ ), .B2(_03007_ ), .ZN(_03194_ ) );
INV_X1 _10790_ ( .A(_03017_ ), .ZN(_03195_ ) );
OAI21_X1 _10791_ ( .A(_02486_ ), .B1(_03194_ ), .B2(_03195_ ), .ZN(_03196_ ) );
NAND2_X1 _10792_ ( .A1(_03196_ ), .A2(_03019_ ), .ZN(_03197_ ) );
XNOR2_X1 _10793_ ( .A(_03197_ ), .B(_02464_ ), .ZN(_03198_ ) );
NOR2_X1 _10794_ ( .A1(_03198_ ), .A2(_03190_ ), .ZN(_00135_ ) );
OR3_X1 _10795_ ( .A1(_03194_ ), .A2(_02486_ ), .A3(_03195_ ), .ZN(_03199_ ) );
AND3_X1 _10796_ ( .A1(_03199_ ), .A2(_03193_ ), .A3(_03196_ ), .ZN(_00136_ ) );
INV_X1 _10797_ ( .A(_02582_ ), .ZN(_03200_ ) );
AOI21_X1 _10798_ ( .A(_03200_ ), .B1(_02989_ ), .B2(_03007_ ), .ZN(_03201_ ) );
AND2_X1 _10799_ ( .A1(_03201_ ), .A2(_02559_ ), .ZN(_03202_ ) );
OAI21_X1 _10800_ ( .A(_02512_ ), .B1(_03202_ ), .B2(_03012_ ), .ZN(_03203_ ) );
INV_X1 _10801_ ( .A(_03014_ ), .ZN(_03204_ ) );
NAND2_X1 _10802_ ( .A1(_03203_ ), .A2(_03204_ ), .ZN(_03205_ ) );
XNOR2_X1 _10803_ ( .A(_03205_ ), .B(_02535_ ), .ZN(_03206_ ) );
NOR2_X1 _10804_ ( .A1(_03206_ ), .A2(_03190_ ), .ZN(_00137_ ) );
NOR2_X1 _10805_ ( .A1(_03202_ ), .A2(_03012_ ), .ZN(_03207_ ) );
XNOR2_X1 _10806_ ( .A(_03207_ ), .B(_02512_ ), .ZN(_03208_ ) );
AND2_X1 _10807_ ( .A1(_03208_ ), .A2(_03193_ ), .ZN(_00138_ ) );
OR2_X1 _10808_ ( .A1(_03201_ ), .A2(_03009_ ), .ZN(_03209_ ) );
XNOR2_X1 _10809_ ( .A(_03209_ ), .B(_02559_ ), .ZN(_03210_ ) );
NOR2_X1 _10810_ ( .A1(_03210_ ), .A2(_03190_ ), .ZN(_00139_ ) );
AND3_X1 _10811_ ( .A1(_02989_ ), .A2(_03007_ ), .A3(_03200_ ), .ZN(_03211_ ) );
NOR3_X1 _10812_ ( .A1(_03211_ ), .A2(_03201_ ), .A3(_03189_ ), .ZN(_00140_ ) );
INV_X1 _10813_ ( .A(_02891_ ), .ZN(_03212_ ) );
INV_X1 _10814_ ( .A(_02987_ ), .ZN(_03213_ ) );
AOI21_X1 _10815_ ( .A(_03213_ ), .B1(_02738_ ), .B2(_02839_ ), .ZN(_03214_ ) );
INV_X1 _10816_ ( .A(_03214_ ), .ZN(_03215_ ) );
AOI21_X1 _10817_ ( .A(_03212_ ), .B1(_03215_ ), .B2(_02998_ ), .ZN(_03216_ ) );
OR2_X1 _10818_ ( .A1(_03216_ ), .A2(_03005_ ), .ZN(_03217_ ) );
AND2_X1 _10819_ ( .A1(_03217_ ), .A2(_02630_ ), .ZN(_03218_ ) );
AND2_X1 _10820_ ( .A1(_02629_ ), .A2(\ID_EX_imm [14] ), .ZN(_03219_ ) );
OR2_X1 _10821_ ( .A1(_03218_ ), .A2(_03219_ ), .ZN(_03220_ ) );
XNOR2_X1 _10822_ ( .A(_03220_ ), .B(_02607_ ), .ZN(_03221_ ) );
NOR2_X1 _10823_ ( .A1(_03221_ ), .A2(_03190_ ), .ZN(_00141_ ) );
XOR2_X1 _10824_ ( .A(_03217_ ), .B(_02630_ ), .Z(_03222_ ) );
AND2_X1 _10825_ ( .A1(_03222_ ), .A2(_03193_ ), .ZN(_00142_ ) );
OAI21_X1 _10826_ ( .A(_02865_ ), .B1(_03214_ ), .B2(_02999_ ), .ZN(_03223_ ) );
NAND2_X1 _10827_ ( .A1(_03223_ ), .A2(_03003_ ), .ZN(_03224_ ) );
XNOR2_X1 _10828_ ( .A(_03224_ ), .B(_02890_ ), .ZN(_03225_ ) );
NOR2_X1 _10829_ ( .A1(_03225_ ), .A2(_03190_ ), .ZN(_00143_ ) );
OR3_X1 _10830_ ( .A1(_03214_ ), .A2(_02999_ ), .A3(_02865_ ), .ZN(_03226_ ) );
AND3_X1 _10831_ ( .A1(_03226_ ), .A2(_03192_ ), .A3(_03223_ ), .ZN(_00144_ ) );
OR2_X1 _10832_ ( .A1(_03129_ ), .A2(_03154_ ), .ZN(_03227_ ) );
XNOR2_X1 _10833_ ( .A(_03227_ ), .B(_03152_ ), .ZN(_03228_ ) );
NOR2_X1 _10834_ ( .A1(_03228_ ), .A2(_03190_ ), .ZN(_00145_ ) );
AND3_X1 _10835_ ( .A1(_03125_ ), .A2(_03128_ ), .A3(_02389_ ), .ZN(_03229_ ) );
NOR3_X1 _10836_ ( .A1(_03229_ ), .A2(_03129_ ), .A3(_03189_ ), .ZN(_00146_ ) );
NAND3_X1 _10837_ ( .A1(_03075_ ), .A2(_03122_ ), .A3(_03124_ ), .ZN(_03230_ ) );
OR2_X1 _10838_ ( .A1(_03126_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03231_ ) );
NAND2_X1 _10839_ ( .A1(_03230_ ), .A2(_03231_ ), .ZN(_03232_ ) );
XNOR2_X1 _10840_ ( .A(_03232_ ), .B(_03099_ ), .ZN(_03233_ ) );
NOR2_X1 _10841_ ( .A1(_03233_ ), .A2(_03190_ ), .ZN(_00147_ ) );
NAND2_X1 _10842_ ( .A1(_03075_ ), .A2(_03124_ ), .ZN(_03234_ ) );
XNOR2_X1 _10843_ ( .A(_03234_ ), .B(_03122_ ), .ZN(_03235_ ) );
AND2_X1 _10844_ ( .A1(_03235_ ), .A2(_03193_ ), .ZN(_00148_ ) );
NAND2_X1 _10845_ ( .A1(_03074_ ), .A2(_03124_ ), .ZN(_03236_ ) );
XNOR2_X1 _10846_ ( .A(_03052_ ), .B(_03236_ ), .ZN(_03237_ ) );
NOR2_X1 _10847_ ( .A1(_03237_ ), .A2(_03190_ ), .ZN(_00149_ ) );
XOR2_X1 _10848_ ( .A(_03025_ ), .B(_03049_ ), .Z(_03238_ ) );
AND2_X1 _10849_ ( .A1(_03238_ ), .A2(_03193_ ), .ZN(_00150_ ) );
OAI211_X1 _10850_ ( .A(_02464_ ), .B(_02486_ ), .C1(_03194_ ), .C2(_03195_ ), .ZN(_03239_ ) );
INV_X1 _10851_ ( .A(_03239_ ), .ZN(_03240_ ) );
OAI21_X1 _10852_ ( .A(_02413_ ), .B1(_03240_ ), .B2(_03021_ ), .ZN(_03241_ ) );
NAND2_X1 _10853_ ( .A1(_02411_ ), .A2(\ID_EX_imm [22] ), .ZN(_03242_ ) );
AND4_X1 _10854_ ( .A1(_02437_ ), .A2(_03241_ ), .A3(_02439_ ), .A4(_03242_ ), .ZN(_03243_ ) );
AOI22_X1 _10855_ ( .A1(_03241_ ), .A2(_03242_ ), .B1(_02437_ ), .B2(_02439_ ), .ZN(_03244_ ) );
NOR2_X1 _10856_ ( .A1(_03243_ ), .A2(_03244_ ), .ZN(_03245_ ) );
NOR2_X1 _10857_ ( .A1(_03245_ ), .A2(_03190_ ), .ZN(_00151_ ) );
OR3_X1 _10858_ ( .A1(_03240_ ), .A2(_02413_ ), .A3(_03021_ ), .ZN(_03246_ ) );
AND3_X1 _10859_ ( .A1(_03246_ ), .A2(_03192_ ), .A3(_03241_ ), .ZN(_00152_ ) );
CLKBUF_X2 _10860_ ( .A(_02278_ ), .Z(_03247_ ) );
AND2_X1 _10861_ ( .A1(_03247_ ), .A2(\ID_EX_rd [4] ), .ZN(_00153_ ) );
AND2_X1 _10862_ ( .A1(_03247_ ), .A2(\ID_EX_rd [3] ), .ZN(_00154_ ) );
AND2_X1 _10863_ ( .A1(_03247_ ), .A2(\ID_EX_rd [2] ), .ZN(_00155_ ) );
AND2_X1 _10864_ ( .A1(_03247_ ), .A2(\ID_EX_rd [1] ), .ZN(_00156_ ) );
AND2_X1 _10865_ ( .A1(_03247_ ), .A2(\ID_EX_rd [0] ), .ZN(_00157_ ) );
INV_X2 _10866_ ( .A(_02277_ ), .ZN(_03248_ ) );
AND3_X1 _10867_ ( .A1(_03191_ ), .A2(fanout_net_8 ), .A3(_03158_ ), .ZN(_03249_ ) );
INV_X2 _10868_ ( .A(fanout_net_8 ), .ZN(_03250_ ) );
BUF_X4 _10869_ ( .A(_03250_ ), .Z(_03251_ ) );
BUF_X4 _10870_ ( .A(_03251_ ), .Z(_03252_ ) );
XNOR2_X1 _10871_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .ZN(_03253_ ) );
AND2_X1 _10872_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_03254_ ) );
NOR2_X1 _10873_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_03255_ ) );
NOR3_X1 _10874_ ( .A1(_03253_ ), .A2(_03254_ ), .A3(_03255_ ), .ZN(_03256_ ) );
XOR2_X1 _10875_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_03257_ ) );
XOR2_X1 _10876_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_03258_ ) );
AND3_X1 _10877_ ( .A1(_03256_ ), .A2(_03257_ ), .A3(_03258_ ), .ZN(_03259_ ) );
XOR2_X1 _10878_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_03260_ ) );
XOR2_X1 _10879_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_03261_ ) );
AND2_X1 _10880_ ( .A1(_03260_ ), .A2(_03261_ ), .ZN(_03262_ ) );
XOR2_X1 _10881_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_03263_ ) );
XOR2_X1 _10882_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_03264_ ) );
AND2_X1 _10883_ ( .A1(_03263_ ), .A2(_03264_ ), .ZN(_03265_ ) );
AND2_X1 _10884_ ( .A1(_03262_ ), .A2(_03265_ ), .ZN(_03266_ ) );
XOR2_X1 _10885_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_03267_ ) );
XOR2_X1 _10886_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_03268_ ) );
AND2_X1 _10887_ ( .A1(_03267_ ), .A2(_03268_ ), .ZN(_03269_ ) );
NOR2_X1 _10888_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_03270_ ) );
XOR2_X1 _10889_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_03271_ ) );
AND2_X1 _10890_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_03272_ ) );
NAND2_X1 _10891_ ( .A1(_03271_ ), .A2(_03272_ ), .ZN(_03273_ ) );
INV_X1 _10892_ ( .A(\ID_EX_pc [1] ), .ZN(_03274_ ) );
OAI21_X1 _10893_ ( .A(_03273_ ), .B1(_03274_ ), .B2(_02761_ ), .ZN(_03275_ ) );
XOR2_X1 _10894_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_03276_ ) );
NAND2_X1 _10895_ ( .A1(_03275_ ), .A2(_03276_ ), .ZN(_03277_ ) );
NAND2_X1 _10896_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_03278_ ) );
NAND2_X1 _10897_ ( .A1(_03277_ ), .A2(_03278_ ), .ZN(_03279_ ) );
OAI21_X1 _10898_ ( .A(_03279_ ), .B1(\ID_EX_pc [3] ), .B2(\ID_EX_imm [3] ), .ZN(_03280_ ) );
NAND2_X1 _10899_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_03281_ ) );
NAND2_X1 _10900_ ( .A1(_03280_ ), .A2(_03281_ ), .ZN(_03282_ ) );
XOR2_X1 _10901_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_03283_ ) );
NAND2_X1 _10902_ ( .A1(_03282_ ), .A2(_03283_ ), .ZN(_03284_ ) );
NAND2_X1 _10903_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_03285_ ) );
AOI21_X1 _10904_ ( .A(_03270_ ), .B1(_03284_ ), .B2(_03285_ ), .ZN(_03286_ ) );
AOI21_X1 _10905_ ( .A(_03286_ ), .B1(\ID_EX_pc [5] ), .B2(\ID_EX_imm [5] ), .ZN(_03287_ ) );
AND2_X1 _10906_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03288_ ) );
NOR2_X1 _10907_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_03289_ ) );
NOR3_X1 _10908_ ( .A1(_03287_ ), .A2(_03288_ ), .A3(_03289_ ), .ZN(_03290_ ) );
NOR2_X1 _10909_ ( .A1(_03290_ ), .A2(_03288_ ), .ZN(_03291_ ) );
NOR2_X1 _10910_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03292_ ) );
NOR2_X1 _10911_ ( .A1(_03291_ ), .A2(_03292_ ), .ZN(_03293_ ) );
AND2_X1 _10912_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_03294_ ) );
OR2_X1 _10913_ ( .A1(_03293_ ), .A2(_03294_ ), .ZN(_03295_ ) );
XOR2_X1 _10914_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_03296_ ) );
XOR2_X1 _10915_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_03297_ ) );
XOR2_X1 _10916_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_03298_ ) );
AND2_X1 _10917_ ( .A1(\ID_EX_pc [9] ), .A2(\ID_EX_imm [9] ), .ZN(_03299_ ) );
NOR2_X1 _10918_ ( .A1(\ID_EX_pc [9] ), .A2(\ID_EX_imm [9] ), .ZN(_03300_ ) );
NOR2_X1 _10919_ ( .A1(_03299_ ), .A2(_03300_ ), .ZN(_03301_ ) );
AND2_X1 _10920_ ( .A1(_03298_ ), .A2(_03301_ ), .ZN(_03302_ ) );
NAND4_X1 _10921_ ( .A1(_03295_ ), .A2(_03296_ ), .A3(_03297_ ), .A4(_03302_ ), .ZN(_03303_ ) );
AND2_X1 _10922_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_03304_ ) );
AOI21_X1 _10923_ ( .A(_03299_ ), .B1(_03301_ ), .B2(_03304_ ), .ZN(_03305_ ) );
INV_X1 _10924_ ( .A(_03305_ ), .ZN(_03306_ ) );
AND3_X1 _10925_ ( .A1(_03306_ ), .A2(_03296_ ), .A3(_03297_ ), .ZN(_03307_ ) );
AND2_X1 _10926_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_imm [11] ), .ZN(_03308_ ) );
AND2_X1 _10927_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_03309_ ) );
AND2_X1 _10928_ ( .A1(_03296_ ), .A2(_03309_ ), .ZN(_03310_ ) );
NOR3_X1 _10929_ ( .A1(_03307_ ), .A2(_03308_ ), .A3(_03310_ ), .ZN(_03311_ ) );
NAND2_X1 _10930_ ( .A1(_03303_ ), .A2(_03311_ ), .ZN(_03312_ ) );
AND2_X1 _10931_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_imm [13] ), .ZN(_03313_ ) );
NOR2_X1 _10932_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_imm [13] ), .ZN(_03314_ ) );
NOR2_X1 _10933_ ( .A1(_03313_ ), .A2(_03314_ ), .ZN(_03315_ ) );
XOR2_X1 _10934_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_03316_ ) );
AND4_X1 _10935_ ( .A1(_03269_ ), .A2(_03312_ ), .A3(_03315_ ), .A4(_03316_ ), .ZN(_03317_ ) );
AND2_X1 _10936_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_03318_ ) );
AND2_X1 _10937_ ( .A1(_03267_ ), .A2(_03318_ ), .ZN(_03319_ ) );
AOI21_X1 _10938_ ( .A(_03319_ ), .B1(\ID_EX_pc [15] ), .B2(\ID_EX_imm [15] ), .ZN(_03320_ ) );
INV_X1 _10939_ ( .A(_03314_ ), .ZN(_03321_ ) );
AND2_X1 _10940_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_03322_ ) );
AOI21_X1 _10941_ ( .A(_03313_ ), .B1(_03321_ ), .B2(_03322_ ), .ZN(_03323_ ) );
INV_X1 _10942_ ( .A(_03269_ ), .ZN(_03324_ ) );
OAI21_X1 _10943_ ( .A(_03320_ ), .B1(_03323_ ), .B2(_03324_ ), .ZN(_03325_ ) );
OAI211_X1 _10944_ ( .A(_03259_ ), .B(_03266_ ), .C1(_03317_ ), .C2(_03325_ ), .ZN(_03326_ ) );
AND2_X1 _10945_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_03327_ ) );
NAND2_X1 _10946_ ( .A1(_03257_ ), .A2(_03327_ ), .ZN(_03328_ ) );
INV_X1 _10947_ ( .A(\ID_EX_pc [23] ), .ZN(_03329_ ) );
AND2_X1 _10948_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_03330_ ) );
NAND2_X1 _10949_ ( .A1(_03260_ ), .A2(_03330_ ), .ZN(_03331_ ) );
INV_X1 _10950_ ( .A(\ID_EX_pc [19] ), .ZN(_03332_ ) );
OAI21_X1 _10951_ ( .A(_03331_ ), .B1(_03332_ ), .B2(_02534_ ), .ZN(_03333_ ) );
NAND3_X1 _10952_ ( .A1(_03263_ ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_imm [16] ), .ZN(_03334_ ) );
INV_X1 _10953_ ( .A(\ID_EX_pc [17] ), .ZN(_03335_ ) );
OAI21_X1 _10954_ ( .A(_03334_ ), .B1(_03335_ ), .B2(_02558_ ), .ZN(_03336_ ) );
AOI21_X1 _10955_ ( .A(_03333_ ), .B1(_03336_ ), .B2(_03262_ ), .ZN(_03337_ ) );
INV_X1 _10956_ ( .A(_03259_ ), .ZN(_03338_ ) );
OAI221_X1 _10957_ ( .A(_03328_ ), .B1(_03329_ ), .B2(_02436_ ), .C1(_03337_ ), .C2(_03338_ ), .ZN(_03339_ ) );
AND2_X1 _10958_ ( .A1(_03257_ ), .A2(_03258_ ), .ZN(_03340_ ) );
INV_X1 _10959_ ( .A(_03255_ ), .ZN(_03341_ ) );
AND2_X1 _10960_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_03342_ ) );
OR2_X1 _10961_ ( .A1(_03254_ ), .A2(_03342_ ), .ZN(_03343_ ) );
AND3_X1 _10962_ ( .A1(_03340_ ), .A2(_03341_ ), .A3(_03343_ ), .ZN(_03344_ ) );
NOR2_X1 _10963_ ( .A1(_03339_ ), .A2(_03344_ ), .ZN(_03345_ ) );
NAND2_X1 _10964_ ( .A1(_03326_ ), .A2(_03345_ ), .ZN(_03346_ ) );
XOR2_X1 _10965_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_03347_ ) );
XOR2_X1 _10966_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_03348_ ) );
AND2_X1 _10967_ ( .A1(_03347_ ), .A2(_03348_ ), .ZN(_03349_ ) );
XOR2_X1 _10968_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_03350_ ) );
AND2_X1 _10969_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_03351_ ) );
NOR2_X1 _10970_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_03352_ ) );
NOR2_X1 _10971_ ( .A1(_03351_ ), .A2(_03352_ ), .ZN(_03353_ ) );
AND2_X1 _10972_ ( .A1(_03350_ ), .A2(_03353_ ), .ZN(_03354_ ) );
NAND3_X1 _10973_ ( .A1(_03346_ ), .A2(_03349_ ), .A3(_03354_ ), .ZN(_03355_ ) );
AND2_X1 _10974_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_03356_ ) );
AND2_X1 _10975_ ( .A1(_03347_ ), .A2(_03356_ ), .ZN(_03357_ ) );
NAND2_X1 _10976_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_03358_ ) );
NOR3_X1 _10977_ ( .A1(_03351_ ), .A2(_03352_ ), .A3(_03358_ ), .ZN(_03359_ ) );
OR2_X1 _10978_ ( .A1(_03359_ ), .A2(_03351_ ), .ZN(_03360_ ) );
AOI221_X4 _10979_ ( .A(_03357_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .C1(_03349_ ), .C2(_03360_ ), .ZN(_03361_ ) );
NAND2_X1 _10980_ ( .A1(_03355_ ), .A2(_03361_ ), .ZN(_03362_ ) );
XOR2_X1 _10981_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_03363_ ) );
NAND2_X1 _10982_ ( .A1(_03362_ ), .A2(_03363_ ), .ZN(_03364_ ) );
NAND2_X1 _10983_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_03365_ ) );
INV_X1 _10984_ ( .A(\ID_EX_pc [29] ), .ZN(_03366_ ) );
OAI211_X1 _10985_ ( .A(_03364_ ), .B(_03365_ ), .C1(_03366_ ), .C2(_03151_ ), .ZN(_03367_ ) );
OAI21_X1 _10986_ ( .A(_03367_ ), .B1(\ID_EX_pc [29] ), .B2(\ID_EX_imm [29] ), .ZN(_03368_ ) );
XNOR2_X1 _10987_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .ZN(_03369_ ) );
XOR2_X1 _10988_ ( .A(_03368_ ), .B(_03369_ ), .Z(_03370_ ) );
AOI211_X1 _10989_ ( .A(_02274_ ), .B(_03249_ ), .C1(_03252_ ), .C2(_03370_ ), .ZN(_03371_ ) );
INV_X2 _10990_ ( .A(fanout_net_10 ), .ZN(_03372_ ) );
INV_X1 _10991_ ( .A(\ID_EX_csr [9] ), .ZN(_03373_ ) );
INV_X1 _10992_ ( .A(\ID_EX_csr [8] ), .ZN(_03374_ ) );
AOI22_X1 _10993_ ( .A1(\EX_LS_dest_csreg_mem [9] ), .A2(_03373_ ), .B1(_03374_ ), .B2(\EX_LS_dest_csreg_mem [8] ), .ZN(_03375_ ) );
XNOR2_X1 _10994_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_03376_ ) );
XNOR2_X1 _10995_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_03377_ ) );
INV_X1 _10996_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_03378_ ) );
INV_X1 _10997_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_03379_ ) );
AOI22_X1 _10998_ ( .A1(_03378_ ), .A2(\ID_EX_csr [9] ), .B1(_03379_ ), .B2(\ID_EX_csr [8] ), .ZN(_03380_ ) );
AND4_X1 _10999_ ( .A1(_03375_ ), .A2(_03376_ ), .A3(_03377_ ), .A4(_03380_ ), .ZN(_03381_ ) );
XNOR2_X1 _11000_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_03382_ ) );
XNOR2_X1 _11001_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_03383_ ) );
AND3_X1 _11002_ ( .A1(_03381_ ), .A2(_03382_ ), .A3(_03383_ ), .ZN(_03384_ ) );
XNOR2_X1 _11003_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_03385_ ) );
XNOR2_X1 _11004_ ( .A(fanout_net_7 ), .B(\ID_EX_csr [0] ), .ZN(_03386_ ) );
XNOR2_X1 _11005_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_03387_ ) );
XNOR2_X1 _11006_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_03388_ ) );
NAND4_X1 _11007_ ( .A1(_03385_ ), .A2(_03386_ ), .A3(_03387_ ), .A4(_03388_ ), .ZN(_03389_ ) );
XOR2_X1 _11008_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .Z(_03390_ ) );
XNOR2_X1 _11009_ ( .A(\EX_LS_dest_csreg_mem [1] ), .B(\ID_EX_csr [1] ), .ZN(_03391_ ) );
INV_X1 _11010_ ( .A(_03391_ ), .ZN(_03392_ ) );
NOR4_X1 _11011_ ( .A1(_03389_ ), .A2(_02332_ ), .A3(_03390_ ), .A4(_03392_ ), .ZN(_03393_ ) );
AND2_X1 _11012_ ( .A1(_03384_ ), .A2(_03393_ ), .ZN(_03394_ ) );
INV_X1 _11013_ ( .A(_03394_ ), .ZN(_03395_ ) );
BUF_X4 _11014_ ( .A(_03395_ ), .Z(_03396_ ) );
AND2_X1 _11015_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_03397_ ) );
NOR2_X1 _11016_ ( .A1(\ID_EX_csr [10] ), .A2(\ID_EX_csr [11] ), .ZN(_03398_ ) );
AND2_X1 _11017_ ( .A1(_03397_ ), .A2(_03398_ ), .ZN(_03399_ ) );
BUF_X4 _11018_ ( .A(_03399_ ), .Z(_03400_ ) );
NOR2_X1 _11019_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_03401_ ) );
NOR2_X1 _11020_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_03402_ ) );
AND2_X1 _11021_ ( .A1(_03401_ ), .A2(_03402_ ), .ZN(_03403_ ) );
AND2_X2 _11022_ ( .A1(_03400_ ), .A2(_03403_ ), .ZN(_03404_ ) );
BUF_X4 _11023_ ( .A(_03404_ ), .Z(_03405_ ) );
BUF_X2 _11024_ ( .A(_03405_ ), .Z(_03406_ ) );
INV_X1 _11025_ ( .A(\ID_EX_csr [0] ), .ZN(_03407_ ) );
NOR2_X1 _11026_ ( .A1(_03407_ ), .A2(\ID_EX_csr [1] ), .ZN(_03408_ ) );
INV_X1 _11027_ ( .A(\ID_EX_csr [3] ), .ZN(_03409_ ) );
AND3_X1 _11028_ ( .A1(_03408_ ), .A2(_03409_ ), .A3(\ID_EX_csr [2] ), .ZN(_03410_ ) );
BUF_X2 _11029_ ( .A(_03410_ ), .Z(_03411_ ) );
AND3_X1 _11030_ ( .A1(_03406_ ), .A2(\mtvec [30] ), .A3(_03411_ ), .ZN(_03412_ ) );
NOR2_X1 _11031_ ( .A1(\ID_EX_csr [3] ), .A2(\ID_EX_csr [2] ), .ZN(_03413_ ) );
INV_X1 _11032_ ( .A(\ID_EX_csr [1] ), .ZN(_03414_ ) );
AND3_X2 _11033_ ( .A1(_03413_ ), .A2(_03414_ ), .A3(_03407_ ), .ZN(_03415_ ) );
BUF_X2 _11034_ ( .A(_03415_ ), .Z(_03416_ ) );
AND3_X1 _11035_ ( .A1(_03406_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_03416_ ), .ZN(_03417_ ) );
NOR2_X1 _11036_ ( .A1(_03412_ ), .A2(_03417_ ), .ZN(_03418_ ) );
NAND2_X1 _11037_ ( .A1(_03413_ ), .A2(\ID_EX_csr [1] ), .ZN(_03419_ ) );
NOR2_X1 _11038_ ( .A1(_03419_ ), .A2(\ID_EX_csr [0] ), .ZN(_03420_ ) );
BUF_X2 _11039_ ( .A(_03420_ ), .Z(_03421_ ) );
INV_X1 _11040_ ( .A(\ID_EX_csr [6] ), .ZN(_03422_ ) );
NOR2_X1 _11041_ ( .A1(_03422_ ), .A2(\ID_EX_csr [7] ), .ZN(_03423_ ) );
AND2_X2 _11042_ ( .A1(_03423_ ), .A2(_03401_ ), .ZN(_03424_ ) );
CLKBUF_X2 _11043_ ( .A(_03424_ ), .Z(_03425_ ) );
CLKBUF_X2 _11044_ ( .A(_03400_ ), .Z(_03426_ ) );
AND4_X1 _11045_ ( .A1(\mycsreg.CSReg[3][30] ), .A2(_03421_ ), .A3(_03425_ ), .A4(_03426_ ), .ZN(_03427_ ) );
AND2_X2 _11046_ ( .A1(_03408_ ), .A2(_03413_ ), .ZN(_03428_ ) );
BUF_X2 _11047_ ( .A(_03428_ ), .Z(_03429_ ) );
AND4_X1 _11048_ ( .A1(\ID_EX_csr [10] ), .A2(_03397_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_03430_ ) );
INV_X1 _11049_ ( .A(\ID_EX_csr [5] ), .ZN(_03431_ ) );
AND2_X1 _11050_ ( .A1(_03402_ ), .A2(_03431_ ), .ZN(_03432_ ) );
AND2_X1 _11051_ ( .A1(_03430_ ), .A2(_03432_ ), .ZN(_03433_ ) );
AOI21_X1 _11052_ ( .A(_03427_ ), .B1(_03429_ ), .B2(_03433_ ), .ZN(_03434_ ) );
BUF_X4 _11053_ ( .A(_03424_ ), .Z(_03435_ ) );
BUF_X4 _11054_ ( .A(_03435_ ), .Z(_03436_ ) );
BUF_X4 _11055_ ( .A(_03436_ ), .Z(_03437_ ) );
BUF_X2 _11056_ ( .A(_03426_ ), .Z(_03438_ ) );
NAND4_X1 _11057_ ( .A1(_03429_ ), .A2(_03437_ ), .A3(\mepc [30] ), .A4(_03438_ ), .ZN(_03439_ ) );
NAND3_X1 _11058_ ( .A1(_03418_ ), .A2(_03434_ ), .A3(_03439_ ), .ZN(_03440_ ) );
NAND2_X1 _11059_ ( .A1(_03396_ ), .A2(_03440_ ), .ZN(_03441_ ) );
BUF_X2 _11060_ ( .A(_03384_ ), .Z(_03442_ ) );
BUF_X2 _11061_ ( .A(_03442_ ), .Z(_03443_ ) );
BUF_X2 _11062_ ( .A(_03393_ ), .Z(_03444_ ) );
BUF_X2 _11063_ ( .A(_03444_ ), .Z(_03445_ ) );
NAND3_X1 _11064_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [30] ), .ZN(_03446_ ) );
AOI21_X1 _11065_ ( .A(_03372_ ), .B1(_03441_ ), .B2(_03446_ ), .ZN(_03447_ ) );
AND2_X1 _11066_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_03448_ ) );
AND2_X1 _11067_ ( .A1(_03448_ ), .A2(\ID_EX_pc [4] ), .ZN(_03449_ ) );
AND2_X1 _11068_ ( .A1(_03449_ ), .A2(\ID_EX_pc [5] ), .ZN(_03450_ ) );
AND2_X1 _11069_ ( .A1(_03450_ ), .A2(\ID_EX_pc [6] ), .ZN(_03451_ ) );
AND2_X1 _11070_ ( .A1(_03451_ ), .A2(\ID_EX_pc [7] ), .ZN(_03452_ ) );
AND2_X1 _11071_ ( .A1(_03452_ ), .A2(\ID_EX_pc [8] ), .ZN(_03453_ ) );
AND2_X2 _11072_ ( .A1(_03453_ ), .A2(\ID_EX_pc [9] ), .ZN(_03454_ ) );
AND2_X1 _11073_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_03455_ ) );
AND2_X1 _11074_ ( .A1(_03454_ ), .A2(_03455_ ), .ZN(_03456_ ) );
AND3_X1 _11075_ ( .A1(_03456_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_03457_ ) );
AND3_X1 _11076_ ( .A1(_03457_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_03458_ ) );
AND3_X1 _11077_ ( .A1(_03458_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_03459_ ) );
AND3_X1 _11078_ ( .A1(_03459_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_03460_ ) );
AND3_X1 _11079_ ( .A1(_03460_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_03461_ ) );
AND3_X1 _11080_ ( .A1(_03461_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_03462_ ) );
AND3_X1 _11081_ ( .A1(_03462_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_03463_ ) );
AND3_X1 _11082_ ( .A1(_03463_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_03464_ ) );
NAND3_X1 _11083_ ( .A1(_03464_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_03465_ ) );
XNOR2_X1 _11084_ ( .A(_03465_ ), .B(\ID_EX_pc [30] ), .ZN(_03466_ ) );
NOR2_X1 _11085_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_8 ), .ZN(_03467_ ) );
AND2_X1 _11086_ ( .A1(_03467_ ), .A2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .ZN(_03468_ ) );
INV_X1 _11087_ ( .A(_03468_ ), .ZN(_03469_ ) );
XNOR2_X1 _11088_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_03470_ ) );
NAND2_X1 _11089_ ( .A1(_02337_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_03471_ ) );
NAND4_X4 _11090_ ( .A1(_02333_ ), .A2(_02336_ ), .A3(_03470_ ), .A4(_03471_ ), .ZN(_03472_ ) );
BUF_X8 _11091_ ( .A(_03472_ ), .Z(_03473_ ) );
XNOR2_X1 _11092_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_03474_ ) );
XNOR2_X1 _11093_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_03475_ ) );
INV_X2 _11094_ ( .A(\ID_EX_rs2 [1] ), .ZN(_03476_ ) );
AOI22_X1 _11095_ ( .A1(_02346_ ), .A2(\ID_EX_rs2 [3] ), .B1(_03476_ ), .B2(\EX_LS_dest_reg [1] ), .ZN(_03477_ ) );
INV_X1 _11096_ ( .A(\ID_EX_rs2 [3] ), .ZN(_03478_ ) );
AOI21_X1 _11097_ ( .A(_02349_ ), .B1(\EX_LS_dest_reg [3] ), .B2(_03478_ ), .ZN(_03479_ ) );
NAND4_X2 _11098_ ( .A1(_03474_ ), .A2(_03475_ ), .A3(_03477_ ), .A4(_03479_ ), .ZN(_03480_ ) );
BUF_X4 _11099_ ( .A(_03480_ ), .Z(_03481_ ) );
NOR2_X4 _11100_ ( .A1(_03473_ ), .A2(_03481_ ), .ZN(_03482_ ) );
INV_X32 _11101_ ( .A(fanout_net_35 ), .ZN(_03483_ ) );
BUF_X2 _11102_ ( .A(_03483_ ), .Z(_03484_ ) );
BUF_X2 _11103_ ( .A(_03484_ ), .Z(_03485_ ) );
CLKBUF_X2 _11104_ ( .A(_03485_ ), .Z(_03486_ ) );
CLKBUF_X2 _11105_ ( .A(_03486_ ), .Z(_03487_ ) );
OR2_X1 _11106_ ( .A1(_03487_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03488_ ) );
INV_X2 _11107_ ( .A(fanout_net_43 ), .ZN(_03489_ ) );
BUF_X4 _11108_ ( .A(_03489_ ), .Z(_03490_ ) );
BUF_X4 _11109_ ( .A(_03490_ ), .Z(_03491_ ) );
BUF_X4 _11110_ ( .A(_03491_ ), .Z(_03492_ ) );
BUF_X4 _11111_ ( .A(_03492_ ), .Z(_03493_ ) );
BUF_X4 _11112_ ( .A(_03493_ ), .Z(_03494_ ) );
OAI211_X1 _11113_ ( .A(_03488_ ), .B(_03494_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03495_ ) );
OR2_X1 _11114_ ( .A1(_03487_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03496_ ) );
OAI211_X1 _11115_ ( .A(_03496_ ), .B(fanout_net_43 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03497_ ) );
INV_X1 _11116_ ( .A(fanout_net_45 ), .ZN(_03498_ ) );
BUF_X4 _11117_ ( .A(_03498_ ), .Z(_03499_ ) );
BUF_X4 _11118_ ( .A(_03499_ ), .Z(_03500_ ) );
BUF_X4 _11119_ ( .A(_03500_ ), .Z(_03501_ ) );
BUF_X4 _11120_ ( .A(_03501_ ), .Z(_03502_ ) );
BUF_X4 _11121_ ( .A(_03502_ ), .Z(_03503_ ) );
BUF_X4 _11122_ ( .A(_03503_ ), .Z(_03504_ ) );
NAND3_X1 _11123_ ( .A1(_03495_ ), .A2(_03497_ ), .A3(_03504_ ), .ZN(_03505_ ) );
MUX2_X1 _11124_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03506_ ) );
MUX2_X1 _11125_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03507_ ) );
BUF_X4 _11126_ ( .A(_03492_ ), .Z(_03508_ ) );
MUX2_X1 _11127_ ( .A(_03506_ ), .B(_03507_ ), .S(_03508_ ), .Z(_03509_ ) );
BUF_X4 _11128_ ( .A(_03503_ ), .Z(_03510_ ) );
OAI211_X1 _11129_ ( .A(fanout_net_46 ), .B(_03505_ ), .C1(_03509_ ), .C2(_03510_ ), .ZN(_03511_ ) );
INV_X1 _11130_ ( .A(fanout_net_46 ), .ZN(_03512_ ) );
BUF_X4 _11131_ ( .A(_03512_ ), .Z(_03513_ ) );
BUF_X4 _11132_ ( .A(_03513_ ), .Z(_03514_ ) );
BUF_X4 _11133_ ( .A(_03514_ ), .Z(_03515_ ) );
CLKBUF_X2 _11134_ ( .A(_03484_ ), .Z(_03516_ ) );
CLKBUF_X2 _11135_ ( .A(_03516_ ), .Z(_03517_ ) );
CLKBUF_X2 _11136_ ( .A(_03517_ ), .Z(_03518_ ) );
BUF_X2 _11137_ ( .A(_03518_ ), .Z(_03519_ ) );
NOR2_X1 _11138_ ( .A1(_03519_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03520_ ) );
OAI21_X1 _11139_ ( .A(fanout_net_43 ), .B1(fanout_net_35 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03521_ ) );
NOR2_X1 _11140_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03522_ ) );
OAI21_X1 _11141_ ( .A(_03508_ ), .B1(_03519_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03523_ ) );
OAI221_X1 _11142_ ( .A(_03503_ ), .B1(_03520_ ), .B2(_03521_ ), .C1(_03522_ ), .C2(_03523_ ), .ZN(_03524_ ) );
MUX2_X1 _11143_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03525_ ) );
MUX2_X1 _11144_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03526_ ) );
MUX2_X1 _11145_ ( .A(_03525_ ), .B(_03526_ ), .S(_03508_ ), .Z(_03527_ ) );
OAI211_X1 _11146_ ( .A(_03515_ ), .B(_03524_ ), .C1(_03527_ ), .C2(_03504_ ), .ZN(_03528_ ) );
AOI21_X1 _11147_ ( .A(_03482_ ), .B1(_03511_ ), .B2(_03528_ ), .ZN(_03529_ ) );
BUF_X16 _11148_ ( .A(_03473_ ), .Z(_03530_ ) );
BUF_X8 _11149_ ( .A(_03530_ ), .Z(_03531_ ) );
BUF_X16 _11150_ ( .A(_03531_ ), .Z(_03532_ ) );
BUF_X4 _11151_ ( .A(_03481_ ), .Z(_03533_ ) );
BUF_X8 _11152_ ( .A(_03533_ ), .Z(_03534_ ) );
BUF_X2 _11153_ ( .A(_03534_ ), .Z(_03535_ ) );
NOR3_X1 _11154_ ( .A1(_03532_ ), .A2(\EX_LS_result_reg [26] ), .A3(_03535_ ), .ZN(_03536_ ) );
NOR2_X1 _11155_ ( .A1(_03529_ ), .A2(_03536_ ), .ZN(_03537_ ) );
XNOR2_X2 _11156_ ( .A(_03537_ ), .B(_03120_ ), .ZN(_03538_ ) );
OR2_X1 _11157_ ( .A1(_03487_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03539_ ) );
OAI211_X1 _11158_ ( .A(_03539_ ), .B(_03494_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03540_ ) );
OR2_X1 _11159_ ( .A1(_03487_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03541_ ) );
OAI211_X1 _11160_ ( .A(_03541_ ), .B(fanout_net_43 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03542_ ) );
NAND3_X1 _11161_ ( .A1(_03540_ ), .A2(_03542_ ), .A3(_03504_ ), .ZN(_03543_ ) );
MUX2_X1 _11162_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03544_ ) );
MUX2_X1 _11163_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03545_ ) );
MUX2_X1 _11164_ ( .A(_03544_ ), .B(_03545_ ), .S(_03508_ ), .Z(_03546_ ) );
OAI211_X1 _11165_ ( .A(fanout_net_46 ), .B(_03543_ ), .C1(_03546_ ), .C2(_03504_ ), .ZN(_03547_ ) );
MUX2_X1 _11166_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03548_ ) );
AND2_X1 _11167_ ( .A1(_03548_ ), .A2(_03493_ ), .ZN(_03549_ ) );
MUX2_X1 _11168_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03550_ ) );
AOI211_X1 _11169_ ( .A(fanout_net_45 ), .B(_03549_ ), .C1(fanout_net_43 ), .C2(_03550_ ), .ZN(_03551_ ) );
MUX2_X1 _11170_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03552_ ) );
MUX2_X1 _11171_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03553_ ) );
MUX2_X1 _11172_ ( .A(_03552_ ), .B(_03553_ ), .S(_03493_ ), .Z(_03554_ ) );
OAI21_X1 _11173_ ( .A(_03515_ ), .B1(_03554_ ), .B2(_03504_ ), .ZN(_03555_ ) );
OAI221_X1 _11174_ ( .A(_03547_ ), .B1(_03551_ ), .B2(_03555_ ), .C1(_03532_ ), .C2(_03535_ ), .ZN(_03556_ ) );
INV_X1 _11175_ ( .A(\EX_LS_result_reg [27] ), .ZN(_03557_ ) );
OR3_X1 _11176_ ( .A1(_03532_ ), .A2(_03557_ ), .A3(_03535_ ), .ZN(_03558_ ) );
NAND2_X1 _11177_ ( .A1(_03556_ ), .A2(_03558_ ), .ZN(_03559_ ) );
NAND2_X1 _11178_ ( .A1(_03076_ ), .A2(_03096_ ), .ZN(_03560_ ) );
XNOR2_X1 _11179_ ( .A(_03559_ ), .B(_03560_ ), .ZN(_03561_ ) );
AND2_X1 _11180_ ( .A1(_03538_ ), .A2(_03561_ ), .ZN(_03562_ ) );
NAND2_X1 _11181_ ( .A1(_03482_ ), .A2(\EX_LS_result_reg [24] ), .ZN(_03563_ ) );
BUF_X2 _11182_ ( .A(_03487_ ), .Z(_03564_ ) );
OR2_X1 _11183_ ( .A1(_03564_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03565_ ) );
OAI211_X1 _11184_ ( .A(_03565_ ), .B(fanout_net_43 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03566_ ) );
OR2_X1 _11185_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03567_ ) );
BUF_X4 _11186_ ( .A(_03508_ ), .Z(_03568_ ) );
OAI211_X1 _11187_ ( .A(_03567_ ), .B(_03568_ ), .C1(_03564_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03569_ ) );
NAND3_X1 _11188_ ( .A1(_03566_ ), .A2(fanout_net_45 ), .A3(_03569_ ), .ZN(_03570_ ) );
MUX2_X1 _11189_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03571_ ) );
MUX2_X1 _11190_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03572_ ) );
MUX2_X1 _11191_ ( .A(_03571_ ), .B(_03572_ ), .S(_03568_ ), .Z(_03573_ ) );
OAI211_X1 _11192_ ( .A(_03515_ ), .B(_03570_ ), .C1(_03573_ ), .C2(fanout_net_45 ), .ZN(_03574_ ) );
NOR2_X1 _11193_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03575_ ) );
OAI21_X1 _11194_ ( .A(_03568_ ), .B1(_03564_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03576_ ) );
MUX2_X1 _11195_ ( .A(_03038_ ), .B(_03039_ ), .S(fanout_net_35 ), .Z(_03577_ ) );
OAI221_X1 _11196_ ( .A(_03510_ ), .B1(_03575_ ), .B2(_03576_ ), .C1(_03577_ ), .C2(_03568_ ), .ZN(_03578_ ) );
MUX2_X1 _11197_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03579_ ) );
MUX2_X1 _11198_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03580_ ) );
MUX2_X1 _11199_ ( .A(_03579_ ), .B(_03580_ ), .S(fanout_net_43 ), .Z(_03581_ ) );
OAI211_X1 _11200_ ( .A(fanout_net_46 ), .B(_03578_ ), .C1(_03581_ ), .C2(_03510_ ), .ZN(_03582_ ) );
BUF_X8 _11201_ ( .A(_03532_ ), .Z(_03583_ ) );
BUF_X2 _11202_ ( .A(_03535_ ), .Z(_03584_ ) );
OAI211_X1 _11203_ ( .A(_03574_ ), .B(_03582_ ), .C1(_03583_ ), .C2(_03584_ ), .ZN(_03585_ ) );
NAND2_X1 _11204_ ( .A1(_03563_ ), .A2(_03585_ ), .ZN(_03586_ ) );
XNOR2_X1 _11205_ ( .A(_03586_ ), .B(_03047_ ), .ZN(_03587_ ) );
INV_X1 _11206_ ( .A(\EX_LS_result_reg [25] ), .ZN(_03588_ ) );
OR3_X2 _11207_ ( .A1(_03583_ ), .A2(_03588_ ), .A3(_03584_ ), .ZN(_03589_ ) );
OR2_X1 _11208_ ( .A1(_03519_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03590_ ) );
OAI211_X1 _11209_ ( .A(_03590_ ), .B(_03568_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03591_ ) );
OR2_X1 _11210_ ( .A1(_03519_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03592_ ) );
OAI211_X1 _11211_ ( .A(_03592_ ), .B(fanout_net_43 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03593_ ) );
NAND3_X1 _11212_ ( .A1(_03591_ ), .A2(_03593_ ), .A3(fanout_net_45 ), .ZN(_03594_ ) );
MUX2_X1 _11213_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03595_ ) );
MUX2_X1 _11214_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_03596_ ) );
MUX2_X1 _11215_ ( .A(_03595_ ), .B(_03596_ ), .S(_03494_ ), .Z(_03597_ ) );
OAI211_X1 _11216_ ( .A(_03515_ ), .B(_03594_ ), .C1(_03597_ ), .C2(fanout_net_45 ), .ZN(_03598_ ) );
NOR2_X1 _11217_ ( .A1(_03564_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03599_ ) );
OAI21_X1 _11218_ ( .A(fanout_net_43 ), .B1(fanout_net_35 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03600_ ) );
NOR2_X1 _11219_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03601_ ) );
OAI21_X1 _11220_ ( .A(_03494_ ), .B1(_03564_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03602_ ) );
OAI221_X1 _11221_ ( .A(_03504_ ), .B1(_03599_ ), .B2(_03600_ ), .C1(_03601_ ), .C2(_03602_ ), .ZN(_03603_ ) );
MUX2_X1 _11222_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03604_ ) );
MUX2_X1 _11223_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03605_ ) );
MUX2_X1 _11224_ ( .A(_03604_ ), .B(_03605_ ), .S(fanout_net_43 ), .Z(_03606_ ) );
OAI211_X1 _11225_ ( .A(fanout_net_46 ), .B(_03603_ ), .C1(_03606_ ), .C2(_03510_ ), .ZN(_03607_ ) );
OAI211_X1 _11226_ ( .A(_03598_ ), .B(_03607_ ), .C1(_03583_ ), .C2(_03584_ ), .ZN(_03608_ ) );
NAND2_X1 _11227_ ( .A1(_03589_ ), .A2(_03608_ ), .ZN(_03609_ ) );
XNOR2_X1 _11228_ ( .A(_03073_ ), .B(_03609_ ), .ZN(_03610_ ) );
AND3_X1 _11229_ ( .A1(_03562_ ), .A2(_03587_ ), .A3(_03610_ ), .ZN(_03611_ ) );
OR3_X1 _11230_ ( .A1(_03532_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_03535_ ), .ZN(_03612_ ) );
OR2_X1 _11231_ ( .A1(_03487_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03613_ ) );
OAI211_X1 _11232_ ( .A(_03613_ ), .B(fanout_net_43 ), .C1(fanout_net_36 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03614_ ) );
OR2_X1 _11233_ ( .A1(fanout_net_36 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03615_ ) );
OAI211_X1 _11234_ ( .A(_03615_ ), .B(_03494_ ), .C1(_03564_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03616_ ) );
NAND3_X1 _11235_ ( .A1(_03614_ ), .A2(fanout_net_45 ), .A3(_03616_ ), .ZN(_03617_ ) );
MUX2_X1 _11236_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03618_ ) );
MUX2_X1 _11237_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03619_ ) );
MUX2_X1 _11238_ ( .A(_03618_ ), .B(_03619_ ), .S(_03508_ ), .Z(_03620_ ) );
OAI211_X1 _11239_ ( .A(_03515_ ), .B(_03617_ ), .C1(_03620_ ), .C2(fanout_net_45 ), .ZN(_03621_ ) );
NOR2_X1 _11240_ ( .A1(fanout_net_36 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03622_ ) );
OAI21_X1 _11241_ ( .A(_03493_ ), .B1(_03519_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03623_ ) );
MUX2_X1 _11242_ ( .A(_02375_ ), .B(_02376_ ), .S(fanout_net_36 ), .Z(_03624_ ) );
OAI221_X1 _11243_ ( .A(_03504_ ), .B1(_03622_ ), .B2(_03623_ ), .C1(_03624_ ), .C2(_03494_ ), .ZN(_03625_ ) );
MUX2_X1 _11244_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03626_ ) );
MUX2_X1 _11245_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03627_ ) );
MUX2_X1 _11246_ ( .A(_03626_ ), .B(_03627_ ), .S(fanout_net_43 ), .Z(_03628_ ) );
OAI211_X1 _11247_ ( .A(fanout_net_46 ), .B(_03625_ ), .C1(_03628_ ), .C2(_03510_ ), .ZN(_03629_ ) );
OAI211_X1 _11248_ ( .A(_03621_ ), .B(_03629_ ), .C1(_03583_ ), .C2(_03584_ ), .ZN(_03630_ ) );
NAND2_X1 _11249_ ( .A1(_03612_ ), .A2(_03630_ ), .ZN(_03631_ ) );
XNOR2_X1 _11250_ ( .A(_03631_ ), .B(_02388_ ), .ZN(_03632_ ) );
OR3_X1 _11251_ ( .A1(_03532_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03535_ ), .ZN(_03633_ ) );
OR2_X1 _11252_ ( .A1(_03518_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03634_ ) );
OAI211_X1 _11253_ ( .A(_03634_ ), .B(_03508_ ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03635_ ) );
OR2_X1 _11254_ ( .A1(_03518_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03636_ ) );
OAI211_X1 _11255_ ( .A(_03636_ ), .B(fanout_net_43 ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03637_ ) );
NAND3_X1 _11256_ ( .A1(_03635_ ), .A2(_03637_ ), .A3(_03503_ ), .ZN(_03638_ ) );
MUX2_X1 _11257_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03639_ ) );
MUX2_X1 _11258_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03640_ ) );
MUX2_X1 _11259_ ( .A(_03639_ ), .B(_03640_ ), .S(_03508_ ), .Z(_03641_ ) );
OAI211_X1 _11260_ ( .A(fanout_net_46 ), .B(_03638_ ), .C1(_03641_ ), .C2(_03504_ ), .ZN(_03642_ ) );
NOR2_X1 _11261_ ( .A1(_03519_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03643_ ) );
OAI21_X1 _11262_ ( .A(fanout_net_43 ), .B1(fanout_net_36 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03644_ ) );
NOR2_X1 _11263_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03645_ ) );
OAI21_X1 _11264_ ( .A(_03508_ ), .B1(_03519_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03646_ ) );
OAI221_X1 _11265_ ( .A(_03503_ ), .B1(_03643_ ), .B2(_03644_ ), .C1(_03645_ ), .C2(_03646_ ), .ZN(_03647_ ) );
MUX2_X1 _11266_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03648_ ) );
MUX2_X1 _11267_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03649_ ) );
MUX2_X1 _11268_ ( .A(_03648_ ), .B(_03649_ ), .S(_03508_ ), .Z(_03650_ ) );
OAI211_X1 _11269_ ( .A(_03515_ ), .B(_03647_ ), .C1(_03650_ ), .C2(_03504_ ), .ZN(_03651_ ) );
OAI211_X1 _11270_ ( .A(_03642_ ), .B(_03651_ ), .C1(_03532_ ), .C2(_03535_ ), .ZN(_03652_ ) );
NAND2_X1 _11271_ ( .A1(_03633_ ), .A2(_03652_ ), .ZN(_03653_ ) );
XNOR2_X1 _11272_ ( .A(_03150_ ), .B(_03653_ ), .ZN(_03654_ ) );
AND2_X1 _11273_ ( .A1(_03632_ ), .A2(_03654_ ), .ZN(_03655_ ) );
OR3_X1 _11274_ ( .A1(_03583_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03584_ ), .ZN(_03656_ ) );
OR2_X1 _11275_ ( .A1(_03564_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03657_ ) );
OAI211_X1 _11276_ ( .A(_03657_ ), .B(_03568_ ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03658_ ) );
NAND2_X1 _11277_ ( .A1(_03164_ ), .A2(fanout_net_36 ), .ZN(_03659_ ) );
OAI211_X1 _11278_ ( .A(_03659_ ), .B(fanout_net_43 ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03660_ ) );
NAND3_X1 _11279_ ( .A1(_03658_ ), .A2(_03510_ ), .A3(_03660_ ), .ZN(_03661_ ) );
MUX2_X1 _11280_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03662_ ) );
MUX2_X1 _11281_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03663_ ) );
MUX2_X1 _11282_ ( .A(_03662_ ), .B(_03663_ ), .S(_03568_ ), .Z(_03664_ ) );
OAI211_X1 _11283_ ( .A(_03515_ ), .B(_03661_ ), .C1(_03664_ ), .C2(_03510_ ), .ZN(_03665_ ) );
OR2_X1 _11284_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03666_ ) );
OAI211_X1 _11285_ ( .A(_03666_ ), .B(_03568_ ), .C1(_03564_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03667_ ) );
NAND2_X1 _11286_ ( .A1(_03174_ ), .A2(fanout_net_36 ), .ZN(_03668_ ) );
OAI211_X1 _11287_ ( .A(_03668_ ), .B(fanout_net_43 ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03669_ ) );
NAND3_X1 _11288_ ( .A1(_03667_ ), .A2(_03669_ ), .A3(fanout_net_45 ), .ZN(_03670_ ) );
MUX2_X1 _11289_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03671_ ) );
MUX2_X1 _11290_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_03672_ ) );
MUX2_X1 _11291_ ( .A(_03671_ ), .B(_03672_ ), .S(fanout_net_43 ), .Z(_03673_ ) );
OAI211_X1 _11292_ ( .A(fanout_net_46 ), .B(_03670_ ), .C1(_03673_ ), .C2(fanout_net_45 ), .ZN(_03674_ ) );
OAI211_X1 _11293_ ( .A(_03665_ ), .B(_03674_ ), .C1(_03583_ ), .C2(_03584_ ), .ZN(_03675_ ) );
NAND2_X1 _11294_ ( .A1(_03656_ ), .A2(_03675_ ), .ZN(_03676_ ) );
XNOR2_X1 _11295_ ( .A(_03184_ ), .B(_03676_ ), .ZN(_03677_ ) );
OR3_X1 _11296_ ( .A1(_03583_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_03584_ ), .ZN(_03678_ ) );
OR2_X1 _11297_ ( .A1(_03519_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03679_ ) );
OAI211_X1 _11298_ ( .A(_03679_ ), .B(_03568_ ), .C1(fanout_net_36 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03680_ ) );
OR2_X1 _11299_ ( .A1(_03519_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03681_ ) );
OAI211_X1 _11300_ ( .A(_03681_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03682_ ) );
NAND3_X1 _11301_ ( .A1(_03680_ ), .A2(_03682_ ), .A3(fanout_net_45 ), .ZN(_03683_ ) );
MUX2_X1 _11302_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_03684_ ) );
MUX2_X1 _11303_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_03685_ ) );
MUX2_X1 _11304_ ( .A(_03684_ ), .B(_03685_ ), .S(_03494_ ), .Z(_03686_ ) );
OAI211_X1 _11305_ ( .A(_03515_ ), .B(_03683_ ), .C1(_03686_ ), .C2(fanout_net_45 ), .ZN(_03687_ ) );
NOR2_X1 _11306_ ( .A1(_03564_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03688_ ) );
OAI21_X1 _11307_ ( .A(fanout_net_43 ), .B1(fanout_net_37 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03689_ ) );
NOR2_X1 _11308_ ( .A1(fanout_net_37 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03690_ ) );
OAI21_X1 _11309_ ( .A(_03494_ ), .B1(_03564_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03691_ ) );
OAI221_X1 _11310_ ( .A(_03504_ ), .B1(_03688_ ), .B2(_03689_ ), .C1(_03690_ ), .C2(_03691_ ), .ZN(_03692_ ) );
MUX2_X1 _11311_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_03693_ ) );
MUX2_X1 _11312_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_03694_ ) );
MUX2_X1 _11313_ ( .A(_03693_ ), .B(_03694_ ), .S(fanout_net_43 ), .Z(_03695_ ) );
OAI211_X1 _11314_ ( .A(fanout_net_46 ), .B(_03692_ ), .C1(_03695_ ), .C2(_03510_ ), .ZN(_03696_ ) );
OAI211_X1 _11315_ ( .A(_03687_ ), .B(_03696_ ), .C1(_03583_ ), .C2(_03584_ ), .ZN(_03697_ ) );
NAND2_X1 _11316_ ( .A1(_03678_ ), .A2(_03697_ ), .ZN(_03698_ ) );
INV_X1 _11317_ ( .A(_03698_ ), .ZN(_03699_ ) );
XNOR2_X1 _11318_ ( .A(_03699_ ), .B(_02358_ ), .ZN(_03700_ ) );
AND3_X1 _11319_ ( .A1(_03655_ ), .A2(_03677_ ), .A3(_03700_ ), .ZN(_03701_ ) );
AND2_X2 _11320_ ( .A1(_03611_ ), .A2(_03701_ ), .ZN(_03702_ ) );
INV_X1 _11321_ ( .A(_02438_ ), .ZN(_03703_ ) );
INV_X1 _11322_ ( .A(\EX_LS_result_reg [23] ), .ZN(_03704_ ) );
OR3_X1 _11323_ ( .A1(_03530_ ), .A2(_03704_ ), .A3(_03533_ ), .ZN(_03705_ ) );
BUF_X2 _11324_ ( .A(_03484_ ), .Z(_03706_ ) );
OR2_X1 _11325_ ( .A1(_03706_ ), .A2(\myreg.Reg[1][23] ), .ZN(_03707_ ) );
BUF_X4 _11326_ ( .A(_03489_ ), .Z(_03708_ ) );
BUF_X4 _11327_ ( .A(_03708_ ), .Z(_03709_ ) );
BUF_X4 _11328_ ( .A(_03709_ ), .Z(_03710_ ) );
OAI211_X1 _11329_ ( .A(_03707_ ), .B(_03710_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[0][23] ), .ZN(_03711_ ) );
OR2_X1 _11330_ ( .A1(_03485_ ), .A2(\myreg.Reg[3][23] ), .ZN(_03712_ ) );
OAI211_X1 _11331_ ( .A(_03712_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[2][23] ), .ZN(_03713_ ) );
NAND3_X1 _11332_ ( .A1(_03711_ ), .A2(_03713_ ), .A3(_03501_ ), .ZN(_03714_ ) );
MUX2_X1 _11333_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_37 ), .Z(_03715_ ) );
MUX2_X1 _11334_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_37 ), .Z(_03716_ ) );
MUX2_X1 _11335_ ( .A(_03715_ ), .B(_03716_ ), .S(_03491_ ), .Z(_03717_ ) );
OAI211_X1 _11336_ ( .A(_03514_ ), .B(_03714_ ), .C1(_03717_ ), .C2(_03501_ ), .ZN(_03718_ ) );
OR2_X1 _11337_ ( .A1(_03485_ ), .A2(\myreg.Reg[15][23] ), .ZN(_03719_ ) );
OAI211_X1 _11338_ ( .A(_03719_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][23] ), .ZN(_03720_ ) );
OR2_X1 _11339_ ( .A1(_03485_ ), .A2(\myreg.Reg[13][23] ), .ZN(_03721_ ) );
OAI211_X1 _11340_ ( .A(_03721_ ), .B(_03710_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[12][23] ), .ZN(_03722_ ) );
NAND3_X1 _11341_ ( .A1(_03720_ ), .A2(_03722_ ), .A3(fanout_net_45 ), .ZN(_03723_ ) );
MUX2_X1 _11342_ ( .A(\myreg.Reg[8][23] ), .B(\myreg.Reg[9][23] ), .S(fanout_net_37 ), .Z(_03724_ ) );
MUX2_X1 _11343_ ( .A(\myreg.Reg[10][23] ), .B(\myreg.Reg[11][23] ), .S(fanout_net_37 ), .Z(_03725_ ) );
MUX2_X1 _11344_ ( .A(_03724_ ), .B(_03725_ ), .S(fanout_net_43 ), .Z(_03726_ ) );
OAI211_X1 _11345_ ( .A(fanout_net_46 ), .B(_03723_ ), .C1(_03726_ ), .C2(fanout_net_45 ), .ZN(_03727_ ) );
NAND2_X1 _11346_ ( .A1(_03718_ ), .A2(_03727_ ), .ZN(_03728_ ) );
OAI21_X1 _11347_ ( .A(_03728_ ), .B1(_03531_ ), .B2(_03534_ ), .ZN(_03729_ ) );
AND2_X2 _11348_ ( .A1(_03705_ ), .A2(_03729_ ), .ZN(_03730_ ) );
XNOR2_X1 _11349_ ( .A(_03703_ ), .B(_03730_ ), .ZN(_03731_ ) );
OR3_X1 _11350_ ( .A1(_03531_ ), .A2(\EX_LS_result_reg [22] ), .A3(_03534_ ), .ZN(_03732_ ) );
OR2_X1 _11351_ ( .A1(_03486_ ), .A2(\myreg.Reg[1][22] ), .ZN(_03733_ ) );
OAI211_X1 _11352_ ( .A(_03733_ ), .B(_03492_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[0][22] ), .ZN(_03734_ ) );
OR2_X1 _11353_ ( .A1(_03486_ ), .A2(\myreg.Reg[3][22] ), .ZN(_03735_ ) );
OAI211_X1 _11354_ ( .A(_03735_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[2][22] ), .ZN(_03736_ ) );
NAND3_X1 _11355_ ( .A1(_03734_ ), .A2(_03736_ ), .A3(_03502_ ), .ZN(_03737_ ) );
MUX2_X1 _11356_ ( .A(\myreg.Reg[6][22] ), .B(\myreg.Reg[7][22] ), .S(fanout_net_37 ), .Z(_03738_ ) );
MUX2_X1 _11357_ ( .A(\myreg.Reg[4][22] ), .B(\myreg.Reg[5][22] ), .S(fanout_net_37 ), .Z(_03739_ ) );
MUX2_X1 _11358_ ( .A(_03738_ ), .B(_03739_ ), .S(_03492_ ), .Z(_03740_ ) );
OAI211_X1 _11359_ ( .A(_03514_ ), .B(_03737_ ), .C1(_03740_ ), .C2(_03503_ ), .ZN(_03741_ ) );
OR2_X1 _11360_ ( .A1(_03486_ ), .A2(\myreg.Reg[15][22] ), .ZN(_03742_ ) );
OAI211_X1 _11361_ ( .A(_03742_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][22] ), .ZN(_03743_ ) );
OR2_X1 _11362_ ( .A1(_03486_ ), .A2(\myreg.Reg[13][22] ), .ZN(_03744_ ) );
OAI211_X1 _11363_ ( .A(_03744_ ), .B(_03492_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[12][22] ), .ZN(_03745_ ) );
NAND3_X1 _11364_ ( .A1(_03743_ ), .A2(_03745_ ), .A3(fanout_net_45 ), .ZN(_03746_ ) );
MUX2_X1 _11365_ ( .A(\myreg.Reg[8][22] ), .B(\myreg.Reg[9][22] ), .S(fanout_net_37 ), .Z(_03747_ ) );
MUX2_X1 _11366_ ( .A(\myreg.Reg[10][22] ), .B(\myreg.Reg[11][22] ), .S(fanout_net_37 ), .Z(_03748_ ) );
MUX2_X1 _11367_ ( .A(_03747_ ), .B(_03748_ ), .S(fanout_net_43 ), .Z(_03749_ ) );
OAI211_X1 _11368_ ( .A(fanout_net_46 ), .B(_03746_ ), .C1(_03749_ ), .C2(fanout_net_45 ), .ZN(_03750_ ) );
OAI211_X1 _11369_ ( .A(_03741_ ), .B(_03750_ ), .C1(_03532_ ), .C2(_03535_ ), .ZN(_03751_ ) );
NAND2_X1 _11370_ ( .A1(_03732_ ), .A2(_03751_ ), .ZN(_03752_ ) );
XOR2_X1 _11371_ ( .A(_02410_ ), .B(_03752_ ), .Z(_03753_ ) );
AND2_X1 _11372_ ( .A1(_03731_ ), .A2(_03753_ ), .ZN(_03754_ ) );
OR2_X1 _11373_ ( .A1(_03518_ ), .A2(\myreg.Reg[1][21] ), .ZN(_03755_ ) );
OAI211_X1 _11374_ ( .A(_03755_ ), .B(_03493_ ), .C1(\myreg.Reg[0][21] ), .C2(fanout_net_37 ), .ZN(_03756_ ) );
OR2_X1 _11375_ ( .A1(_03518_ ), .A2(\myreg.Reg[3][21] ), .ZN(_03757_ ) );
OAI211_X1 _11376_ ( .A(_03757_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[2][21] ), .ZN(_03758_ ) );
NAND3_X1 _11377_ ( .A1(_03756_ ), .A2(_03758_ ), .A3(_03503_ ), .ZN(_03759_ ) );
MUX2_X1 _11378_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_37 ), .Z(_03760_ ) );
MUX2_X1 _11379_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_37 ), .Z(_03761_ ) );
MUX2_X1 _11380_ ( .A(_03760_ ), .B(_03761_ ), .S(_03493_ ), .Z(_03762_ ) );
OAI211_X1 _11381_ ( .A(_03514_ ), .B(_03759_ ), .C1(_03762_ ), .C2(_03503_ ), .ZN(_03763_ ) );
OR2_X1 _11382_ ( .A1(_03518_ ), .A2(\myreg.Reg[15][21] ), .ZN(_03764_ ) );
OAI211_X1 _11383_ ( .A(_03764_ ), .B(fanout_net_43 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][21] ), .ZN(_03765_ ) );
OR2_X1 _11384_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][21] ), .ZN(_03766_ ) );
OAI211_X1 _11385_ ( .A(_03766_ ), .B(_03493_ ), .C1(_03487_ ), .C2(\myreg.Reg[13][21] ), .ZN(_03767_ ) );
NAND3_X1 _11386_ ( .A1(_03765_ ), .A2(fanout_net_45 ), .A3(_03767_ ), .ZN(_03768_ ) );
MUX2_X1 _11387_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_37 ), .Z(_03769_ ) );
MUX2_X1 _11388_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_38 ), .Z(_03770_ ) );
MUX2_X1 _11389_ ( .A(_03769_ ), .B(_03770_ ), .S(fanout_net_43 ), .Z(_03771_ ) );
OAI211_X1 _11390_ ( .A(fanout_net_46 ), .B(_03768_ ), .C1(_03771_ ), .C2(fanout_net_45 ), .ZN(_03772_ ) );
AOI21_X1 _11391_ ( .A(_03482_ ), .B1(_03763_ ), .B2(_03772_ ), .ZN(_03773_ ) );
INV_X1 _11392_ ( .A(\EX_LS_result_reg [21] ), .ZN(_03774_ ) );
NOR3_X1 _11393_ ( .A1(_03532_ ), .A2(_03774_ ), .A3(_03535_ ), .ZN(_03775_ ) );
NOR2_X1 _11394_ ( .A1(_03773_ ), .A2(_03775_ ), .ZN(_03776_ ) );
NAND2_X1 _11395_ ( .A1(_02441_ ), .A2(_02461_ ), .ZN(_03777_ ) );
INV_X1 _11396_ ( .A(_03777_ ), .ZN(_03778_ ) );
XNOR2_X1 _11397_ ( .A(_03776_ ), .B(_03778_ ), .ZN(_03779_ ) );
OR3_X1 _11398_ ( .A1(_03531_ ), .A2(\EX_LS_result_reg [20] ), .A3(_03534_ ), .ZN(_03780_ ) );
OR2_X1 _11399_ ( .A1(_03518_ ), .A2(\myreg.Reg[1][20] ), .ZN(_03781_ ) );
OAI211_X1 _11400_ ( .A(_03781_ ), .B(_03493_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[0][20] ), .ZN(_03782_ ) );
OR2_X1 _11401_ ( .A1(_03518_ ), .A2(\myreg.Reg[3][20] ), .ZN(_03783_ ) );
OAI211_X1 _11402_ ( .A(_03783_ ), .B(fanout_net_43 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[2][20] ), .ZN(_03784_ ) );
NAND3_X1 _11403_ ( .A1(_03782_ ), .A2(_03784_ ), .A3(_03503_ ), .ZN(_03785_ ) );
MUX2_X1 _11404_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_38 ), .Z(_03786_ ) );
MUX2_X1 _11405_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_38 ), .Z(_03787_ ) );
MUX2_X1 _11406_ ( .A(_03786_ ), .B(_03787_ ), .S(_03493_ ), .Z(_03788_ ) );
OAI211_X1 _11407_ ( .A(_03515_ ), .B(_03785_ ), .C1(_03788_ ), .C2(_03503_ ), .ZN(_03789_ ) );
OR2_X1 _11408_ ( .A1(_03518_ ), .A2(\myreg.Reg[15][20] ), .ZN(_03790_ ) );
OAI211_X1 _11409_ ( .A(_03790_ ), .B(fanout_net_44 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[14][20] ), .ZN(_03791_ ) );
OR2_X1 _11410_ ( .A1(_03518_ ), .A2(\myreg.Reg[13][20] ), .ZN(_03792_ ) );
OAI211_X1 _11411_ ( .A(_03792_ ), .B(_03493_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[12][20] ), .ZN(_03793_ ) );
NAND3_X1 _11412_ ( .A1(_03791_ ), .A2(_03793_ ), .A3(fanout_net_45 ), .ZN(_03794_ ) );
MUX2_X1 _11413_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_38 ), .Z(_03795_ ) );
MUX2_X1 _11414_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_38 ), .Z(_03796_ ) );
MUX2_X1 _11415_ ( .A(_03795_ ), .B(_03796_ ), .S(fanout_net_44 ), .Z(_03797_ ) );
OAI211_X1 _11416_ ( .A(fanout_net_46 ), .B(_03794_ ), .C1(_03797_ ), .C2(fanout_net_45 ), .ZN(_03798_ ) );
OAI211_X1 _11417_ ( .A(_03789_ ), .B(_03798_ ), .C1(_03532_ ), .C2(_03535_ ), .ZN(_03799_ ) );
NAND2_X1 _11418_ ( .A1(_03780_ ), .A2(_03799_ ), .ZN(_03800_ ) );
XOR2_X1 _11419_ ( .A(_02485_ ), .B(_03800_ ), .Z(_03801_ ) );
AND3_X1 _11420_ ( .A1(_03754_ ), .A2(_03779_ ), .A3(_03801_ ), .ZN(_03802_ ) );
INV_X1 _11421_ ( .A(_02533_ ), .ZN(_03803_ ) );
INV_X1 _11422_ ( .A(\EX_LS_result_reg [19] ), .ZN(_03804_ ) );
OR3_X4 _11423_ ( .A1(_03531_ ), .A2(_03804_ ), .A3(_03534_ ), .ZN(_03805_ ) );
OR2_X1 _11424_ ( .A1(_03517_ ), .A2(\myreg.Reg[1][19] ), .ZN(_03806_ ) );
OAI211_X1 _11425_ ( .A(_03806_ ), .B(_03492_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[0][19] ), .ZN(_03807_ ) );
OR2_X1 _11426_ ( .A1(_03706_ ), .A2(\myreg.Reg[3][19] ), .ZN(_03808_ ) );
OAI211_X1 _11427_ ( .A(_03808_ ), .B(fanout_net_44 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[2][19] ), .ZN(_03809_ ) );
NAND3_X1 _11428_ ( .A1(_03807_ ), .A2(_03809_ ), .A3(_03502_ ), .ZN(_03810_ ) );
MUX2_X1 _11429_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_38 ), .Z(_03811_ ) );
MUX2_X1 _11430_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_38 ), .Z(_03812_ ) );
MUX2_X1 _11431_ ( .A(_03811_ ), .B(_03812_ ), .S(_03710_ ), .Z(_03813_ ) );
OAI211_X1 _11432_ ( .A(_03514_ ), .B(_03810_ ), .C1(_03813_ ), .C2(_03502_ ), .ZN(_03814_ ) );
OR2_X1 _11433_ ( .A1(_03517_ ), .A2(\myreg.Reg[15][19] ), .ZN(_03815_ ) );
OAI211_X1 _11434_ ( .A(_03815_ ), .B(fanout_net_44 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[14][19] ), .ZN(_03816_ ) );
OR2_X1 _11435_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[12][19] ), .ZN(_03817_ ) );
OAI211_X1 _11436_ ( .A(_03817_ ), .B(_03710_ ), .C1(_03486_ ), .C2(\myreg.Reg[13][19] ), .ZN(_03818_ ) );
NAND3_X1 _11437_ ( .A1(_03816_ ), .A2(fanout_net_45 ), .A3(_03818_ ), .ZN(_03819_ ) );
MUX2_X1 _11438_ ( .A(\myreg.Reg[8][19] ), .B(\myreg.Reg[9][19] ), .S(fanout_net_38 ), .Z(_03820_ ) );
MUX2_X1 _11439_ ( .A(\myreg.Reg[10][19] ), .B(\myreg.Reg[11][19] ), .S(fanout_net_38 ), .Z(_03821_ ) );
MUX2_X1 _11440_ ( .A(_03820_ ), .B(_03821_ ), .S(fanout_net_44 ), .Z(_03822_ ) );
OAI211_X1 _11441_ ( .A(fanout_net_46 ), .B(_03819_ ), .C1(_03822_ ), .C2(fanout_net_45 ), .ZN(_03823_ ) );
NAND2_X1 _11442_ ( .A1(_03814_ ), .A2(_03823_ ), .ZN(_03824_ ) );
OAI21_X1 _11443_ ( .A(_03824_ ), .B1(_03531_ ), .B2(_03534_ ), .ZN(_03825_ ) );
AND2_X1 _11444_ ( .A1(_03805_ ), .A2(_03825_ ), .ZN(_03826_ ) );
XNOR2_X1 _11445_ ( .A(_03803_ ), .B(_03826_ ), .ZN(_03827_ ) );
OR3_X1 _11446_ ( .A1(_03531_ ), .A2(\EX_LS_result_reg [18] ), .A3(_03533_ ), .ZN(_03828_ ) );
OR2_X1 _11447_ ( .A1(_03517_ ), .A2(\myreg.Reg[1][18] ), .ZN(_03829_ ) );
OAI211_X1 _11448_ ( .A(_03829_ ), .B(_03492_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[0][18] ), .ZN(_03830_ ) );
OR2_X1 _11449_ ( .A1(_03517_ ), .A2(\myreg.Reg[3][18] ), .ZN(_03831_ ) );
OAI211_X1 _11450_ ( .A(_03831_ ), .B(fanout_net_44 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[2][18] ), .ZN(_03832_ ) );
NAND3_X1 _11451_ ( .A1(_03830_ ), .A2(_03832_ ), .A3(_03502_ ), .ZN(_03833_ ) );
MUX2_X1 _11452_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_38 ), .Z(_03834_ ) );
MUX2_X1 _11453_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_38 ), .Z(_03835_ ) );
MUX2_X1 _11454_ ( .A(_03834_ ), .B(_03835_ ), .S(_03710_ ), .Z(_03836_ ) );
OAI211_X1 _11455_ ( .A(_03514_ ), .B(_03833_ ), .C1(_03836_ ), .C2(_03502_ ), .ZN(_03837_ ) );
OR2_X1 _11456_ ( .A1(_03517_ ), .A2(\myreg.Reg[15][18] ), .ZN(_03838_ ) );
OAI211_X1 _11457_ ( .A(_03838_ ), .B(fanout_net_44 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[14][18] ), .ZN(_03839_ ) );
OR2_X1 _11458_ ( .A1(_03517_ ), .A2(\myreg.Reg[13][18] ), .ZN(_03840_ ) );
OAI211_X1 _11459_ ( .A(_03840_ ), .B(_03710_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[12][18] ), .ZN(_03841_ ) );
NAND3_X1 _11460_ ( .A1(_03839_ ), .A2(_03841_ ), .A3(fanout_net_45 ), .ZN(_03842_ ) );
MUX2_X1 _11461_ ( .A(\myreg.Reg[8][18] ), .B(\myreg.Reg[9][18] ), .S(fanout_net_38 ), .Z(_03843_ ) );
MUX2_X1 _11462_ ( .A(\myreg.Reg[10][18] ), .B(\myreg.Reg[11][18] ), .S(fanout_net_38 ), .Z(_03844_ ) );
MUX2_X1 _11463_ ( .A(_03843_ ), .B(_03844_ ), .S(fanout_net_44 ), .Z(_03845_ ) );
OAI211_X1 _11464_ ( .A(fanout_net_46 ), .B(_03842_ ), .C1(_03845_ ), .C2(fanout_net_45 ), .ZN(_03846_ ) );
OAI211_X1 _11465_ ( .A(_03837_ ), .B(_03846_ ), .C1(_03531_ ), .C2(_03534_ ), .ZN(_03847_ ) );
NAND2_X2 _11466_ ( .A1(_03828_ ), .A2(_03847_ ), .ZN(_03848_ ) );
XOR2_X2 _11467_ ( .A(_02510_ ), .B(_03848_ ), .Z(_03849_ ) );
AND2_X1 _11468_ ( .A1(_03827_ ), .A2(_03849_ ), .ZN(_03850_ ) );
OR3_X2 _11469_ ( .A1(_03583_ ), .A2(\EX_LS_result_reg [16] ), .A3(_03584_ ), .ZN(_03851_ ) );
OR2_X1 _11470_ ( .A1(_03519_ ), .A2(\myreg.Reg[1][16] ), .ZN(_03852_ ) );
OAI211_X1 _11471_ ( .A(_03852_ ), .B(_03568_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[0][16] ), .ZN(_03853_ ) );
OR2_X1 _11472_ ( .A1(_03487_ ), .A2(\myreg.Reg[3][16] ), .ZN(_03854_ ) );
OAI211_X1 _11473_ ( .A(_03854_ ), .B(fanout_net_44 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[2][16] ), .ZN(_03855_ ) );
NAND3_X1 _11474_ ( .A1(_03853_ ), .A2(_03855_ ), .A3(_03510_ ), .ZN(_03856_ ) );
MUX2_X1 _11475_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_38 ), .Z(_03857_ ) );
MUX2_X1 _11476_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_38 ), .Z(_03858_ ) );
MUX2_X1 _11477_ ( .A(_03857_ ), .B(_03858_ ), .S(_03494_ ), .Z(_03859_ ) );
OAI211_X1 _11478_ ( .A(_03515_ ), .B(_03856_ ), .C1(_03859_ ), .C2(_03510_ ), .ZN(_03860_ ) );
OR2_X1 _11479_ ( .A1(_03487_ ), .A2(\myreg.Reg[15][16] ), .ZN(_03861_ ) );
OAI211_X1 _11480_ ( .A(_03861_ ), .B(fanout_net_44 ), .C1(fanout_net_38 ), .C2(\myreg.Reg[14][16] ), .ZN(_03862_ ) );
OR2_X1 _11481_ ( .A1(_03487_ ), .A2(\myreg.Reg[13][16] ), .ZN(_03863_ ) );
OAI211_X1 _11482_ ( .A(_03863_ ), .B(_03494_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[12][16] ), .ZN(_03864_ ) );
NAND3_X1 _11483_ ( .A1(_03862_ ), .A2(_03864_ ), .A3(fanout_net_45 ), .ZN(_03865_ ) );
MUX2_X1 _11484_ ( .A(\myreg.Reg[8][16] ), .B(\myreg.Reg[9][16] ), .S(fanout_net_39 ), .Z(_03866_ ) );
MUX2_X1 _11485_ ( .A(\myreg.Reg[10][16] ), .B(\myreg.Reg[11][16] ), .S(fanout_net_39 ), .Z(_03867_ ) );
MUX2_X1 _11486_ ( .A(_03866_ ), .B(_03867_ ), .S(fanout_net_44 ), .Z(_03868_ ) );
OAI211_X1 _11487_ ( .A(fanout_net_46 ), .B(_03865_ ), .C1(_03868_ ), .C2(fanout_net_45 ), .ZN(_03869_ ) );
OAI211_X1 _11488_ ( .A(_03860_ ), .B(_03869_ ), .C1(_03583_ ), .C2(_03584_ ), .ZN(_03870_ ) );
NAND2_X2 _11489_ ( .A1(_03851_ ), .A2(_03870_ ), .ZN(_03871_ ) );
XOR2_X2 _11490_ ( .A(_02580_ ), .B(_03871_ ), .Z(_03872_ ) );
INV_X1 _11491_ ( .A(_02557_ ), .ZN(_03873_ ) );
INV_X1 _11492_ ( .A(\EX_LS_result_reg [17] ), .ZN(_03874_ ) );
OR3_X2 _11493_ ( .A1(_03531_ ), .A2(_03874_ ), .A3(_03534_ ), .ZN(_03875_ ) );
OR2_X1 _11494_ ( .A1(_03486_ ), .A2(\myreg.Reg[1][17] ), .ZN(_03876_ ) );
OAI211_X1 _11495_ ( .A(_03876_ ), .B(_03492_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[0][17] ), .ZN(_03877_ ) );
OR2_X1 _11496_ ( .A1(_03517_ ), .A2(\myreg.Reg[3][17] ), .ZN(_03878_ ) );
OAI211_X1 _11497_ ( .A(_03878_ ), .B(fanout_net_44 ), .C1(fanout_net_39 ), .C2(\myreg.Reg[2][17] ), .ZN(_03879_ ) );
NAND3_X1 _11498_ ( .A1(_03877_ ), .A2(_03879_ ), .A3(_03502_ ), .ZN(_03880_ ) );
MUX2_X1 _11499_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_39 ), .Z(_03881_ ) );
MUX2_X1 _11500_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_39 ), .Z(_03882_ ) );
MUX2_X1 _11501_ ( .A(_03881_ ), .B(_03882_ ), .S(_03492_ ), .Z(_03883_ ) );
OAI211_X1 _11502_ ( .A(_03514_ ), .B(_03880_ ), .C1(_03883_ ), .C2(_03502_ ), .ZN(_03884_ ) );
OR2_X1 _11503_ ( .A1(_03517_ ), .A2(\myreg.Reg[15][17] ), .ZN(_03885_ ) );
OAI211_X1 _11504_ ( .A(_03885_ ), .B(fanout_net_44 ), .C1(fanout_net_39 ), .C2(\myreg.Reg[14][17] ), .ZN(_03886_ ) );
OR2_X1 _11505_ ( .A1(_03517_ ), .A2(\myreg.Reg[13][17] ), .ZN(_03887_ ) );
OAI211_X1 _11506_ ( .A(_03887_ ), .B(_03492_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[12][17] ), .ZN(_03888_ ) );
NAND3_X1 _11507_ ( .A1(_03886_ ), .A2(_03888_ ), .A3(fanout_net_45 ), .ZN(_03889_ ) );
MUX2_X1 _11508_ ( .A(\myreg.Reg[8][17] ), .B(\myreg.Reg[9][17] ), .S(fanout_net_39 ), .Z(_03890_ ) );
MUX2_X1 _11509_ ( .A(\myreg.Reg[10][17] ), .B(\myreg.Reg[11][17] ), .S(fanout_net_39 ), .Z(_03891_ ) );
MUX2_X1 _11510_ ( .A(_03890_ ), .B(_03891_ ), .S(fanout_net_44 ), .Z(_03892_ ) );
OAI211_X1 _11511_ ( .A(fanout_net_46 ), .B(_03889_ ), .C1(_03892_ ), .C2(fanout_net_45 ), .ZN(_03893_ ) );
NAND2_X1 _11512_ ( .A1(_03884_ ), .A2(_03893_ ), .ZN(_03894_ ) );
OAI21_X1 _11513_ ( .A(_03894_ ), .B1(_03531_ ), .B2(_03534_ ), .ZN(_03895_ ) );
AND2_X4 _11514_ ( .A1(_03875_ ), .A2(_03895_ ), .ZN(_03896_ ) );
XNOR2_X1 _11515_ ( .A(_03873_ ), .B(_03896_ ), .ZN(_03897_ ) );
AND3_X1 _11516_ ( .A1(_03850_ ), .A2(_03872_ ), .A3(_03897_ ), .ZN(_03898_ ) );
AND2_X2 _11517_ ( .A1(_03802_ ), .A2(_03898_ ), .ZN(_03899_ ) );
INV_X1 _11518_ ( .A(\EX_LS_result_reg [7] ), .ZN(_03900_ ) );
OR3_X1 _11519_ ( .A1(_03472_ ), .A2(_03900_ ), .A3(_03480_ ), .ZN(_03901_ ) );
CLKBUF_X2 _11520_ ( .A(_03483_ ), .Z(_03902_ ) );
OR2_X1 _11521_ ( .A1(_03902_ ), .A2(\myreg.Reg[1][7] ), .ZN(_03903_ ) );
OAI211_X1 _11522_ ( .A(_03903_ ), .B(_03708_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[0][7] ), .ZN(_03904_ ) );
OR2_X1 _11523_ ( .A1(_03902_ ), .A2(\myreg.Reg[3][7] ), .ZN(_03905_ ) );
OAI211_X1 _11524_ ( .A(_03905_ ), .B(fanout_net_44 ), .C1(fanout_net_39 ), .C2(\myreg.Reg[2][7] ), .ZN(_03906_ ) );
NAND3_X1 _11525_ ( .A1(_03904_ ), .A2(_03906_ ), .A3(_03498_ ), .ZN(_03907_ ) );
MUX2_X1 _11526_ ( .A(\myreg.Reg[6][7] ), .B(\myreg.Reg[7][7] ), .S(fanout_net_39 ), .Z(_03908_ ) );
MUX2_X1 _11527_ ( .A(\myreg.Reg[4][7] ), .B(\myreg.Reg[5][7] ), .S(fanout_net_39 ), .Z(_03909_ ) );
MUX2_X1 _11528_ ( .A(_03908_ ), .B(_03909_ ), .S(_03708_ ), .Z(_03910_ ) );
OAI211_X1 _11529_ ( .A(_03512_ ), .B(_03907_ ), .C1(_03910_ ), .C2(_03499_ ), .ZN(_03911_ ) );
OR2_X1 _11530_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[14][7] ), .ZN(_03912_ ) );
OAI211_X1 _11531_ ( .A(_03912_ ), .B(fanout_net_44 ), .C1(_03484_ ), .C2(\myreg.Reg[15][7] ), .ZN(_03913_ ) );
OR2_X1 _11532_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[12][7] ), .ZN(_03914_ ) );
OAI211_X1 _11533_ ( .A(_03914_ ), .B(_03708_ ), .C1(_03484_ ), .C2(\myreg.Reg[13][7] ), .ZN(_03915_ ) );
NAND3_X1 _11534_ ( .A1(_03913_ ), .A2(_03915_ ), .A3(fanout_net_45 ), .ZN(_03916_ ) );
MUX2_X1 _11535_ ( .A(\myreg.Reg[8][7] ), .B(\myreg.Reg[9][7] ), .S(fanout_net_39 ), .Z(_03917_ ) );
MUX2_X1 _11536_ ( .A(\myreg.Reg[10][7] ), .B(\myreg.Reg[11][7] ), .S(fanout_net_39 ), .Z(_03918_ ) );
MUX2_X1 _11537_ ( .A(_03917_ ), .B(_03918_ ), .S(fanout_net_44 ), .Z(_03919_ ) );
OAI211_X1 _11538_ ( .A(fanout_net_46 ), .B(_03916_ ), .C1(_03919_ ), .C2(fanout_net_45 ), .ZN(_03920_ ) );
NAND2_X1 _11539_ ( .A1(_03911_ ), .A2(_03920_ ), .ZN(_03921_ ) );
OAI21_X2 _11540_ ( .A(_03921_ ), .B1(_03473_ ), .B2(_03481_ ), .ZN(_03922_ ) );
AND2_X4 _11541_ ( .A1(_03901_ ), .A2(_03922_ ), .ZN(_03923_ ) );
XOR2_X1 _11542_ ( .A(_02706_ ), .B(_03923_ ), .Z(_03924_ ) );
OR3_X4 _11543_ ( .A1(_03530_ ), .A2(\EX_LS_result_reg [6] ), .A3(_03533_ ), .ZN(_03925_ ) );
OR2_X1 _11544_ ( .A1(_03706_ ), .A2(\myreg.Reg[9][6] ), .ZN(_03926_ ) );
OAI211_X1 _11545_ ( .A(_03926_ ), .B(_03710_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[8][6] ), .ZN(_03927_ ) );
OR2_X1 _11546_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[10][6] ), .ZN(_03928_ ) );
OAI211_X1 _11547_ ( .A(_03928_ ), .B(fanout_net_44 ), .C1(_03486_ ), .C2(\myreg.Reg[11][6] ), .ZN(_03929_ ) );
NAND3_X1 _11548_ ( .A1(_03927_ ), .A2(_03501_ ), .A3(_03929_ ), .ZN(_03930_ ) );
MUX2_X1 _11549_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(fanout_net_39 ), .Z(_03931_ ) );
MUX2_X1 _11550_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(fanout_net_39 ), .Z(_03932_ ) );
MUX2_X1 _11551_ ( .A(_03931_ ), .B(_03932_ ), .S(_03710_ ), .Z(_03933_ ) );
OAI211_X1 _11552_ ( .A(fanout_net_46 ), .B(_03930_ ), .C1(_03933_ ), .C2(_03502_ ), .ZN(_03934_ ) );
NOR2_X1 _11553_ ( .A1(_03486_ ), .A2(\myreg.Reg[3][6] ), .ZN(_03935_ ) );
OAI21_X1 _11554_ ( .A(fanout_net_44 ), .B1(fanout_net_39 ), .B2(\myreg.Reg[2][6] ), .ZN(_03936_ ) );
NOR2_X1 _11555_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[0][6] ), .ZN(_03937_ ) );
OAI21_X1 _11556_ ( .A(_03710_ ), .B1(_03486_ ), .B2(\myreg.Reg[1][6] ), .ZN(_03938_ ) );
OAI221_X1 _11557_ ( .A(_03501_ ), .B1(_03935_ ), .B2(_03936_ ), .C1(_03937_ ), .C2(_03938_ ), .ZN(_03939_ ) );
MUX2_X1 _11558_ ( .A(\myreg.Reg[6][6] ), .B(\myreg.Reg[7][6] ), .S(fanout_net_39 ), .Z(_03940_ ) );
MUX2_X1 _11559_ ( .A(\myreg.Reg[4][6] ), .B(\myreg.Reg[5][6] ), .S(fanout_net_39 ), .Z(_03941_ ) );
MUX2_X1 _11560_ ( .A(_03940_ ), .B(_03941_ ), .S(_03710_ ), .Z(_03942_ ) );
OAI211_X1 _11561_ ( .A(_03514_ ), .B(_03939_ ), .C1(_03942_ ), .C2(_03502_ ), .ZN(_03943_ ) );
OAI211_X1 _11562_ ( .A(_03934_ ), .B(_03943_ ), .C1(_03530_ ), .C2(_03534_ ), .ZN(_03944_ ) );
NAND2_X1 _11563_ ( .A1(_03925_ ), .A2(_03944_ ), .ZN(_03945_ ) );
NAND2_X1 _11564_ ( .A1(_03945_ ), .A2(_02729_ ), .ZN(_03946_ ) );
NAND4_X1 _11565_ ( .A1(_02709_ ), .A2(_03925_ ), .A3(_02728_ ), .A4(_03944_ ), .ZN(_03947_ ) );
AND3_X1 _11566_ ( .A1(_03924_ ), .A2(_03946_ ), .A3(_03947_ ), .ZN(_03948_ ) );
BUF_X4 _11567_ ( .A(_03472_ ), .Z(_03949_ ) );
CLKBUF_X2 _11568_ ( .A(_03480_ ), .Z(_03950_ ) );
OR3_X1 _11569_ ( .A1(_03949_ ), .A2(\EX_LS_result_reg [4] ), .A3(_03950_ ), .ZN(_03951_ ) );
OR2_X1 _11570_ ( .A1(_03516_ ), .A2(\myreg.Reg[7][4] ), .ZN(_03952_ ) );
OAI211_X1 _11571_ ( .A(_03952_ ), .B(fanout_net_44 ), .C1(fanout_net_39 ), .C2(\myreg.Reg[6][4] ), .ZN(_03953_ ) );
OR2_X1 _11572_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[4][4] ), .ZN(_03954_ ) );
OAI211_X1 _11573_ ( .A(_03954_ ), .B(_03491_ ), .C1(_03706_ ), .C2(\myreg.Reg[5][4] ), .ZN(_03955_ ) );
NAND3_X1 _11574_ ( .A1(_03953_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_03955_ ), .ZN(_03956_ ) );
MUX2_X1 _11575_ ( .A(\myreg.Reg[2][4] ), .B(\myreg.Reg[3][4] ), .S(fanout_net_39 ), .Z(_03957_ ) );
MUX2_X1 _11576_ ( .A(\myreg.Reg[0][4] ), .B(\myreg.Reg[1][4] ), .S(fanout_net_40 ), .Z(_03958_ ) );
BUF_X4 _11577_ ( .A(_03490_ ), .Z(_03959_ ) );
MUX2_X1 _11578_ ( .A(_03957_ ), .B(_03958_ ), .S(_03959_ ), .Z(_03960_ ) );
OAI211_X1 _11579_ ( .A(_03513_ ), .B(_03956_ ), .C1(_03960_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03961_ ) );
NOR2_X1 _11580_ ( .A1(_03706_ ), .A2(\myreg.Reg[11][4] ), .ZN(_03962_ ) );
OAI21_X1 _11581_ ( .A(fanout_net_44 ), .B1(fanout_net_40 ), .B2(\myreg.Reg[10][4] ), .ZN(_03963_ ) );
NOR2_X1 _11582_ ( .A1(fanout_net_40 ), .A2(\myreg.Reg[8][4] ), .ZN(_03964_ ) );
OAI21_X1 _11583_ ( .A(_03959_ ), .B1(_03706_ ), .B2(\myreg.Reg[9][4] ), .ZN(_03965_ ) );
OAI221_X1 _11584_ ( .A(_03500_ ), .B1(_03962_ ), .B2(_03963_ ), .C1(_03964_ ), .C2(_03965_ ), .ZN(_03966_ ) );
MUX2_X1 _11585_ ( .A(\myreg.Reg[12][4] ), .B(\myreg.Reg[13][4] ), .S(fanout_net_40 ), .Z(_03967_ ) );
MUX2_X1 _11586_ ( .A(\myreg.Reg[14][4] ), .B(\myreg.Reg[15][4] ), .S(fanout_net_40 ), .Z(_03968_ ) );
MUX2_X1 _11587_ ( .A(_03967_ ), .B(_03968_ ), .S(fanout_net_44 ), .Z(_03969_ ) );
OAI211_X1 _11588_ ( .A(fanout_net_46 ), .B(_03966_ ), .C1(_03969_ ), .C2(_03501_ ), .ZN(_03970_ ) );
OAI211_X1 _11589_ ( .A(_03961_ ), .B(_03970_ ), .C1(_03530_ ), .C2(_03533_ ), .ZN(_03971_ ) );
NAND2_X1 _11590_ ( .A1(_03951_ ), .A2(_03971_ ), .ZN(_03972_ ) );
XOR2_X1 _11591_ ( .A(_03972_ ), .B(_02676_ ), .Z(_03973_ ) );
BUF_X8 _11592_ ( .A(_03902_ ), .Z(_03974_ ) );
OR2_X1 _11593_ ( .A1(_03974_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03975_ ) );
OAI211_X1 _11594_ ( .A(_03975_ ), .B(fanout_net_44 ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03976_ ) );
BUF_X4 _11595_ ( .A(_03499_ ), .Z(_03977_ ) );
NAND2_X1 _11596_ ( .A1(_02641_ ), .A2(fanout_net_40 ), .ZN(_03978_ ) );
OAI211_X1 _11597_ ( .A(_03978_ ), .B(_03491_ ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03979_ ) );
NAND3_X1 _11598_ ( .A1(_03976_ ), .A2(_03977_ ), .A3(_03979_ ), .ZN(_03980_ ) );
MUX2_X1 _11599_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_03981_ ) );
MUX2_X1 _11600_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_03982_ ) );
MUX2_X1 _11601_ ( .A(_03981_ ), .B(_03982_ ), .S(_03959_ ), .Z(_03983_ ) );
OAI211_X1 _11602_ ( .A(fanout_net_46 ), .B(_03980_ ), .C1(_03983_ ), .C2(_03501_ ), .ZN(_03984_ ) );
MUX2_X1 _11603_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_03985_ ) );
AND2_X1 _11604_ ( .A1(_03985_ ), .A2(_03959_ ), .ZN(_03986_ ) );
MUX2_X1 _11605_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_03987_ ) );
AOI211_X1 _11606_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_03986_ ), .C1(fanout_net_44 ), .C2(_03987_ ), .ZN(_03988_ ) );
MUX2_X1 _11607_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_03989_ ) );
MUX2_X1 _11608_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_03990_ ) );
MUX2_X1 _11609_ ( .A(_03989_ ), .B(_03990_ ), .S(_03709_ ), .Z(_03991_ ) );
OAI21_X1 _11610_ ( .A(_03513_ ), .B1(_03991_ ), .B2(_03977_ ), .ZN(_03992_ ) );
OAI221_X2 _11611_ ( .A(_03984_ ), .B1(_03988_ ), .B2(_03992_ ), .C1(_03530_ ), .C2(_03533_ ), .ZN(_03993_ ) );
OR3_X1 _11612_ ( .A1(_03949_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_03950_ ), .ZN(_03994_ ) );
NAND2_X2 _11613_ ( .A1(_03993_ ), .A2(_03994_ ), .ZN(_03995_ ) );
XNOR2_X1 _11614_ ( .A(_02652_ ), .B(_03995_ ), .ZN(_03996_ ) );
AND2_X1 _11615_ ( .A1(_03973_ ), .A2(_03996_ ), .ZN(_03997_ ) );
AND2_X1 _11616_ ( .A1(_03948_ ), .A2(_03997_ ), .ZN(_03998_ ) );
NAND3_X1 _11617_ ( .A1(_03702_ ), .A2(_03899_ ), .A3(_03998_ ), .ZN(_03999_ ) );
OR2_X1 _11618_ ( .A1(_03484_ ), .A2(\myreg.Reg[9][2] ), .ZN(_04000_ ) );
OAI211_X1 _11619_ ( .A(_04000_ ), .B(_03490_ ), .C1(fanout_net_40 ), .C2(\myreg.Reg[8][2] ), .ZN(_04001_ ) );
OR2_X1 _11620_ ( .A1(_03484_ ), .A2(\myreg.Reg[11][2] ), .ZN(_04002_ ) );
OAI211_X1 _11621_ ( .A(_04002_ ), .B(fanout_net_44 ), .C1(fanout_net_40 ), .C2(\myreg.Reg[10][2] ), .ZN(_04003_ ) );
NAND3_X1 _11622_ ( .A1(_04001_ ), .A2(_04003_ ), .A3(_03499_ ), .ZN(_04004_ ) );
MUX2_X1 _11623_ ( .A(\myreg.Reg[14][2] ), .B(\myreg.Reg[15][2] ), .S(fanout_net_40 ), .Z(_04005_ ) );
MUX2_X1 _11624_ ( .A(\myreg.Reg[12][2] ), .B(\myreg.Reg[13][2] ), .S(fanout_net_40 ), .Z(_04006_ ) );
MUX2_X1 _11625_ ( .A(_04005_ ), .B(_04006_ ), .S(_03490_ ), .Z(_04007_ ) );
OAI211_X1 _11626_ ( .A(fanout_net_46 ), .B(_04004_ ), .C1(_04007_ ), .C2(_03500_ ), .ZN(_04008_ ) );
MUX2_X1 _11627_ ( .A(\myreg.Reg[0][2] ), .B(\myreg.Reg[1][2] ), .S(fanout_net_40 ), .Z(_04009_ ) );
AND2_X1 _11628_ ( .A1(_04009_ ), .A2(_03708_ ), .ZN(_04010_ ) );
MUX2_X1 _11629_ ( .A(\myreg.Reg[2][2] ), .B(\myreg.Reg[3][2] ), .S(fanout_net_40 ), .Z(_04011_ ) );
AOI211_X1 _11630_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_04010_ ), .C1(fanout_net_44 ), .C2(_04011_ ), .ZN(_04012_ ) );
MUX2_X1 _11631_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_40 ), .Z(_04013_ ) );
MUX2_X1 _11632_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_40 ), .Z(_04014_ ) );
MUX2_X1 _11633_ ( .A(_04013_ ), .B(_04014_ ), .S(_03708_ ), .Z(_04015_ ) );
OAI21_X1 _11634_ ( .A(_03512_ ), .B1(_04015_ ), .B2(_03499_ ), .ZN(_04016_ ) );
OAI221_X1 _11635_ ( .A(_04008_ ), .B1(_04012_ ), .B2(_04016_ ), .C1(_03473_ ), .C2(_03481_ ), .ZN(_04017_ ) );
OR3_X2 _11636_ ( .A1(_03473_ ), .A2(\EX_LS_result_reg [2] ), .A3(_03480_ ), .ZN(_04018_ ) );
NAND2_X2 _11637_ ( .A1(_04017_ ), .A2(_04018_ ), .ZN(_04019_ ) );
XOR2_X1 _11638_ ( .A(_04019_ ), .B(_02806_ ), .Z(_04020_ ) );
INV_X1 _11639_ ( .A(_04020_ ), .ZN(_04021_ ) );
NAND2_X2 _11640_ ( .A1(_03482_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04022_ ) );
OR2_X1 _11641_ ( .A1(_03902_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04023_ ) );
OAI211_X1 _11642_ ( .A(_04023_ ), .B(_03490_ ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04024_ ) );
OR2_X1 _11643_ ( .A1(_03902_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04025_ ) );
OAI211_X1 _11644_ ( .A(_04025_ ), .B(fanout_net_44 ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04026_ ) );
NAND3_X1 _11645_ ( .A1(_04024_ ), .A2(_04026_ ), .A3(_03499_ ), .ZN(_04027_ ) );
MUX2_X1 _11646_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04028_ ) );
MUX2_X1 _11647_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04029_ ) );
MUX2_X1 _11648_ ( .A(_04028_ ), .B(_04029_ ), .S(_03708_ ), .Z(_04030_ ) );
OAI211_X1 _11649_ ( .A(_03513_ ), .B(_04027_ ), .C1(_04030_ ), .C2(_03500_ ), .ZN(_04031_ ) );
OR2_X1 _11650_ ( .A1(_03902_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04032_ ) );
OAI211_X1 _11651_ ( .A(_04032_ ), .B(fanout_net_44 ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04033_ ) );
OR2_X1 _11652_ ( .A1(_03902_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04034_ ) );
OAI211_X1 _11653_ ( .A(_04034_ ), .B(_03490_ ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04035_ ) );
NAND3_X1 _11654_ ( .A1(_04033_ ), .A2(_04035_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04036_ ) );
MUX2_X1 _11655_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04037_ ) );
MUX2_X1 _11656_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04038_ ) );
MUX2_X1 _11657_ ( .A(_04037_ ), .B(_04038_ ), .S(fanout_net_44 ), .Z(_04039_ ) );
OAI211_X1 _11658_ ( .A(fanout_net_46 ), .B(_04036_ ), .C1(_04039_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04040_ ) );
NAND2_X1 _11659_ ( .A1(_04031_ ), .A2(_04040_ ), .ZN(_04041_ ) );
OAI21_X4 _11660_ ( .A(_04041_ ), .B1(_03949_ ), .B2(_03950_ ), .ZN(_04042_ ) );
AND2_X4 _11661_ ( .A1(_04022_ ), .A2(_04042_ ), .ZN(_04043_ ) );
XNOR2_X1 _11662_ ( .A(_04043_ ), .B(_02829_ ), .ZN(_04044_ ) );
INV_X1 _11663_ ( .A(_04044_ ), .ZN(_04045_ ) );
OR3_X2 _11664_ ( .A1(_03472_ ), .A2(\EX_LS_result_reg [1] ), .A3(_03480_ ), .ZN(_04046_ ) );
OR2_X1 _11665_ ( .A1(_03483_ ), .A2(\myreg.Reg[3][1] ), .ZN(_04047_ ) );
OAI211_X1 _11666_ ( .A(_04047_ ), .B(fanout_net_44 ), .C1(fanout_net_41 ), .C2(\myreg.Reg[2][1] ), .ZN(_04048_ ) );
OR2_X1 _11667_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[0][1] ), .ZN(_04049_ ) );
OAI211_X1 _11668_ ( .A(_04049_ ), .B(_03489_ ), .C1(_03483_ ), .C2(\myreg.Reg[1][1] ), .ZN(_04050_ ) );
NAND3_X1 _11669_ ( .A1(_04048_ ), .A2(_03498_ ), .A3(_04050_ ), .ZN(_04051_ ) );
MUX2_X1 _11670_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(fanout_net_41 ), .Z(_04052_ ) );
MUX2_X1 _11671_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(fanout_net_41 ), .Z(_04053_ ) );
MUX2_X1 _11672_ ( .A(_04052_ ), .B(_04053_ ), .S(_03489_ ), .Z(_04054_ ) );
OAI211_X1 _11673_ ( .A(_03512_ ), .B(_04051_ ), .C1(_04054_ ), .C2(_03498_ ), .ZN(_04055_ ) );
OR2_X1 _11674_ ( .A1(_03483_ ), .A2(\myreg.Reg[15][1] ), .ZN(_04056_ ) );
OAI211_X1 _11675_ ( .A(_04056_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myreg.Reg[14][1] ), .ZN(_04057_ ) );
OR2_X1 _11676_ ( .A1(_03483_ ), .A2(\myreg.Reg[13][1] ), .ZN(_04058_ ) );
OAI211_X1 _11677_ ( .A(_04058_ ), .B(_03489_ ), .C1(fanout_net_41 ), .C2(\myreg.Reg[12][1] ), .ZN(_04059_ ) );
NAND3_X1 _11678_ ( .A1(_04057_ ), .A2(_04059_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04060_ ) );
MUX2_X1 _11679_ ( .A(\myreg.Reg[8][1] ), .B(\myreg.Reg[9][1] ), .S(fanout_net_41 ), .Z(_04061_ ) );
MUX2_X1 _11680_ ( .A(\myreg.Reg[10][1] ), .B(\myreg.Reg[11][1] ), .S(fanout_net_41 ), .Z(_04062_ ) );
MUX2_X1 _11681_ ( .A(_04061_ ), .B(_04062_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04063_ ) );
OAI211_X1 _11682_ ( .A(fanout_net_46 ), .B(_04060_ ), .C1(_04063_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04064_ ) );
OAI211_X1 _11683_ ( .A(_04055_ ), .B(_04064_ ), .C1(_03472_ ), .C2(_03480_ ), .ZN(_04065_ ) );
NAND2_X1 _11684_ ( .A1(_04046_ ), .A2(_04065_ ), .ZN(_04066_ ) );
NAND2_X4 _11685_ ( .A1(_02760_ ), .A2(_04066_ ), .ZN(_04067_ ) );
NAND4_X1 _11686_ ( .A1(_02739_ ), .A2(_04046_ ), .A3(_02758_ ), .A4(_04065_ ), .ZN(_04068_ ) );
AND2_X2 _11687_ ( .A1(_04067_ ), .A2(_04068_ ), .ZN(_04069_ ) );
INV_X2 _11688_ ( .A(_04069_ ), .ZN(_04070_ ) );
NAND2_X4 _11689_ ( .A1(_02764_ ), .A2(_02783_ ), .ZN(_04071_ ) );
OR2_X1 _11690_ ( .A1(_03902_ ), .A2(\myreg.Reg[1][0] ), .ZN(_04072_ ) );
OAI211_X1 _11691_ ( .A(_04072_ ), .B(_03708_ ), .C1(fanout_net_41 ), .C2(\myreg.Reg[0][0] ), .ZN(_04073_ ) );
OR2_X1 _11692_ ( .A1(_03483_ ), .A2(\myreg.Reg[3][0] ), .ZN(_04074_ ) );
OAI211_X1 _11693_ ( .A(_04074_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myreg.Reg[2][0] ), .ZN(_04075_ ) );
NAND3_X1 _11694_ ( .A1(_04073_ ), .A2(_04075_ ), .A3(_03498_ ), .ZN(_04076_ ) );
MUX2_X1 _11695_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_41 ), .Z(_04077_ ) );
MUX2_X1 _11696_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_41 ), .Z(_04078_ ) );
MUX2_X1 _11697_ ( .A(_04077_ ), .B(_04078_ ), .S(_03489_ ), .Z(_04079_ ) );
OAI211_X1 _11698_ ( .A(_03512_ ), .B(_04076_ ), .C1(_04079_ ), .C2(_03499_ ), .ZN(_04080_ ) );
OR2_X1 _11699_ ( .A1(_03483_ ), .A2(\myreg.Reg[15][0] ), .ZN(_04081_ ) );
OAI211_X1 _11700_ ( .A(_04081_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myreg.Reg[14][0] ), .ZN(_04082_ ) );
OR2_X1 _11701_ ( .A1(_03483_ ), .A2(\myreg.Reg[13][0] ), .ZN(_04083_ ) );
OAI211_X1 _11702_ ( .A(_04083_ ), .B(_03489_ ), .C1(fanout_net_41 ), .C2(\myreg.Reg[12][0] ), .ZN(_04084_ ) );
NAND3_X1 _11703_ ( .A1(_04082_ ), .A2(_04084_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04085_ ) );
MUX2_X1 _11704_ ( .A(\myreg.Reg[8][0] ), .B(\myreg.Reg[9][0] ), .S(fanout_net_41 ), .Z(_04086_ ) );
MUX2_X1 _11705_ ( .A(\myreg.Reg[10][0] ), .B(\myreg.Reg[11][0] ), .S(fanout_net_41 ), .Z(_04087_ ) );
MUX2_X1 _11706_ ( .A(_04086_ ), .B(_04087_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04088_ ) );
OAI211_X1 _11707_ ( .A(fanout_net_46 ), .B(_04085_ ), .C1(_04088_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04089_ ) );
NAND2_X1 _11708_ ( .A1(_04080_ ), .A2(_04089_ ), .ZN(_04090_ ) );
OAI21_X1 _11709_ ( .A(_04090_ ), .B1(_03472_ ), .B2(_03481_ ), .ZN(_04091_ ) );
INV_X1 _11710_ ( .A(\EX_LS_result_reg [0] ), .ZN(_04092_ ) );
OR3_X2 _11711_ ( .A1(_03472_ ), .A2(_04092_ ), .A3(_03480_ ), .ZN(_04093_ ) );
AOI21_X4 _11712_ ( .A(_04071_ ), .B1(_04091_ ), .B2(_04093_ ), .ZN(_04094_ ) );
OR4_X1 _11713_ ( .A1(_04021_ ), .A2(_04045_ ), .A3(_04070_ ), .A4(_04094_ ), .ZN(_04095_ ) );
AND3_X1 _11714_ ( .A1(_04071_ ), .A2(_04091_ ), .A3(_04093_ ), .ZN(_04096_ ) );
NOR2_X1 _11715_ ( .A1(_04095_ ), .A2(_04096_ ), .ZN(_04097_ ) );
INV_X1 _11716_ ( .A(\EX_LS_result_reg [11] ), .ZN(_04098_ ) );
OR3_X4 _11717_ ( .A1(_03473_ ), .A2(_04098_ ), .A3(_03481_ ), .ZN(_04099_ ) );
OR2_X1 _11718_ ( .A1(_03902_ ), .A2(\myreg.Reg[1][11] ), .ZN(_04100_ ) );
OAI211_X1 _11719_ ( .A(_04100_ ), .B(_03490_ ), .C1(fanout_net_41 ), .C2(\myreg.Reg[0][11] ), .ZN(_04101_ ) );
OR2_X1 _11720_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[2][11] ), .ZN(_04102_ ) );
OAI211_X1 _11721_ ( .A(_04102_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03974_ ), .C2(\myreg.Reg[3][11] ), .ZN(_04103_ ) );
NAND3_X1 _11722_ ( .A1(_04101_ ), .A2(_03499_ ), .A3(_04103_ ), .ZN(_04104_ ) );
MUX2_X1 _11723_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_41 ), .Z(_04105_ ) );
MUX2_X1 _11724_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_41 ), .Z(_04106_ ) );
MUX2_X1 _11725_ ( .A(_04105_ ), .B(_04106_ ), .S(_03708_ ), .Z(_04107_ ) );
OAI211_X1 _11726_ ( .A(_03513_ ), .B(_04104_ ), .C1(_04107_ ), .C2(_03499_ ), .ZN(_04108_ ) );
OR2_X1 _11727_ ( .A1(_03902_ ), .A2(\myreg.Reg[15][11] ), .ZN(_04109_ ) );
OAI211_X1 _11728_ ( .A(_04109_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myreg.Reg[14][11] ), .ZN(_04110_ ) );
OR2_X1 _11729_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[12][11] ), .ZN(_04111_ ) );
OAI211_X1 _11730_ ( .A(_04111_ ), .B(_03708_ ), .C1(_03974_ ), .C2(\myreg.Reg[13][11] ), .ZN(_04112_ ) );
NAND3_X1 _11731_ ( .A1(_04110_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04112_ ), .ZN(_04113_ ) );
MUX2_X1 _11732_ ( .A(\myreg.Reg[8][11] ), .B(\myreg.Reg[9][11] ), .S(fanout_net_41 ), .Z(_04114_ ) );
MUX2_X1 _11733_ ( .A(\myreg.Reg[10][11] ), .B(\myreg.Reg[11][11] ), .S(fanout_net_41 ), .Z(_04115_ ) );
MUX2_X1 _11734_ ( .A(_04114_ ), .B(_04115_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04116_ ) );
OAI211_X1 _11735_ ( .A(fanout_net_46 ), .B(_04113_ ), .C1(_04116_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04117_ ) );
NAND2_X1 _11736_ ( .A1(_04108_ ), .A2(_04117_ ), .ZN(_04118_ ) );
OAI21_X4 _11737_ ( .A(_04118_ ), .B1(_03949_ ), .B2(_03950_ ), .ZN(_04119_ ) );
AND2_X4 _11738_ ( .A1(_04099_ ), .A2(_04119_ ), .ZN(_04120_ ) );
XNOR2_X1 _11739_ ( .A(_04120_ ), .B(_02936_ ), .ZN(_04121_ ) );
OR3_X2 _11740_ ( .A1(_03949_ ), .A2(\EX_LS_result_reg [10] ), .A3(_03950_ ), .ZN(_04122_ ) );
OR2_X1 _11741_ ( .A1(_03974_ ), .A2(\myreg.Reg[1][10] ), .ZN(_04123_ ) );
OAI211_X1 _11742_ ( .A(_04123_ ), .B(_03959_ ), .C1(fanout_net_41 ), .C2(\myreg.Reg[0][10] ), .ZN(_04124_ ) );
OR2_X1 _11743_ ( .A1(_03974_ ), .A2(\myreg.Reg[3][10] ), .ZN(_04125_ ) );
OAI211_X1 _11744_ ( .A(_04125_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_41 ), .C2(\myreg.Reg[2][10] ), .ZN(_04126_ ) );
NAND3_X1 _11745_ ( .A1(_04124_ ), .A2(_04126_ ), .A3(_03500_ ), .ZN(_04127_ ) );
MUX2_X1 _11746_ ( .A(\myreg.Reg[6][10] ), .B(\myreg.Reg[7][10] ), .S(fanout_net_41 ), .Z(_04128_ ) );
MUX2_X1 _11747_ ( .A(\myreg.Reg[4][10] ), .B(\myreg.Reg[5][10] ), .S(fanout_net_41 ), .Z(_04129_ ) );
MUX2_X1 _11748_ ( .A(_04128_ ), .B(_04129_ ), .S(_03709_ ), .Z(_04130_ ) );
OAI211_X1 _11749_ ( .A(_03513_ ), .B(_04127_ ), .C1(_04130_ ), .C2(_03977_ ), .ZN(_04131_ ) );
OR2_X1 _11750_ ( .A1(_03974_ ), .A2(\myreg.Reg[13][10] ), .ZN(_04132_ ) );
OAI211_X1 _11751_ ( .A(_04132_ ), .B(_03959_ ), .C1(fanout_net_41 ), .C2(\myreg.Reg[12][10] ), .ZN(_04133_ ) );
OR2_X1 _11752_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[14][10] ), .ZN(_04134_ ) );
OAI211_X1 _11753_ ( .A(_04134_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03706_ ), .C2(\myreg.Reg[15][10] ), .ZN(_04135_ ) );
NAND3_X1 _11754_ ( .A1(_04133_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04135_ ), .ZN(_04136_ ) );
MUX2_X1 _11755_ ( .A(\myreg.Reg[8][10] ), .B(\myreg.Reg[9][10] ), .S(fanout_net_42 ), .Z(_04137_ ) );
MUX2_X1 _11756_ ( .A(\myreg.Reg[10][10] ), .B(\myreg.Reg[11][10] ), .S(fanout_net_42 ), .Z(_04138_ ) );
MUX2_X1 _11757_ ( .A(_04137_ ), .B(_04138_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04139_ ) );
OAI211_X1 _11758_ ( .A(fanout_net_46 ), .B(_04136_ ), .C1(_04139_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04140_ ) );
OAI211_X1 _11759_ ( .A(_04131_ ), .B(_04140_ ), .C1(_03949_ ), .C2(_03533_ ), .ZN(_04141_ ) );
NAND2_X1 _11760_ ( .A1(_04122_ ), .A2(_04141_ ), .ZN(_04142_ ) );
AND2_X1 _11761_ ( .A1(_02912_ ), .A2(_04142_ ), .ZN(_04143_ ) );
AND4_X1 _11762_ ( .A1(_02911_ ), .A2(_02892_ ), .A3(_04122_ ), .A4(_04141_ ), .ZN(_04144_ ) );
NOR3_X1 _11763_ ( .A1(_04121_ ), .A2(_04143_ ), .A3(_04144_ ), .ZN(_04145_ ) );
OR3_X1 _11764_ ( .A1(_03949_ ), .A2(\EX_LS_result_reg [8] ), .A3(_03950_ ), .ZN(_04146_ ) );
OR2_X1 _11765_ ( .A1(_03516_ ), .A2(\myreg.Reg[9][8] ), .ZN(_04147_ ) );
OAI211_X1 _11766_ ( .A(_04147_ ), .B(_03491_ ), .C1(fanout_net_42 ), .C2(\myreg.Reg[8][8] ), .ZN(_04148_ ) );
OR2_X1 _11767_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[10][8] ), .ZN(_04149_ ) );
OAI211_X1 _11768_ ( .A(_04149_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03706_ ), .C2(\myreg.Reg[11][8] ), .ZN(_04150_ ) );
NAND3_X1 _11769_ ( .A1(_04148_ ), .A2(_03977_ ), .A3(_04150_ ), .ZN(_04151_ ) );
MUX2_X1 _11770_ ( .A(\myreg.Reg[14][8] ), .B(\myreg.Reg[15][8] ), .S(fanout_net_42 ), .Z(_04152_ ) );
MUX2_X1 _11771_ ( .A(\myreg.Reg[12][8] ), .B(\myreg.Reg[13][8] ), .S(fanout_net_42 ), .Z(_04153_ ) );
MUX2_X1 _11772_ ( .A(_04152_ ), .B(_04153_ ), .S(_03491_ ), .Z(_04154_ ) );
OAI211_X1 _11773_ ( .A(fanout_net_46 ), .B(_04151_ ), .C1(_04154_ ), .C2(_03501_ ), .ZN(_04155_ ) );
OR2_X1 _11774_ ( .A1(_03516_ ), .A2(\myreg.Reg[1][8] ), .ZN(_04156_ ) );
OAI211_X1 _11775_ ( .A(_04156_ ), .B(_03491_ ), .C1(fanout_net_42 ), .C2(\myreg.Reg[0][8] ), .ZN(_04157_ ) );
OR2_X1 _11776_ ( .A1(_03516_ ), .A2(\myreg.Reg[3][8] ), .ZN(_04158_ ) );
OAI211_X1 _11777_ ( .A(_04158_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myreg.Reg[2][8] ), .ZN(_04159_ ) );
NAND3_X1 _11778_ ( .A1(_04157_ ), .A2(_04159_ ), .A3(_03977_ ), .ZN(_04160_ ) );
MUX2_X1 _11779_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_42 ), .Z(_04161_ ) );
MUX2_X1 _11780_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_42 ), .Z(_04162_ ) );
MUX2_X1 _11781_ ( .A(_04161_ ), .B(_04162_ ), .S(_03959_ ), .Z(_04163_ ) );
OAI211_X1 _11782_ ( .A(_03514_ ), .B(_04160_ ), .C1(_04163_ ), .C2(_03501_ ), .ZN(_04164_ ) );
OAI211_X1 _11783_ ( .A(_04155_ ), .B(_04164_ ), .C1(_03530_ ), .C2(_03533_ ), .ZN(_04165_ ) );
NAND2_X1 _11784_ ( .A1(_04146_ ), .A2(_04165_ ), .ZN(_04166_ ) );
XOR2_X1 _11785_ ( .A(_02960_ ), .B(_04166_ ), .Z(_04167_ ) );
OR3_X2 _11786_ ( .A1(_03473_ ), .A2(\EX_LS_result_reg [9] ), .A3(_03481_ ), .ZN(_04168_ ) );
OR2_X1 _11787_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[4][9] ), .ZN(_04169_ ) );
OAI211_X1 _11788_ ( .A(_04169_ ), .B(_03490_ ), .C1(_03516_ ), .C2(\myreg.Reg[5][9] ), .ZN(_04170_ ) );
OR2_X1 _11789_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[6][9] ), .ZN(_04171_ ) );
OAI211_X1 _11790_ ( .A(_04171_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03974_ ), .C2(\myreg.Reg[7][9] ), .ZN(_04172_ ) );
NAND3_X1 _11791_ ( .A1(_04170_ ), .A2(_04172_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04173_ ) );
MUX2_X1 _11792_ ( .A(\myreg.Reg[2][9] ), .B(\myreg.Reg[3][9] ), .S(fanout_net_42 ), .Z(_04174_ ) );
MUX2_X1 _11793_ ( .A(\myreg.Reg[0][9] ), .B(\myreg.Reg[1][9] ), .S(fanout_net_42 ), .Z(_04175_ ) );
MUX2_X1 _11794_ ( .A(_04174_ ), .B(_04175_ ), .S(_03490_ ), .Z(_04176_ ) );
OAI211_X1 _11795_ ( .A(_03513_ ), .B(_04173_ ), .C1(_04176_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04177_ ) );
NOR2_X1 _11796_ ( .A1(_03974_ ), .A2(\myreg.Reg[11][9] ), .ZN(_04178_ ) );
OAI21_X1 _11797_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_42 ), .B2(\myreg.Reg[10][9] ), .ZN(_04179_ ) );
NOR2_X1 _11798_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[8][9] ), .ZN(_04180_ ) );
OAI21_X1 _11799_ ( .A(_03490_ ), .B1(_03974_ ), .B2(\myreg.Reg[9][9] ), .ZN(_04181_ ) );
OAI221_X1 _11800_ ( .A(_03499_ ), .B1(_04178_ ), .B2(_04179_ ), .C1(_04180_ ), .C2(_04181_ ), .ZN(_04182_ ) );
MUX2_X1 _11801_ ( .A(\myreg.Reg[12][9] ), .B(\myreg.Reg[13][9] ), .S(fanout_net_42 ), .Z(_04183_ ) );
MUX2_X1 _11802_ ( .A(\myreg.Reg[14][9] ), .B(\myreg.Reg[15][9] ), .S(fanout_net_42 ), .Z(_04184_ ) );
MUX2_X1 _11803_ ( .A(_04183_ ), .B(_04184_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04185_ ) );
OAI211_X1 _11804_ ( .A(fanout_net_46 ), .B(_04182_ ), .C1(_04185_ ), .C2(_03500_ ), .ZN(_04186_ ) );
OAI211_X1 _11805_ ( .A(_04177_ ), .B(_04186_ ), .C1(_03473_ ), .C2(_03481_ ), .ZN(_04187_ ) );
NAND2_X1 _11806_ ( .A1(_04168_ ), .A2(_04187_ ), .ZN(_04188_ ) );
AND2_X1 _11807_ ( .A1(_04188_ ), .A2(_02983_ ), .ZN(_04189_ ) );
NOR2_X1 _11808_ ( .A1(_04188_ ), .A2(_02983_ ), .ZN(_04190_ ) );
NOR2_X1 _11809_ ( .A1(_04189_ ), .A2(_04190_ ), .ZN(_04191_ ) );
AND3_X1 _11810_ ( .A1(_04145_ ), .A2(_04167_ ), .A3(_04191_ ), .ZN(_04192_ ) );
NAND2_X1 _11811_ ( .A1(_02866_ ), .A2(_02887_ ), .ZN(_04193_ ) );
BUF_X4 _11812_ ( .A(_04193_ ), .Z(_04194_ ) );
OR3_X4 _11813_ ( .A1(_03473_ ), .A2(\EX_LS_result_reg [13] ), .A3(_03481_ ), .ZN(_04195_ ) );
OR2_X1 _11814_ ( .A1(_03484_ ), .A2(\myreg.Reg[9][13] ), .ZN(_04196_ ) );
OAI211_X1 _11815_ ( .A(_04196_ ), .B(_03709_ ), .C1(fanout_net_42 ), .C2(\myreg.Reg[8][13] ), .ZN(_04197_ ) );
OR2_X1 _11816_ ( .A1(_03484_ ), .A2(\myreg.Reg[11][13] ), .ZN(_04198_ ) );
OAI211_X1 _11817_ ( .A(_04198_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myreg.Reg[10][13] ), .ZN(_04199_ ) );
NAND3_X1 _11818_ ( .A1(_04197_ ), .A2(_04199_ ), .A3(_03500_ ), .ZN(_04200_ ) );
MUX2_X1 _11819_ ( .A(\myreg.Reg[14][13] ), .B(\myreg.Reg[15][13] ), .S(fanout_net_42 ), .Z(_04201_ ) );
MUX2_X1 _11820_ ( .A(\myreg.Reg[12][13] ), .B(\myreg.Reg[13][13] ), .S(fanout_net_42 ), .Z(_04202_ ) );
MUX2_X1 _11821_ ( .A(_04201_ ), .B(_04202_ ), .S(_03709_ ), .Z(_04203_ ) );
OAI211_X1 _11822_ ( .A(fanout_net_46 ), .B(_04200_ ), .C1(_04203_ ), .C2(_03977_ ), .ZN(_04204_ ) );
NOR2_X1 _11823_ ( .A1(_03516_ ), .A2(\myreg.Reg[3][13] ), .ZN(_04205_ ) );
OAI21_X1 _11824_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_42 ), .B2(\myreg.Reg[2][13] ), .ZN(_04206_ ) );
NOR2_X1 _11825_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[0][13] ), .ZN(_04207_ ) );
OAI21_X1 _11826_ ( .A(_03709_ ), .B1(_03485_ ), .B2(\myreg.Reg[1][13] ), .ZN(_04208_ ) );
OAI221_X1 _11827_ ( .A(_03500_ ), .B1(_04205_ ), .B2(_04206_ ), .C1(_04207_ ), .C2(_04208_ ), .ZN(_04209_ ) );
MUX2_X1 _11828_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_42 ), .Z(_04210_ ) );
MUX2_X1 _11829_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_42 ), .Z(_04211_ ) );
MUX2_X1 _11830_ ( .A(_04210_ ), .B(_04211_ ), .S(_03709_ ), .Z(_04212_ ) );
OAI211_X1 _11831_ ( .A(_03513_ ), .B(_04209_ ), .C1(_04212_ ), .C2(_03977_ ), .ZN(_04213_ ) );
OAI211_X1 _11832_ ( .A(_04204_ ), .B(_04213_ ), .C1(_03949_ ), .C2(_03950_ ), .ZN(_04214_ ) );
NAND2_X1 _11833_ ( .A1(_04195_ ), .A2(_04214_ ), .ZN(_04215_ ) );
XOR2_X1 _11834_ ( .A(_04194_ ), .B(_04215_ ), .Z(_04216_ ) );
OR3_X1 _11835_ ( .A1(_03949_ ), .A2(\EX_LS_result_reg [12] ), .A3(_03950_ ), .ZN(_04217_ ) );
OR2_X1 _11836_ ( .A1(_03974_ ), .A2(\myreg.Reg[7][12] ), .ZN(_04218_ ) );
OAI211_X1 _11837_ ( .A(_04218_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_42 ), .C2(\myreg.Reg[6][12] ), .ZN(_04219_ ) );
OR2_X1 _11838_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[4][12] ), .ZN(_04220_ ) );
OAI211_X1 _11839_ ( .A(_04220_ ), .B(_03959_ ), .C1(_03706_ ), .C2(\myreg.Reg[5][12] ), .ZN(_04221_ ) );
NAND3_X1 _11840_ ( .A1(_04219_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04221_ ), .ZN(_04222_ ) );
MUX2_X1 _11841_ ( .A(\myreg.Reg[2][12] ), .B(\myreg.Reg[3][12] ), .S(fanout_net_42 ), .Z(_04223_ ) );
MUX2_X1 _11842_ ( .A(\myreg.Reg[0][12] ), .B(\myreg.Reg[1][12] ), .S(fanout_net_42 ), .Z(_04224_ ) );
MUX2_X1 _11843_ ( .A(_04223_ ), .B(_04224_ ), .S(_03959_ ), .Z(_04225_ ) );
OAI211_X1 _11844_ ( .A(_03513_ ), .B(_04222_ ), .C1(_04225_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04226_ ) );
NOR2_X1 _11845_ ( .A1(_03485_ ), .A2(\myreg.Reg[11][12] ), .ZN(_04227_ ) );
OAI21_X1 _11846_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myreg.Reg[10][12] ), .ZN(_04228_ ) );
NOR2_X1 _11847_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[8][12] ), .ZN(_04229_ ) );
OAI21_X1 _11848_ ( .A(_03709_ ), .B1(_03485_ ), .B2(\myreg.Reg[9][12] ), .ZN(_04230_ ) );
OAI221_X1 _11849_ ( .A(_03500_ ), .B1(_04227_ ), .B2(_04228_ ), .C1(_04229_ ), .C2(_04230_ ), .ZN(_04231_ ) );
MUX2_X1 _11850_ ( .A(\myreg.Reg[12][12] ), .B(\myreg.Reg[13][12] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04232_ ) );
MUX2_X1 _11851_ ( .A(\myreg.Reg[14][12] ), .B(\myreg.Reg[15][12] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04233_ ) );
MUX2_X1 _11852_ ( .A(_04232_ ), .B(_04233_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04234_ ) );
OAI211_X1 _11853_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04231_ ), .C1(_04234_ ), .C2(_03977_ ), .ZN(_04235_ ) );
OAI211_X4 _11854_ ( .A(_04226_ ), .B(_04235_ ), .C1(_03530_ ), .C2(_03533_ ), .ZN(_04236_ ) );
NAND2_X1 _11855_ ( .A1(_04217_ ), .A2(_04236_ ), .ZN(_04237_ ) );
XOR2_X1 _11856_ ( .A(_02863_ ), .B(_04237_ ), .Z(_04238_ ) );
AND2_X1 _11857_ ( .A1(_04216_ ), .A2(_04238_ ), .ZN(_04239_ ) );
OR3_X4 _11858_ ( .A1(_03473_ ), .A2(\EX_LS_result_reg [15] ), .A3(_03481_ ), .ZN(_04240_ ) );
OR2_X1 _11859_ ( .A1(_03484_ ), .A2(\myreg.Reg[5][15] ), .ZN(_04241_ ) );
OAI211_X1 _11860_ ( .A(_04241_ ), .B(_03959_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[4][15] ), .ZN(_04242_ ) );
OR2_X1 _11861_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[6][15] ), .ZN(_04243_ ) );
OAI211_X1 _11862_ ( .A(_04243_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03485_ ), .C2(\myreg.Reg[7][15] ), .ZN(_04244_ ) );
NAND3_X1 _11863_ ( .A1(_04242_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04244_ ), .ZN(_04245_ ) );
MUX2_X1 _11864_ ( .A(\myreg.Reg[2][15] ), .B(\myreg.Reg[3][15] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04246_ ) );
MUX2_X1 _11865_ ( .A(\myreg.Reg[0][15] ), .B(\myreg.Reg[1][15] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04247_ ) );
MUX2_X1 _11866_ ( .A(_04246_ ), .B(_04247_ ), .S(_03709_ ), .Z(_04248_ ) );
OAI211_X1 _11867_ ( .A(_03513_ ), .B(_04245_ ), .C1(_04248_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04249_ ) );
NOR2_X1 _11868_ ( .A1(_03485_ ), .A2(\myreg.Reg[11][15] ), .ZN(_04250_ ) );
OAI21_X1 _11869_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myreg.Reg[10][15] ), .ZN(_04251_ ) );
NOR2_X1 _11870_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[8][15] ), .ZN(_04252_ ) );
OAI21_X1 _11871_ ( .A(_03709_ ), .B1(_03485_ ), .B2(\myreg.Reg[9][15] ), .ZN(_04253_ ) );
OAI221_X1 _11872_ ( .A(_03500_ ), .B1(_04250_ ), .B2(_04251_ ), .C1(_04252_ ), .C2(_04253_ ), .ZN(_04254_ ) );
MUX2_X1 _11873_ ( .A(\myreg.Reg[12][15] ), .B(\myreg.Reg[13][15] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04255_ ) );
MUX2_X1 _11874_ ( .A(\myreg.Reg[14][15] ), .B(\myreg.Reg[15][15] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04256_ ) );
MUX2_X1 _11875_ ( .A(_04255_ ), .B(_04256_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04257_ ) );
OAI211_X1 _11876_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04254_ ), .C1(_04257_ ), .C2(_03977_ ), .ZN(_04258_ ) );
OAI211_X1 _11877_ ( .A(_04249_ ), .B(_04258_ ), .C1(_03949_ ), .C2(_03950_ ), .ZN(_04259_ ) );
NAND2_X1 _11878_ ( .A1(_04240_ ), .A2(_04259_ ), .ZN(_04260_ ) );
XOR2_X1 _11879_ ( .A(_02606_ ), .B(_04260_ ), .Z(_04261_ ) );
OR3_X4 _11880_ ( .A1(_03530_ ), .A2(\EX_LS_result_reg [14] ), .A3(_03950_ ), .ZN(_04262_ ) );
OR2_X1 _11881_ ( .A1(_03516_ ), .A2(\myreg.Reg[1][14] ), .ZN(_04263_ ) );
OAI211_X1 _11882_ ( .A(_04263_ ), .B(_03491_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[0][14] ), .ZN(_04264_ ) );
OR2_X1 _11883_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[2][14] ), .ZN(_04265_ ) );
OAI211_X1 _11884_ ( .A(_04265_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03706_ ), .C2(\myreg.Reg[3][14] ), .ZN(_04266_ ) );
NAND3_X1 _11885_ ( .A1(_04264_ ), .A2(_03977_ ), .A3(_04266_ ), .ZN(_04267_ ) );
MUX2_X1 _11886_ ( .A(\myreg.Reg[6][14] ), .B(\myreg.Reg[7][14] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04268_ ) );
MUX2_X1 _11887_ ( .A(\myreg.Reg[4][14] ), .B(\myreg.Reg[5][14] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04269_ ) );
MUX2_X1 _11888_ ( .A(_04268_ ), .B(_04269_ ), .S(_03491_ ), .Z(_04270_ ) );
OAI211_X1 _11889_ ( .A(_03514_ ), .B(_04267_ ), .C1(_04270_ ), .C2(_03501_ ), .ZN(_04271_ ) );
OR2_X1 _11890_ ( .A1(_03516_ ), .A2(\myreg.Reg[15][14] ), .ZN(_04272_ ) );
OAI211_X1 _11891_ ( .A(_04272_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[14][14] ), .ZN(_04273_ ) );
OR2_X1 _11892_ ( .A1(_03516_ ), .A2(\myreg.Reg[13][14] ), .ZN(_04274_ ) );
OAI211_X1 _11893_ ( .A(_04274_ ), .B(_03491_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[12][14] ), .ZN(_04275_ ) );
NAND3_X1 _11894_ ( .A1(_04273_ ), .A2(_04275_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04276_ ) );
MUX2_X1 _11895_ ( .A(\myreg.Reg[8][14] ), .B(\myreg.Reg[9][14] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04277_ ) );
MUX2_X1 _11896_ ( .A(\myreg.Reg[10][14] ), .B(\myreg.Reg[11][14] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04278_ ) );
MUX2_X1 _11897_ ( .A(_04277_ ), .B(_04278_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04279_ ) );
OAI211_X1 _11898_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04276_ ), .C1(_04279_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04280_ ) );
OAI211_X1 _11899_ ( .A(_04271_ ), .B(_04280_ ), .C1(_03530_ ), .C2(_03533_ ), .ZN(_04281_ ) );
NAND2_X1 _11900_ ( .A1(_04262_ ), .A2(_04281_ ), .ZN(_04282_ ) );
XOR2_X1 _11901_ ( .A(_02628_ ), .B(_04282_ ), .Z(_04283_ ) );
AND2_X1 _11902_ ( .A1(_04261_ ), .A2(_04283_ ), .ZN(_04284_ ) );
AND2_X1 _11903_ ( .A1(_04239_ ), .A2(_04284_ ), .ZN(_04285_ ) );
AND2_X1 _11904_ ( .A1(_04192_ ), .A2(_04285_ ), .ZN(_04286_ ) );
NAND2_X1 _11905_ ( .A1(_04097_ ), .A2(_04286_ ), .ZN(_04287_ ) );
NOR2_X1 _11906_ ( .A1(_03999_ ), .A2(_04287_ ), .ZN(_04288_ ) );
NOR2_X1 _11907_ ( .A1(_03250_ ), .A2(\ID_EX_typ [1] ), .ZN(_04289_ ) );
AND2_X1 _11908_ ( .A1(_04289_ ), .A2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .ZN(_04290_ ) );
INV_X1 _11909_ ( .A(_04290_ ), .ZN(_04291_ ) );
INV_X1 _11910_ ( .A(\ID_EX_typ [1] ), .ZN(_04292_ ) );
NOR2_X1 _11911_ ( .A1(_04292_ ), .A2(fanout_net_8 ), .ZN(_04293_ ) );
AND2_X2 _11912_ ( .A1(_04293_ ), .A2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .ZN(_04294_ ) );
INV_X1 _11913_ ( .A(_04294_ ), .ZN(_04295_ ) );
INV_X1 _11914_ ( .A(fanout_net_11 ), .ZN(_04296_ ) );
BUF_X4 _11915_ ( .A(_04296_ ), .Z(_04297_ ) );
BUF_X4 _11916_ ( .A(_04297_ ), .Z(_04298_ ) );
BUF_X2 _11917_ ( .A(_04298_ ), .Z(_04299_ ) );
NAND2_X1 _11918_ ( .A1(_03676_ ), .A2(_04299_ ), .ZN(_04300_ ) );
OR2_X1 _11919_ ( .A1(_04299_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04301_ ) );
AND3_X1 _11920_ ( .A1(_04300_ ), .A2(_03184_ ), .A3(_04301_ ), .ZN(_04302_ ) );
AOI21_X1 _11921_ ( .A(_03184_ ), .B1(_04300_ ), .B2(_04301_ ), .ZN(_04303_ ) );
NOR2_X1 _11922_ ( .A1(_04302_ ), .A2(_04303_ ), .ZN(_04304_ ) );
INV_X1 _11923_ ( .A(_04304_ ), .ZN(_04305_ ) );
NAND3_X1 _11924_ ( .A1(_03678_ ), .A2(_04299_ ), .A3(_03697_ ), .ZN(_04306_ ) );
NAND2_X1 _11925_ ( .A1(fanout_net_11 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04307_ ) );
AND2_X1 _11926_ ( .A1(_04306_ ), .A2(_04307_ ), .ZN(_04308_ ) );
XNOR2_X1 _11927_ ( .A(_04308_ ), .B(_02358_ ), .ZN(_04309_ ) );
NOR2_X1 _11928_ ( .A1(_04305_ ), .A2(_04309_ ), .ZN(_04310_ ) );
NAND3_X1 _11929_ ( .A1(_03633_ ), .A2(_04298_ ), .A3(_03652_ ), .ZN(_04311_ ) );
NAND2_X1 _11930_ ( .A1(fanout_net_11 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04312_ ) );
AND2_X2 _11931_ ( .A1(_04311_ ), .A2(_04312_ ), .ZN(_04313_ ) );
XNOR2_X1 _11932_ ( .A(_04313_ ), .B(_03156_ ), .ZN(_04314_ ) );
INV_X1 _11933_ ( .A(_04314_ ), .ZN(_04315_ ) );
NAND3_X1 _11934_ ( .A1(_03612_ ), .A2(_04299_ ), .A3(_03630_ ), .ZN(_04316_ ) );
NAND2_X1 _11935_ ( .A1(fanout_net_11 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_04317_ ) );
AND2_X2 _11936_ ( .A1(_04316_ ), .A2(_04317_ ), .ZN(_04318_ ) );
INV_X1 _11937_ ( .A(_02388_ ), .ZN(_04319_ ) );
XNOR2_X1 _11938_ ( .A(_04318_ ), .B(_04319_ ), .ZN(_04320_ ) );
INV_X1 _11939_ ( .A(_04320_ ), .ZN(_04321_ ) );
AND3_X1 _11940_ ( .A1(_04310_ ), .A2(_04315_ ), .A3(_04321_ ), .ZN(_04322_ ) );
NAND3_X1 _11941_ ( .A1(_04262_ ), .A2(_04281_ ), .A3(_04297_ ), .ZN(_04323_ ) );
NAND2_X1 _11942_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [14] ), .ZN(_04324_ ) );
AND2_X2 _11943_ ( .A1(_04323_ ), .A2(_04324_ ), .ZN(_04325_ ) );
XNOR2_X2 _11944_ ( .A(_04325_ ), .B(_02628_ ), .ZN(_04326_ ) );
NAND3_X1 _11945_ ( .A1(_04240_ ), .A2(_04296_ ), .A3(_04259_ ), .ZN(_04327_ ) );
NAND2_X1 _11946_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [15] ), .ZN(_04328_ ) );
AND2_X1 _11947_ ( .A1(_04327_ ), .A2(_04328_ ), .ZN(_04329_ ) );
INV_X2 _11948_ ( .A(_02605_ ), .ZN(_04330_ ) );
NOR2_X2 _11949_ ( .A1(_04329_ ), .A2(_04330_ ), .ZN(_04331_ ) );
AND3_X2 _11950_ ( .A1(_04330_ ), .A2(_04328_ ), .A3(_04327_ ), .ZN(_04332_ ) );
NOR2_X4 _11951_ ( .A1(_04331_ ), .A2(_04332_ ), .ZN(_04333_ ) );
OR2_X2 _11952_ ( .A1(_04326_ ), .A2(_04333_ ), .ZN(_04334_ ) );
NAND3_X1 _11953_ ( .A1(_04195_ ), .A2(_04296_ ), .A3(_04214_ ), .ZN(_04335_ ) );
NAND2_X1 _11954_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [13] ), .ZN(_04336_ ) );
AND2_X2 _11955_ ( .A1(_04335_ ), .A2(_04336_ ), .ZN(_04337_ ) );
XNOR2_X1 _11956_ ( .A(_04337_ ), .B(_04193_ ), .ZN(_04338_ ) );
NAND3_X1 _11957_ ( .A1(_04217_ ), .A2(_04236_ ), .A3(_04297_ ), .ZN(_04339_ ) );
NAND2_X1 _11958_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [12] ), .ZN(_04340_ ) );
NAND2_X1 _11959_ ( .A1(_04339_ ), .A2(_04340_ ), .ZN(_04341_ ) );
INV_X1 _11960_ ( .A(_02862_ ), .ZN(_04342_ ) );
XNOR2_X2 _11961_ ( .A(_04341_ ), .B(_04342_ ), .ZN(_04343_ ) );
NOR3_X4 _11962_ ( .A1(_04334_ ), .A2(_04338_ ), .A3(_04343_ ), .ZN(_04344_ ) );
OR2_X4 _11963_ ( .A1(_04120_ ), .A2(fanout_net_11 ), .ZN(_04345_ ) );
NAND2_X1 _11964_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [11] ), .ZN(_04346_ ) );
AND2_X1 _11965_ ( .A1(_04345_ ), .A2(_04346_ ), .ZN(_04347_ ) );
INV_X1 _11966_ ( .A(_02935_ ), .ZN(_04348_ ) );
NOR2_X2 _11967_ ( .A1(_04347_ ), .A2(_04348_ ), .ZN(_04349_ ) );
AND3_X2 _11968_ ( .A1(_04345_ ), .A2(_04348_ ), .A3(_04346_ ), .ZN(_04350_ ) );
NOR2_X4 _11969_ ( .A1(_04349_ ), .A2(_04350_ ), .ZN(_04351_ ) );
NAND3_X1 _11970_ ( .A1(_04122_ ), .A2(_04141_ ), .A3(_04297_ ), .ZN(_04352_ ) );
NAND2_X1 _11971_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [10] ), .ZN(_04353_ ) );
AND2_X1 _11972_ ( .A1(_04352_ ), .A2(_04353_ ), .ZN(_04354_ ) );
XNOR2_X2 _11973_ ( .A(_04354_ ), .B(_02912_ ), .ZN(_04355_ ) );
NOR2_X2 _11974_ ( .A1(_04351_ ), .A2(_04355_ ), .ZN(_04356_ ) );
AND2_X1 _11975_ ( .A1(_04344_ ), .A2(_04356_ ), .ZN(_04357_ ) );
NAND3_X1 _11976_ ( .A1(_04146_ ), .A2(_04297_ ), .A3(_04165_ ), .ZN(_04358_ ) );
NAND2_X1 _11977_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [8] ), .ZN(_04359_ ) );
AND2_X1 _11978_ ( .A1(_04358_ ), .A2(_04359_ ), .ZN(_04360_ ) );
XNOR2_X1 _11979_ ( .A(_04360_ ), .B(_02960_ ), .ZN(_04361_ ) );
INV_X1 _11980_ ( .A(_04361_ ), .ZN(_04362_ ) );
NAND3_X2 _11981_ ( .A1(_04168_ ), .A2(_04296_ ), .A3(_04187_ ), .ZN(_04363_ ) );
NAND2_X1 _11982_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [9] ), .ZN(_04364_ ) );
AND2_X2 _11983_ ( .A1(_04363_ ), .A2(_04364_ ), .ZN(_04365_ ) );
INV_X16 _11984_ ( .A(_02983_ ), .ZN(_04366_ ) );
NOR2_X2 _11985_ ( .A1(_04365_ ), .A2(_04366_ ), .ZN(_04367_ ) );
AND3_X4 _11986_ ( .A1(_04366_ ), .A2(_04364_ ), .A3(_04363_ ), .ZN(_04368_ ) );
OAI211_X1 _11987_ ( .A(_04357_ ), .B(_04362_ ), .C1(_04367_ ), .C2(_04368_ ), .ZN(_04369_ ) );
NAND3_X1 _11988_ ( .A1(_04017_ ), .A2(_04018_ ), .A3(_04297_ ), .ZN(_04370_ ) );
NAND2_X1 _11989_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [2] ), .ZN(_04371_ ) );
AND2_X2 _11990_ ( .A1(_04370_ ), .A2(_04371_ ), .ZN(_04372_ ) );
XNOR2_X1 _11991_ ( .A(_04372_ ), .B(_02806_ ), .ZN(_04373_ ) );
OR2_X4 _11992_ ( .A1(_04043_ ), .A2(fanout_net_11 ), .ZN(_04374_ ) );
NAND2_X1 _11993_ ( .A1(fanout_net_11 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_04375_ ) );
AND2_X4 _11994_ ( .A1(_04374_ ), .A2(_04375_ ), .ZN(_04376_ ) );
XNOR2_X2 _11995_ ( .A(_04376_ ), .B(_02833_ ), .ZN(_04377_ ) );
NAND2_X1 _11996_ ( .A1(_04066_ ), .A2(_04297_ ), .ZN(_04378_ ) );
NAND2_X1 _11997_ ( .A1(_02761_ ), .A2(fanout_net_11 ), .ZN(_04379_ ) );
NAND2_X1 _11998_ ( .A1(_04378_ ), .A2(_04379_ ), .ZN(_04380_ ) );
NAND2_X1 _11999_ ( .A1(_04380_ ), .A2(_02760_ ), .ZN(_04381_ ) );
AND3_X1 _12000_ ( .A1(_04378_ ), .A2(_02760_ ), .A3(_04379_ ), .ZN(_04382_ ) );
AOI21_X1 _12001_ ( .A(_02760_ ), .B1(_04378_ ), .B2(_04379_ ), .ZN(_04383_ ) );
NAND3_X2 _12002_ ( .A1(_04093_ ), .A2(_04296_ ), .A3(_04091_ ), .ZN(_04384_ ) );
NAND2_X1 _12003_ ( .A1(_02763_ ), .A2(fanout_net_11 ), .ZN(_04385_ ) );
NAND2_X4 _12004_ ( .A1(_04384_ ), .A2(_04385_ ), .ZN(_04386_ ) );
OAI22_X1 _12005_ ( .A1(_04382_ ), .A2(_04383_ ), .B1(_04071_ ), .B2(_04386_ ), .ZN(_04387_ ) );
AOI211_X2 _12006_ ( .A(_04373_ ), .B(_04377_ ), .C1(_04381_ ), .C2(_04387_ ), .ZN(_04388_ ) );
INV_X1 _12007_ ( .A(_02806_ ), .ZN(_04389_ ) );
INV_X1 _12008_ ( .A(_04372_ ), .ZN(_04390_ ) );
NOR3_X1 _12009_ ( .A1(_04377_ ), .A2(_04389_ ), .A3(_04390_ ), .ZN(_04391_ ) );
AOI21_X1 _12010_ ( .A(_02833_ ), .B1(_04374_ ), .B2(_04375_ ), .ZN(_04392_ ) );
OR3_X4 _12011_ ( .A1(_04388_ ), .A2(_04391_ ), .A3(_04392_ ), .ZN(_04393_ ) );
OR2_X2 _12012_ ( .A1(_03923_ ), .A2(fanout_net_11 ), .ZN(_04394_ ) );
NAND2_X1 _12013_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [7] ), .ZN(_04395_ ) );
AND2_X1 _12014_ ( .A1(_04394_ ), .A2(_04395_ ), .ZN(_04396_ ) );
NOR2_X2 _12015_ ( .A1(_04396_ ), .A2(_02734_ ), .ZN(_04397_ ) );
AND3_X4 _12016_ ( .A1(_04394_ ), .A2(_02734_ ), .A3(_04395_ ), .ZN(_04398_ ) );
NOR2_X4 _12017_ ( .A1(_04397_ ), .A2(_04398_ ), .ZN(_04399_ ) );
NAND3_X1 _12018_ ( .A1(_03925_ ), .A2(_04297_ ), .A3(_03944_ ), .ZN(_04400_ ) );
NAND2_X1 _12019_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [6] ), .ZN(_04401_ ) );
AND2_X2 _12020_ ( .A1(_04400_ ), .A2(_04401_ ), .ZN(_04402_ ) );
XNOR2_X1 _12021_ ( .A(_04402_ ), .B(_02729_ ), .ZN(_04403_ ) );
NOR2_X1 _12022_ ( .A1(_04399_ ), .A2(_04403_ ), .ZN(_04404_ ) );
NAND2_X1 _12023_ ( .A1(_03995_ ), .A2(_04297_ ), .ZN(_04405_ ) );
NAND2_X1 _12024_ ( .A1(_02681_ ), .A2(fanout_net_11 ), .ZN(_04406_ ) );
NAND2_X2 _12025_ ( .A1(_04405_ ), .A2(_04406_ ), .ZN(_04407_ ) );
INV_X1 _12026_ ( .A(_02652_ ), .ZN(_04408_ ) );
XNOR2_X1 _12027_ ( .A(_04407_ ), .B(_04408_ ), .ZN(_04409_ ) );
INV_X1 _12028_ ( .A(_04409_ ), .ZN(_04410_ ) );
NAND3_X1 _12029_ ( .A1(_03951_ ), .A2(_03971_ ), .A3(_04297_ ), .ZN(_04411_ ) );
NAND2_X1 _12030_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [4] ), .ZN(_04412_ ) );
AND2_X2 _12031_ ( .A1(_04411_ ), .A2(_04412_ ), .ZN(_04413_ ) );
XNOR2_X1 _12032_ ( .A(_04413_ ), .B(_02677_ ), .ZN(_04414_ ) );
INV_X1 _12033_ ( .A(_04414_ ), .ZN(_04415_ ) );
NAND4_X1 _12034_ ( .A1(_04393_ ), .A2(_04404_ ), .A3(_04410_ ), .A4(_04415_ ), .ZN(_04416_ ) );
INV_X1 _12035_ ( .A(_02729_ ), .ZN(_04417_ ) );
INV_X1 _12036_ ( .A(_04402_ ), .ZN(_04418_ ) );
NOR3_X1 _12037_ ( .A1(_04399_ ), .A2(_04417_ ), .A3(_04418_ ), .ZN(_04419_ ) );
AND2_X4 _12038_ ( .A1(_04407_ ), .A2(_02652_ ), .ZN(_04420_ ) );
AND3_X1 _12039_ ( .A1(_04405_ ), .A2(_04408_ ), .A3(_04406_ ), .ZN(_04421_ ) );
OAI211_X2 _12040_ ( .A(_02677_ ), .B(_04413_ ), .C1(_04420_ ), .C2(_04421_ ), .ZN(_04422_ ) );
OAI21_X1 _12041_ ( .A(_04422_ ), .B1(_04408_ ), .B2(_04407_ ), .ZN(_04423_ ) );
AOI221_X1 _12042_ ( .A(_04419_ ), .B1(_02706_ ), .B2(_04396_ ), .C1(_04404_ ), .C2(_04423_ ), .ZN(_04424_ ) );
AOI21_X1 _12043_ ( .A(_04369_ ), .B1(_04416_ ), .B2(_04424_ ), .ZN(_04425_ ) );
AND3_X1 _12044_ ( .A1(_04363_ ), .A2(_02983_ ), .A3(_04364_ ), .ZN(_04426_ ) );
NOR2_X4 _12045_ ( .A1(_04367_ ), .A2(_04368_ ), .ZN(_04427_ ) );
INV_X1 _12046_ ( .A(_02960_ ), .ZN(_04428_ ) );
INV_X1 _12047_ ( .A(_04360_ ), .ZN(_04429_ ) );
NOR3_X4 _12048_ ( .A1(_04427_ ), .A2(_04428_ ), .A3(_04429_ ), .ZN(_04430_ ) );
OAI21_X1 _12049_ ( .A(_04356_ ), .B1(_04426_ ), .B2(_04430_ ), .ZN(_04431_ ) );
INV_X1 _12050_ ( .A(_04347_ ), .ZN(_04432_ ) );
OAI21_X1 _12051_ ( .A(_04431_ ), .B1(_04348_ ), .B2(_04432_ ), .ZN(_04433_ ) );
INV_X1 _12052_ ( .A(_02912_ ), .ZN(_04434_ ) );
INV_X1 _12053_ ( .A(_04354_ ), .ZN(_04435_ ) );
NOR3_X1 _12054_ ( .A1(_04351_ ), .A2(_04434_ ), .A3(_04435_ ), .ZN(_04436_ ) );
OAI21_X2 _12055_ ( .A(_04344_ ), .B1(_04433_ ), .B2(_04436_ ), .ZN(_04437_ ) );
INV_X1 _12056_ ( .A(_04329_ ), .ZN(_04438_ ) );
NOR3_X1 _12057_ ( .A1(_04338_ ), .A2(_04342_ ), .A3(_04341_ ), .ZN(_04439_ ) );
AOI21_X1 _12058_ ( .A(_04439_ ), .B1(_04194_ ), .B2(_04337_ ), .ZN(_04440_ ) );
OAI221_X1 _12059_ ( .A(_04437_ ), .B1(_04330_ ), .B2(_04438_ ), .C1(_04334_ ), .C2(_04440_ ), .ZN(_04441_ ) );
INV_X1 _12060_ ( .A(_02629_ ), .ZN(_04442_ ) );
INV_X1 _12061_ ( .A(_04325_ ), .ZN(_04443_ ) );
NOR3_X1 _12062_ ( .A1(_04333_ ), .A2(_04442_ ), .A3(_04443_ ), .ZN(_04444_ ) );
OR3_X2 _12063_ ( .A1(_04425_ ), .A2(_04441_ ), .A3(_04444_ ), .ZN(_04445_ ) );
OR2_X1 _12064_ ( .A1(_03730_ ), .A2(fanout_net_11 ), .ZN(_04446_ ) );
NAND2_X1 _12065_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [23] ), .ZN(_04447_ ) );
AND2_X1 _12066_ ( .A1(_04446_ ), .A2(_04447_ ), .ZN(_04448_ ) );
NOR2_X1 _12067_ ( .A1(_04448_ ), .A2(_03703_ ), .ZN(_04449_ ) );
AND3_X4 _12068_ ( .A1(_04446_ ), .A2(_03703_ ), .A3(_04447_ ), .ZN(_04450_ ) );
NOR2_X2 _12069_ ( .A1(_04449_ ), .A2(_04450_ ), .ZN(_04451_ ) );
NAND3_X1 _12070_ ( .A1(_03732_ ), .A2(_04298_ ), .A3(_03751_ ), .ZN(_04452_ ) );
NAND2_X1 _12071_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [22] ), .ZN(_04453_ ) );
AND2_X2 _12072_ ( .A1(_04452_ ), .A2(_04453_ ), .ZN(_04454_ ) );
XNOR2_X1 _12073_ ( .A(_04454_ ), .B(_02411_ ), .ZN(_04455_ ) );
NOR2_X2 _12074_ ( .A1(_04451_ ), .A2(_04455_ ), .ZN(_04456_ ) );
OAI21_X1 _12075_ ( .A(_04298_ ), .B1(_03773_ ), .B2(_03775_ ), .ZN(_04457_ ) );
NAND2_X1 _12076_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [21] ), .ZN(_04458_ ) );
AND2_X2 _12077_ ( .A1(_04457_ ), .A2(_04458_ ), .ZN(_04459_ ) );
XNOR2_X1 _12078_ ( .A(_04459_ ), .B(_03777_ ), .ZN(_04460_ ) );
INV_X1 _12079_ ( .A(_04460_ ), .ZN(_04461_ ) );
NAND3_X1 _12080_ ( .A1(_03780_ ), .A2(_03799_ ), .A3(_04298_ ), .ZN(_04462_ ) );
NAND2_X1 _12081_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [20] ), .ZN(_04463_ ) );
AND2_X2 _12082_ ( .A1(_04462_ ), .A2(_04463_ ), .ZN(_04464_ ) );
XNOR2_X1 _12083_ ( .A(_04464_ ), .B(_02485_ ), .ZN(_04465_ ) );
INV_X1 _12084_ ( .A(_04465_ ), .ZN(_04466_ ) );
AND3_X2 _12085_ ( .A1(_04456_ ), .A2(_04461_ ), .A3(_04466_ ), .ZN(_04467_ ) );
INV_X1 _12086_ ( .A(_04467_ ), .ZN(_04468_ ) );
OR2_X1 _12087_ ( .A1(_03896_ ), .A2(fanout_net_11 ), .ZN(_04469_ ) );
NAND2_X1 _12088_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [17] ), .ZN(_04470_ ) );
AND2_X4 _12089_ ( .A1(_04469_ ), .A2(_04470_ ), .ZN(_04471_ ) );
XNOR2_X1 _12090_ ( .A(_04471_ ), .B(_02557_ ), .ZN(_04472_ ) );
NAND3_X1 _12091_ ( .A1(_03828_ ), .A2(_03847_ ), .A3(_04298_ ), .ZN(_04473_ ) );
NAND2_X1 _12092_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [18] ), .ZN(_04474_ ) );
AND2_X2 _12093_ ( .A1(_04473_ ), .A2(_04474_ ), .ZN(_04475_ ) );
XNOR2_X1 _12094_ ( .A(_04475_ ), .B(_02510_ ), .ZN(_04476_ ) );
INV_X1 _12095_ ( .A(_04476_ ), .ZN(_04477_ ) );
OR2_X4 _12096_ ( .A1(_03826_ ), .A2(\ID_EX_typ [4] ), .ZN(_04478_ ) );
NAND2_X1 _12097_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [19] ), .ZN(_04479_ ) );
AND2_X1 _12098_ ( .A1(_04478_ ), .A2(_04479_ ), .ZN(_04480_ ) );
NOR2_X1 _12099_ ( .A1(_04480_ ), .A2(_03803_ ), .ZN(_04481_ ) );
AND3_X1 _12100_ ( .A1(_04478_ ), .A2(_03803_ ), .A3(_04479_ ), .ZN(_04482_ ) );
OAI21_X2 _12101_ ( .A(_04477_ ), .B1(_04481_ ), .B2(_04482_ ), .ZN(_04483_ ) );
NAND3_X1 _12102_ ( .A1(_03851_ ), .A2(_03870_ ), .A3(_04298_ ), .ZN(_04484_ ) );
NAND2_X1 _12103_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [16] ), .ZN(_04485_ ) );
AND2_X2 _12104_ ( .A1(_04484_ ), .A2(_04485_ ), .ZN(_04486_ ) );
XNOR2_X1 _12105_ ( .A(_04486_ ), .B(_02580_ ), .ZN(_04487_ ) );
NOR4_X4 _12106_ ( .A1(_04468_ ), .A2(_04472_ ), .A3(_04483_ ), .A4(_04487_ ), .ZN(_04488_ ) );
AND2_X4 _12107_ ( .A1(_04445_ ), .A2(_04488_ ), .ZN(_04489_ ) );
AND2_X4 _12108_ ( .A1(_04471_ ), .A2(_03873_ ), .ZN(_04490_ ) );
NOR2_X1 _12109_ ( .A1(_04471_ ), .A2(_03873_ ), .ZN(_04491_ ) );
OAI211_X1 _12110_ ( .A(_02580_ ), .B(_04486_ ), .C1(_04490_ ), .C2(_04491_ ), .ZN(_04492_ ) );
OAI211_X1 _12111_ ( .A(_02557_ ), .B(_04470_ ), .C1(_03896_ ), .C2(\ID_EX_typ [4] ), .ZN(_04493_ ) );
AOI21_X1 _12112_ ( .A(_04483_ ), .B1(_04492_ ), .B2(_04493_ ), .ZN(_04494_ ) );
AOI21_X2 _12113_ ( .A(_04494_ ), .B1(_02533_ ), .B2(_04480_ ), .ZN(_04495_ ) );
NOR2_X1 _12114_ ( .A1(_04481_ ), .A2(_04482_ ), .ZN(_04496_ ) );
INV_X1 _12115_ ( .A(_04496_ ), .ZN(_04497_ ) );
NAND3_X1 _12116_ ( .A1(_04497_ ), .A2(_02510_ ), .A3(_04475_ ), .ZN(_04498_ ) );
AOI21_X1 _12117_ ( .A(_04468_ ), .B1(_04495_ ), .B2(_04498_ ), .ZN(_04499_ ) );
INV_X1 _12118_ ( .A(_02411_ ), .ZN(_04500_ ) );
INV_X1 _12119_ ( .A(_04454_ ), .ZN(_04501_ ) );
NOR3_X1 _12120_ ( .A1(_04451_ ), .A2(_04500_ ), .A3(_04501_ ), .ZN(_04502_ ) );
AND3_X1 _12121_ ( .A1(_04461_ ), .A2(_02485_ ), .A3(_04464_ ), .ZN(_04503_ ) );
AND3_X1 _12122_ ( .A1(_04457_ ), .A2(_03777_ ), .A3(_04458_ ), .ZN(_04504_ ) );
OAI21_X1 _12123_ ( .A(_04456_ ), .B1(_04503_ ), .B2(_04504_ ), .ZN(_04505_ ) );
NAND3_X1 _12124_ ( .A1(_04446_ ), .A2(_02438_ ), .A3(_04447_ ), .ZN(_04506_ ) );
NAND2_X1 _12125_ ( .A1(_04505_ ), .A2(_04506_ ), .ZN(_04507_ ) );
NOR4_X4 _12126_ ( .A1(_04489_ ), .A2(_04499_ ), .A3(_04502_ ), .A4(_04507_ ), .ZN(_04508_ ) );
OAI21_X1 _12127_ ( .A(_04298_ ), .B1(_03529_ ), .B2(_03536_ ), .ZN(_04509_ ) );
NAND2_X1 _12128_ ( .A1(_03121_ ), .A2(\ID_EX_typ [4] ), .ZN(_04510_ ) );
NAND2_X1 _12129_ ( .A1(_04509_ ), .A2(_04510_ ), .ZN(_04511_ ) );
NOR2_X1 _12130_ ( .A1(_04511_ ), .A2(_03126_ ), .ZN(_04512_ ) );
AOI21_X1 _12131_ ( .A(_03120_ ), .B1(_04509_ ), .B2(_04510_ ), .ZN(_04513_ ) );
NOR2_X1 _12132_ ( .A1(_04512_ ), .A2(_04513_ ), .ZN(_04514_ ) );
NAND3_X1 _12133_ ( .A1(_03556_ ), .A2(_03558_ ), .A3(_04298_ ), .ZN(_04515_ ) );
NAND2_X1 _12134_ ( .A1(_03077_ ), .A2(\ID_EX_typ [4] ), .ZN(_04516_ ) );
NAND2_X1 _12135_ ( .A1(_04515_ ), .A2(_04516_ ), .ZN(_04517_ ) );
INV_X1 _12136_ ( .A(_03560_ ), .ZN(_04518_ ) );
NOR2_X1 _12137_ ( .A1(_04517_ ), .A2(_04518_ ), .ZN(_04519_ ) );
AOI21_X1 _12138_ ( .A(_03560_ ), .B1(_04515_ ), .B2(_04516_ ), .ZN(_04520_ ) );
NOR2_X1 _12139_ ( .A1(_04519_ ), .A2(_04520_ ), .ZN(_04521_ ) );
NOR2_X1 _12140_ ( .A1(_04514_ ), .A2(_04521_ ), .ZN(_04522_ ) );
INV_X1 _12141_ ( .A(_04522_ ), .ZN(_04523_ ) );
NAND3_X1 _12142_ ( .A1(_03589_ ), .A2(_04298_ ), .A3(_03608_ ), .ZN(_04524_ ) );
NAND2_X1 _12143_ ( .A1(_03123_ ), .A2(\ID_EX_typ [4] ), .ZN(_04525_ ) );
NAND2_X1 _12144_ ( .A1(_04524_ ), .A2(_04525_ ), .ZN(_04526_ ) );
XNOR2_X1 _12145_ ( .A(_04526_ ), .B(_03073_ ), .ZN(_04527_ ) );
NAND3_X1 _12146_ ( .A1(_03563_ ), .A2(_04299_ ), .A3(_03585_ ), .ZN(_04528_ ) );
NAND2_X1 _12147_ ( .A1(_03048_ ), .A2(\ID_EX_typ [4] ), .ZN(_04529_ ) );
NAND2_X1 _12148_ ( .A1(_04528_ ), .A2(_04529_ ), .ZN(_04530_ ) );
INV_X1 _12149_ ( .A(_03047_ ), .ZN(_04531_ ) );
NOR2_X1 _12150_ ( .A1(_04530_ ), .A2(_04531_ ), .ZN(_04532_ ) );
AOI21_X1 _12151_ ( .A(_03047_ ), .B1(_04528_ ), .B2(_04529_ ), .ZN(_04533_ ) );
NOR2_X1 _12152_ ( .A1(_04532_ ), .A2(_04533_ ), .ZN(_04534_ ) );
NOR4_X4 _12153_ ( .A1(_04508_ ), .A2(_04523_ ), .A3(_04527_ ), .A4(_04534_ ), .ZN(_04535_ ) );
NAND2_X1 _12154_ ( .A1(_04526_ ), .A2(_03073_ ), .ZN(_04536_ ) );
INV_X1 _12155_ ( .A(_03073_ ), .ZN(_04537_ ) );
AND2_X1 _12156_ ( .A1(_04526_ ), .A2(_04537_ ), .ZN(_04538_ ) );
NOR2_X1 _12157_ ( .A1(_04526_ ), .A2(_04537_ ), .ZN(_04539_ ) );
OAI211_X1 _12158_ ( .A(_03047_ ), .B(_04530_ ), .C1(_04538_ ), .C2(_04539_ ), .ZN(_04540_ ) );
AOI21_X1 _12159_ ( .A(_04523_ ), .B1(_04536_ ), .B2(_04540_ ), .ZN(_04541_ ) );
INV_X1 _12160_ ( .A(_04521_ ), .ZN(_04542_ ) );
AND3_X1 _12161_ ( .A1(_04542_ ), .A2(_03120_ ), .A3(_04511_ ), .ZN(_04543_ ) );
AOI21_X1 _12162_ ( .A(_04518_ ), .B1(_04515_ ), .B2(_04516_ ), .ZN(_04544_ ) );
OR3_X1 _12163_ ( .A1(_04541_ ), .A2(_04543_ ), .A3(_04544_ ), .ZN(_04545_ ) );
OAI21_X4 _12164_ ( .A(_04322_ ), .B1(_04535_ ), .B2(_04545_ ), .ZN(_04546_ ) );
AOI21_X1 _12165_ ( .A(_02358_ ), .B1(_04307_ ), .B2(_04306_ ), .ZN(_04547_ ) );
AND2_X1 _12166_ ( .A1(_04304_ ), .A2(_04547_ ), .ZN(_04548_ ) );
OR2_X1 _12167_ ( .A1(_04318_ ), .A2(_04319_ ), .ZN(_04549_ ) );
OR2_X1 _12168_ ( .A1(_04314_ ), .A2(_04549_ ), .ZN(_04550_ ) );
OAI21_X1 _12169_ ( .A(_04550_ ), .B1(_03156_ ), .B2(_04313_ ), .ZN(_04551_ ) );
AOI211_X1 _12170_ ( .A(_04303_ ), .B(_04548_ ), .C1(_04551_ ), .C2(_04310_ ), .ZN(_04552_ ) );
AOI21_X2 _12171_ ( .A(_04295_ ), .B1(_04546_ ), .B2(_04552_ ), .ZN(_04553_ ) );
NAND3_X1 _12172_ ( .A1(_03996_ ), .A2(_02677_ ), .A3(_03972_ ), .ZN(_04554_ ) );
OAI21_X1 _12173_ ( .A(_04554_ ), .B1(_04408_ ), .B2(_03995_ ), .ZN(_04555_ ) );
AND2_X1 _12174_ ( .A1(_04019_ ), .A2(_02806_ ), .ZN(_04556_ ) );
INV_X1 _12175_ ( .A(_04556_ ), .ZN(_04557_ ) );
OR2_X4 _12176_ ( .A1(_04070_ ), .A2(_04094_ ), .ZN(_04558_ ) );
AND2_X4 _12177_ ( .A1(_04558_ ), .A2(_04067_ ), .ZN(_04559_ ) );
OAI221_X2 _12178_ ( .A(_04557_ ), .B1(_02833_ ), .B2(_04043_ ), .C1(_04559_ ), .C2(_04021_ ), .ZN(_04560_ ) );
NAND2_X1 _12179_ ( .A1(_02833_ ), .A2(_04043_ ), .ZN(_04561_ ) );
AND2_X2 _12180_ ( .A1(_04560_ ), .A2(_04561_ ), .ZN(_04562_ ) );
AOI21_X2 _12181_ ( .A(_04555_ ), .B1(_04562_ ), .B2(_03997_ ), .ZN(_04563_ ) );
XNOR2_X1 _12182_ ( .A(_02729_ ), .B(_03945_ ), .ZN(_04564_ ) );
OR2_X4 _12183_ ( .A1(_04563_ ), .A2(_04564_ ), .ZN(_04565_ ) );
AND2_X4 _12184_ ( .A1(_04565_ ), .A2(_03946_ ), .ZN(_04566_ ) );
INV_X4 _12185_ ( .A(_04566_ ), .ZN(_04567_ ) );
OAI21_X4 _12186_ ( .A(_04567_ ), .B1(_02706_ ), .B2(_03923_ ), .ZN(_04568_ ) );
NAND2_X1 _12187_ ( .A1(_02706_ ), .A2(_03923_ ), .ZN(_04569_ ) );
AND2_X4 _12188_ ( .A1(_04568_ ), .A2(_04569_ ), .ZN(_04570_ ) );
INV_X8 _12189_ ( .A(_04570_ ), .ZN(_04571_ ) );
NAND2_X4 _12190_ ( .A1(_04571_ ), .A2(_04286_ ), .ZN(_04572_ ) );
AND3_X1 _12191_ ( .A1(_04261_ ), .A2(_02629_ ), .A3(_04282_ ), .ZN(_04573_ ) );
AND2_X1 _12192_ ( .A1(_02863_ ), .A2(_04237_ ), .ZN(_04574_ ) );
AND2_X1 _12193_ ( .A1(_04216_ ), .A2(_04574_ ), .ZN(_04575_ ) );
AOI21_X1 _12194_ ( .A(_04575_ ), .B1(_04194_ ), .B2(_04215_ ), .ZN(_04576_ ) );
INV_X1 _12195_ ( .A(_04576_ ), .ZN(_04577_ ) );
AOI221_X4 _12196_ ( .A(_04573_ ), .B1(_02606_ ), .B2(_04260_ ), .C1(_04577_ ), .C2(_04284_ ), .ZN(_04578_ ) );
NAND2_X1 _12197_ ( .A1(_02960_ ), .A2(_04166_ ), .ZN(_04579_ ) );
NOR3_X1 _12198_ ( .A1(_04189_ ), .A2(_04190_ ), .A3(_04579_ ), .ZN(_04580_ ) );
OAI21_X1 _12199_ ( .A(_04145_ ), .B1(_04189_ ), .B2(_04580_ ), .ZN(_04581_ ) );
NAND3_X1 _12200_ ( .A1(_02936_ ), .A2(_04119_ ), .A3(_04099_ ), .ZN(_04582_ ) );
INV_X1 _12201_ ( .A(_04143_ ), .ZN(_04583_ ) );
OR2_X1 _12202_ ( .A1(_04121_ ), .A2(_04583_ ), .ZN(_04584_ ) );
AND3_X1 _12203_ ( .A1(_04581_ ), .A2(_04582_ ), .A3(_04584_ ), .ZN(_04585_ ) );
INV_X1 _12204_ ( .A(_04285_ ), .ZN(_04586_ ) );
OR2_X1 _12205_ ( .A1(_04585_ ), .A2(_04586_ ), .ZN(_04587_ ) );
AND2_X1 _12206_ ( .A1(_04578_ ), .A2(_04587_ ), .ZN(_04588_ ) );
AND2_X4 _12207_ ( .A1(_04572_ ), .A2(_04588_ ), .ZN(_04589_ ) );
AND2_X1 _12208_ ( .A1(_03702_ ), .A2(_03899_ ), .ZN(_04590_ ) );
INV_X1 _12209_ ( .A(_04590_ ), .ZN(_04591_ ) );
OR2_X4 _12210_ ( .A1(_04589_ ), .A2(_04591_ ), .ZN(_04592_ ) );
NOR2_X1 _12211_ ( .A1(_03896_ ), .A2(_02557_ ), .ZN(_04593_ ) );
INV_X1 _12212_ ( .A(_03850_ ), .ZN(_04594_ ) );
NAND2_X1 _12213_ ( .A1(_02580_ ), .A2(_03871_ ), .ZN(_04595_ ) );
AND2_X1 _12214_ ( .A1(_03896_ ), .A2(_02557_ ), .ZN(_04596_ ) );
INV_X1 _12215_ ( .A(_04596_ ), .ZN(_04597_ ) );
AOI211_X2 _12216_ ( .A(_04593_ ), .B(_04594_ ), .C1(_04595_ ), .C2(_04597_ ), .ZN(_04598_ ) );
AND3_X1 _12217_ ( .A1(_02533_ ), .A2(_03825_ ), .A3(_03805_ ), .ZN(_04599_ ) );
AND3_X1 _12218_ ( .A1(_03827_ ), .A2(_02510_ ), .A3(_03848_ ), .ZN(_04600_ ) );
NOR3_X2 _12219_ ( .A1(_04598_ ), .A2(_04599_ ), .A3(_04600_ ), .ZN(_04601_ ) );
INV_X1 _12220_ ( .A(_03802_ ), .ZN(_04602_ ) );
NOR2_X1 _12221_ ( .A1(_04601_ ), .A2(_04602_ ), .ZN(_04603_ ) );
INV_X1 _12222_ ( .A(_04603_ ), .ZN(_04604_ ) );
AND2_X1 _12223_ ( .A1(_03776_ ), .A2(_03777_ ), .ZN(_04605_ ) );
NOR2_X1 _12224_ ( .A1(_03776_ ), .A2(_03777_ ), .ZN(_04606_ ) );
NAND2_X1 _12225_ ( .A1(_02485_ ), .A2(_03800_ ), .ZN(_04607_ ) );
NOR3_X1 _12226_ ( .A1(_04605_ ), .A2(_04606_ ), .A3(_04607_ ), .ZN(_04608_ ) );
OR2_X1 _12227_ ( .A1(_04608_ ), .A2(_04605_ ), .ZN(_04609_ ) );
AND2_X1 _12228_ ( .A1(_03754_ ), .A2(_04609_ ), .ZN(_04610_ ) );
INV_X1 _12229_ ( .A(_04610_ ), .ZN(_04611_ ) );
AND2_X1 _12230_ ( .A1(_02411_ ), .A2(_03752_ ), .ZN(_04612_ ) );
AND2_X1 _12231_ ( .A1(_03731_ ), .A2(_04612_ ), .ZN(_04613_ ) );
AOI21_X1 _12232_ ( .A(_04613_ ), .B1(_02438_ ), .B2(_03730_ ), .ZN(_04614_ ) );
AND3_X2 _12233_ ( .A1(_04604_ ), .A2(_04611_ ), .A3(_04614_ ), .ZN(_04615_ ) );
INV_X1 _12234_ ( .A(_03702_ ), .ZN(_04616_ ) );
NOR2_X2 _12235_ ( .A1(_04615_ ), .A2(_04616_ ), .ZN(_04617_ ) );
INV_X1 _12236_ ( .A(_04617_ ), .ZN(_04618_ ) );
NOR2_X1 _12237_ ( .A1(_04531_ ), .A2(_03586_ ), .ZN(_04619_ ) );
AND2_X1 _12238_ ( .A1(_03610_ ), .A2(_04619_ ), .ZN(_04620_ ) );
AOI21_X1 _12239_ ( .A(_03609_ ), .B1(_03072_ ), .B2(_03053_ ), .ZN(_04621_ ) );
OAI211_X1 _12240_ ( .A(_03561_ ), .B(_03538_ ), .C1(_04620_ ), .C2(_04621_ ), .ZN(_04622_ ) );
NAND3_X1 _12241_ ( .A1(_03560_ ), .A2(_03558_ ), .A3(_03556_ ), .ZN(_04623_ ) );
NOR2_X1 _12242_ ( .A1(_03537_ ), .A2(_03126_ ), .ZN(_04624_ ) );
NAND2_X1 _12243_ ( .A1(_03561_ ), .A2(_04624_ ), .ZN(_04625_ ) );
AND3_X2 _12244_ ( .A1(_04622_ ), .A2(_04623_ ), .A3(_04625_ ), .ZN(_04626_ ) );
INV_X1 _12245_ ( .A(_03701_ ), .ZN(_04627_ ) );
NOR2_X1 _12246_ ( .A1(_04626_ ), .A2(_04627_ ), .ZN(_04628_ ) );
INV_X2 _12247_ ( .A(_04628_ ), .ZN(_04629_ ) );
NOR2_X1 _12248_ ( .A1(_03156_ ), .A2(_03653_ ), .ZN(_04630_ ) );
NOR2_X1 _12249_ ( .A1(_04319_ ), .A2(_03631_ ), .ZN(_04631_ ) );
AOI21_X1 _12250_ ( .A(_04630_ ), .B1(_03654_ ), .B2(_04631_ ), .ZN(_04632_ ) );
INV_X1 _12251_ ( .A(_03700_ ), .ZN(_04633_ ) );
INV_X1 _12252_ ( .A(_03677_ ), .ZN(_04634_ ) );
NOR3_X1 _12253_ ( .A1(_04632_ ), .A2(_04633_ ), .A3(_04634_ ), .ZN(_04635_ ) );
INV_X1 _12254_ ( .A(_04635_ ), .ZN(_04636_ ) );
NOR2_X1 _12255_ ( .A1(_02358_ ), .A2(_03698_ ), .ZN(_04637_ ) );
AND2_X1 _12256_ ( .A1(_03677_ ), .A2(_04637_ ), .ZN(_04638_ ) );
INV_X1 _12257_ ( .A(_03676_ ), .ZN(_04639_ ) );
AOI21_X1 _12258_ ( .A(_04638_ ), .B1(_03185_ ), .B2(_04639_ ), .ZN(_04640_ ) );
AND4_X4 _12259_ ( .A1(_04618_ ), .A2(_04629_ ), .A3(_04636_ ), .A4(_04640_ ), .ZN(_04641_ ) );
AND2_X2 _12260_ ( .A1(_04289_ ), .A2(\ID_EX_typ [2] ), .ZN(_04642_ ) );
AND3_X4 _12261_ ( .A1(_04592_ ), .A2(_04641_ ), .A3(_04642_ ), .ZN(_04643_ ) );
AND2_X1 _12262_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_8 ), .ZN(_04644_ ) );
AND2_X2 _12263_ ( .A1(_04644_ ), .A2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .ZN(_04645_ ) );
INV_X1 _12264_ ( .A(_04645_ ), .ZN(_04646_ ) );
AOI21_X1 _12265_ ( .A(_04646_ ), .B1(_04592_ ), .B2(_04641_ ), .ZN(_04647_ ) );
OR4_X4 _12266_ ( .A1(_04553_ ), .A2(_04643_ ), .A3(_04647_ ), .A4(_04290_ ), .ZN(_04648_ ) );
INV_X1 _12267_ ( .A(\ID_EX_typ [2] ), .ZN(_04649_ ) );
NOR3_X1 _12268_ ( .A1(_04649_ ), .A2(\ID_EX_typ [1] ), .A3(fanout_net_8 ), .ZN(_04650_ ) );
AND3_X1 _12269_ ( .A1(_04546_ ), .A2(_04552_ ), .A3(_04650_ ), .ZN(_04651_ ) );
OAI221_X2 _12270_ ( .A(_03469_ ), .B1(_04288_ ), .B2(_04291_ ), .C1(_04648_ ), .C2(_04651_ ), .ZN(_04652_ ) );
BUF_X4 _12271_ ( .A(_04652_ ), .Z(_04653_ ) );
OAI21_X2 _12272_ ( .A(_03468_ ), .B1(_03999_ ), .B2(_04287_ ), .ZN(_04654_ ) );
AND2_X4 _12273_ ( .A1(_04653_ ), .A2(_04654_ ), .ZN(_04655_ ) );
BUF_X16 _12274_ ( .A(_04655_ ), .Z(_04656_ ) );
BUF_X32 _12275_ ( .A(_04656_ ), .Z(_04657_ ) );
MUX2_X1 _12276_ ( .A(_03466_ ), .B(_03370_ ), .S(_04657_ ), .Z(_04658_ ) );
BUF_X4 _12277_ ( .A(_03372_ ), .Z(_04659_ ) );
AOI21_X1 _12278_ ( .A(_03447_ ), .B1(_04658_ ), .B2(_04659_ ), .ZN(_04660_ ) );
BUF_X4 _12279_ ( .A(_02273_ ), .Z(_04661_ ) );
BUF_X4 _12280_ ( .A(_04661_ ), .Z(_04662_ ) );
AOI211_X1 _12281_ ( .A(_03248_ ), .B(_03371_ ), .C1(_04660_ ), .C2(_04662_ ), .ZN(_00158_ ) );
BUF_X4 _12282_ ( .A(_03248_ ), .Z(_04663_ ) );
AND3_X1 _12283_ ( .A1(_03455_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_04664_ ) );
AND2_X1 _12284_ ( .A1(\ID_EX_pc [15] ), .A2(\ID_EX_pc [14] ), .ZN(_04665_ ) );
AND4_X1 _12285_ ( .A1(\ID_EX_pc [17] ), .A2(_04664_ ), .A3(\ID_EX_pc [16] ), .A4(_04665_ ), .ZN(_04666_ ) );
AND2_X1 _12286_ ( .A1(_03454_ ), .A2(_04666_ ), .ZN(_04667_ ) );
AND4_X1 _12287_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_04668_ ) );
AND2_X1 _12288_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_04669_ ) );
AND4_X1 _12289_ ( .A1(\ID_EX_pc [21] ), .A2(_04668_ ), .A3(\ID_EX_pc [20] ), .A4(_04669_ ), .ZN(_04670_ ) );
NAND2_X1 _12290_ ( .A1(_04667_ ), .A2(_04670_ ), .ZN(_04671_ ) );
INV_X1 _12291_ ( .A(\ID_EX_pc [27] ), .ZN(_04672_ ) );
INV_X1 _12292_ ( .A(\ID_EX_pc [26] ), .ZN(_04673_ ) );
NOR3_X1 _12293_ ( .A1(_04671_ ), .A2(_04672_ ), .A3(_04673_ ), .ZN(_04674_ ) );
NAND2_X1 _12294_ ( .A1(_04674_ ), .A2(\ID_EX_pc [28] ), .ZN(_04675_ ) );
XNOR2_X1 _12295_ ( .A(_04675_ ), .B(\ID_EX_pc [29] ), .ZN(_04676_ ) );
AOI21_X1 _12296_ ( .A(_04676_ ), .B1(_04653_ ), .B2(_04654_ ), .ZN(_04677_ ) );
BUF_X4 _12297_ ( .A(_04657_ ), .Z(_04678_ ) );
NAND2_X1 _12298_ ( .A1(_03364_ ), .A2(_03365_ ), .ZN(_04679_ ) );
XOR2_X1 _12299_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .Z(_04680_ ) );
XNOR2_X1 _12300_ ( .A(_04679_ ), .B(_04680_ ), .ZN(_04681_ ) );
AOI211_X1 _12301_ ( .A(fanout_net_10 ), .B(_04677_ ), .C1(_04678_ ), .C2(_04681_ ), .ZN(_04682_ ) );
CLKBUF_X2 _12302_ ( .A(_03421_ ), .Z(_04683_ ) );
BUF_X2 _12303_ ( .A(_03436_ ), .Z(_04684_ ) );
CLKBUF_X2 _12304_ ( .A(_03426_ ), .Z(_04685_ ) );
AND4_X1 _12305_ ( .A1(\mycsreg.CSReg[3][29] ), .A2(_04683_ ), .A3(_04684_ ), .A4(_04685_ ), .ZN(_04686_ ) );
AND3_X1 _12306_ ( .A1(_03397_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_04687_ ) );
AND4_X1 _12307_ ( .A1(\ID_EX_csr [4] ), .A2(_03432_ ), .A3(_03408_ ), .A4(_03413_ ), .ZN(_04688_ ) );
AOI21_X1 _12308_ ( .A(_04686_ ), .B1(_04687_ ), .B2(_04688_ ), .ZN(_04689_ ) );
BUF_X2 _12309_ ( .A(_03405_ ), .Z(_04690_ ) );
BUF_X2 _12310_ ( .A(_03411_ ), .Z(_04691_ ) );
AND3_X1 _12311_ ( .A1(_04690_ ), .A2(\mtvec [29] ), .A3(_04691_ ), .ZN(_04692_ ) );
INV_X1 _12312_ ( .A(_04692_ ), .ZN(_04693_ ) );
INV_X1 _12313_ ( .A(_03400_ ), .ZN(_04694_ ) );
NAND4_X1 _12314_ ( .A1(_03408_ ), .A2(_03423_ ), .A3(_03413_ ), .A4(_03401_ ), .ZN(_04695_ ) );
NOR2_X1 _12315_ ( .A1(_04694_ ), .A2(_04695_ ), .ZN(_04696_ ) );
BUF_X2 _12316_ ( .A(_04696_ ), .Z(_04697_ ) );
NAND2_X1 _12317_ ( .A1(_04697_ ), .A2(\mepc [29] ), .ZN(_04698_ ) );
CLKBUF_X2 _12318_ ( .A(_03415_ ), .Z(_04699_ ) );
BUF_X2 _12319_ ( .A(_04699_ ), .Z(_04700_ ) );
BUF_X2 _12320_ ( .A(_03438_ ), .Z(_04701_ ) );
BUF_X2 _12321_ ( .A(_03403_ ), .Z(_04702_ ) );
NAND4_X1 _12322_ ( .A1(_04700_ ), .A2(_04701_ ), .A3(_04702_ ), .A4(\mycsreg.CSReg[0][29] ), .ZN(_04703_ ) );
NAND4_X1 _12323_ ( .A1(_04689_ ), .A2(_04693_ ), .A3(_04698_ ), .A4(_04703_ ), .ZN(_04704_ ) );
AND4_X1 _12324_ ( .A1(_03377_ ), .A2(_03391_ ), .A3(_03386_ ), .A4(_03388_ ), .ZN(_04705_ ) );
AND2_X1 _12325_ ( .A1(_03383_ ), .A2(_03387_ ), .ZN(_04706_ ) );
NAND4_X1 _12326_ ( .A1(_04705_ ), .A2(_03376_ ), .A3(_03385_ ), .A4(_04706_ ), .ZN(_04707_ ) );
INV_X1 _12327_ ( .A(_03382_ ), .ZN(_04708_ ) );
NAND2_X1 _12328_ ( .A1(_03375_ ), .A2(_03380_ ), .ZN(_04709_ ) );
NOR4_X1 _12329_ ( .A1(_04707_ ), .A2(_04708_ ), .A3(_04709_ ), .A4(_03390_ ), .ZN(_04710_ ) );
INV_X1 _12330_ ( .A(_04710_ ), .ZN(_04711_ ) );
BUF_X4 _12331_ ( .A(_02332_ ), .Z(_04712_ ) );
BUF_X4 _12332_ ( .A(_04712_ ), .Z(_04713_ ) );
OAI21_X1 _12333_ ( .A(_04704_ ), .B1(_04711_ ), .B2(_04713_ ), .ZN(_04714_ ) );
BUF_X4 _12334_ ( .A(_02331_ ), .Z(_04715_ ) );
NAND3_X1 _12335_ ( .A1(_04710_ ), .A2(\EX_LS_result_csreg_mem [29] ), .A3(_04715_ ), .ZN(_04716_ ) );
AOI21_X1 _12336_ ( .A(_04659_ ), .B1(_04714_ ), .B2(_04716_ ), .ZN(_04717_ ) );
OAI21_X1 _12337_ ( .A(_04662_ ), .B1(_04682_ ), .B2(_04717_ ), .ZN(_04718_ ) );
MUX2_X1 _12338_ ( .A(_04681_ ), .B(_03228_ ), .S(fanout_net_8 ), .Z(_04719_ ) );
BUF_X2 _12339_ ( .A(_02273_ ), .Z(_04720_ ) );
OR2_X2 _12340_ ( .A1(_04719_ ), .A2(_04720_ ), .ZN(_04721_ ) );
AOI21_X1 _12341_ ( .A(_04663_ ), .B1(_04718_ ), .B2(_04721_ ), .ZN(_00159_ ) );
NAND3_X1 _12342_ ( .A1(_03454_ ), .A2(_04666_ ), .A3(_04669_ ), .ZN(_04722_ ) );
XNOR2_X1 _12343_ ( .A(_04722_ ), .B(\ID_EX_pc [20] ), .ZN(_04723_ ) );
OAI21_X1 _12344_ ( .A(_03266_ ), .B1(_03317_ ), .B2(_03325_ ), .ZN(_04724_ ) );
AND2_X1 _12345_ ( .A1(_04724_ ), .A2(_03337_ ), .ZN(_04725_ ) );
XOR2_X1 _12346_ ( .A(_04725_ ), .B(_03253_ ), .Z(_04726_ ) );
MUX2_X1 _12347_ ( .A(_04723_ ), .B(_04726_ ), .S(_04657_ ), .Z(_04727_ ) );
OR2_X2 _12348_ ( .A1(_04727_ ), .A2(fanout_net_10 ), .ZN(_04728_ ) );
BUF_X4 _12349_ ( .A(_02274_ ), .Z(_04729_ ) );
BUF_X4 _12350_ ( .A(_03372_ ), .Z(_04730_ ) );
BUF_X2 _12351_ ( .A(_03442_ ), .Z(_04731_ ) );
BUF_X2 _12352_ ( .A(_03444_ ), .Z(_04732_ ) );
NAND3_X1 _12353_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [20] ), .ZN(_04733_ ) );
AND2_X1 _12354_ ( .A1(_03433_ ), .A2(_03428_ ), .ZN(_04734_ ) );
AND2_X1 _12355_ ( .A1(_03433_ ), .A2(_03420_ ), .ZN(_04735_ ) );
NOR2_X1 _12356_ ( .A1(_04734_ ), .A2(_04735_ ), .ZN(_04736_ ) );
BUF_X2 _12357_ ( .A(_03421_ ), .Z(_04737_ ) );
BUF_X2 _12358_ ( .A(_04737_ ), .Z(_04738_ ) );
BUF_X4 _12359_ ( .A(_03400_ ), .Z(_04739_ ) );
BUF_X2 _12360_ ( .A(_04739_ ), .Z(_04740_ ) );
BUF_X2 _12361_ ( .A(_04740_ ), .Z(_04741_ ) );
NAND4_X1 _12362_ ( .A1(_04738_ ), .A2(_03437_ ), .A3(\mycsreg.CSReg[3][20] ), .A4(_04741_ ), .ZN(_04742_ ) );
NAND4_X1 _12363_ ( .A1(_03429_ ), .A2(_03437_ ), .A3(\mepc [20] ), .A4(_04741_ ), .ZN(_04743_ ) );
AND2_X1 _12364_ ( .A1(_04742_ ), .A2(_04743_ ), .ZN(_04744_ ) );
BUF_X2 _12365_ ( .A(_03405_ ), .Z(_04745_ ) );
BUF_X2 _12366_ ( .A(_03411_ ), .Z(_04746_ ) );
AND3_X1 _12367_ ( .A1(_04745_ ), .A2(\mtvec [20] ), .A3(_04746_ ), .ZN(_04747_ ) );
BUF_X2 _12368_ ( .A(_03405_ ), .Z(_04748_ ) );
CLKBUF_X2 _12369_ ( .A(_03416_ ), .Z(_04749_ ) );
AND3_X1 _12370_ ( .A1(_04748_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_04749_ ), .ZN(_04750_ ) );
NOR2_X1 _12371_ ( .A1(_04747_ ), .A2(_04750_ ), .ZN(_04751_ ) );
AND3_X1 _12372_ ( .A1(_04736_ ), .A2(_04744_ ), .A3(_04751_ ), .ZN(_04752_ ) );
OAI21_X1 _12373_ ( .A(_04733_ ), .B1(_04752_ ), .B2(_03394_ ), .ZN(_04753_ ) );
OAI211_X1 _12374_ ( .A(_04728_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_04753_ ), .ZN(_04754_ ) );
BUF_X4 _12375_ ( .A(_02272_ ), .Z(_04755_ ) );
BUF_X4 _12376_ ( .A(_04755_ ), .Z(_04756_ ) );
AND3_X1 _12377_ ( .A1(_03199_ ), .A2(fanout_net_8 ), .A3(_03196_ ), .ZN(_04757_ ) );
BUF_X4 _12378_ ( .A(_03250_ ), .Z(_04758_ ) );
BUF_X2 _12379_ ( .A(_04758_ ), .Z(_04759_ ) );
AND2_X1 _12380_ ( .A1(_04726_ ), .A2(_04759_ ), .ZN(_04760_ ) );
OAI21_X1 _12381_ ( .A(_04756_ ), .B1(_04757_ ), .B2(_04760_ ), .ZN(_04761_ ) );
AOI21_X1 _12382_ ( .A(_04663_ ), .B1(_04754_ ), .B2(_04761_ ), .ZN(_00160_ ) );
NAND3_X1 _12383_ ( .A1(_03454_ ), .A2(\ID_EX_pc [18] ), .A3(_04666_ ), .ZN(_04762_ ) );
XNOR2_X1 _12384_ ( .A(_04762_ ), .B(\ID_EX_pc [19] ), .ZN(_04763_ ) );
OR2_X1 _12385_ ( .A1(_03317_ ), .A2(_03325_ ), .ZN(_04764_ ) );
AOI21_X1 _12386_ ( .A(_03336_ ), .B1(_04764_ ), .B2(_03265_ ), .ZN(_04765_ ) );
XNOR2_X1 _12387_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .ZN(_04766_ ) );
NOR2_X1 _12388_ ( .A1(_04765_ ), .A2(_04766_ ), .ZN(_04767_ ) );
NOR2_X1 _12389_ ( .A1(_04767_ ), .A2(_03330_ ), .ZN(_04768_ ) );
XNOR2_X1 _12390_ ( .A(_04768_ ), .B(_03260_ ), .ZN(_04769_ ) );
MUX2_X1 _12391_ ( .A(_04763_ ), .B(_04769_ ), .S(_04656_ ), .Z(_04770_ ) );
OR2_X2 _12392_ ( .A1(_04770_ ), .A2(fanout_net_10 ), .ZN(_04771_ ) );
AND3_X1 _12393_ ( .A1(_04748_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_04749_ ), .ZN(_04772_ ) );
NOR3_X1 _12394_ ( .A1(_02332_ ), .A2(_04709_ ), .A3(_03390_ ), .ZN(_04773_ ) );
AND4_X2 _12395_ ( .A1(_03376_ ), .A2(_03391_ ), .A3(_03385_ ), .A4(_03386_ ), .ZN(_04774_ ) );
AND2_X2 _12396_ ( .A1(_04773_ ), .A2(_04774_ ), .ZN(_04775_ ) );
BUF_X4 _12397_ ( .A(_04775_ ), .Z(_04776_ ) );
AND4_X1 _12398_ ( .A1(_03382_ ), .A2(_04706_ ), .A3(_03377_ ), .A4(_03388_ ), .ZN(_04777_ ) );
BUF_X4 _12399_ ( .A(_04777_ ), .Z(_04778_ ) );
BUF_X2 _12400_ ( .A(_04778_ ), .Z(_04779_ ) );
AOI21_X1 _12401_ ( .A(_04772_ ), .B1(_04776_ ), .B2(_04779_ ), .ZN(_04780_ ) );
BUF_X2 _12402_ ( .A(_04697_ ), .Z(_04781_ ) );
NAND2_X1 _12403_ ( .A1(_04781_ ), .A2(\mepc [19] ), .ZN(_04782_ ) );
AND3_X1 _12404_ ( .A1(_04687_ ), .A2(\ID_EX_csr [4] ), .A3(_03432_ ), .ZN(_04783_ ) );
AND2_X2 _12405_ ( .A1(_04783_ ), .A2(_03420_ ), .ZN(_04784_ ) );
AND3_X1 _12406_ ( .A1(_04748_ ), .A2(\mtvec [19] ), .A3(_04746_ ), .ZN(_04785_ ) );
AND4_X1 _12407_ ( .A1(\mycsreg.CSReg[3][19] ), .A2(_04683_ ), .A3(_04684_ ), .A4(_04685_ ), .ZN(_04786_ ) );
NOR3_X1 _12408_ ( .A1(_04784_ ), .A2(_04785_ ), .A3(_04786_ ), .ZN(_04787_ ) );
NAND3_X1 _12409_ ( .A1(_04780_ ), .A2(_04782_ ), .A3(_04787_ ), .ZN(_04788_ ) );
BUF_X4 _12410_ ( .A(_04778_ ), .Z(_04789_ ) );
INV_X1 _12411_ ( .A(\EX_LS_result_csreg_mem [19] ), .ZN(_04790_ ) );
BUF_X2 _12412_ ( .A(_04774_ ), .Z(_04791_ ) );
BUF_X2 _12413_ ( .A(_04773_ ), .Z(_04792_ ) );
NAND4_X1 _12414_ ( .A1(_04789_ ), .A2(_04790_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_04793_ ) );
NAND2_X1 _12415_ ( .A1(_04788_ ), .A2(_04793_ ), .ZN(_04794_ ) );
INV_X1 _12416_ ( .A(_04794_ ), .ZN(_04795_ ) );
OAI211_X1 _12417_ ( .A(_04771_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_04795_ ), .ZN(_04796_ ) );
NAND2_X1 _12418_ ( .A1(_03206_ ), .A2(fanout_net_8 ), .ZN(_04797_ ) );
OAI211_X1 _12419_ ( .A(_04797_ ), .B(_04756_ ), .C1(fanout_net_8 ), .C2(_04769_ ), .ZN(_04798_ ) );
AOI21_X1 _12420_ ( .A(_04663_ ), .B1(_04796_ ), .B2(_04798_ ), .ZN(_00161_ ) );
NAND2_X1 _12421_ ( .A1(_04696_ ), .A2(\mepc [18] ), .ZN(_04799_ ) );
NAND3_X1 _12422_ ( .A1(_03404_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_03415_ ), .ZN(_04800_ ) );
NAND2_X1 _12423_ ( .A1(_04799_ ), .A2(_04800_ ), .ZN(_04801_ ) );
AOI21_X1 _12424_ ( .A(_04801_ ), .B1(_04775_ ), .B2(_04777_ ), .ZN(_04802_ ) );
AND3_X1 _12425_ ( .A1(_03404_ ), .A2(\mtvec [18] ), .A3(_03410_ ), .ZN(_04803_ ) );
AND4_X1 _12426_ ( .A1(\mycsreg.CSReg[3][18] ), .A2(_03420_ ), .A3(_03424_ ), .A4(_03400_ ), .ZN(_04804_ ) );
NOR3_X1 _12427_ ( .A1(_04784_ ), .A2(_04803_ ), .A3(_04804_ ), .ZN(_04805_ ) );
NAND2_X1 _12428_ ( .A1(_04802_ ), .A2(_04805_ ), .ZN(_04806_ ) );
INV_X1 _12429_ ( .A(\EX_LS_result_csreg_mem [18] ), .ZN(_04807_ ) );
AND4_X1 _12430_ ( .A1(_04807_ ), .A2(_04777_ ), .A3(_04774_ ), .A4(_04773_ ), .ZN(_04808_ ) );
INV_X1 _12431_ ( .A(_04808_ ), .ZN(_04809_ ) );
AND2_X1 _12432_ ( .A1(_04806_ ), .A2(_04809_ ), .ZN(_04810_ ) );
INV_X4 _12433_ ( .A(_04656_ ), .ZN(_04811_ ) );
BUF_X4 _12434_ ( .A(_04811_ ), .Z(_04812_ ) );
XNOR2_X1 _12435_ ( .A(_04765_ ), .B(_03261_ ), .ZN(_04813_ ) );
INV_X1 _12436_ ( .A(_04813_ ), .ZN(_04814_ ) );
OAI21_X1 _12437_ ( .A(_04659_ ), .B1(_04812_ ), .B2(_04814_ ), .ZN(_04815_ ) );
XNOR2_X1 _12438_ ( .A(_04667_ ), .B(\ID_EX_pc [18] ), .ZN(_04816_ ) );
AOI21_X1 _12439_ ( .A(_04816_ ), .B1(_04653_ ), .B2(_04654_ ), .ZN(_04817_ ) );
OAI221_X1 _12440_ ( .A(_02275_ ), .B1(_04659_ ), .B2(_04810_ ), .C1(_04815_ ), .C2(_04817_ ), .ZN(_04818_ ) );
AOI21_X1 _12441_ ( .A(_02274_ ), .B1(_04814_ ), .B2(_03252_ ), .ZN(_04819_ ) );
BUF_X4 _12442_ ( .A(_03251_ ), .Z(_04820_ ) );
OAI21_X1 _12443_ ( .A(_04819_ ), .B1(_03208_ ), .B2(_04820_ ), .ZN(_04821_ ) );
AOI21_X1 _12444_ ( .A(_04663_ ), .B1(_04818_ ), .B2(_04821_ ), .ZN(_00162_ ) );
NAND3_X1 _12445_ ( .A1(_03454_ ), .A2(_04665_ ), .A3(_04664_ ), .ZN(_04822_ ) );
INV_X1 _12446_ ( .A(\ID_EX_pc [16] ), .ZN(_04823_ ) );
NOR2_X1 _12447_ ( .A1(_04822_ ), .A2(_04823_ ), .ZN(_04824_ ) );
XNOR2_X1 _12448_ ( .A(_04824_ ), .B(_03335_ ), .ZN(_04825_ ) );
AOI21_X1 _12449_ ( .A(_04825_ ), .B1(_04653_ ), .B2(_04654_ ), .ZN(_04826_ ) );
OAI21_X1 _12450_ ( .A(_03264_ ), .B1(_03317_ ), .B2(_03325_ ), .ZN(_04827_ ) );
NAND2_X1 _12451_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_04828_ ) );
NAND2_X1 _12452_ ( .A1(_04827_ ), .A2(_04828_ ), .ZN(_04829_ ) );
XOR2_X1 _12453_ ( .A(_04829_ ), .B(_03263_ ), .Z(_04830_ ) );
INV_X1 _12454_ ( .A(_04830_ ), .ZN(_04831_ ) );
AOI211_X1 _12455_ ( .A(fanout_net_10 ), .B(_04826_ ), .C1(_04678_ ), .C2(_04831_ ), .ZN(_04832_ ) );
AND3_X1 _12456_ ( .A1(_03420_ ), .A2(\ID_EX_csr [4] ), .A3(_03432_ ), .ZN(_04833_ ) );
NAND2_X1 _12457_ ( .A1(_04833_ ), .A2(_04687_ ), .ZN(_04834_ ) );
NAND2_X1 _12458_ ( .A1(_04688_ ), .A2(_04687_ ), .ZN(_04835_ ) );
BUF_X2 _12459_ ( .A(_04737_ ), .Z(_04836_ ) );
NAND4_X1 _12460_ ( .A1(_04836_ ), .A2(_03437_ ), .A3(\mycsreg.CSReg[3][17] ), .A4(_03438_ ), .ZN(_04837_ ) );
AND3_X1 _12461_ ( .A1(_04834_ ), .A2(_04835_ ), .A3(_04837_ ), .ZN(_04838_ ) );
BUF_X2 _12462_ ( .A(_03406_ ), .Z(_04839_ ) );
AND3_X1 _12463_ ( .A1(_04839_ ), .A2(\mtvec [17] ), .A3(_04746_ ), .ZN(_04840_ ) );
INV_X1 _12464_ ( .A(_04840_ ), .ZN(_04841_ ) );
NAND2_X1 _12465_ ( .A1(_04697_ ), .A2(\mepc [17] ), .ZN(_04842_ ) );
NAND4_X1 _12466_ ( .A1(_04700_ ), .A2(_04701_ ), .A3(_04702_ ), .A4(\mycsreg.CSReg[0][17] ), .ZN(_04843_ ) );
NAND4_X1 _12467_ ( .A1(_04838_ ), .A2(_04841_ ), .A3(_04842_ ), .A4(_04843_ ), .ZN(_04844_ ) );
OAI21_X1 _12468_ ( .A(_04844_ ), .B1(_04711_ ), .B2(_04713_ ), .ZN(_04845_ ) );
NAND3_X1 _12469_ ( .A1(_04710_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_04715_ ), .ZN(_04846_ ) );
AOI21_X1 _12470_ ( .A(_04659_ ), .B1(_04845_ ), .B2(_04846_ ), .ZN(_04847_ ) );
OAI21_X1 _12471_ ( .A(_04662_ ), .B1(_04832_ ), .B2(_04847_ ), .ZN(_04848_ ) );
NAND2_X1 _12472_ ( .A1(_03210_ ), .A2(fanout_net_8 ), .ZN(_04849_ ) );
OAI211_X1 _12473_ ( .A(_04849_ ), .B(_04756_ ), .C1(fanout_net_8 ), .C2(_04830_ ), .ZN(_04850_ ) );
AOI21_X1 _12474_ ( .A(_04663_ ), .B1(_04848_ ), .B2(_04850_ ), .ZN(_00163_ ) );
XNOR2_X1 _12475_ ( .A(_04822_ ), .B(\ID_EX_pc [16] ), .ZN(_04851_ ) );
NAND2_X1 _12476_ ( .A1(_04812_ ), .A2(_04851_ ), .ZN(_04852_ ) );
XOR2_X1 _12477_ ( .A(_04764_ ), .B(_03264_ ), .Z(_04853_ ) );
NAND3_X1 _12478_ ( .A1(_04653_ ), .A2(_04654_ ), .A3(_04853_ ), .ZN(_04854_ ) );
AOI21_X1 _12479_ ( .A(fanout_net_10 ), .B1(_04852_ ), .B2(_04854_ ), .ZN(_04855_ ) );
BUF_X4 _12480_ ( .A(_03372_ ), .Z(_04856_ ) );
INV_X1 _12481_ ( .A(_04734_ ), .ZN(_04857_ ) );
INV_X1 _12482_ ( .A(_04735_ ), .ZN(_04858_ ) );
NAND4_X1 _12483_ ( .A1(_04737_ ), .A2(_03436_ ), .A3(\mycsreg.CSReg[3][16] ), .A4(_04740_ ), .ZN(_04859_ ) );
BUF_X2 _12484_ ( .A(_03428_ ), .Z(_04860_ ) );
NAND4_X1 _12485_ ( .A1(_04860_ ), .A2(_03436_ ), .A3(\mepc [16] ), .A4(_04740_ ), .ZN(_04861_ ) );
AND2_X1 _12486_ ( .A1(_04859_ ), .A2(_04861_ ), .ZN(_04862_ ) );
NAND3_X1 _12487_ ( .A1(_04857_ ), .A2(_04858_ ), .A3(_04862_ ), .ZN(_04863_ ) );
NAND3_X1 _12488_ ( .A1(_04748_ ), .A2(\mtvec [16] ), .A3(_04746_ ), .ZN(_04864_ ) );
NAND3_X1 _12489_ ( .A1(_04745_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_04699_ ), .ZN(_04865_ ) );
NAND2_X1 _12490_ ( .A1(_04864_ ), .A2(_04865_ ), .ZN(_04866_ ) );
OAI21_X1 _12491_ ( .A(_03395_ ), .B1(_04863_ ), .B2(_04866_ ), .ZN(_04867_ ) );
NAND3_X1 _12492_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [16] ), .ZN(_04868_ ) );
AOI21_X1 _12493_ ( .A(_04856_ ), .B1(_04867_ ), .B2(_04868_ ), .ZN(_04869_ ) );
OAI21_X1 _12494_ ( .A(_04662_ ), .B1(_04855_ ), .B2(_04869_ ), .ZN(_04870_ ) );
OAI21_X1 _12495_ ( .A(fanout_net_8 ), .B1(_03211_ ), .B2(_03201_ ), .ZN(_04871_ ) );
OAI211_X1 _12496_ ( .A(_04871_ ), .B(_04756_ ), .C1(fanout_net_8 ), .C2(_04853_ ), .ZN(_04872_ ) );
AOI21_X1 _12497_ ( .A(_04663_ ), .B1(_04870_ ), .B2(_04872_ ), .ZN(_00164_ ) );
BUF_X16 _12498_ ( .A(_04657_ ), .Z(_04873_ ) );
INV_X1 _12499_ ( .A(_03316_ ), .ZN(_04874_ ) );
AOI21_X1 _12500_ ( .A(_04874_ ), .B1(_03303_ ), .B2(_03311_ ), .ZN(_04875_ ) );
OR2_X1 _12501_ ( .A1(_04875_ ), .A2(_03322_ ), .ZN(_04876_ ) );
AOI21_X1 _12502_ ( .A(_03313_ ), .B1(_04876_ ), .B2(_03321_ ), .ZN(_04877_ ) );
NOR2_X1 _12503_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04878_ ) );
NOR3_X1 _12504_ ( .A1(_04877_ ), .A2(_03318_ ), .A3(_04878_ ), .ZN(_04879_ ) );
NOR2_X1 _12505_ ( .A1(_04879_ ), .A2(_03318_ ), .ZN(_04880_ ) );
XNOR2_X1 _12506_ ( .A(_04880_ ), .B(_03267_ ), .ZN(_04881_ ) );
AOI21_X2 _12507_ ( .A(fanout_net_10 ), .B1(_04873_ ), .B2(_04881_ ), .ZN(_04882_ ) );
NAND3_X1 _12508_ ( .A1(_03454_ ), .A2(\ID_EX_pc [14] ), .A3(_04664_ ), .ZN(_04883_ ) );
INV_X1 _12509_ ( .A(\ID_EX_pc [15] ), .ZN(_04884_ ) );
XNOR2_X1 _12510_ ( .A(_04883_ ), .B(_04884_ ), .ZN(_04885_ ) );
OAI21_X1 _12511_ ( .A(_04882_ ), .B1(_04678_ ), .B2(_04885_ ), .ZN(_04886_ ) );
NAND3_X1 _12512_ ( .A1(_04690_ ), .A2(\mtvec [15] ), .A3(_04691_ ), .ZN(_04887_ ) );
NAND3_X1 _12513_ ( .A1(_03406_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_03416_ ), .ZN(_04888_ ) );
AND2_X1 _12514_ ( .A1(_04887_ ), .A2(_04888_ ), .ZN(_04889_ ) );
AND4_X1 _12515_ ( .A1(\mepc [15] ), .A2(_04860_ ), .A3(_03425_ ), .A4(_03426_ ), .ZN(_04890_ ) );
AOI21_X1 _12516_ ( .A(_04890_ ), .B1(_04836_ ), .B2(_03433_ ), .ZN(_04891_ ) );
NAND4_X1 _12517_ ( .A1(_04836_ ), .A2(_03437_ ), .A3(\mycsreg.CSReg[3][15] ), .A4(_03438_ ), .ZN(_04892_ ) );
NAND3_X1 _12518_ ( .A1(_04889_ ), .A2(_04891_ ), .A3(_04892_ ), .ZN(_04893_ ) );
NAND2_X1 _12519_ ( .A1(_03396_ ), .A2(_04893_ ), .ZN(_04894_ ) );
NAND3_X1 _12520_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [15] ), .ZN(_04895_ ) );
AND2_X1 _12521_ ( .A1(_04894_ ), .A2(_04895_ ), .ZN(_04896_ ) );
INV_X1 _12522_ ( .A(_04896_ ), .ZN(_04897_ ) );
OAI211_X1 _12523_ ( .A(_04886_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_04897_ ), .ZN(_04898_ ) );
NAND2_X1 _12524_ ( .A1(_03221_ ), .A2(fanout_net_8 ), .ZN(_04899_ ) );
OAI211_X1 _12525_ ( .A(_04899_ ), .B(_04756_ ), .C1(fanout_net_8 ), .C2(_04881_ ), .ZN(_04900_ ) );
AOI21_X1 _12526_ ( .A(_04663_ ), .B1(_04898_ ), .B2(_04900_ ), .ZN(_00165_ ) );
XNOR2_X1 _12527_ ( .A(_04877_ ), .B(_03268_ ), .ZN(_04901_ ) );
AOI21_X2 _12528_ ( .A(fanout_net_10 ), .B1(_04873_ ), .B2(_04901_ ), .ZN(_04902_ ) );
NAND2_X1 _12529_ ( .A1(_03454_ ), .A2(_04664_ ), .ZN(_04903_ ) );
INV_X1 _12530_ ( .A(\ID_EX_pc [14] ), .ZN(_04904_ ) );
XNOR2_X1 _12531_ ( .A(_04903_ ), .B(_04904_ ), .ZN(_04905_ ) );
OAI21_X1 _12532_ ( .A(_04902_ ), .B1(_04678_ ), .B2(_04905_ ), .ZN(_04906_ ) );
NAND4_X1 _12533_ ( .A1(_03428_ ), .A2(_03435_ ), .A3(\mepc [14] ), .A4(_04739_ ), .ZN(_04907_ ) );
NAND4_X1 _12534_ ( .A1(_03421_ ), .A2(_03435_ ), .A3(\mycsreg.CSReg[3][14] ), .A4(_04739_ ), .ZN(_04908_ ) );
AND2_X1 _12535_ ( .A1(_04907_ ), .A2(_04908_ ), .ZN(_04909_ ) );
NAND3_X1 _12536_ ( .A1(_03404_ ), .A2(\mtvec [14] ), .A3(_03410_ ), .ZN(_04910_ ) );
NAND3_X1 _12537_ ( .A1(_03404_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_03415_ ), .ZN(_04911_ ) );
AND2_X1 _12538_ ( .A1(_04910_ ), .A2(_04911_ ), .ZN(_04912_ ) );
NAND3_X1 _12539_ ( .A1(_04736_ ), .A2(_04909_ ), .A3(_04912_ ), .ZN(_04913_ ) );
NAND2_X1 _12540_ ( .A1(_04913_ ), .A2(_03395_ ), .ZN(_04914_ ) );
NAND3_X1 _12541_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(\EX_LS_result_csreg_mem [14] ), .ZN(_04915_ ) );
AND2_X1 _12542_ ( .A1(_04914_ ), .A2(_04915_ ), .ZN(_04916_ ) );
INV_X1 _12543_ ( .A(_04916_ ), .ZN(_04917_ ) );
OAI211_X1 _12544_ ( .A(_04906_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_04917_ ), .ZN(_04918_ ) );
OR2_X1 _12545_ ( .A1(_03222_ ), .A2(_03251_ ), .ZN(_04919_ ) );
OAI211_X1 _12546_ ( .A(_04919_ ), .B(_04756_ ), .C1(fanout_net_8 ), .C2(_04901_ ), .ZN(_04920_ ) );
AOI21_X1 _12547_ ( .A(_04663_ ), .B1(_04918_ ), .B2(_04920_ ), .ZN(_00166_ ) );
XOR2_X1 _12548_ ( .A(_04876_ ), .B(_03315_ ), .Z(_04921_ ) );
NOR2_X1 _12549_ ( .A1(_04812_ ), .A2(_04921_ ), .ZN(_04922_ ) );
AND2_X1 _12550_ ( .A1(_03456_ ), .A2(\ID_EX_pc [12] ), .ZN(_04923_ ) );
XNOR2_X1 _12551_ ( .A(_04923_ ), .B(\ID_EX_pc [13] ), .ZN(_04924_ ) );
AOI211_X1 _12552_ ( .A(fanout_net_10 ), .B(_04922_ ), .C1(_04812_ ), .C2(_04924_ ), .ZN(_04925_ ) );
NAND2_X1 _12553_ ( .A1(_04697_ ), .A2(\mepc [13] ), .ZN(_04926_ ) );
NAND3_X1 _12554_ ( .A1(_04748_ ), .A2(\mtvec [13] ), .A3(_04746_ ), .ZN(_04927_ ) );
NAND4_X1 _12555_ ( .A1(_04836_ ), .A2(_03437_ ), .A3(\mycsreg.CSReg[3][13] ), .A4(_03438_ ), .ZN(_04928_ ) );
NAND4_X1 _12556_ ( .A1(_04835_ ), .A2(_04926_ ), .A3(_04927_ ), .A4(_04928_ ), .ZN(_04929_ ) );
AND4_X1 _12557_ ( .A1(\mycsreg.CSReg[0][13] ), .A2(_04749_ ), .A3(_03438_ ), .A4(_04702_ ), .ZN(_04930_ ) );
OAI21_X1 _12558_ ( .A(_03396_ ), .B1(_04929_ ), .B2(_04930_ ), .ZN(_04931_ ) );
NAND3_X1 _12559_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [13] ), .ZN(_04932_ ) );
AOI21_X1 _12560_ ( .A(_04856_ ), .B1(_04931_ ), .B2(_04932_ ), .ZN(_04933_ ) );
OAI21_X1 _12561_ ( .A(_04662_ ), .B1(_04925_ ), .B2(_04933_ ), .ZN(_04934_ ) );
NAND2_X1 _12562_ ( .A1(_03225_ ), .A2(fanout_net_8 ), .ZN(_04935_ ) );
OAI211_X1 _12563_ ( .A(_04935_ ), .B(_04756_ ), .C1(fanout_net_8 ), .C2(_04921_ ), .ZN(_04936_ ) );
AOI21_X1 _12564_ ( .A(_04663_ ), .B1(_04934_ ), .B2(_04936_ ), .ZN(_00167_ ) );
BUF_X4 _12565_ ( .A(_03248_ ), .Z(_04937_ ) );
INV_X1 _12566_ ( .A(\ID_EX_pc [12] ), .ZN(_04938_ ) );
XNOR2_X1 _12567_ ( .A(_03456_ ), .B(_04938_ ), .ZN(_04939_ ) );
XNOR2_X1 _12568_ ( .A(_03312_ ), .B(_04874_ ), .ZN(_04940_ ) );
MUX2_X1 _12569_ ( .A(_04939_ ), .B(_04940_ ), .S(_04656_ ), .Z(_04941_ ) );
OR2_X2 _12570_ ( .A1(_04941_ ), .A2(fanout_net_10 ), .ZN(_04942_ ) );
AND3_X1 _12571_ ( .A1(_04745_ ), .A2(\mtvec [12] ), .A3(_04691_ ), .ZN(_04943_ ) );
AND3_X1 _12572_ ( .A1(_04745_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_04699_ ), .ZN(_04944_ ) );
NOR2_X1 _12573_ ( .A1(_04943_ ), .A2(_04944_ ), .ZN(_04945_ ) );
NAND4_X1 _12574_ ( .A1(_04836_ ), .A2(_04684_ ), .A3(\mycsreg.CSReg[3][12] ), .A4(_04685_ ), .ZN(_04946_ ) );
NAND4_X1 _12575_ ( .A1(_03429_ ), .A2(_04684_ ), .A3(\mepc [12] ), .A4(_04685_ ), .ZN(_04947_ ) );
AND2_X1 _12576_ ( .A1(_04946_ ), .A2(_04947_ ), .ZN(_04948_ ) );
NAND4_X1 _12577_ ( .A1(_04945_ ), .A2(_04857_ ), .A3(_04858_ ), .A4(_04948_ ), .ZN(_04949_ ) );
NAND2_X1 _12578_ ( .A1(_04949_ ), .A2(_03396_ ), .ZN(_04950_ ) );
NAND3_X1 _12579_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [12] ), .ZN(_04951_ ) );
NAND2_X1 _12580_ ( .A1(_04950_ ), .A2(_04951_ ), .ZN(_04952_ ) );
OAI211_X1 _12581_ ( .A(_04942_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_04952_ ), .ZN(_04953_ ) );
OAI21_X1 _12582_ ( .A(_04755_ ), .B1(_04940_ ), .B2(fanout_net_8 ), .ZN(_04954_ ) );
AOI21_X1 _12583_ ( .A(_03251_ ), .B1(_03226_ ), .B2(_03223_ ), .ZN(_04955_ ) );
OR2_X1 _12584_ ( .A1(_04954_ ), .A2(_04955_ ), .ZN(_04956_ ) );
AOI21_X1 _12585_ ( .A(_04937_ ), .B1(_04953_ ), .B2(_04956_ ), .ZN(_00168_ ) );
AND2_X1 _12586_ ( .A1(_03454_ ), .A2(\ID_EX_pc [10] ), .ZN(_04957_ ) );
INV_X1 _12587_ ( .A(\ID_EX_pc [11] ), .ZN(_04958_ ) );
XNOR2_X1 _12588_ ( .A(_04957_ ), .B(_04958_ ), .ZN(_04959_ ) );
AOI21_X1 _12589_ ( .A(_04959_ ), .B1(_04653_ ), .B2(_04654_ ), .ZN(_04960_ ) );
AOI21_X1 _12590_ ( .A(_03306_ ), .B1(_03295_ ), .B2(_03302_ ), .ZN(_04961_ ) );
NOR2_X1 _12591_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_04962_ ) );
NOR3_X1 _12592_ ( .A1(_04961_ ), .A2(_03309_ ), .A3(_04962_ ), .ZN(_04963_ ) );
NOR2_X1 _12593_ ( .A1(_04963_ ), .A2(_03309_ ), .ZN(_04964_ ) );
XNOR2_X1 _12594_ ( .A(_04964_ ), .B(_03296_ ), .ZN(_04965_ ) );
INV_X1 _12595_ ( .A(_04965_ ), .ZN(_04966_ ) );
AOI211_X1 _12596_ ( .A(fanout_net_10 ), .B(_04960_ ), .C1(_04678_ ), .C2(_04966_ ), .ZN(_04967_ ) );
NAND4_X1 _12597_ ( .A1(_04737_ ), .A2(_03436_ ), .A3(\mycsreg.CSReg[3][11] ), .A4(_04740_ ), .ZN(_04968_ ) );
NAND4_X1 _12598_ ( .A1(_04860_ ), .A2(_03436_ ), .A3(\mepc [11] ), .A4(_04740_ ), .ZN(_04969_ ) );
AND2_X1 _12599_ ( .A1(_04968_ ), .A2(_04969_ ), .ZN(_04970_ ) );
NAND3_X1 _12600_ ( .A1(_04690_ ), .A2(\mtvec [11] ), .A3(_03411_ ), .ZN(_04971_ ) );
NAND3_X1 _12601_ ( .A1(_03406_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_03416_ ), .ZN(_04972_ ) );
AND2_X1 _12602_ ( .A1(_04971_ ), .A2(_04972_ ), .ZN(_04973_ ) );
NAND3_X1 _12603_ ( .A1(_04736_ ), .A2(_04970_ ), .A3(_04973_ ), .ZN(_04974_ ) );
NAND2_X1 _12604_ ( .A1(_04974_ ), .A2(_03396_ ), .ZN(_04975_ ) );
NAND3_X1 _12605_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [11] ), .ZN(_04976_ ) );
AOI21_X1 _12606_ ( .A(_04856_ ), .B1(_04975_ ), .B2(_04976_ ), .ZN(_04977_ ) );
OAI21_X1 _12607_ ( .A(_04662_ ), .B1(_04967_ ), .B2(_04977_ ), .ZN(_04978_ ) );
AOI21_X1 _12608_ ( .A(_02274_ ), .B1(_04966_ ), .B2(_03252_ ), .ZN(_04979_ ) );
AOI21_X1 _12609_ ( .A(_02993_ ), .B1(_02841_ ), .B2(_02986_ ), .ZN(_04980_ ) );
AND3_X1 _12610_ ( .A1(_02892_ ), .A2(_02913_ ), .A3(_02911_ ), .ZN(_04981_ ) );
NOR3_X1 _12611_ ( .A1(_04980_ ), .A2(_02996_ ), .A3(_04981_ ), .ZN(_04982_ ) );
NOR2_X1 _12612_ ( .A1(_04982_ ), .A2(_02996_ ), .ZN(_04983_ ) );
XNOR2_X1 _12613_ ( .A(_04983_ ), .B(_02938_ ), .ZN(_04984_ ) );
OAI21_X1 _12614_ ( .A(_04979_ ), .B1(_04984_ ), .B2(_04820_ ), .ZN(_04985_ ) );
AOI21_X1 _12615_ ( .A(_04937_ ), .B1(_04978_ ), .B2(_04985_ ), .ZN(_00169_ ) );
INV_X1 _12616_ ( .A(\ID_EX_pc [28] ), .ZN(_04986_ ) );
XNOR2_X1 _12617_ ( .A(_04674_ ), .B(_04986_ ), .ZN(_04987_ ) );
AOI21_X1 _12618_ ( .A(_04987_ ), .B1(_04653_ ), .B2(_04654_ ), .ZN(_04988_ ) );
XNOR2_X1 _12619_ ( .A(_03362_ ), .B(_03363_ ), .ZN(_04989_ ) );
AOI211_X1 _12620_ ( .A(fanout_net_10 ), .B(_04988_ ), .C1(_04873_ ), .C2(_04989_ ), .ZN(_04990_ ) );
AND4_X1 _12621_ ( .A1(\mycsreg.CSReg[3][28] ), .A2(_04683_ ), .A3(_04684_ ), .A4(_04685_ ), .ZN(_04991_ ) );
AOI21_X1 _12622_ ( .A(_04991_ ), .B1(_04687_ ), .B2(_04688_ ), .ZN(_04992_ ) );
NAND3_X1 _12623_ ( .A1(_04748_ ), .A2(\mtvec [28] ), .A3(_04746_ ), .ZN(_04993_ ) );
NAND2_X1 _12624_ ( .A1(_04781_ ), .A2(\mepc [28] ), .ZN(_04994_ ) );
NAND4_X1 _12625_ ( .A1(_04700_ ), .A2(_04701_ ), .A3(_04702_ ), .A4(\mycsreg.CSReg[0][28] ), .ZN(_04995_ ) );
NAND4_X1 _12626_ ( .A1(_04992_ ), .A2(_04993_ ), .A3(_04994_ ), .A4(_04995_ ), .ZN(_04996_ ) );
OAI21_X1 _12627_ ( .A(_04996_ ), .B1(_04711_ ), .B2(_04713_ ), .ZN(_04997_ ) );
NAND3_X1 _12628_ ( .A1(_04710_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_04715_ ), .ZN(_04998_ ) );
AOI21_X1 _12629_ ( .A(_04856_ ), .B1(_04997_ ), .B2(_04998_ ), .ZN(_04999_ ) );
OAI21_X1 _12630_ ( .A(_04662_ ), .B1(_04990_ ), .B2(_04999_ ), .ZN(_05000_ ) );
OAI21_X1 _12631_ ( .A(fanout_net_8 ), .B1(_03229_ ), .B2(_03129_ ), .ZN(_05001_ ) );
AOI21_X1 _12632_ ( .A(_04661_ ), .B1(_04989_ ), .B2(_03252_ ), .ZN(_05002_ ) );
NAND2_X1 _12633_ ( .A1(_05001_ ), .A2(_05002_ ), .ZN(_05003_ ) );
AOI21_X1 _12634_ ( .A(_04937_ ), .B1(_05000_ ), .B2(_05003_ ), .ZN(_00170_ ) );
BUF_X4 _12635_ ( .A(_02274_ ), .Z(_05004_ ) );
XNOR2_X1 _12636_ ( .A(_03454_ ), .B(\ID_EX_pc [10] ), .ZN(_05005_ ) );
AND2_X2 _12637_ ( .A1(_04811_ ), .A2(_05005_ ), .ZN(_05006_ ) );
XNOR2_X1 _12638_ ( .A(_04961_ ), .B(_03297_ ), .ZN(_05007_ ) );
INV_X1 _12639_ ( .A(_05007_ ), .ZN(_05008_ ) );
AOI211_X2 _12640_ ( .A(fanout_net_10 ), .B(_05006_ ), .C1(_04873_ ), .C2(_05008_ ), .ZN(_05009_ ) );
NAND2_X1 _12641_ ( .A1(_04696_ ), .A2(\mepc [10] ), .ZN(_05010_ ) );
NAND3_X1 _12642_ ( .A1(_04745_ ), .A2(\mtvec [10] ), .A3(_04691_ ), .ZN(_05011_ ) );
BUF_X2 _12643_ ( .A(_03435_ ), .Z(_05012_ ) );
BUF_X2 _12644_ ( .A(_04739_ ), .Z(_05013_ ) );
NAND4_X1 _12645_ ( .A1(_04683_ ), .A2(_05012_ ), .A3(\mycsreg.CSReg[3][10] ), .A4(_05013_ ), .ZN(_05014_ ) );
NAND4_X1 _12646_ ( .A1(_04834_ ), .A2(_05010_ ), .A3(_05011_ ), .A4(_05014_ ), .ZN(_05015_ ) );
AND4_X1 _12647_ ( .A1(\mycsreg.CSReg[0][10] ), .A2(_04699_ ), .A3(_05013_ ), .A4(_03403_ ), .ZN(_05016_ ) );
OAI21_X1 _12648_ ( .A(_03395_ ), .B1(_05015_ ), .B2(_05016_ ), .ZN(_05017_ ) );
NAND3_X1 _12649_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(\EX_LS_result_csreg_mem [10] ), .ZN(_05018_ ) );
AOI21_X1 _12650_ ( .A(_04856_ ), .B1(_05017_ ), .B2(_05018_ ), .ZN(_05019_ ) );
OAI21_X1 _12651_ ( .A(_05004_ ), .B1(_05009_ ), .B2(_05019_ ), .ZN(_05020_ ) );
AOI21_X1 _12652_ ( .A(_02274_ ), .B1(_05008_ ), .B2(_03252_ ), .ZN(_05021_ ) );
XNOR2_X1 _12653_ ( .A(_04980_ ), .B(_02914_ ), .ZN(_05022_ ) );
OAI21_X1 _12654_ ( .A(_05021_ ), .B1(_05022_ ), .B2(_04820_ ), .ZN(_05023_ ) );
AOI21_X1 _12655_ ( .A(_04937_ ), .B1(_05020_ ), .B2(_05023_ ), .ZN(_00171_ ) );
AND2_X1 _12656_ ( .A1(_03295_ ), .A2(_03298_ ), .ZN(_05024_ ) );
NOR2_X1 _12657_ ( .A1(_05024_ ), .A2(_03304_ ), .ZN(_05025_ ) );
XNOR2_X1 _12658_ ( .A(_05025_ ), .B(_03301_ ), .ZN(_05026_ ) );
AOI21_X2 _12659_ ( .A(fanout_net_10 ), .B1(_04873_ ), .B2(_05026_ ), .ZN(_05027_ ) );
XNOR2_X1 _12660_ ( .A(_03453_ ), .B(\ID_EX_pc [9] ), .ZN(_05028_ ) );
OAI21_X1 _12661_ ( .A(_05027_ ), .B1(_04678_ ), .B2(_05028_ ), .ZN(_05029_ ) );
NAND2_X1 _12662_ ( .A1(_04696_ ), .A2(\mepc [9] ), .ZN(_05030_ ) );
NAND3_X1 _12663_ ( .A1(_03405_ ), .A2(\mtvec [9] ), .A3(_03411_ ), .ZN(_05031_ ) );
NAND4_X1 _12664_ ( .A1(_03421_ ), .A2(_03435_ ), .A3(\mycsreg.CSReg[3][9] ), .A4(_04739_ ), .ZN(_05032_ ) );
NAND4_X1 _12665_ ( .A1(_04834_ ), .A2(_05030_ ), .A3(_05031_ ), .A4(_05032_ ), .ZN(_05033_ ) );
AND4_X1 _12666_ ( .A1(\mycsreg.CSReg[0][9] ), .A2(_03416_ ), .A3(_04739_ ), .A4(_03403_ ), .ZN(_05034_ ) );
OAI21_X1 _12667_ ( .A(_03395_ ), .B1(_05033_ ), .B2(_05034_ ), .ZN(_05035_ ) );
NAND3_X1 _12668_ ( .A1(_03384_ ), .A2(_03393_ ), .A3(\EX_LS_result_csreg_mem [9] ), .ZN(_05036_ ) );
AND2_X1 _12669_ ( .A1(_05035_ ), .A2(_05036_ ), .ZN(_05037_ ) );
INV_X1 _12670_ ( .A(_05037_ ), .ZN(_05038_ ) );
OAI211_X1 _12671_ ( .A(_05029_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_05038_ ), .ZN(_05039_ ) );
INV_X1 _12672_ ( .A(_02962_ ), .ZN(_05040_ ) );
AOI21_X1 _12673_ ( .A(_05040_ ), .B1(_02738_ ), .B2(_02839_ ), .ZN(_05041_ ) );
OR2_X1 _12674_ ( .A1(_05041_ ), .A2(_02990_ ), .ZN(_05042_ ) );
XNOR2_X1 _12675_ ( .A(_05042_ ), .B(_02985_ ), .ZN(_05043_ ) );
NAND2_X1 _12676_ ( .A1(_05043_ ), .A2(fanout_net_8 ), .ZN(_05044_ ) );
OAI211_X1 _12677_ ( .A(_05044_ ), .B(_04756_ ), .C1(fanout_net_8 ), .C2(_05026_ ), .ZN(_05045_ ) );
AOI21_X1 _12678_ ( .A(_04937_ ), .B1(_05039_ ), .B2(_05045_ ), .ZN(_00172_ ) );
XOR2_X1 _12679_ ( .A(_03295_ ), .B(_03298_ ), .Z(_05046_ ) );
AOI21_X1 _12680_ ( .A(fanout_net_10 ), .B1(_04657_ ), .B2(_05046_ ), .ZN(_05047_ ) );
XNOR2_X1 _12681_ ( .A(_03452_ ), .B(\ID_EX_pc [8] ), .ZN(_05048_ ) );
OAI21_X1 _12682_ ( .A(_05047_ ), .B1(_04678_ ), .B2(_05048_ ), .ZN(_05049_ ) );
NAND4_X1 _12683_ ( .A1(_03428_ ), .A2(_03435_ ), .A3(\mepc [8] ), .A4(_03400_ ), .ZN(_05050_ ) );
NAND4_X1 _12684_ ( .A1(_03421_ ), .A2(_03435_ ), .A3(\mycsreg.CSReg[3][8] ), .A4(_03400_ ), .ZN(_05051_ ) );
AND2_X1 _12685_ ( .A1(_05050_ ), .A2(_05051_ ), .ZN(_05052_ ) );
NAND3_X1 _12686_ ( .A1(_03404_ ), .A2(\mtvec [8] ), .A3(_03410_ ), .ZN(_05053_ ) );
NAND3_X1 _12687_ ( .A1(_03404_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_03415_ ), .ZN(_05054_ ) );
AND2_X1 _12688_ ( .A1(_05053_ ), .A2(_05054_ ), .ZN(_05055_ ) );
NAND3_X1 _12689_ ( .A1(_04736_ ), .A2(_05052_ ), .A3(_05055_ ), .ZN(_05056_ ) );
NAND2_X1 _12690_ ( .A1(_05056_ ), .A2(_03395_ ), .ZN(_05057_ ) );
NAND3_X1 _12691_ ( .A1(_03384_ ), .A2(_03393_ ), .A3(\EX_LS_result_csreg_mem [8] ), .ZN(_05058_ ) );
AND2_X1 _12692_ ( .A1(_05057_ ), .A2(_05058_ ), .ZN(_05059_ ) );
INV_X1 _12693_ ( .A(_05059_ ), .ZN(_05060_ ) );
OAI211_X1 _12694_ ( .A(_05049_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_05060_ ), .ZN(_05061_ ) );
XNOR2_X1 _12695_ ( .A(_02840_ ), .B(_05040_ ), .ZN(_05062_ ) );
NAND2_X1 _12696_ ( .A1(_05062_ ), .A2(fanout_net_8 ), .ZN(_05063_ ) );
BUF_X4 _12697_ ( .A(_04755_ ), .Z(_05064_ ) );
OAI211_X1 _12698_ ( .A(_05063_ ), .B(_05064_ ), .C1(fanout_net_8 ), .C2(_05046_ ), .ZN(_05065_ ) );
AOI21_X1 _12699_ ( .A(_04937_ ), .B1(_05061_ ), .B2(_05065_ ), .ZN(_00173_ ) );
NOR2_X1 _12700_ ( .A1(_03294_ ), .A2(_03292_ ), .ZN(_05066_ ) );
XNOR2_X1 _12701_ ( .A(_03291_ ), .B(_05066_ ), .ZN(_05067_ ) );
AOI21_X1 _12702_ ( .A(fanout_net_10 ), .B1(_04657_ ), .B2(_05067_ ), .ZN(_05068_ ) );
XNOR2_X1 _12703_ ( .A(_03451_ ), .B(\ID_EX_pc [7] ), .ZN(_05069_ ) );
OAI21_X1 _12704_ ( .A(_05068_ ), .B1(_04678_ ), .B2(_05069_ ), .ZN(_05070_ ) );
NAND3_X1 _12705_ ( .A1(_04690_ ), .A2(\mtvec [7] ), .A3(_04691_ ), .ZN(_05071_ ) );
NAND3_X1 _12706_ ( .A1(_04690_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_03416_ ), .ZN(_05072_ ) );
NAND4_X1 _12707_ ( .A1(_04737_ ), .A2(_03436_ ), .A3(\mycsreg.CSReg[3][7] ), .A4(_04740_ ), .ZN(_05073_ ) );
NAND4_X1 _12708_ ( .A1(_04860_ ), .A2(_03436_ ), .A3(\mepc [7] ), .A4(_04740_ ), .ZN(_05074_ ) );
AND4_X1 _12709_ ( .A1(_05071_ ), .A2(_05072_ ), .A3(_05073_ ), .A4(_05074_ ), .ZN(_05075_ ) );
OR2_X1 _12710_ ( .A1(_03394_ ), .A2(_05075_ ), .ZN(_05076_ ) );
NAND3_X1 _12711_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [7] ), .ZN(_05077_ ) );
AND2_X1 _12712_ ( .A1(_05076_ ), .A2(_05077_ ), .ZN(_05078_ ) );
INV_X1 _12713_ ( .A(_05078_ ), .ZN(_05079_ ) );
OAI211_X1 _12714_ ( .A(_05070_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_05079_ ), .ZN(_05080_ ) );
OAI21_X1 _12715_ ( .A(_02838_ ), .B1(_02831_ ), .B2(_02834_ ), .ZN(_05081_ ) );
NAND2_X1 _12716_ ( .A1(_05081_ ), .A2(_02682_ ), .ZN(_05082_ ) );
NAND2_X1 _12717_ ( .A1(_05082_ ), .A2(_02731_ ), .ZN(_05083_ ) );
NAND2_X1 _12718_ ( .A1(_05083_ ), .A2(_02736_ ), .ZN(_05084_ ) );
XNOR2_X1 _12719_ ( .A(_05084_ ), .B(_02708_ ), .ZN(_05085_ ) );
NAND2_X1 _12720_ ( .A1(_05085_ ), .A2(fanout_net_8 ), .ZN(_05086_ ) );
OAI211_X1 _12721_ ( .A(_05086_ ), .B(_05064_ ), .C1(fanout_net_8 ), .C2(_05067_ ), .ZN(_05087_ ) );
AOI21_X1 _12722_ ( .A(_04937_ ), .B1(_05080_ ), .B2(_05087_ ), .ZN(_00174_ ) );
XOR2_X1 _12723_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_05088_ ) );
XNOR2_X1 _12724_ ( .A(_03287_ ), .B(_05088_ ), .ZN(_05089_ ) );
NAND3_X1 _12725_ ( .A1(_04653_ ), .A2(_04654_ ), .A3(_05089_ ), .ZN(_05090_ ) );
XNOR2_X1 _12726_ ( .A(_03450_ ), .B(\ID_EX_pc [6] ), .ZN(_05091_ ) );
OAI211_X1 _12727_ ( .A(_05090_ ), .B(_04659_ ), .C1(_04873_ ), .C2(_05091_ ), .ZN(_05092_ ) );
AND3_X1 _12728_ ( .A1(_03406_ ), .A2(\mtvec [6] ), .A3(_03411_ ), .ZN(_05093_ ) );
AND3_X1 _12729_ ( .A1(_03406_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_03416_ ), .ZN(_05094_ ) );
NOR2_X1 _12730_ ( .A1(_05093_ ), .A2(_05094_ ), .ZN(_05095_ ) );
AND4_X1 _12731_ ( .A1(\mepc [6] ), .A2(_04860_ ), .A3(_03425_ ), .A4(_03426_ ), .ZN(_05096_ ) );
AOI21_X1 _12732_ ( .A(_05096_ ), .B1(_03429_ ), .B2(_03433_ ), .ZN(_05097_ ) );
NAND4_X1 _12733_ ( .A1(_04836_ ), .A2(_03437_ ), .A3(\mycsreg.CSReg[3][6] ), .A4(_03438_ ), .ZN(_05098_ ) );
NAND3_X1 _12734_ ( .A1(_05095_ ), .A2(_05097_ ), .A3(_05098_ ), .ZN(_05099_ ) );
NAND2_X1 _12735_ ( .A1(_03396_ ), .A2(_05099_ ), .ZN(_05100_ ) );
NAND3_X1 _12736_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [6] ), .ZN(_05101_ ) );
NAND2_X1 _12737_ ( .A1(_05100_ ), .A2(_05101_ ), .ZN(_05102_ ) );
OAI211_X1 _12738_ ( .A(_05092_ ), .B(_04729_ ), .C1(_04730_ ), .C2(_05102_ ), .ZN(_05103_ ) );
XNOR2_X1 _12739_ ( .A(_05082_ ), .B(_02731_ ), .ZN(_05104_ ) );
NAND2_X1 _12740_ ( .A1(_05104_ ), .A2(fanout_net_8 ), .ZN(_05105_ ) );
OAI211_X1 _12741_ ( .A(_05105_ ), .B(_05064_ ), .C1(fanout_net_8 ), .C2(_05089_ ), .ZN(_05106_ ) );
AOI21_X1 _12742_ ( .A(_04937_ ), .B1(_05103_ ), .B2(_05106_ ), .ZN(_00175_ ) );
NAND2_X1 _12743_ ( .A1(_03284_ ), .A2(_03285_ ), .ZN(_05107_ ) );
XNOR2_X1 _12744_ ( .A(\ID_EX_pc [5] ), .B(\ID_EX_imm [5] ), .ZN(_05108_ ) );
XNOR2_X1 _12745_ ( .A(_05107_ ), .B(_05108_ ), .ZN(_05109_ ) );
AOI21_X1 _12746_ ( .A(fanout_net_10 ), .B1(_04657_ ), .B2(_05109_ ), .ZN(_05110_ ) );
XNOR2_X1 _12747_ ( .A(_03449_ ), .B(\ID_EX_pc [5] ), .ZN(_05111_ ) );
OAI21_X1 _12748_ ( .A(_05110_ ), .B1(_04678_ ), .B2(_05111_ ), .ZN(_05112_ ) );
NAND2_X1 _12749_ ( .A1(_04697_ ), .A2(\mepc [5] ), .ZN(_05113_ ) );
NAND3_X1 _12750_ ( .A1(_04748_ ), .A2(\mtvec [5] ), .A3(_04746_ ), .ZN(_05114_ ) );
NAND4_X1 _12751_ ( .A1(_04836_ ), .A2(_03437_ ), .A3(\mycsreg.CSReg[3][5] ), .A4(_03438_ ), .ZN(_05115_ ) );
NAND4_X1 _12752_ ( .A1(_04835_ ), .A2(_05113_ ), .A3(_05114_ ), .A4(_05115_ ), .ZN(_05116_ ) );
AND4_X1 _12753_ ( .A1(\mycsreg.CSReg[0][5] ), .A2(_04749_ ), .A3(_03438_ ), .A4(_04702_ ), .ZN(_05117_ ) );
OAI21_X1 _12754_ ( .A(_03396_ ), .B1(_05116_ ), .B2(_05117_ ), .ZN(_05118_ ) );
NAND3_X1 _12755_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [5] ), .ZN(_05119_ ) );
AND2_X1 _12756_ ( .A1(_05118_ ), .A2(_05119_ ), .ZN(_05120_ ) );
INV_X1 _12757_ ( .A(_05120_ ), .ZN(_05121_ ) );
OAI211_X1 _12758_ ( .A(_05112_ ), .B(_02275_ ), .C1(_04659_ ), .C2(_05121_ ), .ZN(_05122_ ) );
OAI21_X1 _12759_ ( .A(_02837_ ), .B1(_02831_ ), .B2(_02834_ ), .ZN(_05123_ ) );
NAND2_X1 _12760_ ( .A1(_05123_ ), .A2(_02679_ ), .ZN(_05124_ ) );
XNOR2_X1 _12761_ ( .A(_05124_ ), .B(_02836_ ), .ZN(_05125_ ) );
NAND2_X1 _12762_ ( .A1(_05125_ ), .A2(fanout_net_9 ), .ZN(_05126_ ) );
OAI211_X1 _12763_ ( .A(_05126_ ), .B(_05064_ ), .C1(fanout_net_9 ), .C2(_05109_ ), .ZN(_05127_ ) );
AOI21_X1 _12764_ ( .A(_04937_ ), .B1(_05122_ ), .B2(_05127_ ), .ZN(_00176_ ) );
INV_X1 _12765_ ( .A(\ID_EX_pc [4] ), .ZN(_05128_ ) );
XNOR2_X1 _12766_ ( .A(_03448_ ), .B(_05128_ ), .ZN(_05129_ ) );
XOR2_X1 _12767_ ( .A(_03282_ ), .B(_03283_ ), .Z(_05130_ ) );
MUX2_X1 _12768_ ( .A(_05129_ ), .B(_05130_ ), .S(_04656_ ), .Z(_05131_ ) );
OR2_X2 _12769_ ( .A1(_05131_ ), .A2(fanout_net_10 ), .ZN(_05132_ ) );
INV_X1 _12770_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_05133_ ) );
AND4_X1 _12771_ ( .A1(_05133_ ), .A2(_04779_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_05134_ ) );
AND2_X1 _12772_ ( .A1(_04783_ ), .A2(_04860_ ), .ZN(_05135_ ) );
BUF_X4 _12773_ ( .A(_05135_ ), .Z(_05136_ ) );
AND2_X1 _12774_ ( .A1(_04697_ ), .A2(\mepc [4] ), .ZN(_05137_ ) );
AND3_X1 _12775_ ( .A1(_04748_ ), .A2(\mtvec [4] ), .A3(_04746_ ), .ZN(_05138_ ) );
AND4_X1 _12776_ ( .A1(\mycsreg.CSReg[3][4] ), .A2(_04836_ ), .A3(_04684_ ), .A4(_03438_ ), .ZN(_05139_ ) );
NOR4_X1 _12777_ ( .A1(_05136_ ), .A2(_05137_ ), .A3(_05138_ ), .A4(_05139_ ), .ZN(_05140_ ) );
AND3_X1 _12778_ ( .A1(_04839_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_04749_ ), .ZN(_05141_ ) );
AOI21_X1 _12779_ ( .A(_05141_ ), .B1(_04776_ ), .B2(_04789_ ), .ZN(_05142_ ) );
AOI21_X1 _12780_ ( .A(_05134_ ), .B1(_05140_ ), .B2(_05142_ ), .ZN(_05143_ ) );
OAI211_X1 _12781_ ( .A(_05132_ ), .B(_02275_ ), .C1(_04659_ ), .C2(_05143_ ), .ZN(_05144_ ) );
XNOR2_X1 _12782_ ( .A(_02835_ ), .B(_02837_ ), .ZN(_05145_ ) );
NAND2_X1 _12783_ ( .A1(_05145_ ), .A2(fanout_net_9 ), .ZN(_05146_ ) );
OAI211_X1 _12784_ ( .A(_05146_ ), .B(_05064_ ), .C1(fanout_net_9 ), .C2(_05130_ ), .ZN(_05147_ ) );
AOI21_X1 _12785_ ( .A(_04937_ ), .B1(_05144_ ), .B2(_05147_ ), .ZN(_00177_ ) );
BUF_X4 _12786_ ( .A(_03248_ ), .Z(_05148_ ) );
INV_X1 _12787_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_05149_ ) );
AND4_X1 _12788_ ( .A1(_05149_ ), .A2(_04778_ ), .A3(_04774_ ), .A4(_04773_ ), .ZN(_05150_ ) );
AND2_X1 _12789_ ( .A1(_04697_ ), .A2(\mepc [3] ), .ZN(_05151_ ) );
AND3_X1 _12790_ ( .A1(_04690_ ), .A2(\mtvec [3] ), .A3(_04691_ ), .ZN(_05152_ ) );
AND4_X1 _12791_ ( .A1(\mycsreg.CSReg[3][3] ), .A2(_04737_ ), .A3(_03436_ ), .A4(_04740_ ), .ZN(_05153_ ) );
NOR4_X1 _12792_ ( .A1(_05136_ ), .A2(_05151_ ), .A3(_05152_ ), .A4(_05153_ ), .ZN(_05154_ ) );
AND3_X1 _12793_ ( .A1(_04745_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_04749_ ), .ZN(_05155_ ) );
AOI21_X1 _12794_ ( .A(_05155_ ), .B1(_04776_ ), .B2(_04779_ ), .ZN(_05156_ ) );
AOI21_X1 _12795_ ( .A(_05150_ ), .B1(_05154_ ), .B2(_05156_ ), .ZN(_05157_ ) );
XOR2_X1 _12796_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .Z(_05158_ ) );
XNOR2_X1 _12797_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_imm [3] ), .ZN(_05159_ ) );
XNOR2_X1 _12798_ ( .A(_03279_ ), .B(_05159_ ), .ZN(_05160_ ) );
MUX2_X1 _12799_ ( .A(_05158_ ), .B(_05160_ ), .S(_04656_ ), .Z(_05161_ ) );
MUX2_X1 _12800_ ( .A(_05157_ ), .B(_05161_ ), .S(_03372_ ), .Z(_05162_ ) );
NAND2_X1 _12801_ ( .A1(_05162_ ), .A2(_04662_ ), .ZN(_05163_ ) );
OAI21_X1 _12802_ ( .A(_02832_ ), .B1(_02785_ ), .B2(_02808_ ), .ZN(_05164_ ) );
XOR2_X1 _12803_ ( .A(_05164_ ), .B(_02830_ ), .Z(_05165_ ) );
NAND2_X1 _12804_ ( .A1(_05165_ ), .A2(fanout_net_9 ), .ZN(_05166_ ) );
OAI211_X1 _12805_ ( .A(_05166_ ), .B(_05064_ ), .C1(fanout_net_9 ), .C2(_05160_ ), .ZN(_05167_ ) );
AOI21_X1 _12806_ ( .A(_05148_ ), .B1(_05163_ ), .B2(_05167_ ), .ZN(_00178_ ) );
XOR2_X1 _12807_ ( .A(_03275_ ), .B(_03276_ ), .Z(_05168_ ) );
MUX2_X1 _12808_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B(_05168_ ), .S(_04656_ ), .Z(_05169_ ) );
OR2_X2 _12809_ ( .A1(_05169_ ), .A2(fanout_net_10 ), .ZN(_05170_ ) );
AND3_X1 _12810_ ( .A1(_03405_ ), .A2(\mtvec [2] ), .A3(_03411_ ), .ZN(_05171_ ) );
AOI21_X1 _12811_ ( .A(_05171_ ), .B1(_04775_ ), .B2(_04778_ ), .ZN(_05172_ ) );
NAND2_X1 _12812_ ( .A1(_04696_ ), .A2(\mepc [2] ), .ZN(_05173_ ) );
NAND3_X1 _12813_ ( .A1(_03406_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_03416_ ), .ZN(_05174_ ) );
NAND2_X1 _12814_ ( .A1(_05173_ ), .A2(_05174_ ), .ZN(_05175_ ) );
AND4_X1 _12815_ ( .A1(\mycsreg.CSReg[3][2] ), .A2(_03421_ ), .A3(_03425_ ), .A4(_03426_ ), .ZN(_05176_ ) );
NOR3_X1 _12816_ ( .A1(_05175_ ), .A2(_04784_ ), .A3(_05176_ ), .ZN(_05177_ ) );
NAND2_X1 _12817_ ( .A1(_05172_ ), .A2(_05177_ ), .ZN(_05178_ ) );
INV_X1 _12818_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_05179_ ) );
NAND4_X1 _12819_ ( .A1(_04778_ ), .A2(_05179_ ), .A3(_04774_ ), .A4(_04773_ ), .ZN(_05180_ ) );
AND2_X1 _12820_ ( .A1(_05178_ ), .A2(_05180_ ), .ZN(_05181_ ) );
OAI211_X1 _12821_ ( .A(_05170_ ), .B(_02275_ ), .C1(_04659_ ), .C2(_05181_ ), .ZN(_05182_ ) );
XNOR2_X1 _12822_ ( .A(_02785_ ), .B(_02808_ ), .ZN(_05183_ ) );
NAND2_X1 _12823_ ( .A1(_05183_ ), .A2(fanout_net_9 ), .ZN(_05184_ ) );
OAI211_X1 _12824_ ( .A(_05184_ ), .B(_05064_ ), .C1(fanout_net_9 ), .C2(_05168_ ), .ZN(_05185_ ) );
AOI21_X1 _12825_ ( .A(_05148_ ), .B1(_05182_ ), .B2(_05185_ ), .ZN(_00179_ ) );
AOI21_X1 _12826_ ( .A(\ID_EX_pc [1] ), .B1(_04653_ ), .B2(_04654_ ), .ZN(_05186_ ) );
XOR2_X1 _12827_ ( .A(_03271_ ), .B(_03272_ ), .Z(_05187_ ) );
INV_X1 _12828_ ( .A(_05187_ ), .ZN(_05188_ ) );
AOI211_X1 _12829_ ( .A(fanout_net_10 ), .B(_05186_ ), .C1(_04873_ ), .C2(_05188_ ), .ZN(_05189_ ) );
AND3_X1 _12830_ ( .A1(_03404_ ), .A2(\mtvec [1] ), .A3(_03410_ ), .ZN(_05190_ ) );
INV_X1 _12831_ ( .A(_05190_ ), .ZN(_05191_ ) );
NAND2_X1 _12832_ ( .A1(_04781_ ), .A2(\mepc [1] ), .ZN(_05192_ ) );
BUF_X2 _12833_ ( .A(_04684_ ), .Z(_05193_ ) );
NAND4_X1 _12834_ ( .A1(_04738_ ), .A2(_05193_ ), .A3(\mycsreg.CSReg[3][1] ), .A4(_04701_ ), .ZN(_05194_ ) );
NAND4_X1 _12835_ ( .A1(_04700_ ), .A2(_04701_ ), .A3(_04702_ ), .A4(\mycsreg.CSReg[0][1] ), .ZN(_05195_ ) );
NAND4_X1 _12836_ ( .A1(_05191_ ), .A2(_05192_ ), .A3(_05194_ ), .A4(_05195_ ), .ZN(_05196_ ) );
OAI21_X1 _12837_ ( .A(_05196_ ), .B1(_04711_ ), .B2(_04713_ ), .ZN(_05197_ ) );
NAND3_X1 _12838_ ( .A1(_04710_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_04715_ ), .ZN(_05198_ ) );
AOI21_X1 _12839_ ( .A(_04856_ ), .B1(_05197_ ), .B2(_05198_ ), .ZN(_05199_ ) );
OAI21_X1 _12840_ ( .A(_05004_ ), .B1(_05189_ ), .B2(_05199_ ), .ZN(_05200_ ) );
AOI21_X1 _12841_ ( .A(_02274_ ), .B1(_05188_ ), .B2(_03252_ ), .ZN(_05201_ ) );
XOR2_X1 _12842_ ( .A(_02762_ ), .B(_02784_ ), .Z(_05202_ ) );
OAI21_X1 _12843_ ( .A(_05201_ ), .B1(_05202_ ), .B2(_04820_ ), .ZN(_05203_ ) );
AOI21_X1 _12844_ ( .A(_05148_ ), .B1(_05200_ ), .B2(_05203_ ), .ZN(_00180_ ) );
AOI21_X1 _12845_ ( .A(_03360_ ), .B1(_03346_ ), .B2(_03354_ ), .ZN(_05204_ ) );
NOR2_X1 _12846_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_05205_ ) );
NOR3_X1 _12847_ ( .A1(_05204_ ), .A2(_03356_ ), .A3(_05205_ ), .ZN(_05206_ ) );
NOR2_X1 _12848_ ( .A1(_05206_ ), .A2(_03356_ ), .ZN(_05207_ ) );
XNOR2_X1 _12849_ ( .A(_05207_ ), .B(_03347_ ), .ZN(_05208_ ) );
NOR2_X1 _12850_ ( .A1(_04812_ ), .A2(_05208_ ), .ZN(_05209_ ) );
NAND3_X1 _12851_ ( .A1(_04667_ ), .A2(\ID_EX_pc [26] ), .A3(_04670_ ), .ZN(_05210_ ) );
XNOR2_X1 _12852_ ( .A(_05210_ ), .B(_04672_ ), .ZN(_05211_ ) );
AOI211_X1 _12853_ ( .A(fanout_net_10 ), .B(_05209_ ), .C1(_04812_ ), .C2(_05211_ ), .ZN(_05212_ ) );
NAND2_X1 _12854_ ( .A1(_04696_ ), .A2(\mepc [27] ), .ZN(_05213_ ) );
NAND3_X1 _12855_ ( .A1(_04745_ ), .A2(\mtvec [27] ), .A3(_04691_ ), .ZN(_05214_ ) );
NAND4_X1 _12856_ ( .A1(_04683_ ), .A2(_05012_ ), .A3(\mycsreg.CSReg[3][27] ), .A4(_05013_ ), .ZN(_05215_ ) );
NAND4_X1 _12857_ ( .A1(_04835_ ), .A2(_05213_ ), .A3(_05214_ ), .A4(_05215_ ), .ZN(_05216_ ) );
AND4_X1 _12858_ ( .A1(\mycsreg.CSReg[0][27] ), .A2(_04699_ ), .A3(_04685_ ), .A4(_04702_ ), .ZN(_05217_ ) );
OAI21_X1 _12859_ ( .A(_03396_ ), .B1(_05216_ ), .B2(_05217_ ), .ZN(_05218_ ) );
NAND3_X1 _12860_ ( .A1(_04710_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_04715_ ), .ZN(_05219_ ) );
AOI21_X1 _12861_ ( .A(_04856_ ), .B1(_05218_ ), .B2(_05219_ ), .ZN(_05220_ ) );
OAI21_X1 _12862_ ( .A(_05004_ ), .B1(_05212_ ), .B2(_05220_ ), .ZN(_05221_ ) );
NAND2_X1 _12863_ ( .A1(_03233_ ), .A2(fanout_net_9 ), .ZN(_05222_ ) );
OAI211_X1 _12864_ ( .A(_05222_ ), .B(_05064_ ), .C1(fanout_net_9 ), .C2(_05208_ ), .ZN(_05223_ ) );
AOI21_X1 _12865_ ( .A(_05148_ ), .B1(_05221_ ), .B2(_05223_ ), .ZN(_00181_ ) );
CLKBUF_X2 _12866_ ( .A(_02272_ ), .Z(_05224_ ) );
XOR2_X1 _12867_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05225_ ) );
NAND2_X1 _12868_ ( .A1(_05225_ ), .A2(\myexu.pc_jump_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_05226_ ) );
XNOR2_X1 _12869_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .ZN(_05227_ ) );
AOI21_X1 _12870_ ( .A(fanout_net_10 ), .B1(_04657_ ), .B2(_05227_ ), .ZN(_05228_ ) );
OAI21_X1 _12871_ ( .A(_05228_ ), .B1(\ID_EX_pc [0] ), .B2(_04657_ ), .ZN(_05229_ ) );
AND4_X1 _12872_ ( .A1(\mepc [0] ), .A2(_04860_ ), .A3(_03425_ ), .A4(_03426_ ), .ZN(_05230_ ) );
AND4_X1 _12873_ ( .A1(\mycsreg.CSReg[3][0] ), .A2(_03421_ ), .A3(_03425_ ), .A4(_03426_ ), .ZN(_05231_ ) );
NOR3_X1 _12874_ ( .A1(_04735_ ), .A2(_05230_ ), .A3(_05231_ ), .ZN(_05232_ ) );
NAND3_X1 _12875_ ( .A1(_03406_ ), .A2(\mtvec [0] ), .A3(_03411_ ), .ZN(_05233_ ) );
NAND3_X1 _12876_ ( .A1(_03406_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_03416_ ), .ZN(_05234_ ) );
AND2_X1 _12877_ ( .A1(_05233_ ), .A2(_05234_ ), .ZN(_05235_ ) );
AOI21_X1 _12878_ ( .A(_03394_ ), .B1(_05232_ ), .B2(_05235_ ), .ZN(_05236_ ) );
AND3_X1 _12879_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(\EX_LS_result_csreg_mem [0] ), .ZN(_05237_ ) );
OAI21_X1 _12880_ ( .A(fanout_net_10 ), .B1(_05236_ ), .B2(_05237_ ), .ZN(_05238_ ) );
AND2_X1 _12881_ ( .A1(_05238_ ), .A2(_02273_ ), .ZN(_05239_ ) );
AOI221_X1 _12882_ ( .A(_03248_ ), .B1(_05224_ ), .B2(_05226_ ), .C1(_05229_ ), .C2(_05239_ ), .ZN(_00182_ ) );
XNOR2_X1 _12883_ ( .A(_04671_ ), .B(\ID_EX_pc [26] ), .ZN(_05240_ ) );
AOI21_X1 _12884_ ( .A(_05240_ ), .B1(_04653_ ), .B2(_04654_ ), .ZN(_05241_ ) );
XNOR2_X1 _12885_ ( .A(_05204_ ), .B(_03348_ ), .ZN(_05242_ ) );
INV_X1 _12886_ ( .A(_05242_ ), .ZN(_05243_ ) );
AOI211_X1 _12887_ ( .A(fanout_net_10 ), .B(_05241_ ), .C1(_04873_ ), .C2(_05243_ ), .ZN(_05244_ ) );
NAND2_X1 _12888_ ( .A1(_04781_ ), .A2(\mepc [26] ), .ZN(_05245_ ) );
NAND3_X1 _12889_ ( .A1(_04839_ ), .A2(\mtvec [26] ), .A3(_04746_ ), .ZN(_05246_ ) );
NAND4_X1 _12890_ ( .A1(_04738_ ), .A2(_05193_ ), .A3(\mycsreg.CSReg[3][26] ), .A4(_04701_ ), .ZN(_05247_ ) );
NAND4_X1 _12891_ ( .A1(_04700_ ), .A2(_04701_ ), .A3(_04702_ ), .A4(\mycsreg.CSReg[0][26] ), .ZN(_05248_ ) );
NAND4_X1 _12892_ ( .A1(_05245_ ), .A2(_05246_ ), .A3(_05247_ ), .A4(_05248_ ), .ZN(_05249_ ) );
OAI21_X1 _12893_ ( .A(_05249_ ), .B1(_04711_ ), .B2(_04713_ ), .ZN(_05250_ ) );
NAND3_X1 _12894_ ( .A1(_04710_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_04715_ ), .ZN(_05251_ ) );
AOI21_X1 _12895_ ( .A(_04856_ ), .B1(_05250_ ), .B2(_05251_ ), .ZN(_05252_ ) );
OAI21_X1 _12896_ ( .A(_05004_ ), .B1(_05244_ ), .B2(_05252_ ), .ZN(_05253_ ) );
AOI21_X1 _12897_ ( .A(_02274_ ), .B1(_05243_ ), .B2(_03252_ ), .ZN(_05254_ ) );
OAI21_X1 _12898_ ( .A(_05254_ ), .B1(_03235_ ), .B2(_04820_ ), .ZN(_05255_ ) );
AOI21_X1 _12899_ ( .A(_05148_ ), .B1(_05253_ ), .B2(_05255_ ), .ZN(_00183_ ) );
NAND2_X1 _12900_ ( .A1(_03346_ ), .A2(_03350_ ), .ZN(_05256_ ) );
AND2_X1 _12901_ ( .A1(_05256_ ), .A2(_03358_ ), .ZN(_05257_ ) );
XNOR2_X1 _12902_ ( .A(_05257_ ), .B(_03353_ ), .ZN(_05258_ ) );
NOR2_X1 _12903_ ( .A1(_04812_ ), .A2(_05258_ ), .ZN(_05259_ ) );
AND3_X1 _12904_ ( .A1(_04669_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05260_ ) );
AND2_X1 _12905_ ( .A1(_04667_ ), .A2(_05260_ ), .ZN(_05261_ ) );
NAND3_X1 _12906_ ( .A1(_05261_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05262_ ) );
INV_X1 _12907_ ( .A(\ID_EX_pc [24] ), .ZN(_05263_ ) );
NOR2_X1 _12908_ ( .A1(_05262_ ), .A2(_05263_ ), .ZN(_05264_ ) );
XNOR2_X1 _12909_ ( .A(_05264_ ), .B(\ID_EX_pc [25] ), .ZN(_05265_ ) );
AOI211_X1 _12910_ ( .A(fanout_net_10 ), .B(_05259_ ), .C1(_04812_ ), .C2(_05265_ ), .ZN(_05266_ ) );
NAND4_X1 _12911_ ( .A1(_03420_ ), .A2(_03424_ ), .A3(\mycsreg.CSReg[3][25] ), .A4(_03400_ ), .ZN(_05267_ ) );
NAND4_X1 _12912_ ( .A1(_03428_ ), .A2(_03424_ ), .A3(\mepc [25] ), .A4(_03400_ ), .ZN(_05268_ ) );
AND2_X1 _12913_ ( .A1(_05267_ ), .A2(_05268_ ), .ZN(_05269_ ) );
NAND3_X1 _12914_ ( .A1(_03405_ ), .A2(\mtvec [25] ), .A3(_03411_ ), .ZN(_05270_ ) );
NAND3_X1 _12915_ ( .A1(_03405_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_03415_ ), .ZN(_05271_ ) );
NAND3_X1 _12916_ ( .A1(_05269_ ), .A2(_05270_ ), .A3(_05271_ ), .ZN(_05272_ ) );
AOI21_X1 _12917_ ( .A(_05272_ ), .B1(_04775_ ), .B2(_04778_ ), .ZN(_05273_ ) );
INV_X1 _12918_ ( .A(\EX_LS_result_csreg_mem [25] ), .ZN(_05274_ ) );
AND4_X1 _12919_ ( .A1(_05274_ ), .A2(_04777_ ), .A3(_04774_ ), .A4(_04773_ ), .ZN(_05275_ ) );
NOR3_X1 _12920_ ( .A1(_05273_ ), .A2(_04856_ ), .A3(_05275_ ), .ZN(_05276_ ) );
OAI21_X1 _12921_ ( .A(_05004_ ), .B1(_05266_ ), .B2(_05276_ ), .ZN(_05277_ ) );
NAND2_X1 _12922_ ( .A1(_03237_ ), .A2(fanout_net_9 ), .ZN(_05278_ ) );
OAI211_X1 _12923_ ( .A(_05278_ ), .B(_05064_ ), .C1(fanout_net_9 ), .C2(_05258_ ), .ZN(_05279_ ) );
AOI21_X1 _12924_ ( .A(_05148_ ), .B1(_05277_ ), .B2(_05279_ ), .ZN(_00184_ ) );
AND3_X1 _12925_ ( .A1(_04690_ ), .A2(\mtvec [24] ), .A3(_04691_ ), .ZN(_05280_ ) );
AND3_X1 _12926_ ( .A1(_04690_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_04699_ ), .ZN(_05281_ ) );
NOR2_X1 _12927_ ( .A1(_05280_ ), .A2(_05281_ ), .ZN(_05282_ ) );
NAND4_X1 _12928_ ( .A1(_04683_ ), .A2(_05012_ ), .A3(\mycsreg.CSReg[3][24] ), .A4(_05013_ ), .ZN(_05283_ ) );
NAND4_X1 _12929_ ( .A1(_03429_ ), .A2(_05012_ ), .A3(\mepc [24] ), .A4(_05013_ ), .ZN(_05284_ ) );
AND2_X1 _12930_ ( .A1(_05283_ ), .A2(_05284_ ), .ZN(_05285_ ) );
NAND4_X1 _12931_ ( .A1(_05282_ ), .A2(_04857_ ), .A3(_04858_ ), .A4(_05285_ ), .ZN(_05286_ ) );
NAND2_X1 _12932_ ( .A1(_05286_ ), .A2(_03396_ ), .ZN(_05287_ ) );
NAND3_X1 _12933_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [24] ), .ZN(_05288_ ) );
NAND2_X1 _12934_ ( .A1(_05287_ ), .A2(_05288_ ), .ZN(_05289_ ) );
XNOR2_X1 _12935_ ( .A(_05262_ ), .B(\ID_EX_pc [24] ), .ZN(_05290_ ) );
XOR2_X1 _12936_ ( .A(_03346_ ), .B(_03350_ ), .Z(_05291_ ) );
MUX2_X1 _12937_ ( .A(_05290_ ), .B(_05291_ ), .S(_04656_ ), .Z(_05292_ ) );
MUX2_X1 _12938_ ( .A(_05289_ ), .B(_05292_ ), .S(_03372_ ), .Z(_05293_ ) );
NAND2_X1 _12939_ ( .A1(_05293_ ), .A2(_04662_ ), .ZN(_05294_ ) );
OR2_X1 _12940_ ( .A1(_03238_ ), .A2(_03251_ ), .ZN(_05295_ ) );
OAI211_X1 _12941_ ( .A(_05295_ ), .B(_05064_ ), .C1(fanout_net_9 ), .C2(_05291_ ), .ZN(_05296_ ) );
AOI21_X1 _12942_ ( .A(_05148_ ), .B1(_05294_ ), .B2(_05296_ ), .ZN(_00185_ ) );
AOI21_X1 _12943_ ( .A(_03253_ ), .B1(_04724_ ), .B2(_03337_ ), .ZN(_05297_ ) );
OAI21_X1 _12944_ ( .A(_03341_ ), .B1(_05297_ ), .B2(_03343_ ), .ZN(_05298_ ) );
XNOR2_X1 _12945_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .ZN(_05299_ ) );
NOR2_X1 _12946_ ( .A1(_05298_ ), .A2(_05299_ ), .ZN(_05300_ ) );
NOR2_X1 _12947_ ( .A1(_05300_ ), .A2(_03327_ ), .ZN(_05301_ ) );
XNOR2_X1 _12948_ ( .A(_05301_ ), .B(_03257_ ), .ZN(_05302_ ) );
NOR2_X1 _12949_ ( .A1(_04812_ ), .A2(_05302_ ), .ZN(_05303_ ) );
NAND3_X1 _12950_ ( .A1(_04667_ ), .A2(\ID_EX_pc [22] ), .A3(_05260_ ), .ZN(_05304_ ) );
XNOR2_X1 _12951_ ( .A(_05304_ ), .B(_03329_ ), .ZN(_05305_ ) );
AOI211_X1 _12952_ ( .A(fanout_net_10 ), .B(_05303_ ), .C1(_04812_ ), .C2(_05305_ ), .ZN(_05306_ ) );
NAND4_X1 _12953_ ( .A1(_04737_ ), .A2(_03425_ ), .A3(\mycsreg.CSReg[3][23] ), .A4(_03426_ ), .ZN(_05307_ ) );
NAND4_X1 _12954_ ( .A1(_04860_ ), .A2(_03425_ ), .A3(\mepc [23] ), .A4(_03426_ ), .ZN(_05308_ ) );
AND2_X1 _12955_ ( .A1(_05307_ ), .A2(_05308_ ), .ZN(_05309_ ) );
NAND3_X1 _12956_ ( .A1(_04690_ ), .A2(\mtvec [23] ), .A3(_04691_ ), .ZN(_05310_ ) );
NAND3_X1 _12957_ ( .A1(_04690_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_04699_ ), .ZN(_05311_ ) );
NAND3_X1 _12958_ ( .A1(_05309_ ), .A2(_05310_ ), .A3(_05311_ ), .ZN(_05312_ ) );
AOI21_X1 _12959_ ( .A(_05312_ ), .B1(_04776_ ), .B2(_04779_ ), .ZN(_05313_ ) );
INV_X1 _12960_ ( .A(\EX_LS_result_csreg_mem [23] ), .ZN(_05314_ ) );
AND4_X1 _12961_ ( .A1(_05314_ ), .A2(_04778_ ), .A3(_04774_ ), .A4(_04773_ ), .ZN(_05315_ ) );
NOR3_X1 _12962_ ( .A1(_05313_ ), .A2(_03372_ ), .A3(_05315_ ), .ZN(_05316_ ) );
OAI21_X1 _12963_ ( .A(_05004_ ), .B1(_05306_ ), .B2(_05316_ ), .ZN(_05317_ ) );
OR3_X1 _12964_ ( .A1(_03243_ ), .A2(_03251_ ), .A3(_03244_ ), .ZN(_05318_ ) );
CLKBUF_X2 _12965_ ( .A(_02272_ ), .Z(_05319_ ) );
BUF_X4 _12966_ ( .A(_05319_ ), .Z(_05320_ ) );
OAI211_X1 _12967_ ( .A(_05318_ ), .B(_05320_ ), .C1(fanout_net_9 ), .C2(_05302_ ), .ZN(_05321_ ) );
AOI21_X1 _12968_ ( .A(_05148_ ), .B1(_05317_ ), .B2(_05321_ ), .ZN(_00186_ ) );
XNOR2_X1 _12969_ ( .A(_05261_ ), .B(\ID_EX_pc [22] ), .ZN(_05322_ ) );
AND2_X2 _12970_ ( .A1(_04811_ ), .A2(_05322_ ), .ZN(_05323_ ) );
XNOR2_X1 _12971_ ( .A(_05298_ ), .B(_03258_ ), .ZN(_05324_ ) );
INV_X1 _12972_ ( .A(_05324_ ), .ZN(_05325_ ) );
AOI211_X2 _12973_ ( .A(fanout_net_10 ), .B(_05323_ ), .C1(_04873_ ), .C2(_05325_ ), .ZN(_05326_ ) );
NAND4_X1 _12974_ ( .A1(_03421_ ), .A2(_03435_ ), .A3(\mycsreg.CSReg[3][22] ), .A4(_04739_ ), .ZN(_05327_ ) );
NAND4_X1 _12975_ ( .A1(_04860_ ), .A2(_03435_ ), .A3(\mepc [22] ), .A4(_04739_ ), .ZN(_05328_ ) );
AND2_X1 _12976_ ( .A1(_05327_ ), .A2(_05328_ ), .ZN(_05329_ ) );
NAND3_X1 _12977_ ( .A1(_03405_ ), .A2(\mtvec [22] ), .A3(_03411_ ), .ZN(_05330_ ) );
NAND3_X1 _12978_ ( .A1(_03405_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_03416_ ), .ZN(_05331_ ) );
AND2_X1 _12979_ ( .A1(_05330_ ), .A2(_05331_ ), .ZN(_05332_ ) );
NAND3_X1 _12980_ ( .A1(_04736_ ), .A2(_05329_ ), .A3(_05332_ ), .ZN(_05333_ ) );
NAND2_X1 _12981_ ( .A1(_05333_ ), .A2(_03395_ ), .ZN(_05334_ ) );
NAND3_X1 _12982_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(\EX_LS_result_csreg_mem [22] ), .ZN(_05335_ ) );
AOI21_X1 _12983_ ( .A(_04856_ ), .B1(_05334_ ), .B2(_05335_ ), .ZN(_05336_ ) );
OAI21_X1 _12984_ ( .A(_05004_ ), .B1(_05326_ ), .B2(_05336_ ), .ZN(_05337_ ) );
AOI21_X1 _12985_ ( .A(_02274_ ), .B1(_05325_ ), .B2(_03252_ ), .ZN(_05338_ ) );
AND2_X1 _12986_ ( .A1(_03246_ ), .A2(_03241_ ), .ZN(_05339_ ) );
OAI21_X1 _12987_ ( .A(_05338_ ), .B1(_05339_ ), .B2(_04820_ ), .ZN(_05340_ ) );
AOI21_X1 _12988_ ( .A(_05148_ ), .B1(_05337_ ), .B2(_05340_ ), .ZN(_00187_ ) );
NOR2_X1 _12989_ ( .A1(_05297_ ), .A2(_03342_ ), .ZN(_05341_ ) );
NOR2_X1 _12990_ ( .A1(_03254_ ), .A2(_03255_ ), .ZN(_05342_ ) );
XNOR2_X1 _12991_ ( .A(_05341_ ), .B(_05342_ ), .ZN(_05343_ ) );
AOI21_X1 _12992_ ( .A(fanout_net_10 ), .B1(_04657_ ), .B2(_05343_ ), .ZN(_05344_ ) );
INV_X1 _12993_ ( .A(\ID_EX_pc [20] ), .ZN(_05345_ ) );
NOR2_X1 _12994_ ( .A1(_04722_ ), .A2(_05345_ ), .ZN(_05346_ ) );
XNOR2_X1 _12995_ ( .A(_05346_ ), .B(\ID_EX_pc [21] ), .ZN(_05347_ ) );
OAI21_X1 _12996_ ( .A(_05344_ ), .B1(_04678_ ), .B2(_05347_ ), .ZN(_05348_ ) );
NAND2_X1 _12997_ ( .A1(_04696_ ), .A2(\mepc [21] ), .ZN(_05349_ ) );
NAND3_X1 _12998_ ( .A1(_04745_ ), .A2(\mtvec [21] ), .A3(_04691_ ), .ZN(_05350_ ) );
NAND4_X1 _12999_ ( .A1(_04683_ ), .A2(_05012_ ), .A3(\mycsreg.CSReg[3][21] ), .A4(_05013_ ), .ZN(_05351_ ) );
NAND4_X1 _13000_ ( .A1(_04835_ ), .A2(_05349_ ), .A3(_05350_ ), .A4(_05351_ ), .ZN(_05352_ ) );
AND4_X1 _13001_ ( .A1(\mycsreg.CSReg[0][21] ), .A2(_04699_ ), .A3(_04685_ ), .A4(_04702_ ), .ZN(_05353_ ) );
OAI21_X1 _13002_ ( .A(_03395_ ), .B1(_05352_ ), .B2(_05353_ ), .ZN(_05354_ ) );
NAND3_X1 _13003_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [21] ), .ZN(_05355_ ) );
AND2_X1 _13004_ ( .A1(_05354_ ), .A2(_05355_ ), .ZN(_05356_ ) );
INV_X1 _13005_ ( .A(_05356_ ), .ZN(_05357_ ) );
OAI211_X1 _13006_ ( .A(_05348_ ), .B(_02275_ ), .C1(_04659_ ), .C2(_05357_ ), .ZN(_05358_ ) );
NAND2_X1 _13007_ ( .A1(_03198_ ), .A2(fanout_net_9 ), .ZN(_05359_ ) );
OAI211_X1 _13008_ ( .A(_05359_ ), .B(_05320_ ), .C1(fanout_net_9 ), .C2(_05343_ ), .ZN(_05360_ ) );
AOI21_X1 _13009_ ( .A(_05148_ ), .B1(_05358_ ), .B2(_05360_ ), .ZN(_00188_ ) );
INV_X1 _13010_ ( .A(\ID_EX_pc [30] ), .ZN(_05361_ ) );
NOR2_X1 _13011_ ( .A1(_03465_ ), .A2(_05361_ ), .ZN(_05362_ ) );
XNOR2_X1 _13012_ ( .A(_05362_ ), .B(\ID_EX_pc [31] ), .ZN(_05363_ ) );
AND2_X2 _13013_ ( .A1(_04811_ ), .A2(_05363_ ), .ZN(_05364_ ) );
NOR2_X1 _13014_ ( .A1(_03368_ ), .A2(_03369_ ), .ZN(_05365_ ) );
AND2_X1 _13015_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_05366_ ) );
NOR2_X1 _13016_ ( .A1(_05365_ ), .A2(_05366_ ), .ZN(_05367_ ) );
XNOR2_X1 _13017_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_05368_ ) );
XOR2_X1 _13018_ ( .A(_05367_ ), .B(_05368_ ), .Z(_05369_ ) );
INV_X1 _13019_ ( .A(_05369_ ), .ZN(_05370_ ) );
AOI211_X2 _13020_ ( .A(fanout_net_10 ), .B(_05364_ ), .C1(_04873_ ), .C2(_05370_ ), .ZN(_05371_ ) );
NAND2_X1 _13021_ ( .A1(_04781_ ), .A2(\mepc [31] ), .ZN(_05372_ ) );
NAND3_X1 _13022_ ( .A1(_04839_ ), .A2(\mtvec [31] ), .A3(_04746_ ), .ZN(_05373_ ) );
NAND4_X1 _13023_ ( .A1(_04738_ ), .A2(_05193_ ), .A3(\mycsreg.CSReg[3][31] ), .A4(_04741_ ), .ZN(_05374_ ) );
NAND4_X1 _13024_ ( .A1(_04700_ ), .A2(_04741_ ), .A3(_04702_ ), .A4(\mycsreg.CSReg[0][31] ), .ZN(_05375_ ) );
NAND4_X1 _13025_ ( .A1(_05372_ ), .A2(_05373_ ), .A3(_05374_ ), .A4(_05375_ ), .ZN(_05376_ ) );
BUF_X4 _13026_ ( .A(_04712_ ), .Z(_05377_ ) );
OAI21_X1 _13027_ ( .A(_05376_ ), .B1(_04711_ ), .B2(_05377_ ), .ZN(_05378_ ) );
NAND3_X1 _13028_ ( .A1(_04710_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_04715_ ), .ZN(_05379_ ) );
AOI21_X1 _13029_ ( .A(_03372_ ), .B1(_05378_ ), .B2(_05379_ ), .ZN(_05380_ ) );
OAI21_X1 _13030_ ( .A(_02275_ ), .B1(_05371_ ), .B2(_05380_ ), .ZN(_05381_ ) );
MUX2_X1 _13031_ ( .A(_05370_ ), .B(_03187_ ), .S(fanout_net_9 ), .Z(_05382_ ) );
OAI211_X1 _13032_ ( .A(_05381_ ), .B(_03247_ ), .C1(_04662_ ), .C2(_05382_ ), .ZN(_00189_ ) );
AND2_X1 _13033_ ( .A1(_03247_ ), .A2(\ID_EX_pc [31] ), .ZN(_00190_ ) );
NOR3_X1 _13034_ ( .A1(_05361_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00191_ ) );
INV_X1 _13035_ ( .A(\ID_EX_pc [21] ), .ZN(_05383_ ) );
NOR3_X1 _13036_ ( .A1(_05383_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00192_ ) );
NOR3_X1 _13037_ ( .A1(_05345_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00193_ ) );
NOR3_X1 _13038_ ( .A1(_03332_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00194_ ) );
INV_X1 _13039_ ( .A(\ID_EX_pc [18] ), .ZN(_05384_ ) );
NOR3_X1 _13040_ ( .A1(_05384_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00195_ ) );
NOR3_X1 _13041_ ( .A1(_03335_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00196_ ) );
NOR3_X1 _13042_ ( .A1(_04823_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00197_ ) );
NOR3_X1 _13043_ ( .A1(_04884_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00198_ ) );
NOR3_X1 _13044_ ( .A1(_04904_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00199_ ) );
AND2_X1 _13045_ ( .A1(_03247_ ), .A2(\ID_EX_pc [13] ), .ZN(_00200_ ) );
NOR3_X1 _13046_ ( .A1(_04938_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00201_ ) );
NOR3_X1 _13047_ ( .A1(_03366_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00202_ ) );
NOR3_X1 _13048_ ( .A1(_04958_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00203_ ) );
INV_X1 _13049_ ( .A(\ID_EX_pc [10] ), .ZN(_05385_ ) );
NOR3_X1 _13050_ ( .A1(_05385_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00204_ ) );
INV_X1 _13051_ ( .A(\ID_EX_pc [9] ), .ZN(_05386_ ) );
NOR3_X1 _13052_ ( .A1(_05386_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00205_ ) );
INV_X1 _13053_ ( .A(\ID_EX_pc [8] ), .ZN(_05387_ ) );
NOR3_X1 _13054_ ( .A1(_05387_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00206_ ) );
AND2_X1 _13055_ ( .A1(_03247_ ), .A2(\ID_EX_pc [7] ), .ZN(_00207_ ) );
INV_X1 _13056_ ( .A(\ID_EX_pc [6] ), .ZN(_05388_ ) );
NOR3_X1 _13057_ ( .A1(_05388_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00208_ ) );
AND2_X1 _13058_ ( .A1(_03247_ ), .A2(\ID_EX_pc [5] ), .ZN(_00209_ ) );
NOR3_X1 _13059_ ( .A1(_05128_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00210_ ) );
INV_X1 _13060_ ( .A(\ID_EX_pc [3] ), .ZN(_05389_ ) );
NOR3_X1 _13061_ ( .A1(_05389_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00211_ ) );
AND2_X1 _13062_ ( .A1(_02279_ ), .A2(\ID_EX_pc [2] ), .ZN(_00212_ ) );
NOR3_X1 _13063_ ( .A1(_04986_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00213_ ) );
NOR3_X1 _13064_ ( .A1(_03274_ ), .A2(fanout_net_4 ), .A3(fanout_net_20 ), .ZN(_00214_ ) );
AND2_X1 _13065_ ( .A1(_02279_ ), .A2(\ID_EX_pc [0] ), .ZN(_00215_ ) );
NOR3_X1 _13066_ ( .A1(_04672_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00216_ ) );
NOR3_X1 _13067_ ( .A1(_04673_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00217_ ) );
AND2_X1 _13068_ ( .A1(_02279_ ), .A2(\ID_EX_pc [25] ), .ZN(_00218_ ) );
NOR3_X1 _13069_ ( .A1(_05263_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00219_ ) );
NOR3_X1 _13070_ ( .A1(_03329_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00220_ ) );
AND2_X1 _13071_ ( .A1(_02279_ ), .A2(\ID_EX_pc [22] ), .ZN(_00221_ ) );
NOR3_X1 _13072_ ( .A1(_02270_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00222_ ) );
MUX2_X1 _13073_ ( .A(io_master_arready ), .B(_02212_ ), .S(_02207_ ), .Z(_05390_ ) );
BUF_X2 _13074_ ( .A(_02150_ ), .Z(_05391_ ) );
AND2_X1 _13075_ ( .A1(_05390_ ), .A2(_05391_ ), .ZN(_05392_ ) );
BUF_X4 _13076_ ( .A(_02120_ ), .Z(_05393_ ) );
INV_X1 _13077_ ( .A(_05393_ ), .ZN(_05394_ ) );
NOR3_X1 _13078_ ( .A1(_05392_ ), .A2(_02186_ ), .A3(_05394_ ), .ZN(_05395_ ) );
INV_X1 _13079_ ( .A(_05395_ ), .ZN(_05396_ ) );
BUF_X4 _13080_ ( .A(_02131_ ), .Z(_05397_ ) );
INV_X1 _13081_ ( .A(io_master_awready ), .ZN(_05398_ ) );
NAND3_X1 _13082_ ( .A1(_05397_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A3(_05398_ ), .ZN(_05399_ ) );
OAI21_X1 _13083_ ( .A(_05399_ ), .B1(\mylsu.state [4] ), .B2(\mylsu.state [0] ), .ZN(_05400_ ) );
AOI21_X1 _13084_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .B1(_05400_ ), .B2(EXU_valid_LSU ), .ZN(_05401_ ) );
AOI21_X1 _13085_ ( .A(_03248_ ), .B1(_05396_ ), .B2(_05401_ ), .ZN(_00223_ ) );
NOR3_X1 _13086_ ( .A1(_02267_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00224_ ) );
NOR3_X1 _13087_ ( .A1(_02262_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00225_ ) );
NOR3_X1 _13088_ ( .A1(_04299_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00226_ ) );
NOR3_X1 _13089_ ( .A1(_04730_ ), .A2(fanout_net_5 ), .A3(fanout_net_20 ), .ZN(_00227_ ) );
BUF_X4 _13090_ ( .A(_04649_ ), .Z(_05402_ ) );
NOR3_X1 _13091_ ( .A1(_05402_ ), .A2(fanout_net_5 ), .A3(excp_written ), .ZN(_00228_ ) );
NOR3_X1 _13092_ ( .A1(_04292_ ), .A2(fanout_net_5 ), .A3(excp_written ), .ZN(_00229_ ) );
NOR3_X1 _13093_ ( .A1(_04820_ ), .A2(fanout_net_5 ), .A3(excp_written ), .ZN(_00230_ ) );
AND2_X1 _13094_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_05403_ ) );
NOR2_X1 _13095_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_05404_ ) );
AND2_X2 _13096_ ( .A1(_05403_ ), .A2(_05404_ ), .ZN(_05405_ ) );
CLKBUF_X2 _13097_ ( .A(_05405_ ), .Z(_05406_ ) );
AND3_X1 _13098_ ( .A1(_05406_ ), .A2(\IF_ID_inst [12] ), .A3(\IF_ID_inst [6] ), .ZN(_05407_ ) );
AND2_X2 _13099_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05408_ ) );
AND2_X2 _13100_ ( .A1(_05407_ ), .A2(_05408_ ), .ZN(_05409_ ) );
INV_X1 _13101_ ( .A(\IF_ID_inst [6] ), .ZN(_05410_ ) );
NOR2_X1 _13102_ ( .A1(_05410_ ), .A2(\IF_ID_inst [12] ), .ZN(_05411_ ) );
AND3_X1 _13103_ ( .A1(_05411_ ), .A2(\IF_ID_inst [13] ), .A3(_05408_ ), .ZN(_05412_ ) );
AND2_X1 _13104_ ( .A1(_05412_ ), .A2(_05406_ ), .ZN(_05413_ ) );
NOR2_X1 _13105_ ( .A1(_05409_ ), .A2(_05413_ ), .ZN(_05414_ ) );
BUF_X4 _13106_ ( .A(_05414_ ), .Z(_05415_ ) );
INV_X1 _13107_ ( .A(\IF_ID_inst [31] ), .ZN(_05416_ ) );
AND2_X1 _13108_ ( .A1(_02249_ ), .A2(_02277_ ), .ZN(_05417_ ) );
INV_X1 _13109_ ( .A(_05417_ ), .ZN(_05418_ ) );
BUF_X4 _13110_ ( .A(_05418_ ), .Z(_05419_ ) );
BUF_X4 _13111_ ( .A(_05419_ ), .Z(_05420_ ) );
NOR3_X1 _13112_ ( .A1(_05415_ ), .A2(_05416_ ), .A3(_05420_ ), .ZN(_00231_ ) );
INV_X1 _13113_ ( .A(\IF_ID_inst [30] ), .ZN(_05421_ ) );
NOR3_X1 _13114_ ( .A1(_05415_ ), .A2(_05421_ ), .A3(_05420_ ), .ZN(_00232_ ) );
INV_X1 _13115_ ( .A(\IF_ID_inst [21] ), .ZN(_05422_ ) );
NOR3_X1 _13116_ ( .A1(_05415_ ), .A2(_05422_ ), .A3(_05420_ ), .ZN(_00233_ ) );
BUF_X4 _13117_ ( .A(_05419_ ), .Z(_05423_ ) );
INV_X1 _13118_ ( .A(_05414_ ), .ZN(_05424_ ) );
INV_X1 _13119_ ( .A(\IF_ID_inst [20] ), .ZN(_05425_ ) );
AOI21_X1 _13120_ ( .A(_05423_ ), .B1(_05424_ ), .B2(_05425_ ), .ZN(_00234_ ) );
INV_X1 _13121_ ( .A(\IF_ID_inst [29] ), .ZN(_05426_ ) );
AOI21_X1 _13122_ ( .A(_05423_ ), .B1(_05424_ ), .B2(_05426_ ), .ZN(_00235_ ) );
INV_X1 _13123_ ( .A(\IF_ID_inst [28] ), .ZN(_05427_ ) );
AOI21_X1 _13124_ ( .A(_05423_ ), .B1(_05424_ ), .B2(_05427_ ), .ZN(_00236_ ) );
INV_X1 _13125_ ( .A(\IF_ID_inst [27] ), .ZN(_05428_ ) );
NOR3_X1 _13126_ ( .A1(_05415_ ), .A2(_05428_ ), .A3(_05420_ ), .ZN(_00237_ ) );
INV_X1 _13127_ ( .A(\IF_ID_inst [26] ), .ZN(_05429_ ) );
AOI21_X1 _13128_ ( .A(_05423_ ), .B1(_05424_ ), .B2(_05429_ ), .ZN(_00238_ ) );
INV_X1 _13129_ ( .A(\IF_ID_inst [25] ), .ZN(_05430_ ) );
BUF_X4 _13130_ ( .A(_05418_ ), .Z(_05431_ ) );
NOR3_X1 _13131_ ( .A1(_05415_ ), .A2(_05430_ ), .A3(_05431_ ), .ZN(_00239_ ) );
INV_X1 _13132_ ( .A(\IF_ID_inst [24] ), .ZN(_05432_ ) );
NOR3_X1 _13133_ ( .A1(_05415_ ), .A2(_05432_ ), .A3(_05431_ ), .ZN(_00240_ ) );
INV_X1 _13134_ ( .A(\IF_ID_inst [23] ), .ZN(_05433_ ) );
NOR3_X1 _13135_ ( .A1(_05415_ ), .A2(_05433_ ), .A3(_05431_ ), .ZN(_00241_ ) );
INV_X1 _13136_ ( .A(\IF_ID_inst [22] ), .ZN(_05434_ ) );
NOR3_X1 _13137_ ( .A1(_05415_ ), .A2(_05434_ ), .A3(_05431_ ), .ZN(_00242_ ) );
AND3_X1 _13138_ ( .A1(_02249_ ), .A2(_02279_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00243_ ) );
AND3_X1 _13139_ ( .A1(_02249_ ), .A2(_02278_ ), .A3(\myidu.state [2] ), .ZN(_00244_ ) );
INV_X1 _13140_ ( .A(\IF_ID_inst [12] ), .ZN(_05435_ ) );
INV_X1 _13141_ ( .A(\IF_ID_inst [7] ), .ZN(_05436_ ) );
INV_X1 _13142_ ( .A(\IF_ID_inst [15] ), .ZN(_05437_ ) );
AND4_X1 _13143_ ( .A1(_05435_ ), .A2(_05436_ ), .A3(_05437_ ), .A4(\IF_ID_inst [6] ), .ZN(_05438_ ) );
NOR2_X1 _13144_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_05439_ ) );
BUF_X2 _13145_ ( .A(_05439_ ), .Z(_05440_ ) );
AND3_X1 _13146_ ( .A1(_05438_ ), .A2(_05408_ ), .A3(_05440_ ), .ZN(_05441_ ) );
INV_X1 _13147_ ( .A(\IF_ID_inst [11] ), .ZN(_05442_ ) );
INV_X1 _13148_ ( .A(\IF_ID_inst [10] ), .ZN(_05443_ ) );
INV_X1 _13149_ ( .A(\IF_ID_inst [9] ), .ZN(_05444_ ) );
NAND3_X1 _13150_ ( .A1(_05442_ ), .A2(_05443_ ), .A3(_05444_ ), .ZN(_05445_ ) );
NOR2_X1 _13151_ ( .A1(_05445_ ), .A2(\IF_ID_inst [8] ), .ZN(_05446_ ) );
AND3_X1 _13152_ ( .A1(_05441_ ), .A2(_05406_ ), .A3(_05446_ ), .ZN(_05447_ ) );
NOR4_X1 _13153_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .A4(\IF_ID_inst [31] ), .ZN(_05448_ ) );
NOR2_X1 _13154_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_05449_ ) );
NOR2_X1 _13155_ ( .A1(\IF_ID_inst [27] ), .A2(\IF_ID_inst [24] ), .ZN(_05450_ ) );
AND2_X1 _13156_ ( .A1(_05449_ ), .A2(_05450_ ), .ZN(_05451_ ) );
AND2_X1 _13157_ ( .A1(_05448_ ), .A2(_05451_ ), .ZN(_05452_ ) );
NAND2_X1 _13158_ ( .A1(_05447_ ), .A2(_05452_ ), .ZN(_05453_ ) );
NOR2_X1 _13159_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [18] ), .ZN(_05454_ ) );
NOR2_X1 _13160_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_05455_ ) );
AND2_X1 _13161_ ( .A1(_05454_ ), .A2(_05455_ ), .ZN(_05456_ ) );
NOR2_X1 _13162_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_05457_ ) );
NAND4_X1 _13163_ ( .A1(_05456_ ), .A2(_05422_ ), .A3(\IF_ID_inst [20] ), .A4(_05457_ ), .ZN(_05458_ ) );
NOR2_X1 _13164_ ( .A1(_05453_ ), .A2(_05458_ ), .ZN(_05459_ ) );
INV_X1 _13165_ ( .A(_05459_ ), .ZN(_05460_ ) );
INV_X1 _13166_ ( .A(\IF_ID_inst [5] ), .ZN(_05461_ ) );
NOR2_X1 _13167_ ( .A1(_05461_ ), .A2(\IF_ID_inst [4] ), .ZN(_05462_ ) );
NOR2_X1 _13168_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_05463_ ) );
AND3_X1 _13169_ ( .A1(_05405_ ), .A2(_05462_ ), .A3(_05463_ ), .ZN(_05464_ ) );
NAND2_X1 _13170_ ( .A1(_05464_ ), .A2(_05439_ ), .ZN(_05465_ ) );
NOR2_X1 _13171_ ( .A1(_05435_ ), .A2(\IF_ID_inst [6] ), .ZN(_05466_ ) );
AND3_X1 _13172_ ( .A1(_05466_ ), .A2(_05403_ ), .A3(_05404_ ), .ZN(_05467_ ) );
NAND3_X1 _13173_ ( .A1(_05467_ ), .A2(_05439_ ), .A3(_05462_ ), .ZN(_05468_ ) );
AND2_X1 _13174_ ( .A1(_05465_ ), .A2(_05468_ ), .ZN(_05469_ ) );
INV_X1 _13175_ ( .A(\IF_ID_inst [13] ), .ZN(_05470_ ) );
NOR2_X1 _13176_ ( .A1(_05470_ ), .A2(\IF_ID_inst [14] ), .ZN(_05471_ ) );
AND2_X1 _13177_ ( .A1(_05464_ ), .A2(_05471_ ), .ZN(_05472_ ) );
INV_X1 _13178_ ( .A(_05472_ ), .ZN(_05473_ ) );
AND2_X1 _13179_ ( .A1(_05469_ ), .A2(_05473_ ), .ZN(_05474_ ) );
NOR2_X1 _13180_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_05475_ ) );
AND4_X1 _13181_ ( .A1(\IF_ID_inst [12] ), .A2(_05440_ ), .A3(_05475_ ), .A4(_05410_ ), .ZN(_05476_ ) );
AND3_X2 _13182_ ( .A1(_05403_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_05477_ ) );
CLKBUF_X2 _13183_ ( .A(_05477_ ), .Z(_05478_ ) );
AND2_X1 _13184_ ( .A1(_05476_ ), .A2(_05478_ ), .ZN(_05479_ ) );
AND2_X1 _13185_ ( .A1(_05411_ ), .A2(_05462_ ), .ZN(_05480_ ) );
AND2_X1 _13186_ ( .A1(_05480_ ), .A2(_05406_ ), .ZN(_05481_ ) );
AND3_X1 _13187_ ( .A1(_05457_ ), .A2(\IF_ID_inst [21] ), .A3(_05425_ ), .ZN(_05482_ ) );
NAND2_X1 _13188_ ( .A1(\IF_ID_inst [29] ), .A2(\IF_ID_inst [28] ), .ZN(_05483_ ) );
NOR3_X1 _13189_ ( .A1(_05483_ ), .A2(\IF_ID_inst [30] ), .A3(\IF_ID_inst [31] ), .ZN(_05484_ ) );
AND4_X1 _13190_ ( .A1(_05451_ ), .A2(_05482_ ), .A3(_05456_ ), .A4(_05484_ ), .ZN(_05485_ ) );
AOI221_X4 _13191_ ( .A(_05479_ ), .B1(_05440_ ), .B2(_05481_ ), .C1(_05447_ ), .C2(_05485_ ), .ZN(_05486_ ) );
NAND3_X1 _13192_ ( .A1(_05460_ ), .A2(_05474_ ), .A3(_05486_ ), .ZN(_05487_ ) );
AND4_X1 _13193_ ( .A1(\IF_ID_inst [14] ), .A2(_05407_ ), .A3(\IF_ID_inst [13] ), .A4(_05462_ ), .ZN(_05488_ ) );
AND2_X1 _13194_ ( .A1(_05481_ ), .A2(\IF_ID_inst [14] ), .ZN(_05489_ ) );
AND3_X1 _13195_ ( .A1(_05407_ ), .A2(_05470_ ), .A3(_05462_ ), .ZN(_05490_ ) );
OR3_X1 _13196_ ( .A1(_05488_ ), .A2(_05489_ ), .A3(_05490_ ), .ZN(_05491_ ) );
NOR4_X1 _13197_ ( .A1(_05487_ ), .A2(_05442_ ), .A3(_05431_ ), .A4(_05491_ ), .ZN(_00245_ ) );
NOR4_X1 _13198_ ( .A1(_05487_ ), .A2(_05443_ ), .A3(_05431_ ), .A4(_05491_ ), .ZN(_00246_ ) );
NOR4_X1 _13199_ ( .A1(_05487_ ), .A2(_05444_ ), .A3(_05431_ ), .A4(_05491_ ), .ZN(_00247_ ) );
AND3_X1 _13200_ ( .A1(_05460_ ), .A2(_05474_ ), .A3(_05486_ ), .ZN(_05492_ ) );
CLKBUF_X2 _13201_ ( .A(_05417_ ), .Z(_05493_ ) );
NOR3_X1 _13202_ ( .A1(_05488_ ), .A2(_05490_ ), .A3(_05489_ ), .ZN(_05494_ ) );
AND4_X1 _13203_ ( .A1(\IF_ID_inst [8] ), .A2(_05492_ ), .A3(_05493_ ), .A4(_05494_ ), .ZN(_00248_ ) );
NOR4_X1 _13204_ ( .A1(_05487_ ), .A2(_05436_ ), .A3(_05431_ ), .A4(_05491_ ), .ZN(_00249_ ) );
NAND4_X1 _13205_ ( .A1(_05406_ ), .A2(\IF_ID_inst [6] ), .A3(_05436_ ), .A4(_05408_ ), .ZN(_05495_ ) );
NOR4_X1 _13206_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_05496_ ) );
NAND2_X1 _13207_ ( .A1(_05446_ ), .A2(_05496_ ), .ZN(_05497_ ) );
NOR2_X1 _13208_ ( .A1(_05495_ ), .A2(_05497_ ), .ZN(_05498_ ) );
AND4_X1 _13209_ ( .A1(_05451_ ), .A2(_05482_ ), .A3(_05456_ ), .A4(_05484_ ), .ZN(_05499_ ) );
AND2_X1 _13210_ ( .A1(_05498_ ), .A2(_05499_ ), .ZN(_05500_ ) );
INV_X1 _13211_ ( .A(_05500_ ), .ZN(_05501_ ) );
INV_X1 _13212_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_05502_ ) );
AND2_X1 _13213_ ( .A1(_05462_ ), .A2(_05502_ ), .ZN(_05503_ ) );
AND2_X2 _13214_ ( .A1(_05503_ ), .A2(_05477_ ), .ZN(_05504_ ) );
INV_X1 _13215_ ( .A(_05504_ ), .ZN(_05505_ ) );
NAND3_X1 _13216_ ( .A1(\IF_ID_inst [2] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [1] ), .ZN(_05506_ ) );
NOR2_X1 _13217_ ( .A1(_05506_ ), .A2(\IF_ID_inst [3] ), .ZN(_05507_ ) );
AND3_X1 _13218_ ( .A1(_05410_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_05508_ ) );
NAND2_X1 _13219_ ( .A1(_05507_ ), .A2(_05508_ ), .ZN(_05509_ ) );
INV_X1 _13220_ ( .A(\IF_ID_inst [4] ), .ZN(_05510_ ) );
NOR2_X1 _13221_ ( .A1(_05510_ ), .A2(\IF_ID_inst [5] ), .ZN(_05511_ ) );
NAND3_X1 _13222_ ( .A1(_05507_ ), .A2(_05410_ ), .A3(_05511_ ), .ZN(_05512_ ) );
NAND4_X1 _13223_ ( .A1(_05501_ ), .A2(_05505_ ), .A3(_05509_ ), .A4(_05512_ ), .ZN(_05513_ ) );
AND4_X1 _13224_ ( .A1(_05422_ ), .A2(_05433_ ), .A3(_05434_ ), .A4(\IF_ID_inst [20] ), .ZN(_05514_ ) );
AND4_X1 _13225_ ( .A1(_05451_ ), .A2(_05448_ ), .A3(_05456_ ), .A4(_05514_ ), .ZN(_05515_ ) );
AOI21_X1 _13226_ ( .A(_05479_ ), .B1(_05498_ ), .B2(_05515_ ), .ZN(_05516_ ) );
INV_X1 _13227_ ( .A(_05516_ ), .ZN(_05517_ ) );
INV_X1 _13228_ ( .A(\IF_ID_inst [19] ), .ZN(_05518_ ) );
NOR4_X1 _13229_ ( .A1(_05513_ ), .A2(_05517_ ), .A3(_05518_ ), .A4(_05419_ ), .ZN(_00250_ ) );
INV_X1 _13230_ ( .A(\IF_ID_inst [18] ), .ZN(_05519_ ) );
NOR4_X1 _13231_ ( .A1(_05513_ ), .A2(_05517_ ), .A3(_05519_ ), .A4(_05419_ ), .ZN(_00251_ ) );
INV_X1 _13232_ ( .A(\IF_ID_inst [17] ), .ZN(_05520_ ) );
NOR4_X1 _13233_ ( .A1(_05513_ ), .A2(_05517_ ), .A3(_05520_ ), .A4(_05419_ ), .ZN(_00252_ ) );
AND2_X2 _13234_ ( .A1(_05405_ ), .A2(_05463_ ), .ZN(_05521_ ) );
AND2_X1 _13235_ ( .A1(_05521_ ), .A2(_05475_ ), .ZN(_05522_ ) );
AND2_X1 _13236_ ( .A1(_05522_ ), .A2(_05471_ ), .ZN(_05523_ ) );
INV_X1 _13237_ ( .A(_05523_ ), .ZN(_05524_ ) );
NAND2_X1 _13238_ ( .A1(_05481_ ), .A2(_05440_ ), .ZN(_05525_ ) );
AND3_X1 _13239_ ( .A1(_05411_ ), .A2(_05462_ ), .A3(_05440_ ), .ZN(_05526_ ) );
AND2_X1 _13240_ ( .A1(_05526_ ), .A2(_05507_ ), .ZN(_05527_ ) );
INV_X1 _13241_ ( .A(_05527_ ), .ZN(_05528_ ) );
NAND3_X1 _13242_ ( .A1(_05524_ ), .A2(_05525_ ), .A3(_05528_ ), .ZN(_05529_ ) );
INV_X1 _13243_ ( .A(_05474_ ), .ZN(_05530_ ) );
AND2_X1 _13244_ ( .A1(_05467_ ), .A2(_05511_ ), .ZN(_05531_ ) );
NOR3_X1 _13245_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_05532_ ) );
AND3_X1 _13246_ ( .A1(_05532_ ), .A2(_05428_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05533_ ) );
INV_X1 _13247_ ( .A(\IF_ID_inst [14] ), .ZN(_05534_ ) );
NOR2_X1 _13248_ ( .A1(_05534_ ), .A2(\IF_ID_inst [13] ), .ZN(_05535_ ) );
AND2_X1 _13249_ ( .A1(_05535_ ), .A2(_05449_ ), .ZN(_05536_ ) );
AND2_X2 _13250_ ( .A1(_05533_ ), .A2(_05536_ ), .ZN(_05537_ ) );
NAND3_X1 _13251_ ( .A1(_05427_ ), .A2(_05428_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05538_ ) );
NOR3_X1 _13252_ ( .A1(_05538_ ), .A2(_05421_ ), .A3(\IF_ID_inst [29] ), .ZN(_05539_ ) );
AND2_X1 _13253_ ( .A1(_05539_ ), .A2(_05536_ ), .ZN(_05540_ ) );
OAI21_X1 _13254_ ( .A(_05531_ ), .B1(_05537_ ), .B2(_05540_ ), .ZN(_05541_ ) );
INV_X1 _13255_ ( .A(_05541_ ), .ZN(_05542_ ) );
OR4_X1 _13256_ ( .A1(_05424_ ), .A2(_05529_ ), .A3(_05530_ ), .A4(_05542_ ), .ZN(_05543_ ) );
AND2_X1 _13257_ ( .A1(_05532_ ), .A2(_05428_ ), .ZN(_05544_ ) );
AND4_X1 _13258_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A2(_05449_ ), .A3(_05534_ ), .A4(\IF_ID_inst [13] ), .ZN(_05545_ ) );
AND2_X1 _13259_ ( .A1(_05544_ ), .A2(_05545_ ), .ZN(_05546_ ) );
NAND3_X1 _13260_ ( .A1(_05546_ ), .A2(_05408_ ), .A3(_05521_ ), .ZN(_05547_ ) );
AND2_X1 _13261_ ( .A1(_05439_ ), .A2(_05449_ ), .ZN(_05548_ ) );
NAND4_X1 _13262_ ( .A1(_05521_ ), .A2(_05408_ ), .A3(_05539_ ), .A4(_05548_ ), .ZN(_05549_ ) );
AND2_X1 _13263_ ( .A1(_05547_ ), .A2(_05549_ ), .ZN(_05550_ ) );
INV_X1 _13264_ ( .A(_05550_ ), .ZN(_05551_ ) );
AND3_X1 _13265_ ( .A1(_05406_ ), .A2(_05466_ ), .A3(_05475_ ), .ZN(_05552_ ) );
AND2_X1 _13266_ ( .A1(_05552_ ), .A2(_05470_ ), .ZN(_05553_ ) );
AND3_X1 _13267_ ( .A1(_05521_ ), .A2(_05470_ ), .A3(_05475_ ), .ZN(_05554_ ) );
AND2_X1 _13268_ ( .A1(_05533_ ), .A2(_05548_ ), .ZN(_05555_ ) );
AND2_X1 _13269_ ( .A1(_05555_ ), .A2(_05531_ ), .ZN(_05556_ ) );
OR4_X1 _13270_ ( .A1(_05551_ ), .A2(_05553_ ), .A3(_05554_ ), .A4(_05556_ ), .ZN(_05557_ ) );
AND3_X1 _13271_ ( .A1(_05467_ ), .A2(\IF_ID_inst [13] ), .A3(_05511_ ), .ZN(_05558_ ) );
AND2_X1 _13272_ ( .A1(_05558_ ), .A2(_05534_ ), .ZN(_05559_ ) );
AND2_X1 _13273_ ( .A1(_05521_ ), .A2(_05511_ ), .ZN(_05560_ ) );
AND4_X1 _13274_ ( .A1(\IF_ID_inst [14] ), .A2(_05467_ ), .A3(\IF_ID_inst [13] ), .A4(_05511_ ), .ZN(_05561_ ) );
OR3_X1 _13275_ ( .A1(_05559_ ), .A2(_05560_ ), .A3(_05561_ ), .ZN(_05562_ ) );
NOR4_X1 _13276_ ( .A1(_05543_ ), .A2(_05491_ ), .A3(_05557_ ), .A4(_05562_ ), .ZN(_05563_ ) );
AND2_X1 _13277_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_05564_ ) );
AND3_X1 _13278_ ( .A1(_05544_ ), .A2(_05564_ ), .A3(_05449_ ), .ZN(_05565_ ) );
AND2_X1 _13279_ ( .A1(_05565_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05566_ ) );
AND4_X1 _13280_ ( .A1(\IF_ID_inst [4] ), .A2(_05410_ ), .A3(\IF_ID_inst [5] ), .A4(\IF_ID_inst [12] ), .ZN(_05567_ ) );
AND2_X2 _13281_ ( .A1(_05406_ ), .A2(_05567_ ), .ZN(_05568_ ) );
AND2_X1 _13282_ ( .A1(_05566_ ), .A2(_05568_ ), .ZN(_05569_ ) );
AND2_X2 _13283_ ( .A1(_05521_ ), .A2(_05408_ ), .ZN(_05570_ ) );
OR2_X1 _13284_ ( .A1(_05537_ ), .A2(_05555_ ), .ZN(_05571_ ) );
OAI22_X1 _13285_ ( .A1(_05569_ ), .A2(_05570_ ), .B1(_05571_ ), .B2(_05566_ ), .ZN(_05572_ ) );
AND2_X1 _13286_ ( .A1(_05540_ ), .A2(_05568_ ), .ZN(_05573_ ) );
INV_X1 _13287_ ( .A(_05573_ ), .ZN(_05574_ ) );
NOR3_X1 _13288_ ( .A1(_05537_ ), .A2(_05555_ ), .A3(_05546_ ), .ZN(_05575_ ) );
INV_X1 _13289_ ( .A(_05568_ ), .ZN(_05576_ ) );
NOR2_X1 _13290_ ( .A1(_05575_ ), .A2(_05576_ ), .ZN(_05577_ ) );
INV_X1 _13291_ ( .A(_05577_ ), .ZN(_05578_ ) );
AND3_X1 _13292_ ( .A1(_05572_ ), .A2(_05574_ ), .A3(_05578_ ), .ZN(_05579_ ) );
NAND2_X1 _13293_ ( .A1(_05563_ ), .A2(_05579_ ), .ZN(_05580_ ) );
NOR2_X1 _13294_ ( .A1(_05513_ ), .A2(_05517_ ), .ZN(_05581_ ) );
INV_X1 _13295_ ( .A(_05581_ ), .ZN(_05582_ ) );
NOR2_X2 _13296_ ( .A1(_05580_ ), .A2(_05582_ ), .ZN(_05583_ ) );
INV_X1 _13297_ ( .A(_05583_ ), .ZN(_05584_ ) );
XNOR2_X1 _13298_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_05585_ ) );
XNOR2_X1 _13299_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_05586_ ) );
XNOR2_X1 _13300_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_05587_ ) );
XNOR2_X1 _13301_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_05588_ ) );
AND4_X1 _13302_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(_05587_ ), .A4(_05588_ ), .ZN(_05589_ ) );
XNOR2_X1 _13303_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_05590_ ) );
XNOR2_X1 _13304_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_05591_ ) );
XNOR2_X1 _13305_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_05592_ ) );
XNOR2_X1 _13306_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_05593_ ) );
AND4_X1 _13307_ ( .A1(_05590_ ), .A2(_05591_ ), .A3(_05592_ ), .A4(_05593_ ), .ZN(_05594_ ) );
XNOR2_X1 _13308_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_05595_ ) );
XNOR2_X1 _13309_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_05596_ ) );
XNOR2_X1 _13310_ ( .A(\IF_ID_pc [21] ), .B(\myexu.pc_jump [21] ), .ZN(_05597_ ) );
XNOR2_X1 _13311_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_05598_ ) );
AND4_X1 _13312_ ( .A1(_05595_ ), .A2(_05596_ ), .A3(_05597_ ), .A4(_05598_ ), .ZN(_05599_ ) );
XNOR2_X1 _13313_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_05600_ ) );
XNOR2_X1 _13314_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_05601_ ) );
XNOR2_X1 _13315_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_05602_ ) );
XNOR2_X1 _13316_ ( .A(fanout_net_16 ), .B(\myexu.pc_jump [4] ), .ZN(_05603_ ) );
AND4_X1 _13317_ ( .A1(_05600_ ), .A2(_05601_ ), .A3(_05602_ ), .A4(_05603_ ), .ZN(_05604_ ) );
XNOR2_X1 _13318_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_05605_ ) );
XNOR2_X1 _13319_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_05606_ ) );
XNOR2_X1 _13320_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_05607_ ) );
XNOR2_X1 _13321_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_05608_ ) );
AND4_X1 _13322_ ( .A1(_05605_ ), .A2(_05606_ ), .A3(_05607_ ), .A4(_05608_ ), .ZN(_05609_ ) );
AND4_X1 _13323_ ( .A1(_05594_ ), .A2(_05599_ ), .A3(_05604_ ), .A4(_05609_ ), .ZN(_05610_ ) );
XNOR2_X1 _13324_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_05611_ ) );
XNOR2_X1 _13325_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_05612_ ) );
XNOR2_X1 _13326_ ( .A(fanout_net_12 ), .B(\myexu.pc_jump [3] ), .ZN(_05613_ ) );
XNOR2_X1 _13327_ ( .A(\myexu.pc_jump [2] ), .B(\IF_ID_pc [2] ), .ZN(_05614_ ) );
AND4_X1 _13328_ ( .A1(_05611_ ), .A2(_05612_ ), .A3(_05613_ ), .A4(_05614_ ), .ZN(_05615_ ) );
XNOR2_X1 _13329_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_05616_ ) );
XNOR2_X1 _13330_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_05617_ ) );
XNOR2_X1 _13331_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_05618_ ) );
XNOR2_X1 _13332_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_05619_ ) );
XNOR2_X1 _13333_ ( .A(\IF_ID_pc [25] ), .B(\myexu.pc_jump [25] ), .ZN(_05620_ ) );
AND4_X1 _13334_ ( .A1(_05617_ ), .A2(_05618_ ), .A3(_05619_ ), .A4(_05620_ ), .ZN(_05621_ ) );
XNOR2_X1 _13335_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_05622_ ) );
XOR2_X1 _13336_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .Z(_05623_ ) );
XOR2_X1 _13337_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .Z(_05624_ ) );
NOR2_X1 _13338_ ( .A1(_05623_ ), .A2(_05624_ ), .ZN(_05625_ ) );
AND4_X1 _13339_ ( .A1(_05616_ ), .A2(_05621_ ), .A3(_05622_ ), .A4(_05625_ ), .ZN(_05626_ ) );
AND4_X1 _13340_ ( .A1(_05589_ ), .A2(_05610_ ), .A3(_05615_ ), .A4(_05626_ ), .ZN(_05627_ ) );
NOR2_X1 _13341_ ( .A1(_05627_ ), .A2(_02265_ ), .ZN(_05628_ ) );
INV_X1 _13342_ ( .A(\myifu.state [1] ), .ZN(_05629_ ) );
NOR2_X1 _13343_ ( .A1(_05629_ ), .A2(fanout_net_48 ), .ZN(_05630_ ) );
INV_X1 _13344_ ( .A(_05630_ ), .ZN(_05631_ ) );
NOR2_X1 _13345_ ( .A1(_05628_ ), .A2(_05631_ ), .ZN(_05632_ ) );
AND2_X1 _13346_ ( .A1(_05632_ ), .A2(IDU_ready_IFU ), .ZN(_05633_ ) );
BUF_X4 _13347_ ( .A(_05633_ ), .Z(_05634_ ) );
OAI211_X1 _13348_ ( .A(_05584_ ), .B(_05634_ ), .C1(_05519_ ), .C2(_05582_ ), .ZN(_05635_ ) );
INV_X1 _13349_ ( .A(_05635_ ), .ZN(_05636_ ) );
INV_X1 _13350_ ( .A(_05634_ ), .ZN(_05637_ ) );
NOR2_X1 _13351_ ( .A1(_05583_ ), .A2(_05637_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _13352_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_05638_ ) );
AOI211_X1 _13353_ ( .A(_05431_ ), .B(_05636_ ), .C1(_02350_ ), .C2(_05638_ ), .ZN(_00253_ ) );
INV_X1 _13354_ ( .A(\IF_ID_inst [16] ), .ZN(_05639_ ) );
NOR4_X1 _13355_ ( .A1(_05513_ ), .A2(_05517_ ), .A3(_05639_ ), .A4(_05419_ ), .ZN(_00254_ ) );
OAI21_X1 _13356_ ( .A(\ID_EX_rs1 [2] ), .B1(_05583_ ), .B2(_05637_ ), .ZN(_05640_ ) );
NAND4_X1 _13357_ ( .A1(_05580_ ), .A2(\IF_ID_inst [17] ), .A3(_05581_ ), .A4(_05634_ ), .ZN(_05641_ ) );
AOI21_X1 _13358_ ( .A(_05423_ ), .B1(_05640_ ), .B2(_05641_ ), .ZN(_00255_ ) );
NOR4_X1 _13359_ ( .A1(_05513_ ), .A2(_05517_ ), .A3(_05437_ ), .A4(_05419_ ), .ZN(_00256_ ) );
OAI211_X1 _13360_ ( .A(_05584_ ), .B(_05634_ ), .C1(_05639_ ), .C2(_05582_ ), .ZN(_05642_ ) );
INV_X1 _13361_ ( .A(_05642_ ), .ZN(_05643_ ) );
AOI211_X1 _13362_ ( .A(_05419_ ), .B(_05643_ ), .C1(_02347_ ), .C2(_05638_ ), .ZN(_00257_ ) );
NOR2_X1 _13363_ ( .A1(_05459_ ), .A2(_05424_ ), .ZN(_05644_ ) );
NOR4_X1 _13364_ ( .A1(_05500_ ), .A2(_05553_ ), .A3(_05554_ ), .A4(_05479_ ), .ZN(_05645_ ) );
NOR2_X1 _13365_ ( .A1(_05527_ ), .A2(_05504_ ), .ZN(_05646_ ) );
INV_X1 _13366_ ( .A(_05646_ ), .ZN(_05647_ ) );
NOR2_X1 _13367_ ( .A1(_05523_ ), .A2(_05647_ ), .ZN(_05648_ ) );
INV_X1 _13368_ ( .A(_05471_ ), .ZN(_05649_ ) );
AND3_X1 _13369_ ( .A1(_05521_ ), .A2(_05649_ ), .A3(_05511_ ), .ZN(_05650_ ) );
NOR2_X1 _13370_ ( .A1(_05650_ ), .A2(_05558_ ), .ZN(_05651_ ) );
AND4_X1 _13371_ ( .A1(_05644_ ), .A2(_05645_ ), .A3(_05648_ ), .A4(_05651_ ), .ZN(_05652_ ) );
AND2_X1 _13372_ ( .A1(_05560_ ), .A2(_05471_ ), .ZN(_05653_ ) );
NOR2_X1 _13373_ ( .A1(_05510_ ), .A2(\IF_ID_inst [6] ), .ZN(_05654_ ) );
AND2_X1 _13374_ ( .A1(_05507_ ), .A2(_05654_ ), .ZN(_05655_ ) );
NOR2_X1 _13375_ ( .A1(_05653_ ), .A2(_05655_ ), .ZN(_05656_ ) );
NOR2_X1 _13376_ ( .A1(_05542_ ), .A2(_05556_ ), .ZN(_05657_ ) );
AND2_X2 _13377_ ( .A1(_05656_ ), .A2(_05657_ ), .ZN(_05658_ ) );
AND4_X1 _13378_ ( .A1(\IF_ID_inst [24] ), .A2(_05652_ ), .A3(_05493_ ), .A4(_05658_ ), .ZN(_00258_ ) );
OAI21_X1 _13379_ ( .A(\ID_EX_rs1 [0] ), .B1(_05583_ ), .B2(_05637_ ), .ZN(_05659_ ) );
NAND4_X1 _13380_ ( .A1(_05580_ ), .A2(\IF_ID_inst [15] ), .A3(_05581_ ), .A4(_05634_ ), .ZN(_05660_ ) );
AOI21_X1 _13381_ ( .A(_05423_ ), .B1(_05659_ ), .B2(_05660_ ), .ZN(_00259_ ) );
AND4_X1 _13382_ ( .A1(\IF_ID_inst [23] ), .A2(_05652_ ), .A3(_05493_ ), .A4(_05658_ ), .ZN(_00260_ ) );
AND4_X1 _13383_ ( .A1(\IF_ID_inst [22] ), .A2(_05652_ ), .A3(_05493_ ), .A4(_05658_ ), .ZN(_00261_ ) );
AND2_X1 _13384_ ( .A1(_05652_ ), .A2(_05658_ ), .ZN(_05661_ ) );
INV_X1 _13385_ ( .A(_05661_ ), .ZN(_05662_ ) );
OAI221_X1 _13386_ ( .A(_05634_ ), .B1(_05433_ ), .B2(_05662_ ), .C1(_05580_ ), .C2(_05582_ ), .ZN(_05663_ ) );
INV_X1 _13387_ ( .A(_05663_ ), .ZN(_05664_ ) );
AOI211_X1 _13388_ ( .A(_05419_ ), .B(_05664_ ), .C1(_03478_ ), .C2(_05638_ ), .ZN(_00262_ ) );
AND4_X1 _13389_ ( .A1(\IF_ID_inst [21] ), .A2(_05652_ ), .A3(_05493_ ), .A4(_05658_ ), .ZN(_00263_ ) );
NAND4_X1 _13390_ ( .A1(_05584_ ), .A2(\IF_ID_inst [22] ), .A3(_05634_ ), .A4(_05661_ ), .ZN(_05665_ ) );
OAI21_X1 _13391_ ( .A(\ID_EX_rs2 [2] ), .B1(_05583_ ), .B2(_05637_ ), .ZN(_05666_ ) );
AOI21_X1 _13392_ ( .A(_05423_ ), .B1(_05665_ ), .B2(_05666_ ), .ZN(_00264_ ) );
AND4_X1 _13393_ ( .A1(\IF_ID_inst [20] ), .A2(_05652_ ), .A3(_05493_ ), .A4(_05658_ ), .ZN(_00265_ ) );
OAI221_X1 _13394_ ( .A(_05634_ ), .B1(_05422_ ), .B2(_05662_ ), .C1(_05580_ ), .C2(_05582_ ), .ZN(_05667_ ) );
INV_X1 _13395_ ( .A(_05667_ ), .ZN(_05668_ ) );
AOI211_X1 _13396_ ( .A(_05419_ ), .B(_05668_ ), .C1(_03476_ ), .C2(_05638_ ), .ZN(_00266_ ) );
AND4_X1 _13397_ ( .A1(_02260_ ), .A2(_05476_ ), .A3(_05493_ ), .A4(_05478_ ), .ZN(_00267_ ) );
NAND4_X1 _13398_ ( .A1(_05584_ ), .A2(\IF_ID_inst [20] ), .A3(_05634_ ), .A4(_05661_ ), .ZN(_05669_ ) );
OAI21_X1 _13399_ ( .A(\ID_EX_rs2 [0] ), .B1(_05583_ ), .B2(_05637_ ), .ZN(_05670_ ) );
AOI21_X1 _13400_ ( .A(_05423_ ), .B1(_05669_ ), .B2(_05670_ ), .ZN(_00268_ ) );
INV_X1 _13401_ ( .A(IDU_ready_IFU ), .ZN(_05671_ ) );
OR2_X1 _13402_ ( .A1(_05523_ ), .A2(_05554_ ), .ZN(_05672_ ) );
OR3_X1 _13403_ ( .A1(_05672_ ), .A2(_05553_ ), .A3(_05527_ ), .ZN(_05673_ ) );
NOR3_X1 _13404_ ( .A1(_05673_ ), .A2(_05424_ ), .A3(_05562_ ), .ZN(_05674_ ) );
NOR2_X1 _13405_ ( .A1(_05500_ ), .A2(_05479_ ), .ZN(_05675_ ) );
XNOR2_X1 _13406_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_05676_ ) );
XNOR2_X1 _13407_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_05677_ ) );
XNOR2_X1 _13408_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_05678_ ) );
XNOR2_X1 _13409_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_05679_ ) );
AND4_X1 _13410_ ( .A1(_05676_ ), .A2(_05677_ ), .A3(_05678_ ), .A4(_05679_ ), .ZN(_05680_ ) );
AND2_X1 _13411_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_05681_ ) );
AND2_X1 _13412_ ( .A1(_05681_ ), .A2(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A ), .ZN(_05682_ ) );
XNOR2_X1 _13413_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_05683_ ) );
AND3_X1 _13414_ ( .A1(_05680_ ), .A2(_05682_ ), .A3(_05683_ ), .ZN(_05684_ ) );
XNOR2_X1 _13415_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_05685_ ) );
XNOR2_X1 _13416_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_05686_ ) );
XNOR2_X1 _13417_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_05687_ ) );
NAND4_X1 _13418_ ( .A1(_05682_ ), .A2(_05685_ ), .A3(_05686_ ), .A4(_05687_ ), .ZN(_05688_ ) );
XOR2_X1 _13419_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .Z(_05689_ ) );
XOR2_X1 _13420_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .Z(_05690_ ) );
NOR3_X1 _13421_ ( .A1(_05688_ ), .A2(_05689_ ), .A3(_05690_ ), .ZN(_05691_ ) );
OR2_X1 _13422_ ( .A1(_05684_ ), .A2(_05691_ ), .ZN(_05692_ ) );
NOR2_X1 _13423_ ( .A1(_05504_ ), .A2(_05655_ ), .ZN(_05693_ ) );
NAND4_X1 _13424_ ( .A1(_05460_ ), .A2(_05675_ ), .A3(_05692_ ), .A4(_05693_ ), .ZN(_05694_ ) );
AOI211_X1 _13425_ ( .A(_05671_ ), .B(_05418_ ), .C1(_05674_ ), .C2(_05694_ ), .ZN(_05695_ ) );
OR2_X1 _13426_ ( .A1(_05674_ ), .A2(_05684_ ), .ZN(_05696_ ) );
AND2_X1 _13427_ ( .A1(_05695_ ), .A2(_05696_ ), .ZN(_00269_ ) );
AND2_X1 _13428_ ( .A1(_05407_ ), .A2(_05462_ ), .ZN(_05697_ ) );
AOI22_X1 _13429_ ( .A1(_05697_ ), .A2(_05440_ ), .B1(\IF_ID_inst [14] ), .B2(_05481_ ), .ZN(_05698_ ) );
AOI22_X1 _13430_ ( .A1(_05697_ ), .A2(\IF_ID_inst [14] ), .B1(_05406_ ), .B2(_05526_ ), .ZN(_05699_ ) );
AND4_X1 _13431_ ( .A1(_05675_ ), .A2(_05646_ ), .A3(_05698_ ), .A4(_05699_ ), .ZN(_05700_ ) );
NAND3_X1 _13432_ ( .A1(_05441_ ), .A2(_05406_ ), .A3(_05446_ ), .ZN(_05701_ ) );
NAND4_X1 _13433_ ( .A1(_05448_ ), .A2(_05451_ ), .A3(_05422_ ), .A4(_05425_ ), .ZN(_05702_ ) );
NOR2_X1 _13434_ ( .A1(_05701_ ), .A2(_05702_ ), .ZN(_05703_ ) );
NAND3_X1 _13435_ ( .A1(_05703_ ), .A2(_05456_ ), .A3(_05457_ ), .ZN(_05704_ ) );
AND2_X1 _13436_ ( .A1(_05704_ ), .A2(_05414_ ), .ZN(_05705_ ) );
AOI21_X1 _13437_ ( .A(_05423_ ), .B1(_05700_ ), .B2(_05705_ ), .ZN(_00270_ ) );
AND2_X1 _13438_ ( .A1(_05552_ ), .A2(_05440_ ), .ZN(_05706_ ) );
AND3_X1 _13439_ ( .A1(_05552_ ), .A2(\IF_ID_inst [14] ), .A3(_05470_ ), .ZN(_05707_ ) );
NOR4_X1 _13440_ ( .A1(_05530_ ), .A2(_05672_ ), .A3(_05706_ ), .A4(_05707_ ), .ZN(_05708_ ) );
AOI21_X1 _13441_ ( .A(_05423_ ), .B1(_05708_ ), .B2(_05705_ ), .ZN(_00271_ ) );
NAND4_X1 _13442_ ( .A1(_05570_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_05544_ ), .A4(_05548_ ), .ZN(_05709_ ) );
NAND2_X1 _13443_ ( .A1(_05570_ ), .A2(_05537_ ), .ZN(_05710_ ) );
AND2_X1 _13444_ ( .A1(_05709_ ), .A2(_05710_ ), .ZN(_05711_ ) );
OAI211_X1 _13445_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B(_05565_ ), .C1(_05570_ ), .C2(_05568_ ), .ZN(_05712_ ) );
AND4_X1 _13446_ ( .A1(_05578_ ), .A2(_05711_ ), .A3(_05712_ ), .A4(_05651_ ), .ZN(_05713_ ) );
AND2_X1 _13447_ ( .A1(_05704_ ), .A2(_05574_ ), .ZN(_05714_ ) );
NAND2_X1 _13448_ ( .A1(_05539_ ), .A2(_05548_ ), .ZN(_05715_ ) );
NAND2_X1 _13449_ ( .A1(_05544_ ), .A2(_05545_ ), .ZN(_05716_ ) );
NAND2_X1 _13450_ ( .A1(_05715_ ), .A2(_05716_ ), .ZN(_05717_ ) );
AND2_X1 _13451_ ( .A1(_05570_ ), .A2(_05717_ ), .ZN(_05718_ ) );
NOR3_X1 _13452_ ( .A1(_05718_ ), .A2(_05553_ ), .A3(_05554_ ), .ZN(_05719_ ) );
AND4_X1 _13453_ ( .A1(_05648_ ), .A2(_05713_ ), .A3(_05714_ ), .A4(_05719_ ), .ZN(_05720_ ) );
AOI21_X1 _13454_ ( .A(_05420_ ), .B1(_05720_ ), .B2(_05658_ ), .ZN(_00272_ ) );
NOR3_X1 _13455_ ( .A1(_05650_ ), .A2(_05479_ ), .A3(_05558_ ), .ZN(_05721_ ) );
AOI21_X1 _13456_ ( .A(_05420_ ), .B1(_05658_ ), .B2(_05721_ ), .ZN(_00273_ ) );
AND2_X1 _13457_ ( .A1(_05447_ ), .A2(_05485_ ), .ZN(_05722_ ) );
AND3_X1 _13458_ ( .A1(_05546_ ), .A2(_05408_ ), .A3(_05521_ ), .ZN(_05723_ ) );
AND4_X1 _13459_ ( .A1(_05408_ ), .A2(_05521_ ), .A3(_05539_ ), .A4(_05548_ ), .ZN(_05724_ ) );
NOR4_X1 _13460_ ( .A1(_05722_ ), .A2(_05472_ ), .A3(_05723_ ), .A4(_05724_ ), .ZN(_05725_ ) );
AOI21_X1 _13461_ ( .A(_05420_ ), .B1(_05725_ ), .B2(_05656_ ), .ZN(_00274_ ) );
AOI221_X4 _13462_ ( .A(_05559_ ), .B1(\IF_ID_inst [14] ), .B2(_05697_ ), .C1(\IF_ID_inst [13] ), .C2(_05409_ ), .ZN(_05726_ ) );
INV_X1 _13463_ ( .A(_05655_ ), .ZN(_05727_ ) );
AOI22_X1 _13464_ ( .A1(_05522_ ), .A2(_05471_ ), .B1(_05568_ ), .B2(_05540_ ), .ZN(_05728_ ) );
AND4_X1 _13465_ ( .A1(_05473_ ), .A2(_05726_ ), .A3(_05727_ ), .A4(_05728_ ), .ZN(_05729_ ) );
NOR3_X1 _13466_ ( .A1(_05577_ ), .A2(_05542_ ), .A3(_05556_ ), .ZN(_05730_ ) );
AOI21_X1 _13467_ ( .A(_05420_ ), .B1(_05729_ ), .B2(_05730_ ), .ZN(_00275_ ) );
AOI221_X4 _13468_ ( .A(_05413_ ), .B1(_05464_ ), .B2(_05471_ ), .C1(\IF_ID_inst [14] ), .C2(_05481_ ), .ZN(_05731_ ) );
AND3_X1 _13469_ ( .A1(_05467_ ), .A2(_05440_ ), .A3(_05462_ ), .ZN(_05732_ ) );
AOI21_X1 _13470_ ( .A(_05732_ ), .B1(_05440_ ), .B2(_05552_ ), .ZN(_05733_ ) );
OAI21_X1 _13471_ ( .A(\IF_ID_inst [14] ), .B1(_05553_ ), .B2(_05560_ ), .ZN(_05734_ ) );
AND4_X1 _13472_ ( .A1(_05509_ ), .A2(_05731_ ), .A3(_05733_ ), .A4(_05734_ ), .ZN(_05735_ ) );
OAI21_X1 _13473_ ( .A(_05570_ ), .B1(_05566_ ), .B2(_05537_ ), .ZN(_05736_ ) );
OAI22_X1 _13474_ ( .A1(_05537_ ), .A2(_05540_ ), .B1(_05531_ ), .B2(_05568_ ), .ZN(_05737_ ) );
AND2_X1 _13475_ ( .A1(_05736_ ), .A2(_05737_ ), .ZN(_05738_ ) );
AOI21_X1 _13476_ ( .A(_05420_ ), .B1(_05735_ ), .B2(_05738_ ), .ZN(_00276_ ) );
NAND2_X1 _13477_ ( .A1(_05560_ ), .A2(_05535_ ), .ZN(_05739_ ) );
NAND4_X1 _13478_ ( .A1(_05539_ ), .A2(_05467_ ), .A3(_05511_ ), .A4(_05536_ ), .ZN(_05740_ ) );
NAND2_X1 _13479_ ( .A1(_05739_ ), .A2(_05740_ ), .ZN(_05741_ ) );
AND3_X1 _13480_ ( .A1(_05412_ ), .A2(\IF_ID_inst [14] ), .A3(_05406_ ), .ZN(_05742_ ) );
NOR3_X1 _13481_ ( .A1(_05741_ ), .A2(_05707_ ), .A3(_05742_ ), .ZN(_05743_ ) );
AOI22_X1 _13482_ ( .A1(_05566_ ), .A2(_05568_ ), .B1(_05546_ ), .B2(_05570_ ), .ZN(_05744_ ) );
AND3_X1 _13483_ ( .A1(_05744_ ), .A2(_05473_ ), .A3(_05528_ ), .ZN(_05745_ ) );
OAI21_X1 _13484_ ( .A(_05568_ ), .B1(_05555_ ), .B2(_05540_ ), .ZN(_05746_ ) );
OAI21_X1 _13485_ ( .A(_05535_ ), .B1(_05409_ ), .B2(_05522_ ), .ZN(_05747_ ) );
AND4_X1 _13486_ ( .A1(_05743_ ), .A2(_05745_ ), .A3(_05746_ ), .A4(_05747_ ), .ZN(_05748_ ) );
OR3_X1 _13487_ ( .A1(_05409_ ), .A2(_05481_ ), .A3(_05531_ ), .ZN(_05749_ ) );
OAI22_X1 _13488_ ( .A1(_05749_ ), .A2(_05697_ ), .B1(_05564_ ), .B2(_05556_ ), .ZN(_05750_ ) );
AOI22_X1 _13489_ ( .A1(_05697_ ), .A2(_05440_ ), .B1(_05570_ ), .B2(_05537_ ), .ZN(_05751_ ) );
AND4_X1 _13490_ ( .A1(_05469_ ), .A2(_05750_ ), .A3(_05460_ ), .A4(_05751_ ), .ZN(_05752_ ) );
AOI21_X1 _13491_ ( .A(_05420_ ), .B1(_05748_ ), .B2(_05752_ ), .ZN(_00277_ ) );
INV_X1 _13492_ ( .A(_05627_ ), .ZN(_05753_ ) );
INV_X1 _13493_ ( .A(fanout_net_48 ), .ZN(_05754_ ) );
BUF_X4 _13494_ ( .A(_05754_ ), .Z(_05755_ ) );
NAND4_X1 _13495_ ( .A1(_05753_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_05755_ ), .ZN(_05756_ ) );
NAND2_X1 _13496_ ( .A1(\mtvec [0] ), .A2(fanout_net_48 ), .ZN(_05757_ ) );
AOI21_X1 _13497_ ( .A(fanout_net_5 ), .B1(_05756_ ), .B2(_05757_ ), .ZN(_00281_ ) );
BUF_X2 _13498_ ( .A(_05628_ ), .Z(_05758_ ) );
AND4_X2 _13499_ ( .A1(\IF_ID_inst [31] ), .A2(_05510_ ), .A3(_05502_ ), .A4(\IF_ID_inst [5] ), .ZN(_05759_ ) );
AND2_X1 _13500_ ( .A1(_05405_ ), .A2(_05759_ ), .ZN(_05760_ ) );
AND2_X1 _13501_ ( .A1(_05760_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05761_ ) );
CLKBUF_X2 _13502_ ( .A(_05503_ ), .Z(_05762_ ) );
OAI211_X1 _13503_ ( .A(_05762_ ), .B(\IF_ID_inst [31] ), .C1(_05478_ ), .C2(_05405_ ), .ZN(_05763_ ) );
NOR2_X1 _13504_ ( .A1(_05761_ ), .A2(_05763_ ), .ZN(_05764_ ) );
XNOR2_X1 _13505_ ( .A(_05764_ ), .B(_02197_ ), .ZN(_05765_ ) );
AND2_X1 _13506_ ( .A1(_05504_ ), .A2(\IF_ID_inst [27] ), .ZN(_05766_ ) );
INV_X1 _13507_ ( .A(_05766_ ), .ZN(_05767_ ) );
INV_X1 _13508_ ( .A(_05760_ ), .ZN(_05768_ ) );
OAI21_X1 _13509_ ( .A(_05767_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_05768_ ), .ZN(_05769_ ) );
XNOR2_X1 _13510_ ( .A(_05769_ ), .B(_01962_ ), .ZN(_05770_ ) );
NAND3_X1 _13511_ ( .A1(_05503_ ), .A2(_05477_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_05771_ ) );
NAND3_X1 _13512_ ( .A1(_05405_ ), .A2(_05759_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_05772_ ) );
AND3_X1 _13513_ ( .A1(_05771_ ), .A2(\IF_ID_pc [2] ), .A3(_05772_ ), .ZN(_05773_ ) );
AOI21_X1 _13514_ ( .A(\IF_ID_pc [2] ), .B1(_05771_ ), .B2(_05772_ ), .ZN(_05774_ ) );
NOR2_X1 _13515_ ( .A1(_05773_ ), .A2(_05774_ ), .ZN(_05775_ ) );
NAND3_X1 _13516_ ( .A1(_05503_ ), .A2(_05477_ ), .A3(\IF_ID_inst [21] ), .ZN(_05776_ ) );
INV_X1 _13517_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_05777_ ) );
NAND3_X1 _13518_ ( .A1(_05405_ ), .A2(_05759_ ), .A3(_05777_ ), .ZN(_05778_ ) );
NAND2_X1 _13519_ ( .A1(_05776_ ), .A2(_05778_ ), .ZN(_05779_ ) );
AND2_X1 _13520_ ( .A1(_05779_ ), .A2(\IF_ID_pc [1] ), .ZN(_05780_ ) );
AND2_X1 _13521_ ( .A1(_05775_ ), .A2(_05780_ ), .ZN(_05781_ ) );
NOR2_X1 _13522_ ( .A1(_05781_ ), .A2(_05773_ ), .ZN(_05782_ ) );
NAND3_X1 _13523_ ( .A1(_05762_ ), .A2(_05477_ ), .A3(\IF_ID_inst [23] ), .ZN(_05783_ ) );
INV_X1 _13524_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_05784_ ) );
NAND3_X1 _13525_ ( .A1(_05405_ ), .A2(_05759_ ), .A3(_05784_ ), .ZN(_05785_ ) );
NAND2_X1 _13526_ ( .A1(_05783_ ), .A2(_05785_ ), .ZN(_05786_ ) );
XNOR2_X1 _13527_ ( .A(_05786_ ), .B(fanout_net_12 ), .ZN(_05787_ ) );
NAND3_X1 _13528_ ( .A1(_05503_ ), .A2(_05477_ ), .A3(\IF_ID_inst [24] ), .ZN(_05788_ ) );
INV_X1 _13529_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05789_ ) );
NAND3_X1 _13530_ ( .A1(_05405_ ), .A2(_05759_ ), .A3(_05789_ ), .ZN(_05790_ ) );
NAND2_X1 _13531_ ( .A1(_05788_ ), .A2(_05790_ ), .ZN(_05791_ ) );
NAND2_X1 _13532_ ( .A1(_05791_ ), .A2(fanout_net_16 ), .ZN(_05792_ ) );
INV_X1 _13533_ ( .A(fanout_net_16 ), .ZN(_05793_ ) );
NAND3_X1 _13534_ ( .A1(_05788_ ), .A2(_05793_ ), .A3(_05790_ ), .ZN(_05794_ ) );
AND2_X1 _13535_ ( .A1(_05792_ ), .A2(_05794_ ), .ZN(_05795_ ) );
INV_X1 _13536_ ( .A(_05795_ ), .ZN(_05796_ ) );
NOR3_X1 _13537_ ( .A1(_05782_ ), .A2(_05787_ ), .A3(_05796_ ), .ZN(_05797_ ) );
INV_X1 _13538_ ( .A(_05786_ ), .ZN(_05798_ ) );
OR2_X1 _13539_ ( .A1(_05798_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05799_ ) );
OAI21_X1 _13540_ ( .A(_05792_ ), .B1(_05796_ ), .B2(_05799_ ), .ZN(_05800_ ) );
NOR2_X1 _13541_ ( .A1(_05797_ ), .A2(_05800_ ), .ZN(_05801_ ) );
INV_X1 _13542_ ( .A(_05801_ ), .ZN(_05802_ ) );
NOR2_X1 _13543_ ( .A1(_05768_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_05803_ ) );
AND2_X1 _13544_ ( .A1(_05504_ ), .A2(\IF_ID_inst [25] ), .ZN(_05804_ ) );
NOR2_X1 _13545_ ( .A1(_05803_ ), .A2(_05804_ ), .ZN(_05805_ ) );
XNOR2_X1 _13546_ ( .A(_05805_ ), .B(\IF_ID_pc [5] ), .ZN(_05806_ ) );
AND2_X1 _13547_ ( .A1(_05504_ ), .A2(\IF_ID_inst [26] ), .ZN(_05807_ ) );
INV_X1 _13548_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05808_ ) );
AOI21_X1 _13549_ ( .A(_05807_ ), .B1(_05808_ ), .B2(_05760_ ), .ZN(_05809_ ) );
XNOR2_X1 _13550_ ( .A(_05809_ ), .B(\IF_ID_pc [6] ), .ZN(_05810_ ) );
AND3_X1 _13551_ ( .A1(_05802_ ), .A2(_05806_ ), .A3(_05810_ ), .ZN(_05811_ ) );
AND2_X1 _13552_ ( .A1(_05809_ ), .A2(_02033_ ), .ZN(_05812_ ) );
OR2_X1 _13553_ ( .A1(_05805_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05813_ ) );
NOR2_X1 _13554_ ( .A1(_05809_ ), .A2(_02033_ ), .ZN(_05814_ ) );
OR3_X1 _13555_ ( .A1(_05812_ ), .A2(_05813_ ), .A3(_05814_ ), .ZN(_05815_ ) );
OAI21_X1 _13556_ ( .A(_05815_ ), .B1(_02033_ ), .B2(_05809_ ), .ZN(_05816_ ) );
OAI21_X1 _13557_ ( .A(_05770_ ), .B1(_05811_ ), .B2(_05816_ ), .ZN(_05817_ ) );
INV_X1 _13558_ ( .A(_05817_ ), .ZN(_05818_ ) );
AND2_X1 _13559_ ( .A1(_05769_ ), .A2(\IF_ID_pc [7] ), .ZN(_05819_ ) );
AND2_X1 _13560_ ( .A1(_05504_ ), .A2(\IF_ID_inst [28] ), .ZN(_05820_ ) );
INV_X1 _13561_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05821_ ) );
BUF_X4 _13562_ ( .A(_05760_ ), .Z(_05822_ ) );
AOI21_X1 _13563_ ( .A(_05820_ ), .B1(_05821_ ), .B2(_05822_ ), .ZN(_05823_ ) );
INV_X1 _13564_ ( .A(_05823_ ), .ZN(_05824_ ) );
OAI22_X1 _13565_ ( .A1(_05818_ ), .A2(_05819_ ), .B1(\IF_ID_pc [8] ), .B2(_05824_ ), .ZN(_05825_ ) );
INV_X1 _13566_ ( .A(\IF_ID_pc [8] ), .ZN(_05826_ ) );
OR2_X1 _13567_ ( .A1(_05823_ ), .A2(_05826_ ), .ZN(_05827_ ) );
NAND2_X1 _13568_ ( .A1(_05825_ ), .A2(_05827_ ), .ZN(_05828_ ) );
NAND3_X1 _13569_ ( .A1(_05762_ ), .A2(_05478_ ), .A3(\IF_ID_inst [16] ), .ZN(_05829_ ) );
MUX2_X1 _13570_ ( .A(_05829_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .S(_05822_ ), .Z(_05830_ ) );
XNOR2_X1 _13571_ ( .A(_05830_ ), .B(\IF_ID_pc [16] ), .ZN(_05831_ ) );
AND3_X1 _13572_ ( .A1(_05762_ ), .A2(_05478_ ), .A3(\IF_ID_inst [15] ), .ZN(_05832_ ) );
INV_X1 _13573_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_05833_ ) );
MUX2_X1 _13574_ ( .A(_05832_ ), .B(_05833_ ), .S(_05822_ ), .Z(_05834_ ) );
XNOR2_X1 _13575_ ( .A(_05834_ ), .B(_02049_ ), .ZN(_05835_ ) );
AND2_X1 _13576_ ( .A1(_05831_ ), .A2(_05835_ ), .ZN(_05836_ ) );
OAI21_X1 _13577_ ( .A(_05768_ ), .B1(_05505_ ), .B2(_05534_ ), .ZN(_05837_ ) );
INV_X1 _13578_ ( .A(_05761_ ), .ZN(_05838_ ) );
NAND2_X1 _13579_ ( .A1(_05837_ ), .A2(_05838_ ), .ZN(_05839_ ) );
XNOR2_X1 _13580_ ( .A(_05839_ ), .B(\IF_ID_pc [14] ), .ZN(_05840_ ) );
AND3_X1 _13581_ ( .A1(_05762_ ), .A2(_05478_ ), .A3(\IF_ID_inst [13] ), .ZN(_05841_ ) );
MUX2_X1 _13582_ ( .A(_05841_ ), .B(_05833_ ), .S(_05822_ ), .Z(_05842_ ) );
XNOR2_X1 _13583_ ( .A(_05842_ ), .B(_02038_ ), .ZN(_05843_ ) );
AND3_X1 _13584_ ( .A1(_05836_ ), .A2(_05840_ ), .A3(_05843_ ), .ZN(_05844_ ) );
AND3_X1 _13585_ ( .A1(_05762_ ), .A2(_05477_ ), .A3(\IF_ID_inst [12] ), .ZN(_05845_ ) );
MUX2_X1 _13586_ ( .A(_05845_ ), .B(_05833_ ), .S(_05822_ ), .Z(_05846_ ) );
XNOR2_X1 _13587_ ( .A(_05846_ ), .B(_02023_ ), .ZN(_05847_ ) );
INV_X1 _13588_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05848_ ) );
AND3_X1 _13589_ ( .A1(_05405_ ), .A2(_05759_ ), .A3(_05848_ ), .ZN(_05849_ ) );
AOI21_X1 _13590_ ( .A(_05849_ ), .B1(\IF_ID_inst [20] ), .B2(_05504_ ), .ZN(_05850_ ) );
XNOR2_X1 _13591_ ( .A(_05850_ ), .B(\IF_ID_pc [11] ), .ZN(_05851_ ) );
AND2_X1 _13592_ ( .A1(_05847_ ), .A2(_05851_ ), .ZN(_05852_ ) );
AND2_X1 _13593_ ( .A1(_05504_ ), .A2(\IF_ID_inst [29] ), .ZN(_05853_ ) );
INV_X1 _13594_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_05854_ ) );
AOI21_X1 _13595_ ( .A(_05853_ ), .B1(_05854_ ), .B2(_05822_ ), .ZN(_05855_ ) );
XNOR2_X1 _13596_ ( .A(_05855_ ), .B(\IF_ID_pc [9] ), .ZN(_05856_ ) );
AND2_X1 _13597_ ( .A1(_05504_ ), .A2(\IF_ID_inst [30] ), .ZN(_05857_ ) );
INV_X1 _13598_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_05858_ ) );
AOI21_X1 _13599_ ( .A(_05857_ ), .B1(_05858_ ), .B2(_05822_ ), .ZN(_05859_ ) );
XNOR2_X1 _13600_ ( .A(_05859_ ), .B(\IF_ID_pc [10] ), .ZN(_05860_ ) );
AND3_X1 _13601_ ( .A1(_05852_ ), .A2(_05856_ ), .A3(_05860_ ), .ZN(_05861_ ) );
NAND3_X1 _13602_ ( .A1(_05828_ ), .A2(_05844_ ), .A3(_05861_ ), .ZN(_05862_ ) );
AND2_X1 _13603_ ( .A1(_05842_ ), .A2(\IF_ID_pc [13] ), .ZN(_05863_ ) );
NAND2_X1 _13604_ ( .A1(_05840_ ), .A2(_05863_ ), .ZN(_05864_ ) );
OAI21_X1 _13605_ ( .A(_05864_ ), .B1(_02016_ ), .B2(_05839_ ), .ZN(_05865_ ) );
AND2_X1 _13606_ ( .A1(_05865_ ), .A2(_05836_ ), .ZN(_05866_ ) );
NOR2_X1 _13607_ ( .A1(_05830_ ), .A2(_01944_ ), .ZN(_05867_ ) );
AND2_X1 _13608_ ( .A1(_05834_ ), .A2(\IF_ID_pc [15] ), .ZN(_05868_ ) );
AND2_X1 _13609_ ( .A1(_05831_ ), .A2(_05868_ ), .ZN(_05869_ ) );
OR3_X1 _13610_ ( .A1(_05866_ ), .A2(_05867_ ), .A3(_05869_ ), .ZN(_05870_ ) );
INV_X1 _13611_ ( .A(\IF_ID_pc [11] ), .ZN(_05871_ ) );
NOR2_X1 _13612_ ( .A1(_05850_ ), .A2(_05871_ ), .ZN(_05872_ ) );
AND2_X1 _13613_ ( .A1(_05847_ ), .A2(_05872_ ), .ZN(_05873_ ) );
AOI21_X1 _13614_ ( .A(_05873_ ), .B1(\IF_ID_pc [12] ), .B2(_05846_ ), .ZN(_05874_ ) );
INV_X1 _13615_ ( .A(\IF_ID_pc [10] ), .ZN(_05875_ ) );
NOR2_X1 _13616_ ( .A1(_05859_ ), .A2(_05875_ ), .ZN(_05876_ ) );
AND2_X1 _13617_ ( .A1(_05859_ ), .A2(_05875_ ), .ZN(_05877_ ) );
INV_X1 _13618_ ( .A(_05877_ ), .ZN(_05878_ ) );
INV_X1 _13619_ ( .A(\IF_ID_pc [9] ), .ZN(_05879_ ) );
NOR2_X1 _13620_ ( .A1(_05855_ ), .A2(_05879_ ), .ZN(_05880_ ) );
AOI21_X1 _13621_ ( .A(_05876_ ), .B1(_05878_ ), .B2(_05880_ ), .ZN(_05881_ ) );
INV_X1 _13622_ ( .A(_05852_ ), .ZN(_05882_ ) );
OAI21_X1 _13623_ ( .A(_05874_ ), .B1(_05881_ ), .B2(_05882_ ), .ZN(_05883_ ) );
AND2_X1 _13624_ ( .A1(_05883_ ), .A2(_05844_ ), .ZN(_05884_ ) );
NOR2_X1 _13625_ ( .A1(_05870_ ), .A2(_05884_ ), .ZN(_05885_ ) );
AND2_X1 _13626_ ( .A1(_05862_ ), .A2(_05885_ ), .ZN(_05886_ ) );
INV_X1 _13627_ ( .A(_05886_ ), .ZN(_05887_ ) );
AND3_X1 _13628_ ( .A1(_05762_ ), .A2(_05478_ ), .A3(\IF_ID_inst [19] ), .ZN(_05888_ ) );
MUX2_X1 _13629_ ( .A(_05888_ ), .B(_05833_ ), .S(_05822_ ), .Z(_05889_ ) );
XNOR2_X1 _13630_ ( .A(_05889_ ), .B(_02194_ ), .ZN(_05890_ ) );
AND3_X1 _13631_ ( .A1(_05762_ ), .A2(_05478_ ), .A3(\IF_ID_inst [18] ), .ZN(_05891_ ) );
MUX2_X1 _13632_ ( .A(_05891_ ), .B(_05833_ ), .S(_05822_ ), .Z(_05892_ ) );
XNOR2_X1 _13633_ ( .A(_05892_ ), .B(_02185_ ), .ZN(_05893_ ) );
AND3_X1 _13634_ ( .A1(_05762_ ), .A2(_05478_ ), .A3(\IF_ID_inst [17] ), .ZN(_05894_ ) );
MUX2_X1 _13635_ ( .A(_05894_ ), .B(_05833_ ), .S(_05822_ ), .Z(_05895_ ) );
XNOR2_X1 _13636_ ( .A(_05895_ ), .B(_02200_ ), .ZN(_05896_ ) );
AND2_X1 _13637_ ( .A1(_05893_ ), .A2(_05896_ ), .ZN(_05897_ ) );
AND4_X1 _13638_ ( .A1(_05765_ ), .A2(_05887_ ), .A3(_05890_ ), .A4(_05897_ ), .ZN(_05898_ ) );
AND2_X1 _13639_ ( .A1(_05892_ ), .A2(\IF_ID_pc [18] ), .ZN(_05899_ ) );
AND2_X1 _13640_ ( .A1(_05895_ ), .A2(\IF_ID_pc [17] ), .ZN(_05900_ ) );
OR2_X1 _13641_ ( .A1(_05899_ ), .A2(_05900_ ), .ZN(_05901_ ) );
NOR2_X1 _13642_ ( .A1(_05892_ ), .A2(\IF_ID_pc [18] ), .ZN(_05902_ ) );
INV_X1 _13643_ ( .A(_05902_ ), .ZN(_05903_ ) );
AND4_X1 _13644_ ( .A1(_05765_ ), .A2(_05901_ ), .A3(_05890_ ), .A4(_05903_ ), .ZN(_05904_ ) );
NOR3_X1 _13645_ ( .A1(_05761_ ), .A2(_02197_ ), .A3(_05763_ ), .ZN(_05905_ ) );
AND2_X1 _13646_ ( .A1(_05889_ ), .A2(\IF_ID_pc [19] ), .ZN(_05906_ ) );
AND2_X1 _13647_ ( .A1(_05765_ ), .A2(_05906_ ), .ZN(_05907_ ) );
OR3_X1 _13648_ ( .A1(_05904_ ), .A2(_05905_ ), .A3(_05907_ ), .ZN(_05908_ ) );
OR2_X1 _13649_ ( .A1(_05898_ ), .A2(_05908_ ), .ZN(_05909_ ) );
XNOR2_X1 _13650_ ( .A(_05764_ ), .B(_01932_ ), .ZN(_05910_ ) );
XNOR2_X1 _13651_ ( .A(_05764_ ), .B(_01939_ ), .ZN(_05911_ ) );
AND2_X1 _13652_ ( .A1(_05910_ ), .A2(_05911_ ), .ZN(_05912_ ) );
BUF_X4 _13653_ ( .A(_05764_ ), .Z(_05913_ ) );
XNOR2_X1 _13654_ ( .A(_05913_ ), .B(\IF_ID_pc [22] ), .ZN(_05914_ ) );
AND2_X1 _13655_ ( .A1(_05764_ ), .A2(\IF_ID_pc [21] ), .ZN(_05915_ ) );
NOR2_X1 _13656_ ( .A1(_05913_ ), .A2(\IF_ID_pc [21] ), .ZN(_05916_ ) );
NOR3_X1 _13657_ ( .A1(_05914_ ), .A2(_05915_ ), .A3(_05916_ ), .ZN(_05917_ ) );
AND3_X1 _13658_ ( .A1(_05909_ ), .A2(_05912_ ), .A3(_05917_ ), .ZN(_05918_ ) );
AND2_X1 _13659_ ( .A1(_05913_ ), .A2(\IF_ID_pc [22] ), .ZN(_05919_ ) );
OAI21_X1 _13660_ ( .A(_05912_ ), .B1(_05919_ ), .B2(_05915_ ), .ZN(_05920_ ) );
NAND2_X1 _13661_ ( .A1(_05913_ ), .A2(\IF_ID_pc [24] ), .ZN(_05921_ ) );
NAND2_X1 _13662_ ( .A1(_05913_ ), .A2(\IF_ID_pc [23] ), .ZN(_05922_ ) );
NAND3_X1 _13663_ ( .A1(_05920_ ), .A2(_05921_ ), .A3(_05922_ ), .ZN(_05923_ ) );
NOR2_X1 _13664_ ( .A1(_05918_ ), .A2(_05923_ ), .ZN(_05924_ ) );
XNOR2_X1 _13665_ ( .A(_05913_ ), .B(_02182_ ), .ZN(_05925_ ) );
XNOR2_X1 _13666_ ( .A(_05913_ ), .B(_01927_ ), .ZN(_05926_ ) );
AND2_X1 _13667_ ( .A1(_05925_ ), .A2(_05926_ ), .ZN(_05927_ ) );
INV_X1 _13668_ ( .A(_05927_ ), .ZN(_05928_ ) );
XNOR2_X1 _13669_ ( .A(_05913_ ), .B(_01987_ ), .ZN(_05929_ ) );
XNOR2_X1 _13670_ ( .A(_05913_ ), .B(_02171_ ), .ZN(_05930_ ) );
NAND2_X1 _13671_ ( .A1(_05929_ ), .A2(_05930_ ), .ZN(_05931_ ) );
NOR3_X1 _13672_ ( .A1(_05924_ ), .A2(_05928_ ), .A3(_05931_ ), .ZN(_05932_ ) );
BUF_X4 _13673_ ( .A(_05913_ ), .Z(_05933_ ) );
OAI21_X1 _13674_ ( .A(_05933_ ), .B1(\IF_ID_pc [28] ), .B2(\IF_ID_pc [27] ), .ZN(_05934_ ) );
OAI21_X1 _13675_ ( .A(_05933_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_05935_ ) );
OAI21_X1 _13676_ ( .A(_05934_ ), .B1(_05928_ ), .B2(_05935_ ), .ZN(_05936_ ) );
NOR2_X1 _13677_ ( .A1(_05932_ ), .A2(_05936_ ), .ZN(_05937_ ) );
XNOR2_X1 _13678_ ( .A(_05933_ ), .B(\IF_ID_pc [29] ), .ZN(_05938_ ) );
NOR2_X1 _13679_ ( .A1(_05937_ ), .A2(_05938_ ), .ZN(_05939_ ) );
NOR3_X1 _13680_ ( .A1(_05761_ ), .A2(_02161_ ), .A3(_05763_ ), .ZN(_05940_ ) );
NOR2_X1 _13681_ ( .A1(_05939_ ), .A2(_05940_ ), .ZN(_05941_ ) );
XNOR2_X1 _13682_ ( .A(_05933_ ), .B(\IF_ID_pc [30] ), .ZN(_05942_ ) );
OR2_X1 _13683_ ( .A1(_05941_ ), .A2(_05942_ ), .ZN(_05943_ ) );
AOI21_X1 _13684_ ( .A(_05758_ ), .B1(_05941_ ), .B2(_05942_ ), .ZN(_05944_ ) );
AOI221_X4 _13685_ ( .A(fanout_net_48 ), .B1(\myexu.pc_jump [30] ), .B2(_05758_ ), .C1(_05943_ ), .C2(_05944_ ), .ZN(_05945_ ) );
BUF_X4 _13686_ ( .A(_05754_ ), .Z(_05946_ ) );
NOR2_X1 _13687_ ( .A1(_05946_ ), .A2(\mtvec [30] ), .ZN(_05947_ ) );
NOR3_X1 _13688_ ( .A1(_05945_ ), .A2(fanout_net_5 ), .A3(_05947_ ), .ZN(_00282_ ) );
XNOR2_X1 _13689_ ( .A(_05933_ ), .B(_02062_ ), .ZN(_05948_ ) );
AND2_X1 _13690_ ( .A1(_05909_ ), .A2(_05948_ ), .ZN(_05949_ ) );
BUF_X4 _13691_ ( .A(_05758_ ), .Z(_05950_ ) );
NOR3_X1 _13692_ ( .A1(_05898_ ), .A2(_05948_ ), .A3(_05908_ ), .ZN(_05951_ ) );
NOR3_X1 _13693_ ( .A1(_05949_ ), .A2(_05950_ ), .A3(_05951_ ), .ZN(_05952_ ) );
BUF_X4 _13694_ ( .A(_05950_ ), .Z(_05953_ ) );
AOI211_X1 _13695_ ( .A(fanout_net_48 ), .B(_05952_ ), .C1(\myexu.pc_jump [21] ), .C2(_05953_ ), .ZN(_05954_ ) );
NOR2_X1 _13696_ ( .A1(_05946_ ), .A2(\mtvec [21] ), .ZN(_05955_ ) );
NOR3_X1 _13697_ ( .A1(_05954_ ), .A2(fanout_net_5 ), .A3(_05955_ ), .ZN(_00283_ ) );
AND2_X1 _13698_ ( .A1(_05828_ ), .A2(_05861_ ), .ZN(_05956_ ) );
OR2_X1 _13699_ ( .A1(_05956_ ), .A2(_05883_ ), .ZN(_05957_ ) );
AND2_X1 _13700_ ( .A1(_05957_ ), .A2(_05844_ ), .ZN(_05958_ ) );
OAI21_X1 _13701_ ( .A(_05896_ ), .B1(_05958_ ), .B2(_05870_ ), .ZN(_05959_ ) );
INV_X1 _13702_ ( .A(_05893_ ), .ZN(_05960_ ) );
NOR2_X1 _13703_ ( .A1(_05959_ ), .A2(_05960_ ), .ZN(_05961_ ) );
NAND2_X1 _13704_ ( .A1(_05901_ ), .A2(_05903_ ), .ZN(_05962_ ) );
INV_X1 _13705_ ( .A(_05962_ ), .ZN(_05963_ ) );
OAI21_X1 _13706_ ( .A(_05890_ ), .B1(_05961_ ), .B2(_05963_ ), .ZN(_05964_ ) );
INV_X1 _13707_ ( .A(_05906_ ), .ZN(_05965_ ) );
AND3_X1 _13708_ ( .A1(_05964_ ), .A2(_05965_ ), .A3(_05765_ ), .ZN(_05966_ ) );
AOI21_X1 _13709_ ( .A(_05765_ ), .B1(_05964_ ), .B2(_05965_ ), .ZN(_05967_ ) );
OR3_X1 _13710_ ( .A1(_05966_ ), .A2(_05967_ ), .A3(_05758_ ), .ZN(_05968_ ) );
BUF_X4 _13711_ ( .A(_05754_ ), .Z(_05969_ ) );
INV_X1 _13712_ ( .A(_05628_ ), .ZN(_05970_ ) );
BUF_X4 _13713_ ( .A(_05970_ ), .Z(_05971_ ) );
BUF_X4 _13714_ ( .A(_05971_ ), .Z(_05972_ ) );
OAI211_X1 _13715_ ( .A(_05968_ ), .B(_05969_ ), .C1(\myexu.pc_jump [20] ), .C2(_05972_ ), .ZN(_05973_ ) );
NAND2_X1 _13716_ ( .A1(\mtvec [20] ), .A2(fanout_net_48 ), .ZN(_05974_ ) );
AOI21_X1 _13717_ ( .A(fanout_net_5 ), .B1(_05973_ ), .B2(_05974_ ), .ZN(_00284_ ) );
NOR2_X1 _13718_ ( .A1(_05961_ ), .A2(_05963_ ), .ZN(_05975_ ) );
XOR2_X1 _13719_ ( .A(_05975_ ), .B(_05890_ ), .Z(_05976_ ) );
BUF_X4 _13720_ ( .A(_05971_ ), .Z(_05977_ ) );
NAND2_X1 _13721_ ( .A1(_05976_ ), .A2(_05977_ ), .ZN(_05978_ ) );
OAI211_X1 _13722_ ( .A(_05978_ ), .B(_05969_ ), .C1(\myexu.pc_jump [19] ), .C2(_05972_ ), .ZN(_05979_ ) );
NAND2_X1 _13723_ ( .A1(\mtvec [19] ), .A2(fanout_net_48 ), .ZN(_05980_ ) );
AOI21_X1 _13724_ ( .A(fanout_net_5 ), .B1(_05979_ ), .B2(_05980_ ), .ZN(_00285_ ) );
INV_X1 _13725_ ( .A(_05900_ ), .ZN(_05981_ ) );
AND3_X1 _13726_ ( .A1(_05959_ ), .A2(_05960_ ), .A3(_05981_ ), .ZN(_05982_ ) );
AOI21_X1 _13727_ ( .A(_05960_ ), .B1(_05959_ ), .B2(_05981_ ), .ZN(_05983_ ) );
NOR3_X1 _13728_ ( .A1(_05982_ ), .A2(_05983_ ), .A3(_05950_ ), .ZN(_05984_ ) );
AOI211_X1 _13729_ ( .A(fanout_net_48 ), .B(_05984_ ), .C1(\myexu.pc_jump [18] ), .C2(_05953_ ), .ZN(_05985_ ) );
NOR2_X1 _13730_ ( .A1(_05946_ ), .A2(\mtvec [18] ), .ZN(_05986_ ) );
NOR3_X1 _13731_ ( .A1(_05985_ ), .A2(fanout_net_5 ), .A3(_05986_ ), .ZN(_00286_ ) );
XOR2_X1 _13732_ ( .A(_05886_ ), .B(_05896_ ), .Z(_05987_ ) );
NAND2_X1 _13733_ ( .A1(_05987_ ), .A2(_05977_ ), .ZN(_05988_ ) );
OAI211_X1 _13734_ ( .A(_05988_ ), .B(_05969_ ), .C1(\myexu.pc_jump [17] ), .C2(_05972_ ), .ZN(_05989_ ) );
NAND2_X1 _13735_ ( .A1(\mtvec [17] ), .A2(fanout_net_48 ), .ZN(_05990_ ) );
AOI21_X1 _13736_ ( .A(fanout_net_5 ), .B1(_05989_ ), .B2(_05990_ ), .ZN(_00287_ ) );
AND3_X1 _13737_ ( .A1(_05957_ ), .A2(_05840_ ), .A3(_05843_ ), .ZN(_05991_ ) );
OAI21_X1 _13738_ ( .A(_05835_ ), .B1(_05991_ ), .B2(_05865_ ), .ZN(_05992_ ) );
INV_X1 _13739_ ( .A(_05868_ ), .ZN(_05993_ ) );
NAND2_X1 _13740_ ( .A1(_05992_ ), .A2(_05993_ ), .ZN(_05994_ ) );
XNOR2_X1 _13741_ ( .A(_05994_ ), .B(_05831_ ), .ZN(_05995_ ) );
NOR2_X1 _13742_ ( .A1(_05995_ ), .A2(_05950_ ), .ZN(_05996_ ) );
AOI211_X1 _13743_ ( .A(fanout_net_48 ), .B(_05996_ ), .C1(\myexu.pc_jump [16] ), .C2(_05953_ ), .ZN(_05997_ ) );
NOR2_X1 _13744_ ( .A1(_05946_ ), .A2(\mtvec [16] ), .ZN(_05998_ ) );
NOR3_X1 _13745_ ( .A1(_05997_ ), .A2(fanout_net_5 ), .A3(_05998_ ), .ZN(_00288_ ) );
OR3_X1 _13746_ ( .A1(_05991_ ), .A2(_05835_ ), .A3(_05865_ ), .ZN(_05999_ ) );
AND3_X1 _13747_ ( .A1(_05999_ ), .A2(_05970_ ), .A3(_05992_ ), .ZN(_06000_ ) );
AOI211_X1 _13748_ ( .A(fanout_net_48 ), .B(_06000_ ), .C1(\myexu.pc_jump [15] ), .C2(_05953_ ), .ZN(_06001_ ) );
NOR2_X1 _13749_ ( .A1(_05946_ ), .A2(\mtvec [15] ), .ZN(_06002_ ) );
NOR3_X1 _13750_ ( .A1(_06001_ ), .A2(fanout_net_5 ), .A3(_06002_ ), .ZN(_00289_ ) );
AND2_X1 _13751_ ( .A1(_05957_ ), .A2(_05843_ ), .ZN(_06003_ ) );
OR3_X1 _13752_ ( .A1(_06003_ ), .A2(_05863_ ), .A3(_05840_ ), .ZN(_06004_ ) );
OAI21_X1 _13753_ ( .A(_05840_ ), .B1(_06003_ ), .B2(_05863_ ), .ZN(_06005_ ) );
AND3_X1 _13754_ ( .A1(_06004_ ), .A2(_05970_ ), .A3(_06005_ ), .ZN(_06006_ ) );
AOI211_X1 _13755_ ( .A(fanout_net_48 ), .B(_06006_ ), .C1(\myexu.pc_jump [14] ), .C2(_05953_ ), .ZN(_06007_ ) );
NOR2_X1 _13756_ ( .A1(_05946_ ), .A2(\mtvec [14] ), .ZN(_06008_ ) );
NOR3_X1 _13757_ ( .A1(_06007_ ), .A2(fanout_net_5 ), .A3(_06008_ ), .ZN(_00290_ ) );
NOR3_X1 _13758_ ( .A1(_05956_ ), .A2(_05843_ ), .A3(_05883_ ), .ZN(_06009_ ) );
NOR3_X1 _13759_ ( .A1(_06003_ ), .A2(_05950_ ), .A3(_06009_ ), .ZN(_06010_ ) );
AOI211_X1 _13760_ ( .A(fanout_net_48 ), .B(_06010_ ), .C1(\myexu.pc_jump [13] ), .C2(_05953_ ), .ZN(_06011_ ) );
NOR2_X1 _13761_ ( .A1(_05946_ ), .A2(\mtvec [13] ), .ZN(_06012_ ) );
NOR3_X1 _13762_ ( .A1(_06011_ ), .A2(fanout_net_5 ), .A3(_06012_ ), .ZN(_00291_ ) );
AND2_X1 _13763_ ( .A1(_05856_ ), .A2(_05860_ ), .ZN(_06013_ ) );
NAND2_X1 _13764_ ( .A1(_05828_ ), .A2(_06013_ ), .ZN(_06014_ ) );
AND2_X1 _13765_ ( .A1(_06014_ ), .A2(_05881_ ), .ZN(_06015_ ) );
INV_X1 _13766_ ( .A(_05851_ ), .ZN(_06016_ ) );
OR2_X1 _13767_ ( .A1(_06015_ ), .A2(_06016_ ), .ZN(_06017_ ) );
INV_X1 _13768_ ( .A(_05872_ ), .ZN(_06018_ ) );
AND3_X1 _13769_ ( .A1(_06017_ ), .A2(_06018_ ), .A3(_05847_ ), .ZN(_06019_ ) );
AOI21_X1 _13770_ ( .A(_05847_ ), .B1(_06017_ ), .B2(_06018_ ), .ZN(_06020_ ) );
OR3_X1 _13771_ ( .A1(_06019_ ), .A2(_06020_ ), .A3(_05758_ ), .ZN(_06021_ ) );
OAI211_X1 _13772_ ( .A(_06021_ ), .B(_05969_ ), .C1(\myexu.pc_jump [12] ), .C2(_05972_ ), .ZN(_06022_ ) );
NAND2_X1 _13773_ ( .A1(\mtvec [12] ), .A2(fanout_net_48 ), .ZN(_06023_ ) );
AOI21_X1 _13774_ ( .A(fanout_net_5 ), .B1(_06022_ ), .B2(_06023_ ), .ZN(_00292_ ) );
AND2_X1 _13775_ ( .A1(_05937_ ), .A2(_05938_ ), .ZN(_06024_ ) );
OAI21_X1 _13776_ ( .A(_05971_ ), .B1(_06024_ ), .B2(_05939_ ), .ZN(_06025_ ) );
OAI211_X1 _13777_ ( .A(_06025_ ), .B(_05969_ ), .C1(\myexu.pc_jump [29] ), .C2(_05972_ ), .ZN(_06026_ ) );
NAND2_X1 _13778_ ( .A1(\mtvec [29] ), .A2(fanout_net_48 ), .ZN(_06027_ ) );
AOI21_X1 _13779_ ( .A(fanout_net_5 ), .B1(_06026_ ), .B2(_06027_ ), .ZN(_00293_ ) );
OAI21_X1 _13780_ ( .A(_05970_ ), .B1(_06015_ ), .B2(_06016_ ), .ZN(_06028_ ) );
AOI21_X1 _13781_ ( .A(_06028_ ), .B1(_06016_ ), .B2(_06015_ ), .ZN(_06029_ ) );
AOI211_X1 _13782_ ( .A(fanout_net_48 ), .B(_06029_ ), .C1(\myexu.pc_jump [11] ), .C2(_05953_ ), .ZN(_06030_ ) );
NOR2_X1 _13783_ ( .A1(_05946_ ), .A2(\mtvec [11] ), .ZN(_06031_ ) );
NOR3_X1 _13784_ ( .A1(_06030_ ), .A2(fanout_net_5 ), .A3(_06031_ ), .ZN(_00294_ ) );
INV_X1 _13785_ ( .A(_05856_ ), .ZN(_06032_ ) );
AOI21_X1 _13786_ ( .A(_06032_ ), .B1(_05825_ ), .B2(_05827_ ), .ZN(_06033_ ) );
NOR2_X1 _13787_ ( .A1(_06033_ ), .A2(_05880_ ), .ZN(_06034_ ) );
INV_X1 _13788_ ( .A(_06034_ ), .ZN(_06035_ ) );
OAI21_X1 _13789_ ( .A(_05970_ ), .B1(_06035_ ), .B2(_05860_ ), .ZN(_06036_ ) );
AOI21_X1 _13790_ ( .A(_06036_ ), .B1(_06035_ ), .B2(_05860_ ), .ZN(_06037_ ) );
AOI211_X1 _13791_ ( .A(fanout_net_48 ), .B(_06037_ ), .C1(\myexu.pc_jump [10] ), .C2(_05953_ ), .ZN(_06038_ ) );
NOR2_X1 _13792_ ( .A1(_05946_ ), .A2(\mtvec [10] ), .ZN(_06039_ ) );
NOR3_X1 _13793_ ( .A1(_06038_ ), .A2(fanout_net_5 ), .A3(_06039_ ), .ZN(_00295_ ) );
AND3_X1 _13794_ ( .A1(_05825_ ), .A2(_05827_ ), .A3(_06032_ ), .ZN(_06040_ ) );
NOR3_X1 _13795_ ( .A1(_06040_ ), .A2(_06033_ ), .A3(_05950_ ), .ZN(_06041_ ) );
AOI211_X1 _13796_ ( .A(fanout_net_48 ), .B(_06041_ ), .C1(\myexu.pc_jump [9] ), .C2(_05953_ ), .ZN(_06042_ ) );
NOR2_X1 _13797_ ( .A1(_05969_ ), .A2(\mtvec [9] ), .ZN(_06043_ ) );
NOR3_X1 _13798_ ( .A1(_06042_ ), .A2(fanout_net_5 ), .A3(_06043_ ), .ZN(_00296_ ) );
NOR2_X1 _13799_ ( .A1(_05818_ ), .A2(_05819_ ), .ZN(_06044_ ) );
XNOR2_X1 _13800_ ( .A(_05823_ ), .B(_05826_ ), .ZN(_06045_ ) );
OR2_X1 _13801_ ( .A1(_06044_ ), .A2(_06045_ ), .ZN(_06046_ ) );
AOI21_X1 _13802_ ( .A(_05758_ ), .B1(_06044_ ), .B2(_06045_ ), .ZN(_06047_ ) );
AOI221_X4 _13803_ ( .A(fanout_net_48 ), .B1(\myexu.pc_jump [8] ), .B2(_05758_ ), .C1(_06046_ ), .C2(_06047_ ), .ZN(_06048_ ) );
NOR2_X1 _13804_ ( .A1(_05969_ ), .A2(\mtvec [8] ), .ZN(_06049_ ) );
NOR3_X1 _13805_ ( .A1(_06048_ ), .A2(fanout_net_5 ), .A3(_06049_ ), .ZN(_00297_ ) );
NOR3_X1 _13806_ ( .A1(_05811_ ), .A2(_05770_ ), .A3(_05816_ ), .ZN(_06050_ ) );
OAI21_X1 _13807_ ( .A(_05971_ ), .B1(_05818_ ), .B2(_06050_ ), .ZN(_06051_ ) );
OAI211_X1 _13808_ ( .A(_06051_ ), .B(_05969_ ), .C1(\myexu.pc_jump [7] ), .C2(_05972_ ), .ZN(_06052_ ) );
NAND2_X1 _13809_ ( .A1(\mtvec [7] ), .A2(fanout_net_48 ), .ZN(_06053_ ) );
AOI21_X1 _13810_ ( .A(fanout_net_5 ), .B1(_06052_ ), .B2(_06053_ ), .ZN(_00298_ ) );
OAI21_X1 _13811_ ( .A(_05806_ ), .B1(_05797_ ), .B2(_05800_ ), .ZN(_06054_ ) );
AND3_X1 _13812_ ( .A1(_06054_ ), .A2(_05813_ ), .A3(_05810_ ), .ZN(_06055_ ) );
AOI21_X1 _13813_ ( .A(_05810_ ), .B1(_06054_ ), .B2(_05813_ ), .ZN(_06056_ ) );
OR3_X1 _13814_ ( .A1(_06055_ ), .A2(_06056_ ), .A3(_05758_ ), .ZN(_06057_ ) );
OAI211_X1 _13815_ ( .A(_06057_ ), .B(_05755_ ), .C1(\myexu.pc_jump [6] ), .C2(_05972_ ), .ZN(_06058_ ) );
NAND2_X1 _13816_ ( .A1(\mtvec [6] ), .A2(fanout_net_48 ), .ZN(_06059_ ) );
AOI21_X1 _13817_ ( .A(fanout_net_6 ), .B1(_06058_ ), .B2(_06059_ ), .ZN(_00299_ ) );
XOR2_X1 _13818_ ( .A(_05801_ ), .B(_05806_ ), .Z(_06060_ ) );
NAND2_X1 _13819_ ( .A1(_06060_ ), .A2(_05977_ ), .ZN(_06061_ ) );
OAI211_X1 _13820_ ( .A(_06061_ ), .B(_05755_ ), .C1(\myexu.pc_jump [5] ), .C2(_05972_ ), .ZN(_06062_ ) );
NAND2_X1 _13821_ ( .A1(\mtvec [5] ), .A2(fanout_net_48 ), .ZN(_06063_ ) );
AOI21_X1 _13822_ ( .A(fanout_net_6 ), .B1(_06062_ ), .B2(_06063_ ), .ZN(_00300_ ) );
OR2_X1 _13823_ ( .A1(_05782_ ), .A2(_05787_ ), .ZN(_06064_ ) );
AND3_X1 _13824_ ( .A1(_06064_ ), .A2(_05799_ ), .A3(_05795_ ), .ZN(_06065_ ) );
AOI21_X1 _13825_ ( .A(_05795_ ), .B1(_06064_ ), .B2(_05799_ ), .ZN(_06066_ ) );
OR3_X1 _13826_ ( .A1(_06065_ ), .A2(_06066_ ), .A3(_05758_ ), .ZN(_06067_ ) );
OAI211_X1 _13827_ ( .A(_06067_ ), .B(_05754_ ), .C1(\myexu.pc_jump [4] ), .C2(_05970_ ), .ZN(_06068_ ) );
NAND2_X1 _13828_ ( .A1(\mtvec [4] ), .A2(fanout_net_48 ), .ZN(_06069_ ) );
AOI21_X1 _13829_ ( .A(fanout_net_6 ), .B1(_06068_ ), .B2(_06069_ ), .ZN(_00301_ ) );
AND2_X1 _13830_ ( .A1(\mtvec [3] ), .A2(fanout_net_48 ), .ZN(_06070_ ) );
XOR2_X1 _13831_ ( .A(_05782_ ), .B(_05787_ ), .Z(_06071_ ) );
MUX2_X1 _13832_ ( .A(\myexu.pc_jump [3] ), .B(_06071_ ), .S(_05970_ ), .Z(_06072_ ) );
AOI21_X1 _13833_ ( .A(_06070_ ), .B1(_06072_ ), .B2(_05946_ ), .ZN(_06073_ ) );
NOR2_X1 _13834_ ( .A1(_06073_ ), .A2(fanout_net_6 ), .ZN(_00302_ ) );
AND2_X1 _13835_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
NOR2_X1 _13836_ ( .A1(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A2(fanout_net_6 ), .ZN(_06074_ ) );
NOR2_X1 _13837_ ( .A1(_00301_ ), .A2(_06074_ ), .ZN(_06075_ ) );
BUF_X4 _13838_ ( .A(_05793_ ), .Z(_06076_ ) );
BUF_X4 _13839_ ( .A(_06076_ ), .Z(_06077_ ) );
BUF_X2 _13840_ ( .A(_06077_ ), .Z(_06078_ ) );
INV_X1 _13841_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_06079_ ) );
AOI21_X1 _13842_ ( .A(_06075_ ), .B1(_06078_ ), .B2(_06079_ ), .ZN(_00303_ ) );
NOR2_X1 _13843_ ( .A1(_05775_ ), .A2(_05780_ ), .ZN(_06080_ ) );
NOR3_X1 _13844_ ( .A1(_05950_ ), .A2(_05781_ ), .A3(_06080_ ), .ZN(_06081_ ) );
AOI211_X1 _13845_ ( .A(fanout_net_48 ), .B(_06081_ ), .C1(\myexu.pc_jump [2] ), .C2(_05950_ ), .ZN(_06082_ ) );
NOR2_X1 _13846_ ( .A1(_05969_ ), .A2(\mtvec [2] ), .ZN(_06083_ ) );
NOR3_X1 _13847_ ( .A1(_06082_ ), .A2(fanout_net_6 ), .A3(_06083_ ), .ZN(_00304_ ) );
AOI211_X1 _13848_ ( .A(_06070_ ), .B(_06079_ ), .C1(_06072_ ), .C2(_05754_ ), .ZN(_06084_ ) );
INV_X1 _13849_ ( .A(fanout_net_12 ), .ZN(_06085_ ) );
BUF_X4 _13850_ ( .A(_06085_ ), .Z(_06086_ ) );
BUF_X2 _13851_ ( .A(_06086_ ), .Z(_06087_ ) );
AOI211_X1 _13852_ ( .A(fanout_net_6 ), .B(_06084_ ), .C1(_06087_ ), .C2(_06079_ ), .ZN(_00305_ ) );
NOR2_X1 _13853_ ( .A1(_05924_ ), .A2(_05931_ ), .ZN(_06088_ ) );
INV_X1 _13854_ ( .A(_05935_ ), .ZN(_06089_ ) );
OAI21_X1 _13855_ ( .A(_05926_ ), .B1(_06088_ ), .B2(_06089_ ), .ZN(_06090_ ) );
NAND2_X1 _13856_ ( .A1(_05933_ ), .A2(\IF_ID_pc [27] ), .ZN(_06091_ ) );
NAND2_X1 _13857_ ( .A1(_06090_ ), .A2(_06091_ ), .ZN(_06092_ ) );
XNOR2_X1 _13858_ ( .A(_06092_ ), .B(_05925_ ), .ZN(_06093_ ) );
NAND2_X1 _13859_ ( .A1(_06093_ ), .A2(_05971_ ), .ZN(_06094_ ) );
OAI211_X1 _13860_ ( .A(_06094_ ), .B(_05755_ ), .C1(\myexu.pc_jump [28] ), .C2(_05977_ ), .ZN(_06095_ ) );
NAND2_X1 _13861_ ( .A1(\mtvec [28] ), .A2(fanout_net_48 ), .ZN(_06096_ ) );
AOI21_X1 _13862_ ( .A(fanout_net_6 ), .B1(_06095_ ), .B2(_06096_ ), .ZN(_00306_ ) );
XNOR2_X1 _13863_ ( .A(_05779_ ), .B(\IF_ID_pc [1] ), .ZN(_06097_ ) );
AOI21_X1 _13864_ ( .A(_06097_ ), .B1(_05753_ ), .B2(check_quest ), .ZN(_06098_ ) );
AOI211_X1 _13865_ ( .A(fanout_net_48 ), .B(_06098_ ), .C1(\myexu.pc_jump [1] ), .C2(_05950_ ), .ZN(_06099_ ) );
NOR2_X1 _13866_ ( .A1(_05969_ ), .A2(\mtvec [1] ), .ZN(_06100_ ) );
NOR3_X1 _13867_ ( .A1(_06099_ ), .A2(fanout_net_6 ), .A3(_06100_ ), .ZN(_00307_ ) );
NOR2_X1 _13868_ ( .A1(_06088_ ), .A2(_06089_ ), .ZN(_06101_ ) );
XOR2_X1 _13869_ ( .A(_06101_ ), .B(_05926_ ), .Z(_06102_ ) );
NAND2_X1 _13870_ ( .A1(_06102_ ), .A2(_05971_ ), .ZN(_06103_ ) );
OAI211_X1 _13871_ ( .A(_06103_ ), .B(_05755_ ), .C1(\myexu.pc_jump [27] ), .C2(_05977_ ), .ZN(_06104_ ) );
NAND2_X1 _13872_ ( .A1(\mtvec [27] ), .A2(fanout_net_48 ), .ZN(_06105_ ) );
AOI21_X1 _13873_ ( .A(fanout_net_6 ), .B1(_06104_ ), .B2(_06105_ ), .ZN(_00308_ ) );
OAI21_X1 _13874_ ( .A(_05930_ ), .B1(_05918_ ), .B2(_05923_ ), .ZN(_06106_ ) );
NAND2_X1 _13875_ ( .A1(_05933_ ), .A2(\IF_ID_pc [25] ), .ZN(_06107_ ) );
AND3_X1 _13876_ ( .A1(_06106_ ), .A2(_06107_ ), .A3(_05929_ ), .ZN(_06108_ ) );
AOI21_X1 _13877_ ( .A(_05929_ ), .B1(_06106_ ), .B2(_06107_ ), .ZN(_06109_ ) );
OR3_X1 _13878_ ( .A1(_06108_ ), .A2(_06109_ ), .A3(_05758_ ), .ZN(_06110_ ) );
OAI211_X1 _13879_ ( .A(_06110_ ), .B(_05755_ ), .C1(\myexu.pc_jump [26] ), .C2(_05977_ ), .ZN(_06111_ ) );
NAND2_X1 _13880_ ( .A1(\mtvec [26] ), .A2(fanout_net_48 ), .ZN(_06112_ ) );
AOI21_X1 _13881_ ( .A(fanout_net_6 ), .B1(_06111_ ), .B2(_06112_ ), .ZN(_00309_ ) );
XOR2_X1 _13882_ ( .A(_05924_ ), .B(_05930_ ), .Z(_06113_ ) );
NAND2_X1 _13883_ ( .A1(_06113_ ), .A2(_05971_ ), .ZN(_06114_ ) );
OAI211_X1 _13884_ ( .A(_06114_ ), .B(_05755_ ), .C1(\myexu.pc_jump [25] ), .C2(_05977_ ), .ZN(_06115_ ) );
NAND2_X1 _13885_ ( .A1(\mtvec [25] ), .A2(fanout_net_48 ), .ZN(_06116_ ) );
AOI21_X1 _13886_ ( .A(fanout_net_6 ), .B1(_06115_ ), .B2(_06116_ ), .ZN(_00310_ ) );
OAI21_X1 _13887_ ( .A(_05917_ ), .B1(_05898_ ), .B2(_05908_ ), .ZN(_06117_ ) );
OAI21_X1 _13888_ ( .A(_05933_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_06118_ ) );
NAND2_X1 _13889_ ( .A1(_06117_ ), .A2(_06118_ ), .ZN(_06119_ ) );
NAND2_X1 _13890_ ( .A1(_06119_ ), .A2(_05911_ ), .ZN(_06120_ ) );
NAND2_X1 _13891_ ( .A1(_06120_ ), .A2(_05922_ ), .ZN(_06121_ ) );
XNOR2_X1 _13892_ ( .A(_06121_ ), .B(_05910_ ), .ZN(_06122_ ) );
NAND2_X1 _13893_ ( .A1(_06122_ ), .A2(_05971_ ), .ZN(_06123_ ) );
OAI211_X1 _13894_ ( .A(_06123_ ), .B(_05755_ ), .C1(\myexu.pc_jump [24] ), .C2(_05977_ ), .ZN(_06124_ ) );
NAND2_X1 _13895_ ( .A1(\mtvec [24] ), .A2(\myifu.to_reset ), .ZN(_06125_ ) );
AOI21_X1 _13896_ ( .A(fanout_net_6 ), .B1(_06124_ ), .B2(_06125_ ), .ZN(_00311_ ) );
XNOR2_X1 _13897_ ( .A(_06119_ ), .B(_05911_ ), .ZN(_06126_ ) );
NAND2_X1 _13898_ ( .A1(_06126_ ), .A2(_05971_ ), .ZN(_06127_ ) );
OAI211_X1 _13899_ ( .A(_06127_ ), .B(_05755_ ), .C1(\myexu.pc_jump [23] ), .C2(_05977_ ), .ZN(_06128_ ) );
NAND2_X1 _13900_ ( .A1(\mtvec [23] ), .A2(\myifu.to_reset ), .ZN(_06129_ ) );
AOI21_X1 _13901_ ( .A(fanout_net_6 ), .B1(_06128_ ), .B2(_06129_ ), .ZN(_00312_ ) );
OR3_X1 _13902_ ( .A1(_05949_ ), .A2(_05915_ ), .A3(_05914_ ), .ZN(_06130_ ) );
OAI21_X1 _13903_ ( .A(_05914_ ), .B1(_05949_ ), .B2(_05915_ ), .ZN(_06131_ ) );
NAND3_X1 _13904_ ( .A1(_06130_ ), .A2(_05971_ ), .A3(_06131_ ), .ZN(_06132_ ) );
OAI211_X1 _13905_ ( .A(_06132_ ), .B(_05755_ ), .C1(\myexu.pc_jump [22] ), .C2(_05977_ ), .ZN(_06133_ ) );
NAND2_X1 _13906_ ( .A1(\mtvec [22] ), .A2(\myifu.to_reset ), .ZN(_06134_ ) );
AOI21_X1 _13907_ ( .A(fanout_net_6 ), .B1(_06133_ ), .B2(_06134_ ), .ZN(_00313_ ) );
NAND2_X1 _13908_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_06135_ ) );
OR3_X1 _13909_ ( .A1(_05937_ ), .A2(_05938_ ), .A3(_05942_ ), .ZN(_06136_ ) );
OAI21_X1 _13910_ ( .A(_05933_ ), .B1(\IF_ID_pc [30] ), .B2(\IF_ID_pc [29] ), .ZN(_06137_ ) );
AND2_X1 _13911_ ( .A1(_06136_ ), .A2(_06137_ ), .ZN(_06138_ ) );
XOR2_X1 _13912_ ( .A(_05933_ ), .B(\IF_ID_pc [31] ), .Z(_06139_ ) );
OR2_X1 _13913_ ( .A1(_06138_ ), .A2(_06139_ ), .ZN(_06140_ ) );
AOI21_X1 _13914_ ( .A(_05950_ ), .B1(_06138_ ), .B2(_06139_ ), .ZN(_06141_ ) );
AND2_X1 _13915_ ( .A1(_06140_ ), .A2(_06141_ ), .ZN(_06142_ ) );
OAI21_X1 _13916_ ( .A(_05754_ ), .B1(_05972_ ), .B2(\myexu.pc_jump [31] ), .ZN(_06143_ ) );
OAI211_X1 _13917_ ( .A(_01794_ ), .B(_06135_ ), .C1(_06142_ ), .C2(_06143_ ), .ZN(_00314_ ) );
OR2_X1 _13918_ ( .A1(_02208_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .ZN(_06144_ ) );
NAND2_X1 _13919_ ( .A1(_02208_ ), .A2(io_master_rvalid ), .ZN(_06145_ ) );
NAND2_X2 _13920_ ( .A1(_06144_ ), .A2(_06145_ ), .ZN(_06146_ ) );
NOR2_X1 _13921_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_06147_ ) );
NOR2_X1 _13922_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_06148_ ) );
INV_X1 _13923_ ( .A(\io_master_rid [1] ), .ZN(_06149_ ) );
NAND4_X1 _13924_ ( .A1(_06147_ ), .A2(_06148_ ), .A3(_06149_ ), .A4(\io_master_rid [0] ), .ZN(_06150_ ) );
AOI21_X1 _13925_ ( .A(_02156_ ), .B1(_02208_ ), .B2(_06150_ ), .ZN(_06151_ ) );
AND2_X1 _13926_ ( .A1(_06146_ ), .A2(_06151_ ), .ZN(_06152_ ) );
BUF_X4 _13927_ ( .A(_06152_ ), .Z(_06153_ ) );
OR2_X1 _13928_ ( .A1(_02207_ ), .A2(io_master_rlast ), .ZN(_06154_ ) );
NAND2_X1 _13929_ ( .A1(_06153_ ), .A2(_06154_ ), .ZN(_06155_ ) );
INV_X1 _13930_ ( .A(\myifu.tmp_offset [2] ), .ZN(_06156_ ) );
NAND3_X1 _13931_ ( .A1(_06155_ ), .A2(_01794_ ), .A3(_06156_ ), .ZN(_06157_ ) );
INV_X1 _13932_ ( .A(_06157_ ), .ZN(_00315_ ) );
NOR3_X1 _13933_ ( .A1(fanout_net_6 ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00316_ ) );
AND3_X1 _13934_ ( .A1(_02249_ ), .A2(_05629_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_06158_ ) );
INV_X1 _13935_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_06159_ ) );
MUX2_X1 _13936_ ( .A(_02249_ ), .B(_06159_ ), .S(\myifu.to_reset ), .Z(_06160_ ) );
AOI211_X1 _13937_ ( .A(fanout_net_6 ), .B(_06158_ ), .C1(_06160_ ), .C2(\myifu.state [1] ), .ZN(_00317_ ) );
AND2_X1 _13938_ ( .A1(_02279_ ), .A2(\EX_LS_pc [2] ), .ZN(_00318_ ) );
INV_X1 _13939_ ( .A(\mylsu.state [3] ), .ZN(_06161_ ) );
BUF_X4 _13940_ ( .A(_06161_ ), .Z(_06162_ ) );
NOR3_X1 _13941_ ( .A1(_06162_ ), .A2(fanout_net_6 ), .A3(excp_written ), .ZN(_00319_ ) );
AOI21_X1 _13942_ ( .A(\LS_WB_waddr_csreg [11] ), .B1(_05397_ ), .B2(\EX_LS_flag [2] ), .ZN(_06163_ ) );
INV_X1 _13943_ ( .A(_02132_ ), .ZN(_06164_ ) );
NOR2_X1 _13944_ ( .A1(_02141_ ), .A2(_06164_ ), .ZN(_06165_ ) );
NOR2_X1 _13945_ ( .A1(\EX_LS_flag [2] ), .A2(\EX_LS_flag [1] ), .ZN(_06166_ ) );
NOR2_X1 _13946_ ( .A1(_02131_ ), .A2(_06166_ ), .ZN(_06167_ ) );
NOR2_X1 _13947_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_06168_ ) );
AND2_X2 _13948_ ( .A1(_06168_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_06169_ ) );
NOR2_X1 _13949_ ( .A1(_06167_ ), .A2(_06169_ ), .ZN(_06170_ ) );
INV_X1 _13950_ ( .A(_06170_ ), .ZN(_06171_ ) );
OR2_X2 _13951_ ( .A1(_06165_ ), .A2(_06171_ ), .ZN(_06172_ ) );
BUF_X4 _13952_ ( .A(_06172_ ), .Z(_06173_ ) );
INV_X1 _13953_ ( .A(\EX_LS_dest_csreg_mem [11] ), .ZN(_06174_ ) );
AOI211_X1 _13954_ ( .A(_06163_ ), .B(_06173_ ), .C1(_06174_ ), .C2(_04715_ ), .ZN(_00320_ ) );
NOR2_X1 _13955_ ( .A1(_06165_ ), .A2(_06169_ ), .ZN(_06175_ ) );
INV_X1 _13956_ ( .A(_06175_ ), .ZN(_06176_ ) );
NAND3_X1 _13957_ ( .A1(_05397_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_06177_ ) );
BUF_X4 _13958_ ( .A(_02105_ ), .Z(_06178_ ) );
NAND2_X1 _13959_ ( .A1(_06178_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06179_ ) );
AOI211_X1 _13960_ ( .A(_05393_ ), .B(_06176_ ), .C1(_06177_ ), .C2(_06179_ ), .ZN(_00321_ ) );
NAND3_X1 _13961_ ( .A1(_05397_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_06180_ ) );
NAND2_X1 _13962_ ( .A1(_06178_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06181_ ) );
AOI211_X1 _13963_ ( .A(_05393_ ), .B(_06176_ ), .C1(_06180_ ), .C2(_06181_ ), .ZN(_00322_ ) );
NAND3_X1 _13964_ ( .A1(_05397_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_06182_ ) );
NAND2_X1 _13965_ ( .A1(_06178_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_06183_ ) );
AOI211_X1 _13966_ ( .A(_05393_ ), .B(_06176_ ), .C1(_06182_ ), .C2(_06183_ ), .ZN(_00323_ ) );
NAND3_X1 _13967_ ( .A1(_05397_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_06184_ ) );
NAND2_X1 _13968_ ( .A1(_06178_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06185_ ) );
AOI211_X1 _13969_ ( .A(_05393_ ), .B(_06176_ ), .C1(_06184_ ), .C2(_06185_ ), .ZN(_00324_ ) );
NAND3_X1 _13970_ ( .A1(_05397_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_06186_ ) );
NAND2_X1 _13971_ ( .A1(_06178_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_06187_ ) );
AOI211_X1 _13972_ ( .A(_05393_ ), .B(_06176_ ), .C1(_06186_ ), .C2(_06187_ ), .ZN(_00325_ ) );
NAND3_X1 _13973_ ( .A1(_05397_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_06188_ ) );
NAND2_X1 _13974_ ( .A1(_06178_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_06189_ ) );
AOI211_X1 _13975_ ( .A(_05393_ ), .B(_06176_ ), .C1(_06188_ ), .C2(_06189_ ), .ZN(_00326_ ) );
NAND3_X1 _13976_ ( .A1(_05397_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_flag [2] ), .ZN(_06190_ ) );
NAND2_X1 _13977_ ( .A1(_06178_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_06191_ ) );
AOI211_X1 _13978_ ( .A(_05393_ ), .B(_06176_ ), .C1(_06190_ ), .C2(_06191_ ), .ZN(_00327_ ) );
AND4_X1 _13979_ ( .A1(_03378_ ), .A2(_02327_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06192_ ) );
NOR2_X1 _13980_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_06193_ ) );
OAI211_X1 _13981_ ( .A(_06175_ ), .B(_05394_ ), .C1(_06192_ ), .C2(_06193_ ), .ZN(_00328_ ) );
AND4_X1 _13982_ ( .A1(_03379_ ), .A2(_02327_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06194_ ) );
NOR2_X1 _13983_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06195_ ) );
OAI211_X1 _13984_ ( .A(_06175_ ), .B(_05394_ ), .C1(_06194_ ), .C2(_06195_ ), .ZN(_00329_ ) );
INV_X1 _13985_ ( .A(\EX_LS_dest_csreg_mem [6] ), .ZN(_06196_ ) );
AND4_X1 _13986_ ( .A1(_06196_ ), .A2(_02327_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06197_ ) );
NOR2_X1 _13987_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06198_ ) );
OAI211_X1 _13988_ ( .A(_06175_ ), .B(_05394_ ), .C1(_06197_ ), .C2(_06198_ ), .ZN(_00330_ ) );
INV_X1 _13989_ ( .A(fanout_net_7 ), .ZN(_06199_ ) );
AND4_X1 _13990_ ( .A1(_06199_ ), .A2(_02327_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_06200_ ) );
NOR2_X1 _13991_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_06201_ ) );
OAI211_X1 _13992_ ( .A(_06175_ ), .B(_05394_ ), .C1(_06200_ ), .C2(_06201_ ), .ZN(_00331_ ) );
NOR4_X1 _13993_ ( .A1(fanout_net_6 ), .A2(\mylsu.state [3] ), .A3(\mylsu.state [1] ), .A4(excp_written ), .ZN(_06202_ ) );
INV_X1 _13994_ ( .A(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06203_ ) );
NAND2_X1 _13995_ ( .A1(_06202_ ), .A2(_06203_ ), .ZN(_06204_ ) );
OAI21_X1 _13996_ ( .A(_02130_ ), .B1(_02251_ ), .B2(_02252_ ), .ZN(_06205_ ) );
INV_X1 _13997_ ( .A(_02255_ ), .ZN(_06206_ ) );
OR2_X1 _13998_ ( .A1(_06205_ ), .A2(_06206_ ), .ZN(_06207_ ) );
AOI221_X4 _13999_ ( .A(_06169_ ), .B1(_06207_ ), .B2(\EX_LS_flag [2] ), .C1(_02258_ ), .C2(_02132_ ), .ZN(_06208_ ) );
AOI21_X1 _14000_ ( .A(_06204_ ), .B1(_06208_ ), .B2(_02129_ ), .ZN(_00332_ ) );
INV_X1 _14001_ ( .A(_02129_ ), .ZN(_06209_ ) );
NOR2_X1 _14002_ ( .A1(_02131_ ), .A2(_02105_ ), .ZN(_06210_ ) );
AOI21_X1 _14003_ ( .A(_06209_ ), .B1(_06210_ ), .B2(_06207_ ), .ZN(_06211_ ) );
AOI21_X1 _14004_ ( .A(_06204_ ), .B1(_06211_ ), .B2(_06175_ ), .ZN(_00333_ ) );
NOR2_X1 _14005_ ( .A1(_02253_ ), .A2(_06206_ ), .ZN(_06212_ ) );
AND2_X1 _14006_ ( .A1(_02119_ ), .A2(\EX_LS_flag [2] ), .ZN(_06213_ ) );
AND4_X1 _14007_ ( .A1(_06203_ ), .A2(_06212_ ), .A3(_06213_ ), .A4(_06202_ ), .ZN(_00334_ ) );
INV_X1 _14008_ ( .A(_06165_ ), .ZN(_06214_ ) );
BUF_X4 _14009_ ( .A(_06214_ ), .Z(_06215_ ) );
AOI21_X1 _14010_ ( .A(_06204_ ), .B1(_06215_ ), .B2(_02129_ ), .ZN(_00335_ ) );
NAND2_X1 _14011_ ( .A1(_06212_ ), .A2(_06213_ ), .ZN(_06216_ ) );
AOI21_X1 _14012_ ( .A(_06204_ ), .B1(_06175_ ), .B2(_06216_ ), .ZN(_00336_ ) );
NOR2_X1 _14013_ ( .A1(_06169_ ), .A2(_03248_ ), .ZN(_06217_ ) );
BUF_X2 _14014_ ( .A(_02186_ ), .Z(_06218_ ) );
NOR3_X1 _14015_ ( .A1(_06218_ ), .A2(\mylsu.state [3] ), .A3(\mylsu.state [1] ), .ZN(_06219_ ) );
OAI211_X1 _14016_ ( .A(_06217_ ), .B(_06219_ ), .C1(_02136_ ), .C2(_02139_ ), .ZN(_06220_ ) );
INV_X1 _14017_ ( .A(_02128_ ), .ZN(_06221_ ) );
OR2_X1 _14018_ ( .A1(_02123_ ), .A2(_06221_ ), .ZN(_06222_ ) );
AND3_X1 _14019_ ( .A1(_06205_ ), .A2(_02255_ ), .A3(_06210_ ), .ZN(_06223_ ) );
NOR2_X1 _14020_ ( .A1(_06223_ ), .A2(_02133_ ), .ZN(_06224_ ) );
AOI21_X1 _14021_ ( .A(_06220_ ), .B1(_06222_ ), .B2(_06224_ ), .ZN(_00337_ ) );
INV_X1 _14022_ ( .A(_00319_ ), .ZN(_06225_ ) );
OAI211_X1 _14023_ ( .A(_02278_ ), .B(_06219_ ), .C1(_04715_ ), .C2(_02328_ ), .ZN(_06226_ ) );
OAI21_X1 _14024_ ( .A(_06225_ ), .B1(_02133_ ), .B2(_06226_ ), .ZN(_00338_ ) );
INV_X1 _14025_ ( .A(\mysc.state [2] ), .ZN(_06227_ ) );
NOR2_X1 _14026_ ( .A1(_06227_ ), .A2(fanout_net_6 ), .ZN(_00339_ ) );
AND2_X1 _14027_ ( .A1(_02144_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_06228_ ) );
CLKBUF_X2 _14028_ ( .A(_06228_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _14029_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .ZN(_06229_ ) );
BUF_X2 _14030_ ( .A(_06229_ ), .Z(_06230_ ) );
AND3_X1 _14031_ ( .A1(_02144_ ), .A2(_06230_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00278_ ) );
AND3_X1 _14032_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06078_ ), .A3(fanout_net_12 ), .ZN(_00279_ ) );
AND3_X1 _14033_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_16 ), .A3(_06087_ ), .ZN(_00280_ ) );
CLKBUF_X2 _14034_ ( .A(_02104_ ), .Z(_06231_ ) );
CLKBUF_X2 _14035_ ( .A(_06231_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _14036_ ( .A(_02151_ ), .Z(_06232_ ) );
NOR3_X1 _14037_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(_06218_ ), .ZN(_06233_ ) );
INV_X1 _14038_ ( .A(_02150_ ), .ZN(_06234_ ) );
BUF_X4 _14039_ ( .A(_06234_ ), .Z(_06235_ ) );
BUF_X4 _14040_ ( .A(_06235_ ), .Z(_06236_ ) );
BUF_X4 _14041_ ( .A(_06236_ ), .Z(_06237_ ) );
INV_X1 _14042_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06238_ ) );
INV_X1 _14043_ ( .A(_02110_ ), .ZN(_06239_ ) );
AOI211_X1 _14044_ ( .A(_06233_ ), .B(_06237_ ), .C1(_06238_ ), .C2(_06239_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _14045_ ( .A1(_06232_ ), .A2(fanout_net_7 ), .A3(_06218_ ), .ZN(_06240_ ) );
INV_X1 _14046_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06241_ ) );
AOI211_X1 _14047_ ( .A(_06240_ ), .B(_06237_ ), .C1(_06241_ ), .C2(_06239_ ), .ZN(\io_master_araddr [0] ) );
OAI221_X1 _14048_ ( .A(\IF_ID_pc [15] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_06242_ ) );
INV_X1 _14049_ ( .A(_02148_ ), .ZN(_06243_ ) );
OR3_X1 _14050_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(_02186_ ), .ZN(_06244_ ) );
BUF_X4 _14051_ ( .A(_02110_ ), .Z(_06245_ ) );
OAI211_X1 _14052_ ( .A(_06243_ ), .B(_06244_ ), .C1(\mylsu.araddr_tmp [15] ), .C2(_06245_ ), .ZN(_06246_ ) );
OAI21_X1 _14053_ ( .A(_06242_ ), .B1(\io_master_arburst [0] ), .B2(_06246_ ), .ZN(\io_master_araddr [15] ) );
OR3_X1 _14054_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(_06218_ ), .ZN(_06247_ ) );
OAI21_X1 _14055_ ( .A(_06247_ ), .B1(_06245_ ), .B2(\mylsu.araddr_tmp [14] ), .ZN(_06248_ ) );
BUF_X4 _14056_ ( .A(_02156_ ), .Z(_06249_ ) );
BUF_X2 _14057_ ( .A(_06249_ ), .Z(_06250_ ) );
OAI22_X1 _14058_ ( .A1(_06237_ ), .A2(_06248_ ), .B1(_02016_ ), .B2(_06250_ ), .ZN(\io_master_araddr [14] ) );
MUX2_X1 _14059_ ( .A(\mylsu.araddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_02110_ ), .Z(_06251_ ) );
AND2_X1 _14060_ ( .A1(_06251_ ), .A2(_06243_ ), .ZN(_06252_ ) );
MUX2_X1 _14061_ ( .A(_06252_ ), .B(\IF_ID_pc [5] ), .S(_06231_ ), .Z(\io_master_araddr [5] ) );
OAI221_X1 _14062_ ( .A(fanout_net_16 ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_06253_ ) );
OR3_X1 _14063_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(_02186_ ), .ZN(_06254_ ) );
OAI211_X1 _14064_ ( .A(_06243_ ), .B(_06254_ ), .C1(\mylsu.araddr_tmp [4] ), .C2(_06245_ ), .ZN(_06255_ ) );
OAI21_X1 _14065_ ( .A(_06253_ ), .B1(\io_master_arburst [0] ), .B2(_06255_ ), .ZN(\io_master_araddr [4] ) );
OR3_X1 _14066_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(_06218_ ), .ZN(_06256_ ) );
OAI21_X1 _14067_ ( .A(_06256_ ), .B1(_06245_ ), .B2(\mylsu.araddr_tmp [3] ), .ZN(_06257_ ) );
OAI22_X1 _14068_ ( .A1(_06237_ ), .A2(_06257_ ), .B1(_06087_ ), .B2(_06250_ ), .ZN(\io_master_araddr [3] ) );
OAI221_X1 _14069_ ( .A(\IF_ID_pc [13] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_06258_ ) );
OR3_X1 _14070_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(_02186_ ), .ZN(_06259_ ) );
OAI211_X1 _14071_ ( .A(_06243_ ), .B(_06259_ ), .C1(\mylsu.araddr_tmp [13] ), .C2(_06245_ ), .ZN(_06260_ ) );
OAI21_X1 _14072_ ( .A(_06258_ ), .B1(\io_master_arburst [0] ), .B2(_06260_ ), .ZN(\io_master_araddr [13] ) );
INV_X1 _14073_ ( .A(_02168_ ), .ZN(\io_master_araddr [22] ) );
AND2_X1 _14074_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _14075_ ( .A1(\EX_LS_dest_csreg_mem [12] ), .A2(_02119_ ), .A3(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A4(_02105_ ), .ZN(_06261_ ) );
AOI21_X1 _14076_ ( .A(_06261_ ), .B1(_06239_ ), .B2(\mylsu.araddr_tmp [12] ), .ZN(_06262_ ) );
OAI22_X1 _14077_ ( .A1(_06237_ ), .A2(_06262_ ), .B1(_02023_ ), .B2(_06250_ ), .ZN(\io_master_araddr [12] ) );
NOR3_X1 _14078_ ( .A1(_06232_ ), .A2(_06174_ ), .A3(_06218_ ), .ZN(_06263_ ) );
AOI21_X1 _14079_ ( .A(_06263_ ), .B1(_06239_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_06264_ ) );
OAI22_X1 _14080_ ( .A1(_06237_ ), .A2(_06264_ ), .B1(_05871_ ), .B2(_06250_ ), .ZN(\io_master_araddr [11] ) );
OAI221_X1 _14081_ ( .A(\IF_ID_pc [10] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02097_ ), .C2(_02098_ ), .ZN(_06265_ ) );
OR3_X1 _14082_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(_02186_ ), .ZN(_06266_ ) );
OAI211_X1 _14083_ ( .A(_06243_ ), .B(_06266_ ), .C1(\mylsu.araddr_tmp [10] ), .C2(_06245_ ), .ZN(_06267_ ) );
OAI21_X1 _14084_ ( .A(_06265_ ), .B1(\io_master_arburst [0] ), .B2(_06267_ ), .ZN(\io_master_araddr [10] ) );
NAND4_X1 _14085_ ( .A1(_02119_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_03378_ ), .A4(_06178_ ), .ZN(_06268_ ) );
OAI21_X1 _14086_ ( .A(_06268_ ), .B1(_06245_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06269_ ) );
OAI22_X1 _14087_ ( .A1(_06237_ ), .A2(_06269_ ), .B1(_05879_ ), .B2(_06250_ ), .ZN(\io_master_araddr [9] ) );
NAND4_X1 _14088_ ( .A1(_02119_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_03379_ ), .A4(_06178_ ), .ZN(_06270_ ) );
OAI21_X1 _14089_ ( .A(_06270_ ), .B1(_06245_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_06271_ ) );
OAI22_X1 _14090_ ( .A1(_06237_ ), .A2(_06271_ ), .B1(_05826_ ), .B2(_06250_ ), .ZN(\io_master_araddr [8] ) );
OR3_X1 _14091_ ( .A1(_06232_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(_06218_ ), .ZN(_06272_ ) );
OAI21_X1 _14092_ ( .A(_06272_ ), .B1(_06245_ ), .B2(\mylsu.araddr_tmp [7] ), .ZN(_06273_ ) );
OAI22_X1 _14093_ ( .A1(_06237_ ), .A2(_06273_ ), .B1(_01962_ ), .B2(_06250_ ), .ZN(\io_master_araddr [7] ) );
NAND4_X1 _14094_ ( .A1(_02119_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A3(_06196_ ), .A4(_06178_ ), .ZN(_06274_ ) );
OAI21_X1 _14095_ ( .A(_06274_ ), .B1(_06245_ ), .B2(\mylsu.araddr_tmp [6] ), .ZN(_06275_ ) );
OAI22_X1 _14096_ ( .A1(_06237_ ), .A2(_06275_ ), .B1(_02033_ ), .B2(_06250_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _14097_ ( .A1(_02151_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(_02186_ ), .ZN(_06276_ ) );
OAI211_X1 _14098_ ( .A(_06243_ ), .B(_06276_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_02110_ ), .ZN(_06277_ ) );
NOR2_X1 _14099_ ( .A1(_02101_ ), .A2(_06277_ ), .ZN(_06278_ ) );
BUF_X4 _14100_ ( .A(_06278_ ), .Z(_06279_ ) );
BUF_X4 _14101_ ( .A(_06279_ ), .Z(_06280_ ) );
BUF_X2 _14102_ ( .A(_06280_ ), .Z(\io_master_araddr [2] ) );
BUF_X2 _14103_ ( .A(_05391_ ), .Z(_06281_ ) );
BUF_X2 _14104_ ( .A(_06281_ ), .Z(\io_master_arid [1] ) );
AND3_X1 _14105_ ( .A1(_06250_ ), .A2(\EX_LS_typ [3] ), .A3(_06243_ ), .ZN(\io_master_arsize [2] ) );
BUF_X4 _14106_ ( .A(_06249_ ), .Z(_06282_ ) );
AND3_X1 _14107_ ( .A1(_06282_ ), .A2(\EX_LS_typ [1] ), .A3(_06243_ ), .ZN(\io_master_arsize [0] ) );
OAI22_X1 _14108_ ( .A1(_02099_ ), .A2(_02100_ ), .B1(_02115_ ), .B2(_02148_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _14109_ ( .A(_02209_ ), .B(_02210_ ), .C1(_02179_ ), .C2(_02205_ ), .ZN(io_master_arvalid ) );
AND2_X1 _14110_ ( .A1(_02132_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_06283_ ) );
BUF_X4 _14111_ ( .A(_06283_ ), .Z(_06284_ ) );
BUF_X4 _14112_ ( .A(_06284_ ), .Z(_06285_ ) );
MUX2_X1 _14113_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06285_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _14114_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06285_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _14115_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06285_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _14116_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06285_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _14117_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06285_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _14118_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06285_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _14119_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06285_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _14120_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06285_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _14121_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06285_ ), .Z(\io_master_awaddr [15] ) );
BUF_X4 _14122_ ( .A(_06284_ ), .Z(_06286_ ) );
MUX2_X1 _14123_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06286_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _14124_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06286_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _14125_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06286_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _14126_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06286_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _14127_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06286_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _14128_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06286_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _14129_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06286_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _14130_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06286_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _14131_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06286_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _14132_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06286_ ), .Z(\io_master_awaddr [6] ) );
BUF_X4 _14133_ ( .A(_06284_ ), .Z(_06287_ ) );
MUX2_X1 _14134_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06287_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _14135_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06287_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _14136_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06287_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _14137_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06287_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _14138_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06287_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _14139_ ( .A(\mylsu.awaddr_tmp [1] ), .B(\EX_LS_dest_csreg_mem [1] ), .S(_06287_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _14140_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_7 ), .S(_06287_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _14141_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06287_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _14142_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06287_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _14143_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06287_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _14144_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06284_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _14145_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06284_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _14146_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06284_ ), .Z(\io_master_awaddr [22] ) );
AND3_X1 _14147_ ( .A1(_02135_ ), .A2(\EX_LS_typ [1] ), .A3(_02112_ ), .ZN(\io_master_awsize [0] ) );
NAND2_X1 _14148_ ( .A1(_02135_ ), .A2(_02112_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _14149_ ( .A1(_02129_ ), .A2(_02141_ ), .A3(_06285_ ), .ZN(_06288_ ) );
INV_X1 _14150_ ( .A(\mylsu.state [4] ), .ZN(_06289_ ) );
NAND2_X1 _14151_ ( .A1(_06288_ ), .A2(_06289_ ), .ZN(io_master_awvalid ) );
INV_X1 _14152_ ( .A(\mylsu.state [2] ), .ZN(_06290_ ) );
INV_X1 _14153_ ( .A(\mylsu.state [1] ), .ZN(_06291_ ) );
NAND4_X1 _14154_ ( .A1(_06288_ ), .A2(_06290_ ), .A3(_06289_ ), .A4(_06291_ ), .ZN(io_master_bready ) );
NOR3_X1 _14155_ ( .A1(_01910_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_06292_ ) );
NAND3_X1 _14156_ ( .A1(_02179_ ), .A2(_05391_ ), .A3(_02205_ ), .ZN(_06293_ ) );
NOR2_X1 _14157_ ( .A1(_06149_ ), .A2(\io_master_rid [0] ), .ZN(_06294_ ) );
NAND4_X1 _14158_ ( .A1(_06294_ ), .A2(io_master_rlast ), .A3(_06147_ ), .A4(_06148_ ), .ZN(_06295_ ) );
OAI21_X1 _14159_ ( .A(_06293_ ), .B1(_06236_ ), .B2(_06295_ ), .ZN(_06296_ ) );
AOI21_X1 _14160_ ( .A(_06162_ ), .B1(_06146_ ), .B2(_06296_ ), .ZN(_06297_ ) );
NOR2_X1 _14161_ ( .A1(\io_master_bid [3] ), .A2(\io_master_bid [2] ), .ZN(_06298_ ) );
AND3_X1 _14162_ ( .A1(_06298_ ), .A2(\io_master_bid [1] ), .A3(\io_master_bid [0] ), .ZN(_06299_ ) );
NOR2_X1 _14163_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_06300_ ) );
AND2_X1 _14164_ ( .A1(_06300_ ), .A2(io_master_bvalid ), .ZN(_06301_ ) );
AND2_X1 _14165_ ( .A1(_06299_ ), .A2(_06301_ ), .ZN(_06302_ ) );
INV_X1 _14166_ ( .A(_06302_ ), .ZN(_06303_ ) );
AOI211_X1 _14167_ ( .A(_06292_ ), .B(_06297_ ), .C1(\mylsu.state [1] ), .C2(_06303_ ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _14168_ ( .A(_02143_ ), .B(_02146_ ), .C1(_02179_ ), .C2(_02205_ ), .ZN(io_master_rready ) );
MUX2_X1 _14169_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_7 ), .Z(_06304_ ) );
INV_X1 _14170_ ( .A(\EX_LS_dest_csreg_mem [1] ), .ZN(_06305_ ) );
CLKBUF_X2 _14171_ ( .A(_06305_ ), .Z(_06306_ ) );
AND2_X1 _14172_ ( .A1(_06304_ ), .A2(_06306_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _14173_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_7 ), .Z(_06307_ ) );
AND2_X1 _14174_ ( .A1(_06307_ ), .A2(_06306_ ), .ZN(\io_master_wdata [14] ) );
INV_X1 _14175_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_06308_ ) );
NOR3_X1 _14176_ ( .A1(_06308_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _14177_ ( .A1(_05133_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [4] ) );
NOR3_X1 _14178_ ( .A1(_05149_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [3] ) );
NOR3_X1 _14179_ ( .A1(_05179_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14180_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06309_ ) );
NOR3_X1 _14181_ ( .A1(_06309_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14182_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06310_ ) );
NOR3_X1 _14183_ ( .A1(_06310_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14184_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_7 ), .Z(_06311_ ) );
AND2_X1 _14185_ ( .A1(_06311_ ), .A2(_06306_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14186_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_7 ), .Z(_06312_ ) );
AND2_X1 _14187_ ( .A1(_06312_ ), .A2(_06306_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14188_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_7 ), .Z(_06313_ ) );
AND2_X1 _14189_ ( .A1(_06313_ ), .A2(_06306_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14190_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_7 ), .Z(_06314_ ) );
AND2_X1 _14191_ ( .A1(_06314_ ), .A2(_06306_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14192_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_7 ), .Z(_06315_ ) );
AND2_X1 _14193_ ( .A1(_06315_ ), .A2(_06306_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14194_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_7 ), .Z(_06316_ ) );
AND2_X1 _14195_ ( .A1(_06316_ ), .A2(_06306_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14196_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06317_ ) );
NOR3_X1 _14197_ ( .A1(_06317_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [7] ) );
INV_X1 _14198_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_06318_ ) );
NOR3_X1 _14199_ ( .A1(_06318_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14200_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_7 ), .Z(_06319_ ) );
MUX2_X1 _14201_ ( .A(_06319_ ), .B(_06304_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14202_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_7 ), .Z(_06320_ ) );
MUX2_X1 _14203_ ( .A(_06320_ ), .B(_06307_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [30] ) );
NOR2_X1 _14204_ ( .A1(_06305_ ), .A2(fanout_net_7 ), .ZN(_06321_ ) );
INV_X1 _14205_ ( .A(_06321_ ), .ZN(_06322_ ) );
OAI21_X1 _14206_ ( .A(_06305_ ), .B1(_06199_ ), .B2(\EX_LS_result_csreg_mem [13] ), .ZN(_06323_ ) );
NOR2_X1 _14207_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [21] ), .ZN(_06324_ ) );
OAI22_X1 _14208_ ( .A1(_06322_ ), .A2(_06308_ ), .B1(_06323_ ), .B2(_06324_ ), .ZN(\io_master_wdata [21] ) );
INV_X1 _14209_ ( .A(\EX_LS_result_csreg_mem [20] ), .ZN(_06325_ ) );
INV_X1 _14210_ ( .A(\EX_LS_result_csreg_mem [12] ), .ZN(_06326_ ) );
MUX2_X1 _14211_ ( .A(_06325_ ), .B(_06326_ ), .S(fanout_net_7 ), .Z(_06327_ ) );
OAI22_X1 _14212_ ( .A1(_06327_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06322_ ), .B2(_05133_ ), .ZN(\io_master_wdata [20] ) );
OAI21_X1 _14213_ ( .A(_06305_ ), .B1(_06199_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_06328_ ) );
NOR2_X1 _14214_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_06329_ ) );
OAI22_X1 _14215_ ( .A1(_06322_ ), .A2(_05149_ ), .B1(_06328_ ), .B2(_06329_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _14216_ ( .A(_06305_ ), .B1(_06199_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_06330_ ) );
NOR2_X1 _14217_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_06331_ ) );
OAI22_X1 _14218_ ( .A1(_06322_ ), .A2(_05179_ ), .B1(_06330_ ), .B2(_06331_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _14219_ ( .A(_06305_ ), .B1(_06199_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_06332_ ) );
NOR2_X1 _14220_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_06333_ ) );
OAI22_X1 _14221_ ( .A1(_06322_ ), .A2(_06309_ ), .B1(_06332_ ), .B2(_06333_ ), .ZN(\io_master_wdata [17] ) );
OAI21_X1 _14222_ ( .A(_06305_ ), .B1(_06199_ ), .B2(\EX_LS_result_csreg_mem [8] ), .ZN(_06334_ ) );
NOR2_X1 _14223_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [16] ), .ZN(_06335_ ) );
OAI22_X1 _14224_ ( .A1(_06322_ ), .A2(_06310_ ), .B1(_06334_ ), .B2(_06335_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14225_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06336_ ) );
MUX2_X1 _14226_ ( .A(_06336_ ), .B(_06311_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14227_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06337_ ) );
MUX2_X1 _14228_ ( .A(_06337_ ), .B(_06312_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14229_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06338_ ) );
MUX2_X1 _14230_ ( .A(_06338_ ), .B(_06313_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14231_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06339_ ) );
MUX2_X1 _14232_ ( .A(_06339_ ), .B(_06314_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14233_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06340_ ) );
MUX2_X1 _14234_ ( .A(_06340_ ), .B(_06315_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14235_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06341_ ) );
MUX2_X1 _14236_ ( .A(_06341_ ), .B(_06316_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [24] ) );
INV_X1 _14237_ ( .A(\EX_LS_result_csreg_mem [15] ), .ZN(_06342_ ) );
MUX2_X1 _14238_ ( .A(_05314_ ), .B(_06342_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06343_ ) );
OAI22_X1 _14239_ ( .A1(_06343_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_06322_ ), .B2(_06317_ ), .ZN(\io_master_wdata [23] ) );
OAI21_X1 _14240_ ( .A(_06305_ ), .B1(_06199_ ), .B2(\EX_LS_result_csreg_mem [14] ), .ZN(_06344_ ) );
NOR2_X1 _14241_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [22] ), .ZN(_06345_ ) );
OAI22_X1 _14242_ ( .A1(_06322_ ), .A2(_06318_ ), .B1(_06344_ ), .B2(_06345_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14243_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06346_ ) );
AND2_X1 _14244_ ( .A1(_06346_ ), .A2(_06306_ ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _14245_ ( .A1(_06199_ ), .A2(_06306_ ), .A3(\EX_LS_typ [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14246_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06347_ ) );
MUX2_X1 _14247_ ( .A(_06347_ ), .B(_06346_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14248_ ( .A1(_06305_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_06348_ ) );
NAND3_X1 _14249_ ( .A1(_06199_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_typ [0] ), .ZN(_06349_ ) );
OAI211_X1 _14250_ ( .A(_06348_ ), .B(_06349_ ), .C1(_02137_ ), .C2(_02115_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _14251_ ( .A1(_06288_ ), .A2(_06290_ ), .ZN(io_master_wvalid ) );
AND2_X1 _14252_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06350_ ) );
NOR2_X1 _14253_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06351_ ) );
AND2_X1 _14254_ ( .A1(_06350_ ), .A2(_06351_ ), .ZN(_06352_ ) );
NOR4_X1 _14255_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .A3(\LS_WB_waddr_csreg [5] ), .A4(\LS_WB_waddr_csreg [4] ), .ZN(_06353_ ) );
NAND2_X1 _14256_ ( .A1(_06352_ ), .A2(_06353_ ), .ZN(_06354_ ) );
INV_X1 _14257_ ( .A(\LS_WB_wen_csreg [7] ), .ZN(_06355_ ) );
NOR2_X1 _14258_ ( .A1(_06355_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_06356_ ) );
INV_X1 _14259_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_06357_ ) );
INV_X1 _14260_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_06358_ ) );
INV_X1 _14261_ ( .A(\LS_WB_waddr_csreg [2] ), .ZN(_06359_ ) );
NAND4_X1 _14262_ ( .A1(_06356_ ), .A2(_06357_ ), .A3(_06358_ ), .A4(_06359_ ), .ZN(_06360_ ) );
NOR2_X1 _14263_ ( .A1(_06354_ ), .A2(_06360_ ), .ZN(\mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _14264_ ( .A1(_06356_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(_06358_ ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_06361_ ) );
NOR2_X1 _14265_ ( .A1(_06354_ ), .A2(_06361_ ), .ZN(\mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _14266_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06362_ ) );
NAND2_X1 _14267_ ( .A1(_06362_ ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06363_ ) );
NOR2_X1 _14268_ ( .A1(_06363_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06364_ ) );
AND4_X1 _14269_ ( .A1(\LS_WB_waddr_csreg [0] ), .A2(_06364_ ), .A3(_06358_ ), .A4(_06356_ ), .ZN(_06365_ ) );
AND3_X1 _14270_ ( .A1(_06365_ ), .A2(_06359_ ), .A3(_06352_ ), .ZN(\mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14271_ ( .A(_06364_ ), .ZN(_06366_ ) );
NOR4_X1 _14272_ ( .A1(_06366_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(_06358_ ), .A4(\LS_WB_waddr_csreg [3] ), .ZN(_06367_ ) );
NAND3_X1 _14273_ ( .A1(_06367_ ), .A2(_06359_ ), .A3(_06352_ ), .ZN(_06368_ ) );
AOI21_X1 _14274_ ( .A(_06355_ ), .B1(_06368_ ), .B2(_02244_ ), .ZN(\mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ) );
NOR4_X1 _14275_ ( .A1(_02260_ ), .A2(fanout_net_6 ), .A3(excp_written ), .A4(EXU_valid_LSU ), .ZN(\mycsreg.excp_written_$_NOR__A_Y_$_ANDNOT__A_Y ) );
INV_X1 _14276_ ( .A(_02142_ ), .ZN(_06369_ ) );
OR2_X2 _14277_ ( .A1(_06369_ ), .A2(_02256_ ), .ZN(_06370_ ) );
BUF_X4 _14278_ ( .A(_06370_ ), .Z(_06371_ ) );
MUX2_X1 _14279_ ( .A(\ID_EX_pc [21] ), .B(\EX_LS_pc [21] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14280_ ( .A(\ID_EX_pc [20] ), .B(\EX_LS_pc [20] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14281_ ( .A(\ID_EX_pc [19] ), .B(\EX_LS_pc [19] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14282_ ( .A(\ID_EX_pc [18] ), .B(\EX_LS_pc [18] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14283_ ( .A(\ID_EX_pc [17] ), .B(\EX_LS_pc [17] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14284_ ( .A(\ID_EX_pc [16] ), .B(\EX_LS_pc [16] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14285_ ( .A(\ID_EX_pc [15] ), .B(\EX_LS_pc [15] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14286_ ( .A(\ID_EX_pc [14] ), .B(\EX_LS_pc [14] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14287_ ( .A(\ID_EX_pc [13] ), .B(\EX_LS_pc [13] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14288_ ( .A(\ID_EX_pc [12] ), .B(\EX_LS_pc [12] ), .S(_06371_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14289_ ( .A(_06370_ ), .Z(_06372_ ) );
MUX2_X1 _14290_ ( .A(\ID_EX_pc [30] ), .B(\EX_LS_pc [30] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14291_ ( .A(\ID_EX_pc [11] ), .B(\EX_LS_pc [11] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14292_ ( .A(\ID_EX_pc [10] ), .B(\EX_LS_pc [10] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14293_ ( .A(\ID_EX_pc [9] ), .B(\EX_LS_pc [9] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14294_ ( .A(\ID_EX_pc [8] ), .B(\EX_LS_pc [8] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14295_ ( .A(\ID_EX_pc [7] ), .B(\EX_LS_pc [7] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14296_ ( .A(\ID_EX_pc [6] ), .B(\EX_LS_pc [6] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14297_ ( .A(\ID_EX_pc [5] ), .B(\EX_LS_pc [5] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14298_ ( .A(\ID_EX_pc [4] ), .B(\EX_LS_pc [4] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14299_ ( .A(\ID_EX_pc [3] ), .B(\EX_LS_pc [3] ), .S(_06372_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14300_ ( .A(_06370_ ), .Z(_06373_ ) );
MUX2_X1 _14301_ ( .A(\ID_EX_pc [2] ), .B(\EX_LS_pc [2] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14302_ ( .A(\ID_EX_pc [29] ), .B(\EX_LS_pc [29] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14303_ ( .A(\ID_EX_pc [1] ), .B(\EX_LS_pc [1] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14304_ ( .A(\ID_EX_pc [0] ), .B(\EX_LS_pc [0] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14305_ ( .A(\ID_EX_pc [28] ), .B(\EX_LS_pc [28] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14306_ ( .A(\ID_EX_pc [27] ), .B(\EX_LS_pc [27] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14307_ ( .A(\ID_EX_pc [26] ), .B(\EX_LS_pc [26] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14308_ ( .A(\ID_EX_pc [25] ), .B(\EX_LS_pc [25] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14309_ ( .A(\ID_EX_pc [24] ), .B(\EX_LS_pc [24] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14310_ ( .A(\ID_EX_pc [23] ), .B(\EX_LS_pc [23] ), .S(_06373_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14311_ ( .A(\ID_EX_pc [22] ), .B(\EX_LS_pc [22] ), .S(_06370_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14312_ ( .A(\ID_EX_pc [31] ), .B(\EX_LS_pc [31] ), .S(_06370_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
NOR4_X1 _14313_ ( .A1(_06369_ ), .A2(exception_quest_IDU ), .A3(_02256_ ), .A4(_02259_ ), .ZN(_06374_ ) );
XNOR2_X1 _14314_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06375_ ) );
XNOR2_X1 _14315_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06376_ ) );
XNOR2_X1 _14316_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06377_ ) );
XNOR2_X1 _14317_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06378_ ) );
AND4_X1 _14318_ ( .A1(_06375_ ), .A2(_06376_ ), .A3(_06377_ ), .A4(_06378_ ), .ZN(_06379_ ) );
XNOR2_X1 _14319_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06380_ ) );
XNOR2_X1 _14320_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06381_ ) );
XNOR2_X1 _14321_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06382_ ) );
XNOR2_X1 _14322_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06383_ ) );
AND4_X1 _14323_ ( .A1(_06380_ ), .A2(_06381_ ), .A3(_06382_ ), .A4(_06383_ ), .ZN(_06384_ ) );
XNOR2_X1 _14324_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_06385_ ) );
XNOR2_X1 _14325_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_06386_ ) );
XNOR2_X1 _14326_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_06387_ ) );
XNOR2_X1 _14327_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_06388_ ) );
AND4_X1 _14328_ ( .A1(_06385_ ), .A2(_06386_ ), .A3(_06387_ ), .A4(_06388_ ), .ZN(_06389_ ) );
XNOR2_X1 _14329_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06390_ ) );
XNOR2_X1 _14330_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06391_ ) );
XNOR2_X1 _14331_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06392_ ) );
XNOR2_X1 _14332_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06393_ ) );
AND4_X1 _14333_ ( .A1(_06390_ ), .A2(_06391_ ), .A3(_06392_ ), .A4(_06393_ ), .ZN(_06394_ ) );
AND4_X1 _14334_ ( .A1(_06379_ ), .A2(_06384_ ), .A3(_06389_ ), .A4(_06394_ ), .ZN(_06395_ ) );
XNOR2_X1 _14335_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06396_ ) );
XNOR2_X1 _14336_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06397_ ) );
XNOR2_X1 _14337_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06398_ ) );
XNOR2_X1 _14338_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06399_ ) );
NAND4_X1 _14339_ ( .A1(_06396_ ), .A2(_06397_ ), .A3(_06398_ ), .A4(_06399_ ), .ZN(_06400_ ) );
XNOR2_X1 _14340_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06401_ ) );
XNOR2_X1 _14341_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06402_ ) );
XNOR2_X1 _14342_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06403_ ) );
XNOR2_X1 _14343_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06404_ ) );
NAND4_X1 _14344_ ( .A1(_06401_ ), .A2(_06402_ ), .A3(_06403_ ), .A4(_06404_ ), .ZN(_06405_ ) );
NOR2_X1 _14345_ ( .A1(_06400_ ), .A2(_06405_ ), .ZN(_06406_ ) );
XNOR2_X1 _14346_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06407_ ) );
XNOR2_X1 _14347_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06408_ ) );
XNOR2_X1 _14348_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06409_ ) );
XNOR2_X1 _14349_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06410_ ) );
NAND4_X1 _14350_ ( .A1(_06407_ ), .A2(_06408_ ), .A3(_06409_ ), .A4(_06410_ ), .ZN(_06411_ ) );
XNOR2_X1 _14351_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06412_ ) );
XNOR2_X1 _14352_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06413_ ) );
NAND2_X1 _14353_ ( .A1(_06412_ ), .A2(_06413_ ), .ZN(_06414_ ) );
XOR2_X1 _14354_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .Z(_06415_ ) );
XOR2_X1 _14355_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .Z(_06416_ ) );
NOR4_X1 _14356_ ( .A1(_06411_ ), .A2(_06414_ ), .A3(_06415_ ), .A4(_06416_ ), .ZN(_06417_ ) );
NAND4_X1 _14357_ ( .A1(_06395_ ), .A2(_06406_ ), .A3(excp_written ), .A4(_06417_ ), .ZN(_06418_ ) );
AOI21_X1 _14358_ ( .A(_06374_ ), .B1(_02259_ ), .B2(_06418_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _14359_ ( .A1(_05202_ ), .A2(_03192_ ), .ZN(_06419_ ) );
AND2_X1 _14360_ ( .A1(_03189_ ), .A2(_02262_ ), .ZN(_06420_ ) );
BUF_X4 _14361_ ( .A(_06420_ ), .Z(_06421_ ) );
INV_X2 _14362_ ( .A(_06421_ ), .ZN(_06422_ ) );
BUF_X4 _14363_ ( .A(_06422_ ), .Z(_06423_ ) );
BUF_X4 _14364_ ( .A(_06423_ ), .Z(_06424_ ) );
OAI21_X1 _14365_ ( .A(_06419_ ), .B1(_03414_ ), .B2(_06424_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _14366_ ( .A(_04071_ ), .B(\ID_EX_imm [0] ), .ZN(_06425_ ) );
BUF_X4 _14367_ ( .A(_06421_ ), .Z(_06426_ ) );
BUF_X4 _14368_ ( .A(_06426_ ), .Z(_06427_ ) );
AOI22_X1 _14369_ ( .A1(_06425_ ), .A2(_03193_ ), .B1(_03407_ ), .B2(_06427_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND2_X1 _14370_ ( .A1(_05681_ ), .A2(\ID_EX_typ [7] ), .ZN(_06428_ ) );
INV_X1 _14371_ ( .A(_06428_ ), .ZN(_06429_ ) );
BUF_X4 _14372_ ( .A(_06429_ ), .Z(_06430_ ) );
AND2_X1 _14373_ ( .A1(_05022_ ), .A2(_06430_ ), .ZN(_06431_ ) );
BUF_X4 _14374_ ( .A(_06422_ ), .Z(_06432_ ) );
MUX2_X1 _14375_ ( .A(\ID_EX_csr [10] ), .B(_06431_ ), .S(_06432_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
AOI22_X1 _14376_ ( .A1(_05043_ ), .A2(_03193_ ), .B1(_03373_ ), .B2(_06427_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
AOI22_X1 _14377_ ( .A1(_05062_ ), .A2(_03193_ ), .B1(_03374_ ), .B2(_06427_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND4_X1 _14378_ ( .A1(_02262_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_csr [7] ), .ZN(_06433_ ) );
OAI21_X1 _14379_ ( .A(_06433_ ), .B1(_05085_ ), .B2(_03189_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
BUF_X4 _14380_ ( .A(_06421_ ), .Z(_06434_ ) );
BUF_X4 _14381_ ( .A(_06434_ ), .Z(_06435_ ) );
AOI22_X1 _14382_ ( .A1(_05104_ ), .A2(_03193_ ), .B1(_03422_ ), .B2(_06435_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
OAI22_X1 _14383_ ( .A1(_05125_ ), .A2(_03189_ ), .B1(_03431_ ), .B2(_06424_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND4_X1 _14384_ ( .A1(_02262_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_csr [4] ), .ZN(_06436_ ) );
OAI21_X1 _14385_ ( .A(_06436_ ), .B1(_05145_ ), .B2(_03189_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
OAI22_X1 _14386_ ( .A1(_05165_ ), .A2(_03189_ ), .B1(_03409_ ), .B2(_06424_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND4_X1 _14387_ ( .A1(_02262_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_csr [2] ), .ZN(_06437_ ) );
OAI21_X1 _14388_ ( .A(_06437_ ), .B1(_05183_ ), .B2(_03189_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
AND2_X1 _14389_ ( .A1(_04984_ ), .A2(_06430_ ), .ZN(_06438_ ) );
MUX2_X1 _14390_ ( .A(\ID_EX_csr [11] ), .B(_06438_ ), .S(_06432_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
NOR2_X1 _14391_ ( .A1(_04292_ ), .A2(\ID_EX_typ [2] ), .ZN(_06439_ ) );
INV_X1 _14392_ ( .A(_06439_ ), .ZN(_06440_ ) );
BUF_X4 _14393_ ( .A(_06440_ ), .Z(_06441_ ) );
AOI21_X1 _14394_ ( .A(_06441_ ), .B1(_05354_ ), .B2(_05355_ ), .ZN(_06442_ ) );
AOI22_X1 _14395_ ( .A1(_05356_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02442_ ), .ZN(_06443_ ) );
NAND3_X1 _14396_ ( .A1(_02441_ ), .A2(_02461_ ), .A3(_04759_ ), .ZN(_06444_ ) );
AOI211_X1 _14397_ ( .A(_06423_ ), .B(_06442_ ), .C1(_06443_ ), .C2(_06444_ ), .ZN(_06445_ ) );
BUF_X4 _14398_ ( .A(_06429_ ), .Z(_06446_ ) );
MUX2_X1 _14399_ ( .A(_05383_ ), .B(_03776_ ), .S(_06446_ ), .Z(_06447_ ) );
AOI21_X1 _14400_ ( .A(_06445_ ), .B1(_06424_ ), .B2(_06447_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
AND4_X1 _14401_ ( .A1(_06325_ ), .A2(_04779_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_06448_ ) );
AND2_X1 _14402_ ( .A1(_04697_ ), .A2(\mepc [20] ), .ZN(_06449_ ) );
AOI211_X1 _14403_ ( .A(_04750_ ), .B(_06449_ ), .C1(_04776_ ), .C2(_04789_ ), .ZN(_06450_ ) );
AND4_X1 _14404_ ( .A1(\mycsreg.CSReg[3][20] ), .A2(_04683_ ), .A3(_05012_ ), .A4(_05013_ ), .ZN(_06451_ ) );
NOR4_X1 _14405_ ( .A1(_05136_ ), .A2(_04784_ ), .A3(_04747_ ), .A4(_06451_ ), .ZN(_06452_ ) );
AOI21_X1 _14406_ ( .A(_06448_ ), .B1(_06450_ ), .B2(_06452_ ), .ZN(_06453_ ) );
AOI21_X1 _14407_ ( .A(fanout_net_9 ), .B1(_02465_ ), .B2(_02484_ ), .ZN(_06454_ ) );
AND2_X1 _14408_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [20] ), .ZN(_06455_ ) );
OAI221_X1 _14409_ ( .A(_06426_ ), .B1(_05402_ ), .B2(_06453_ ), .C1(_06454_ ), .C2(_06455_ ), .ZN(_06456_ ) );
BUF_X4 _14410_ ( .A(_06434_ ), .Z(_06457_ ) );
BUF_X4 _14411_ ( .A(_06439_ ), .Z(_06458_ ) );
BUF_X4 _14412_ ( .A(_06458_ ), .Z(_06459_ ) );
NAND3_X1 _14413_ ( .A1(_06453_ ), .A2(_06457_ ), .A3(_06459_ ), .ZN(_06460_ ) );
BUF_X4 _14414_ ( .A(_06421_ ), .Z(_06461_ ) );
BUF_X4 _14415_ ( .A(_06461_ ), .Z(_06462_ ) );
MUX2_X1 _14416_ ( .A(_05345_ ), .B(_03800_ ), .S(_06430_ ), .Z(_06463_ ) );
OAI211_X1 _14417_ ( .A(_06456_ ), .B(_06460_ ), .C1(_06462_ ), .C2(_06463_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
AOI21_X1 _14418_ ( .A(fanout_net_9 ), .B1(_02513_ ), .B2(_02532_ ), .ZN(_06464_ ) );
AND2_X1 _14419_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [19] ), .ZN(_06465_ ) );
OAI221_X1 _14420_ ( .A(_06426_ ), .B1(_06464_ ), .B2(_06465_ ), .C1(_04795_ ), .C2(_05402_ ), .ZN(_06466_ ) );
AND3_X1 _14421_ ( .A1(_04788_ ), .A2(_04793_ ), .A3(_06421_ ), .ZN(_06467_ ) );
NAND2_X1 _14422_ ( .A1(_06467_ ), .A2(_06459_ ), .ZN(_06468_ ) );
MUX2_X1 _14423_ ( .A(_03332_ ), .B(_03826_ ), .S(_06430_ ), .Z(_06469_ ) );
OAI211_X1 _14424_ ( .A(_06466_ ), .B(_06468_ ), .C1(_06462_ ), .C2(_06469_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
NOR2_X1 _14425_ ( .A1(_04758_ ), .A2(\ID_EX_imm [18] ), .ZN(_06470_ ) );
INV_X1 _14426_ ( .A(_04810_ ), .ZN(_06471_ ) );
INV_X1 _14427_ ( .A(_02510_ ), .ZN(_06472_ ) );
AOI221_X4 _14428_ ( .A(_06470_ ), .B1(_06471_ ), .B2(\ID_EX_typ [2] ), .C1(_04758_ ), .C2(_06472_ ), .ZN(_06473_ ) );
AOI211_X1 _14429_ ( .A(_06441_ ), .B(_04808_ ), .C1(_04802_ ), .C2(_04805_ ), .ZN(_06474_ ) );
OAI21_X1 _14430_ ( .A(_06435_ ), .B1(_06473_ ), .B2(_06474_ ), .ZN(_06475_ ) );
MUX2_X1 _14431_ ( .A(_05384_ ), .B(_03848_ ), .S(_06430_ ), .Z(_06476_ ) );
OAI21_X1 _14432_ ( .A(_06475_ ), .B1(_06462_ ), .B2(_06476_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
INV_X1 _14433_ ( .A(\EX_LS_result_csreg_mem [17] ), .ZN(_06477_ ) );
AND4_X1 _14434_ ( .A1(_06477_ ), .A2(_04779_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_06478_ ) );
NAND3_X1 _14435_ ( .A1(_04839_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_04700_ ), .ZN(_06479_ ) );
NAND2_X1 _14436_ ( .A1(_04842_ ), .A2(_06479_ ), .ZN(_06480_ ) );
AND4_X1 _14437_ ( .A1(\mycsreg.CSReg[3][17] ), .A2(_04683_ ), .A3(_04684_ ), .A4(_04685_ ), .ZN(_06481_ ) );
NOR4_X1 _14438_ ( .A1(_06480_ ), .A2(_05136_ ), .A3(_04784_ ), .A4(_06481_ ), .ZN(_06482_ ) );
AOI21_X1 _14439_ ( .A(_04840_ ), .B1(_04776_ ), .B2(_04789_ ), .ZN(_06483_ ) );
AOI21_X1 _14440_ ( .A(_06478_ ), .B1(_06482_ ), .B2(_06483_ ), .ZN(_06484_ ) );
AOI21_X1 _14441_ ( .A(fanout_net_9 ), .B1(_02537_ ), .B2(_02556_ ), .ZN(_06485_ ) );
AND2_X1 _14442_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [17] ), .ZN(_06486_ ) );
OAI221_X1 _14443_ ( .A(_06457_ ), .B1(_05402_ ), .B2(_06484_ ), .C1(_06485_ ), .C2(_06486_ ), .ZN(_06487_ ) );
BUF_X4 _14444_ ( .A(_06423_ ), .Z(_06488_ ) );
AOI21_X1 _14445_ ( .A(_06428_ ), .B1(_03875_ ), .B2(_03895_ ), .ZN(_06489_ ) );
CLKBUF_X2 _14446_ ( .A(_05681_ ), .Z(_06490_ ) );
AND3_X1 _14447_ ( .A1(_06490_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_typ [7] ), .ZN(_06491_ ) );
OAI21_X1 _14448_ ( .A(_06488_ ), .B1(_06489_ ), .B2(_06491_ ), .ZN(_06492_ ) );
NAND3_X1 _14449_ ( .A1(_06484_ ), .A2(_06435_ ), .A3(_06459_ ), .ZN(_06493_ ) );
NAND3_X1 _14450_ ( .A1(_06487_ ), .A2(_06492_ ), .A3(_06493_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _14451_ ( .A(_06441_ ), .B1(_04867_ ), .B2(_04868_ ), .ZN(_06494_ ) );
AND2_X1 _14452_ ( .A1(_04867_ ), .A2(_04868_ ), .ZN(_06495_ ) );
AOI22_X1 _14453_ ( .A1(_06495_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02581_ ), .ZN(_06496_ ) );
NAND3_X1 _14454_ ( .A1(_02560_ ), .A2(_04759_ ), .A3(_02579_ ), .ZN(_06497_ ) );
AOI211_X1 _14455_ ( .A(_06423_ ), .B(_06494_ ), .C1(_06496_ ), .C2(_06497_ ), .ZN(_06498_ ) );
MUX2_X1 _14456_ ( .A(_04823_ ), .B(_03871_ ), .S(_06446_ ), .Z(_06499_ ) );
AOI21_X1 _14457_ ( .A(_06498_ ), .B1(_06424_ ), .B2(_06499_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
AOI21_X1 _14458_ ( .A(_06441_ ), .B1(_04894_ ), .B2(_04895_ ), .ZN(_06500_ ) );
NOR2_X1 _14459_ ( .A1(_03251_ ), .A2(\ID_EX_imm [15] ), .ZN(_06501_ ) );
AOI21_X1 _14460_ ( .A(_06501_ ), .B1(_04896_ ), .B2(\ID_EX_typ [2] ), .ZN(_06502_ ) );
NAND3_X1 _14461_ ( .A1(_02584_ ), .A2(_02604_ ), .A3(_04759_ ), .ZN(_06503_ ) );
AOI211_X1 _14462_ ( .A(_06423_ ), .B(_06500_ ), .C1(_06502_ ), .C2(_06503_ ), .ZN(_06504_ ) );
MUX2_X1 _14463_ ( .A(_04884_ ), .B(_04260_ ), .S(_06446_ ), .Z(_06505_ ) );
AOI21_X1 _14464_ ( .A(_06504_ ), .B1(_06424_ ), .B2(_06505_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
NOR2_X1 _14465_ ( .A1(_04758_ ), .A2(\ID_EX_imm [14] ), .ZN(_06506_ ) );
AOI221_X4 _14466_ ( .A(_06506_ ), .B1(_04916_ ), .B2(\ID_EX_typ [2] ), .C1(_04442_ ), .C2(_04758_ ), .ZN(_06507_ ) );
AOI21_X1 _14467_ ( .A(_06441_ ), .B1(_04914_ ), .B2(_04915_ ), .ZN(_06508_ ) );
OAI21_X1 _14468_ ( .A(_06435_ ), .B1(_06507_ ), .B2(_06508_ ), .ZN(_06509_ ) );
MUX2_X1 _14469_ ( .A(_04904_ ), .B(_04282_ ), .S(_06430_ ), .Z(_06510_ ) );
OAI21_X1 _14470_ ( .A(_06509_ ), .B1(_06462_ ), .B2(_06510_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
AND2_X1 _14471_ ( .A1(_04931_ ), .A2(_04932_ ), .ZN(_06511_ ) );
AOI22_X1 _14472_ ( .A1(_06511_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02867_ ), .ZN(_06512_ ) );
OAI211_X1 _14473_ ( .A(_06512_ ), .B(_06457_ ), .C1(fanout_net_9 ), .C2(_04194_ ), .ZN(_06513_ ) );
AOI21_X1 _14474_ ( .A(_06423_ ), .B1(_04931_ ), .B2(_04932_ ), .ZN(_06514_ ) );
NAND2_X1 _14475_ ( .A1(_06514_ ), .A2(_06459_ ), .ZN(_06515_ ) );
AND3_X1 _14476_ ( .A1(_04195_ ), .A2(_04214_ ), .A3(_06429_ ), .ZN(_06516_ ) );
AND3_X1 _14477_ ( .A1(_06490_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_typ [7] ), .ZN(_06517_ ) );
OAI21_X1 _14478_ ( .A(_06488_ ), .B1(_06516_ ), .B2(_06517_ ), .ZN(_06518_ ) );
NAND3_X1 _14479_ ( .A1(_06513_ ), .A2(_06515_ ), .A3(_06518_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AND3_X1 _14480_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(\EX_LS_result_csreg_mem [12] ), .ZN(_06519_ ) );
AOI21_X1 _14481_ ( .A(_06519_ ), .B1(_04949_ ), .B2(_03396_ ), .ZN(_06520_ ) );
AOI22_X1 _14482_ ( .A1(_06520_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02864_ ), .ZN(_06521_ ) );
OAI211_X1 _14483_ ( .A(_06521_ ), .B(_06461_ ), .C1(fanout_net_9 ), .C2(_02863_ ), .ZN(_06522_ ) );
AND2_X1 _14484_ ( .A1(_04781_ ), .A2(\mepc [12] ), .ZN(_06523_ ) );
AOI211_X1 _14485_ ( .A(_04944_ ), .B(_06523_ ), .C1(_04776_ ), .C2(_04789_ ), .ZN(_06524_ ) );
AND4_X1 _14486_ ( .A1(\mycsreg.CSReg[3][12] ), .A2(_04738_ ), .A3(_05193_ ), .A4(_04741_ ), .ZN(_06525_ ) );
NOR3_X1 _14487_ ( .A1(_05136_ ), .A2(_04784_ ), .A3(_06525_ ), .ZN(_06526_ ) );
INV_X1 _14488_ ( .A(_04943_ ), .ZN(_06527_ ) );
NAND3_X1 _14489_ ( .A1(_06524_ ), .A2(_06526_ ), .A3(_06527_ ), .ZN(_06528_ ) );
NAND4_X1 _14490_ ( .A1(_04789_ ), .A2(_06326_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_06529_ ) );
NAND4_X1 _14491_ ( .A1(_06528_ ), .A2(_06529_ ), .A3(_06426_ ), .A4(_06458_ ), .ZN(_06530_ ) );
MUX2_X1 _14492_ ( .A(_04938_ ), .B(_04237_ ), .S(_06446_ ), .Z(_06531_ ) );
OAI211_X1 _14493_ ( .A(_06522_ ), .B(_06530_ ), .C1(_06531_ ), .C2(_06427_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
NAND3_X1 _14494_ ( .A1(_02356_ ), .A2(_02357_ ), .A3(_04758_ ), .ZN(_06532_ ) );
NAND2_X1 _14495_ ( .A1(_03441_ ), .A2(_03446_ ), .ZN(_06533_ ) );
OAI221_X1 _14496_ ( .A(_06532_ ), .B1(_03251_ ), .B2(\ID_EX_imm [30] ), .C1(_04649_ ), .C2(_06533_ ), .ZN(_06534_ ) );
AOI21_X1 _14497_ ( .A(_03412_ ), .B1(_04776_ ), .B2(_04779_ ), .ZN(_06535_ ) );
NAND2_X1 _14498_ ( .A1(_04697_ ), .A2(\mepc [30] ), .ZN(_06536_ ) );
NAND3_X1 _14499_ ( .A1(_04839_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_04749_ ), .ZN(_06537_ ) );
NAND2_X1 _14500_ ( .A1(_06536_ ), .A2(_06537_ ), .ZN(_06538_ ) );
AND4_X1 _14501_ ( .A1(\mycsreg.CSReg[3][30] ), .A2(_04683_ ), .A3(_05012_ ), .A4(_05013_ ), .ZN(_06539_ ) );
NOR3_X1 _14502_ ( .A1(_06538_ ), .A2(_05136_ ), .A3(_06539_ ), .ZN(_06540_ ) );
NAND2_X1 _14503_ ( .A1(_06535_ ), .A2(_06540_ ), .ZN(_06541_ ) );
AND2_X2 _14504_ ( .A1(_04775_ ), .A2(_04778_ ), .ZN(_06542_ ) );
INV_X1 _14505_ ( .A(_06542_ ), .ZN(_06543_ ) );
OAI211_X1 _14506_ ( .A(_06541_ ), .B(_06458_ ), .C1(_06543_ ), .C2(\EX_LS_result_csreg_mem [30] ), .ZN(_06544_ ) );
AND3_X1 _14507_ ( .A1(_06534_ ), .A2(_06434_ ), .A3(_06544_ ), .ZN(_06545_ ) );
MUX2_X1 _14508_ ( .A(_05361_ ), .B(_03699_ ), .S(_06446_ ), .Z(_06546_ ) );
AOI21_X1 _14509_ ( .A(_06545_ ), .B1(_06424_ ), .B2(_06546_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
AND2_X1 _14510_ ( .A1(_04975_ ), .A2(_04976_ ), .ZN(_06547_ ) );
AOI22_X1 _14511_ ( .A1(_06547_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02937_ ), .ZN(_06548_ ) );
OAI211_X1 _14512_ ( .A(_06548_ ), .B(_06461_ ), .C1(\ID_EX_typ [0] ), .C2(_02936_ ), .ZN(_06549_ ) );
AOI21_X1 _14513_ ( .A(_06422_ ), .B1(_04975_ ), .B2(_04976_ ), .ZN(_06550_ ) );
NAND2_X1 _14514_ ( .A1(_06550_ ), .A2(_06459_ ), .ZN(_06551_ ) );
MUX2_X1 _14515_ ( .A(_04958_ ), .B(_04120_ ), .S(_06429_ ), .Z(_06552_ ) );
OAI211_X1 _14516_ ( .A(_06549_ ), .B(_06551_ ), .C1(_06462_ ), .C2(_06552_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _14517_ ( .A(_06440_ ), .B1(_05017_ ), .B2(_05018_ ), .ZN(_06553_ ) );
AND2_X1 _14518_ ( .A1(_05017_ ), .A2(_05018_ ), .ZN(_06554_ ) );
AOI22_X1 _14519_ ( .A1(_06554_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02913_ ), .ZN(_06555_ ) );
NAND3_X1 _14520_ ( .A1(_02892_ ), .A2(_04759_ ), .A3(_02911_ ), .ZN(_06556_ ) );
AOI211_X1 _14521_ ( .A(_06423_ ), .B(_06553_ ), .C1(_06555_ ), .C2(_06556_ ), .ZN(_06557_ ) );
MUX2_X1 _14522_ ( .A(_05385_ ), .B(_04142_ ), .S(_06446_ ), .Z(_06558_ ) );
AOI21_X1 _14523_ ( .A(_06557_ ), .B1(_06424_ ), .B2(_06558_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
BUF_X4 _14524_ ( .A(_06434_ ), .Z(_06559_ ) );
NOR2_X1 _14525_ ( .A1(_03250_ ), .A2(\ID_EX_imm [9] ), .ZN(_06560_ ) );
AOI221_X4 _14526_ ( .A(_06560_ ), .B1(_05037_ ), .B2(\ID_EX_typ [2] ), .C1(_04366_ ), .C2(_04758_ ), .ZN(_06561_ ) );
AOI21_X1 _14527_ ( .A(_06441_ ), .B1(_05035_ ), .B2(_05036_ ), .ZN(_06562_ ) );
OAI21_X1 _14528_ ( .A(_06559_ ), .B1(_06561_ ), .B2(_06562_ ), .ZN(_06563_ ) );
MUX2_X1 _14529_ ( .A(_05386_ ), .B(_04188_ ), .S(_06430_ ), .Z(_06564_ ) );
OAI21_X1 _14530_ ( .A(_06563_ ), .B1(_06462_ ), .B2(_06564_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
NOR2_X1 _14531_ ( .A1(_03250_ ), .A2(\ID_EX_imm [8] ), .ZN(_06565_ ) );
AOI221_X4 _14532_ ( .A(_06565_ ), .B1(_05059_ ), .B2(\ID_EX_typ [2] ), .C1(_04428_ ), .C2(_04758_ ), .ZN(_06566_ ) );
AOI21_X1 _14533_ ( .A(_06441_ ), .B1(_05057_ ), .B2(_05058_ ), .ZN(_06567_ ) );
OAI21_X1 _14534_ ( .A(_06559_ ), .B1(_06566_ ), .B2(_06567_ ), .ZN(_06568_ ) );
MUX2_X1 _14535_ ( .A(_05387_ ), .B(_04166_ ), .S(_06430_ ), .Z(_06569_ ) );
OAI21_X1 _14536_ ( .A(_06568_ ), .B1(_06462_ ), .B2(_06569_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
NAND4_X1 _14537_ ( .A1(_04789_ ), .A2(_06317_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_06570_ ) );
NAND2_X1 _14538_ ( .A1(_04781_ ), .A2(\mepc [7] ), .ZN(_06571_ ) );
NAND4_X1 _14539_ ( .A1(_04738_ ), .A2(_05193_ ), .A3(\mycsreg.CSReg[3][7] ), .A4(_04741_ ), .ZN(_06572_ ) );
NAND4_X1 _14540_ ( .A1(_06571_ ), .A2(_05071_ ), .A3(_05072_ ), .A4(_06572_ ), .ZN(_06573_ ) );
OAI211_X1 _14541_ ( .A(_06570_ ), .B(_06458_ ), .C1(_06542_ ), .C2(_06573_ ), .ZN(_06574_ ) );
AOI21_X1 _14542_ ( .A(\ID_EX_typ [0] ), .B1(_02684_ ), .B2(_02704_ ), .ZN(_06575_ ) );
AND2_X1 _14543_ ( .A1(\ID_EX_typ [0] ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_06576_ ) );
OAI21_X1 _14544_ ( .A(_06574_ ), .B1(_06575_ ), .B2(_06576_ ), .ZN(_06577_ ) );
OAI211_X1 _14545_ ( .A(_06577_ ), .B(_06435_ ), .C1(_05402_ ), .C2(_05079_ ), .ZN(_06578_ ) );
NAND3_X1 _14546_ ( .A1(_03901_ ), .A2(_03922_ ), .A3(_06446_ ), .ZN(_06579_ ) );
BUF_X4 _14547_ ( .A(_06430_ ), .Z(_06580_ ) );
OAI211_X1 _14548_ ( .A(_06579_ ), .B(_06488_ ), .C1(\ID_EX_pc [7] ), .C2(_06580_ ), .ZN(_06581_ ) );
NAND2_X1 _14549_ ( .A1(_06578_ ), .A2(_06581_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
INV_X1 _14550_ ( .A(_05102_ ), .ZN(_06582_ ) );
AOI22_X1 _14551_ ( .A1(_06582_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02730_ ), .ZN(_06583_ ) );
OAI211_X1 _14552_ ( .A(_06583_ ), .B(_06461_ ), .C1(\ID_EX_typ [0] ), .C2(_02729_ ), .ZN(_06584_ ) );
NAND3_X1 _14553_ ( .A1(_05102_ ), .A2(_06457_ ), .A3(_06459_ ), .ZN(_06585_ ) );
MUX2_X1 _14554_ ( .A(_05388_ ), .B(_03945_ ), .S(_06429_ ), .Z(_06586_ ) );
OAI211_X1 _14555_ ( .A(_06584_ ), .B(_06585_ ), .C1(_06462_ ), .C2(_06586_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
AOI21_X1 _14556_ ( .A(_06441_ ), .B1(_05118_ ), .B2(_05119_ ), .ZN(_06587_ ) );
NOR2_X1 _14557_ ( .A1(_03251_ ), .A2(\ID_EX_imm [5] ), .ZN(_06588_ ) );
AOI21_X1 _14558_ ( .A(_06588_ ), .B1(_05120_ ), .B2(\ID_EX_typ [2] ), .ZN(_06589_ ) );
NAND3_X1 _14559_ ( .A1(_02650_ ), .A2(_02651_ ), .A3(_03252_ ), .ZN(_06590_ ) );
AOI211_X1 _14560_ ( .A(_06432_ ), .B(_06587_ ), .C1(_06589_ ), .C2(_06590_ ), .ZN(_06591_ ) );
AND4_X1 _14561_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06592_ ) );
AOI211_X1 _14562_ ( .A(_06426_ ), .B(_06592_ ), .C1(_03995_ ), .C2(_06580_ ), .ZN(_06593_ ) );
NOR2_X1 _14563_ ( .A1(_06591_ ), .A2(_06593_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
AOI21_X1 _14564_ ( .A(\ID_EX_typ [0] ), .B1(_02655_ ), .B2(_02675_ ), .ZN(_06594_ ) );
AND2_X1 _14565_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [4] ), .ZN(_06595_ ) );
OAI221_X1 _14566_ ( .A(_06457_ ), .B1(_05402_ ), .B2(_05143_ ), .C1(_06594_ ), .C2(_06595_ ), .ZN(_06596_ ) );
AND3_X1 _14567_ ( .A1(_03951_ ), .A2(_03971_ ), .A3(_06429_ ), .ZN(_06597_ ) );
AND3_X1 _14568_ ( .A1(_06490_ ), .A2(\ID_EX_pc [4] ), .A3(\ID_EX_typ [7] ), .ZN(_06598_ ) );
OAI21_X1 _14569_ ( .A(_06488_ ), .B1(_06597_ ), .B2(_06598_ ), .ZN(_06599_ ) );
NAND2_X1 _14570_ ( .A1(_04781_ ), .A2(\mepc [4] ), .ZN(_06600_ ) );
NOR3_X1 _14571_ ( .A1(_05136_ ), .A2(_05138_ ), .A3(_05139_ ), .ZN(_06601_ ) );
NAND3_X1 _14572_ ( .A1(_05142_ ), .A2(_06600_ ), .A3(_06601_ ), .ZN(_06602_ ) );
INV_X1 _14573_ ( .A(_05134_ ), .ZN(_06603_ ) );
NAND4_X1 _14574_ ( .A1(_06602_ ), .A2(_06603_ ), .A3(_06461_ ), .A4(_06459_ ), .ZN(_06604_ ) );
NAND3_X1 _14575_ ( .A1(_06596_ ), .A2(_06599_ ), .A3(_06604_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
AOI21_X1 _14576_ ( .A(\ID_EX_typ [0] ), .B1(_02809_ ), .B2(_02828_ ), .ZN(_06605_ ) );
AND2_X1 _14577_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [3] ), .ZN(_06606_ ) );
OAI221_X1 _14578_ ( .A(_06426_ ), .B1(_05402_ ), .B2(_05157_ ), .C1(_06605_ ), .C2(_06606_ ), .ZN(_06607_ ) );
NAND2_X1 _14579_ ( .A1(_04781_ ), .A2(\mepc [3] ), .ZN(_06608_ ) );
NOR3_X1 _14580_ ( .A1(_05136_ ), .A2(_05152_ ), .A3(_05153_ ), .ZN(_06609_ ) );
NAND3_X1 _14581_ ( .A1(_05156_ ), .A2(_06608_ ), .A3(_06609_ ), .ZN(_06610_ ) );
INV_X1 _14582_ ( .A(_05150_ ), .ZN(_06611_ ) );
NAND4_X1 _14583_ ( .A1(_06610_ ), .A2(_06611_ ), .A3(_06426_ ), .A4(_06458_ ), .ZN(_06612_ ) );
AND3_X1 _14584_ ( .A1(_06490_ ), .A2(\ID_EX_pc [3] ), .A3(\ID_EX_typ [7] ), .ZN(_06613_ ) );
AOI21_X1 _14585_ ( .A(_06613_ ), .B1(_04043_ ), .B2(_06580_ ), .ZN(_06614_ ) );
OAI211_X1 _14586_ ( .A(_06607_ ), .B(_06612_ ), .C1(_06427_ ), .C2(_06614_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
INV_X1 _14587_ ( .A(_05181_ ), .ZN(_06615_ ) );
AOI22_X1 _14588_ ( .A1(_04389_ ), .A2(_04759_ ), .B1(_06615_ ), .B2(\ID_EX_typ [2] ), .ZN(_06616_ ) );
OAI211_X1 _14589_ ( .A(_06616_ ), .B(_06457_ ), .C1(_04820_ ), .C2(\ID_EX_imm [2] ), .ZN(_06617_ ) );
AND3_X1 _14590_ ( .A1(_05178_ ), .A2(_05180_ ), .A3(_06434_ ), .ZN(_06618_ ) );
NAND2_X1 _14591_ ( .A1(_06618_ ), .A2(_06459_ ), .ZN(_06619_ ) );
AND3_X1 _14592_ ( .A1(_04017_ ), .A2(_04018_ ), .A3(_06429_ ), .ZN(_06620_ ) );
AND3_X1 _14593_ ( .A1(_06490_ ), .A2(\ID_EX_pc [2] ), .A3(\ID_EX_typ [7] ), .ZN(_06621_ ) );
OAI21_X1 _14594_ ( .A(_06488_ ), .B1(_06620_ ), .B2(_06621_ ), .ZN(_06622_ ) );
NAND3_X1 _14595_ ( .A1(_06617_ ), .A2(_06619_ ), .A3(_06622_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
AOI21_X1 _14596_ ( .A(_04692_ ), .B1(_04776_ ), .B2(_04779_ ), .ZN(_06623_ ) );
NAND3_X1 _14597_ ( .A1(_04745_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_04699_ ), .ZN(_06624_ ) );
NAND2_X1 _14598_ ( .A1(_04698_ ), .A2(_06624_ ), .ZN(_06625_ ) );
AND4_X1 _14599_ ( .A1(\mycsreg.CSReg[3][29] ), .A2(_04737_ ), .A3(_05012_ ), .A4(_05013_ ), .ZN(_06626_ ) );
NOR3_X1 _14600_ ( .A1(_06625_ ), .A2(_05135_ ), .A3(_06626_ ), .ZN(_06627_ ) );
NAND2_X1 _14601_ ( .A1(_06623_ ), .A2(_06627_ ), .ZN(_06628_ ) );
INV_X1 _14602_ ( .A(\EX_LS_result_csreg_mem [29] ), .ZN(_06629_ ) );
NAND4_X1 _14603_ ( .A1(_04779_ ), .A2(_06629_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_06630_ ) );
NAND2_X1 _14604_ ( .A1(_06628_ ), .A2(_06630_ ), .ZN(_06631_ ) );
AOI22_X1 _14605_ ( .A1(_03156_ ), .A2(_04759_ ), .B1(\ID_EX_typ [2] ), .B2(_06631_ ), .ZN(_06632_ ) );
OAI211_X1 _14606_ ( .A(_06632_ ), .B(_06461_ ), .C1(_04820_ ), .C2(\ID_EX_imm [29] ), .ZN(_06633_ ) );
NAND4_X1 _14607_ ( .A1(_06628_ ), .A2(_06630_ ), .A3(_06426_ ), .A4(_06458_ ), .ZN(_06634_ ) );
AND3_X1 _14608_ ( .A1(_06490_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_typ [7] ), .ZN(_06635_ ) );
AOI21_X1 _14609_ ( .A(_06635_ ), .B1(_03653_ ), .B2(_06580_ ), .ZN(_06636_ ) );
OAI211_X1 _14610_ ( .A(_06633_ ), .B(_06634_ ), .C1(_06427_ ), .C2(_06636_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
AND3_X1 _14611_ ( .A1(_03404_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_03415_ ), .ZN(_06637_ ) );
NAND4_X1 _14612_ ( .A1(_03421_ ), .A2(_03425_ ), .A3(\mycsreg.CSReg[3][1] ), .A4(_04739_ ), .ZN(_06638_ ) );
NAND4_X1 _14613_ ( .A1(_04860_ ), .A2(_03425_ ), .A3(\mepc [1] ), .A4(_04739_ ), .ZN(_06639_ ) );
NAND2_X1 _14614_ ( .A1(_06638_ ), .A2(_06639_ ), .ZN(_06640_ ) );
NOR2_X1 _14615_ ( .A1(_06637_ ), .A2(_06640_ ), .ZN(_06641_ ) );
AOI22_X1 _14616_ ( .A1(_06641_ ), .A2(_05191_ ), .B1(_03442_ ), .B2(_03444_ ), .ZN(_06642_ ) );
AND3_X1 _14617_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(\EX_LS_result_csreg_mem [1] ), .ZN(_06643_ ) );
NOR2_X1 _14618_ ( .A1(_06642_ ), .A2(_06643_ ), .ZN(_06644_ ) );
NAND4_X1 _14619_ ( .A1(_04778_ ), .A2(_06309_ ), .A3(_04774_ ), .A4(_04773_ ), .ZN(_06645_ ) );
AND4_X1 _14620_ ( .A1(\mycsreg.CSReg[3][1] ), .A2(_03420_ ), .A3(_03435_ ), .A4(_03400_ ), .ZN(_06646_ ) );
AOI21_X1 _14621_ ( .A(_06646_ ), .B1(\mepc [1] ), .B2(_04696_ ), .ZN(_06647_ ) );
INV_X1 _14622_ ( .A(_06637_ ), .ZN(_06648_ ) );
NAND3_X1 _14623_ ( .A1(_06647_ ), .A2(_05191_ ), .A3(_06648_ ), .ZN(_06649_ ) );
OAI211_X1 _14624_ ( .A(_06645_ ), .B(_06439_ ), .C1(_06542_ ), .C2(_06649_ ), .ZN(_06650_ ) );
INV_X1 _14625_ ( .A(_06650_ ), .ZN(_06651_ ) );
AOI21_X1 _14626_ ( .A(_06651_ ), .B1(_02760_ ), .B2(_04758_ ), .ZN(_06652_ ) );
OR2_X1 _14627_ ( .A1(_03250_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_06653_ ) );
AOI221_X4 _14628_ ( .A(_06422_ ), .B1(\ID_EX_typ [2] ), .B2(_06644_ ), .C1(_06652_ ), .C2(_06653_ ), .ZN(_06654_ ) );
AND4_X1 _14629_ ( .A1(_03274_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06655_ ) );
AOI211_X1 _14630_ ( .A(_06434_ ), .B(_06655_ ), .C1(_04066_ ), .C2(_06446_ ), .ZN(_06656_ ) );
OR2_X1 _14631_ ( .A1(_06654_ ), .A2(_06656_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
NAND3_X1 _14632_ ( .A1(_04093_ ), .A2(_04091_ ), .A3(_06446_ ), .ZN(_06657_ ) );
OAI211_X1 _14633_ ( .A(_06657_ ), .B(_06432_ ), .C1(\ID_EX_pc [0] ), .C2(_06580_ ), .ZN(_06658_ ) );
NOR2_X1 _14634_ ( .A1(_05236_ ), .A2(_05237_ ), .ZN(_06659_ ) );
OAI22_X1 _14635_ ( .A1(_06659_ ), .A2(_06441_ ), .B1(_04759_ ), .B2(_02763_ ), .ZN(_06660_ ) );
AOI21_X1 _14636_ ( .A(_06660_ ), .B1(_04820_ ), .B2(_04071_ ), .ZN(_06661_ ) );
INV_X1 _14637_ ( .A(_06659_ ), .ZN(_06662_ ) );
OAI21_X1 _14638_ ( .A(_06457_ ), .B1(_06662_ ), .B2(_05402_ ), .ZN(_06663_ ) );
OAI21_X1 _14639_ ( .A(_06658_ ), .B1(_06661_ ), .B2(_06663_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
AND4_X1 _14640_ ( .A1(\mepc [28] ), .A2(_03429_ ), .A3(_05012_ ), .A4(_05013_ ), .ZN(_06664_ ) );
AND4_X1 _14641_ ( .A1(\mycsreg.CSReg[3][28] ), .A2(_04737_ ), .A3(_05012_ ), .A4(_04740_ ), .ZN(_06665_ ) );
NOR3_X1 _14642_ ( .A1(_04734_ ), .A2(_06664_ ), .A3(_06665_ ), .ZN(_06666_ ) );
NAND3_X1 _14643_ ( .A1(_04748_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_04749_ ), .ZN(_06667_ ) );
AND2_X1 _14644_ ( .A1(_04993_ ), .A2(_06667_ ), .ZN(_06668_ ) );
AOI22_X1 _14645_ ( .A1(_06666_ ), .A2(_06668_ ), .B1(_03443_ ), .B2(_03445_ ), .ZN(_06669_ ) );
AND3_X1 _14646_ ( .A1(_03442_ ), .A2(_03444_ ), .A3(\EX_LS_result_csreg_mem [28] ), .ZN(_06670_ ) );
OR2_X1 _14647_ ( .A1(_06669_ ), .A2(_06670_ ), .ZN(_06671_ ) );
OAI21_X1 _14648_ ( .A(_06458_ ), .B1(_06669_ ), .B2(_06670_ ), .ZN(_06672_ ) );
NAND2_X1 _14649_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [28] ), .ZN(_06673_ ) );
NAND2_X1 _14650_ ( .A1(_06672_ ), .A2(_06673_ ), .ZN(_06674_ ) );
AOI21_X1 _14651_ ( .A(\ID_EX_typ [0] ), .B1(_02362_ ), .B2(_02387_ ), .ZN(_06675_ ) );
OAI221_X1 _14652_ ( .A(_06435_ ), .B1(_05402_ ), .B2(_06671_ ), .C1(_06674_ ), .C2(_06675_ ), .ZN(_06676_ ) );
NAND4_X1 _14653_ ( .A1(_04986_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06677_ ) );
OAI211_X1 _14654_ ( .A(_06488_ ), .B(_06677_ ), .C1(_03631_ ), .C2(_06428_ ), .ZN(_06678_ ) );
NAND2_X1 _14655_ ( .A1(_06676_ ), .A2(_06678_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND3_X1 _14656_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [27] ), .ZN(_06679_ ) );
AND2_X1 _14657_ ( .A1(_05218_ ), .A2(_06679_ ), .ZN(_06680_ ) );
AOI22_X1 _14658_ ( .A1(_06680_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_03077_ ), .ZN(_06681_ ) );
OAI211_X1 _14659_ ( .A(_06681_ ), .B(_06461_ ), .C1(\ID_EX_typ [0] ), .C2(_03560_ ), .ZN(_06682_ ) );
AOI21_X1 _14660_ ( .A(_06423_ ), .B1(_05218_ ), .B2(_06679_ ), .ZN(_06683_ ) );
NAND2_X1 _14661_ ( .A1(_06683_ ), .A2(_06459_ ), .ZN(_06684_ ) );
AND3_X1 _14662_ ( .A1(_06490_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_06685_ ) );
AOI21_X1 _14663_ ( .A(_06685_ ), .B1(_03559_ ), .B2(_06580_ ), .ZN(_06686_ ) );
OAI211_X1 _14664_ ( .A(_06682_ ), .B(_06684_ ), .C1(_06427_ ), .C2(_06686_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
AND3_X1 _14665_ ( .A1(_04745_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_04699_ ), .ZN(_06687_ ) );
NAND4_X1 _14666_ ( .A1(_04836_ ), .A2(_04684_ ), .A3(\mycsreg.CSReg[3][26] ), .A4(_04685_ ), .ZN(_06688_ ) );
NAND4_X1 _14667_ ( .A1(_03429_ ), .A2(_04684_ ), .A3(\mepc [26] ), .A4(_04685_ ), .ZN(_06689_ ) );
NAND2_X1 _14668_ ( .A1(_06688_ ), .A2(_06689_ ), .ZN(_06690_ ) );
NOR2_X1 _14669_ ( .A1(_06687_ ), .A2(_06690_ ), .ZN(_06691_ ) );
AOI22_X1 _14670_ ( .A1(_06691_ ), .A2(_05246_ ), .B1(_03443_ ), .B2(_03445_ ), .ZN(_06692_ ) );
AND3_X1 _14671_ ( .A1(_03443_ ), .A2(_03445_ ), .A3(\EX_LS_result_csreg_mem [26] ), .ZN(_06693_ ) );
NOR2_X1 _14672_ ( .A1(_06692_ ), .A2(_06693_ ), .ZN(_06694_ ) );
AOI22_X1 _14673_ ( .A1(_06694_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06695_ ) );
OAI211_X1 _14674_ ( .A(_06695_ ), .B(_06461_ ), .C1(\ID_EX_typ [0] ), .C2(_03120_ ), .ZN(_06696_ ) );
OR2_X1 _14675_ ( .A1(_06543_ ), .A2(\EX_LS_result_csreg_mem [26] ), .ZN(_06697_ ) );
INV_X1 _14676_ ( .A(_06687_ ), .ZN(_06698_ ) );
NAND4_X1 _14677_ ( .A1(_04738_ ), .A2(_05193_ ), .A3(\mycsreg.CSReg[3][26] ), .A4(_04701_ ), .ZN(_06699_ ) );
NAND4_X1 _14678_ ( .A1(_06698_ ), .A2(_05246_ ), .A3(_05245_ ), .A4(_06699_ ), .ZN(_06700_ ) );
OR2_X1 _14679_ ( .A1(_06542_ ), .A2(_06700_ ), .ZN(_06701_ ) );
NAND4_X1 _14680_ ( .A1(_06697_ ), .A2(_06701_ ), .A3(_06426_ ), .A4(_06458_ ), .ZN(_06702_ ) );
AND3_X1 _14681_ ( .A1(_06490_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_06703_ ) );
AOI21_X1 _14682_ ( .A(_06703_ ), .B1(_03537_ ), .B2(_06580_ ), .ZN(_06704_ ) );
OAI211_X1 _14683_ ( .A(_06696_ ), .B(_06702_ ), .C1(_06704_ ), .C2(_06427_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
NOR2_X1 _14684_ ( .A1(_03250_ ), .A2(\ID_EX_imm [25] ), .ZN(_06705_ ) );
OR2_X1 _14685_ ( .A1(_05273_ ), .A2(_05275_ ), .ZN(_06706_ ) );
AOI221_X4 _14686_ ( .A(_06705_ ), .B1(_06706_ ), .B2(\ID_EX_typ [2] ), .C1(_04537_ ), .C2(_04758_ ), .ZN(_06707_ ) );
NOR3_X1 _14687_ ( .A1(_05273_ ), .A2(_05275_ ), .A3(_06441_ ), .ZN(_06708_ ) );
OAI21_X1 _14688_ ( .A(_06559_ ), .B1(_06707_ ), .B2(_06708_ ), .ZN(_06709_ ) );
AND4_X1 _14689_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06710_ ) );
AOI21_X1 _14690_ ( .A(_06710_ ), .B1(_03609_ ), .B2(_06580_ ), .ZN(_06711_ ) );
OAI21_X1 _14691_ ( .A(_06709_ ), .B1(_06462_ ), .B2(_06711_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _14692_ ( .A(_05280_ ), .B1(_04775_ ), .B2(_04778_ ), .ZN(_06712_ ) );
AND4_X1 _14693_ ( .A1(\mycsreg.CSReg[3][24] ), .A2(_04737_ ), .A3(_03436_ ), .A4(_04740_ ), .ZN(_06713_ ) );
NOR3_X1 _14694_ ( .A1(_05136_ ), .A2(_04784_ ), .A3(_06713_ ), .ZN(_06714_ ) );
NAND2_X1 _14695_ ( .A1(_04697_ ), .A2(\mepc [24] ), .ZN(_06715_ ) );
NAND3_X1 _14696_ ( .A1(_04748_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_04749_ ), .ZN(_06716_ ) );
AND2_X1 _14697_ ( .A1(_06715_ ), .A2(_06716_ ), .ZN(_06717_ ) );
NAND3_X1 _14698_ ( .A1(_06712_ ), .A2(_06714_ ), .A3(_06717_ ), .ZN(_06718_ ) );
INV_X1 _14699_ ( .A(\EX_LS_result_csreg_mem [24] ), .ZN(_06719_ ) );
NAND4_X1 _14700_ ( .A1(_04779_ ), .A2(_06719_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_06720_ ) );
NAND2_X1 _14701_ ( .A1(_06718_ ), .A2(_06720_ ), .ZN(_06721_ ) );
AOI22_X1 _14702_ ( .A1(_04531_ ), .A2(_04759_ ), .B1(\ID_EX_typ [2] ), .B2(_06721_ ), .ZN(_06722_ ) );
OAI211_X1 _14703_ ( .A(_06722_ ), .B(_06461_ ), .C1(_03252_ ), .C2(\ID_EX_imm [24] ), .ZN(_06723_ ) );
NAND4_X1 _14704_ ( .A1(_06718_ ), .A2(_06720_ ), .A3(_06426_ ), .A4(_06458_ ), .ZN(_06724_ ) );
AND3_X1 _14705_ ( .A1(_06490_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_typ [7] ), .ZN(_06725_ ) );
AOI21_X1 _14706_ ( .A(_06725_ ), .B1(_03586_ ), .B2(_06580_ ), .ZN(_06726_ ) );
OAI211_X1 _14707_ ( .A(_06723_ ), .B(_06724_ ), .C1(_06427_ ), .C2(_06726_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
OR2_X1 _14708_ ( .A1(_05313_ ), .A2(_05315_ ), .ZN(_06727_ ) );
AOI22_X1 _14709_ ( .A1(_06727_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02436_ ), .ZN(_06728_ ) );
OAI211_X1 _14710_ ( .A(_06728_ ), .B(_06461_ ), .C1(\ID_EX_typ [0] ), .C2(_02438_ ), .ZN(_06729_ ) );
NOR3_X1 _14711_ ( .A1(_05313_ ), .A2(_05315_ ), .A3(_06423_ ), .ZN(_06730_ ) );
NAND2_X1 _14712_ ( .A1(_06730_ ), .A2(_06459_ ), .ZN(_06731_ ) );
MUX2_X1 _14713_ ( .A(_03329_ ), .B(_03730_ ), .S(_06430_ ), .Z(_06732_ ) );
OAI211_X1 _14714_ ( .A(_06729_ ), .B(_06731_ ), .C1(_06732_ ), .C2(_06427_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
AND2_X1 _14715_ ( .A1(_05334_ ), .A2(_05335_ ), .ZN(_06733_ ) );
OAI22_X1 _14716_ ( .A1(_06733_ ), .A2(_06440_ ), .B1(_03251_ ), .B2(_02412_ ), .ZN(_06734_ ) );
AOI21_X1 _14717_ ( .A(_06734_ ), .B1(_04759_ ), .B2(_02411_ ), .ZN(_06735_ ) );
INV_X1 _14718_ ( .A(_06733_ ), .ZN(_06736_ ) );
OAI21_X1 _14719_ ( .A(_06434_ ), .B1(_06736_ ), .B2(_04649_ ), .ZN(_06737_ ) );
NOR2_X1 _14720_ ( .A1(_06735_ ), .A2(_06737_ ), .ZN(_06738_ ) );
NOR4_X1 _14721_ ( .A1(_02270_ ), .A2(_02267_ ), .A3(_02262_ ), .A4(\ID_EX_pc [22] ), .ZN(_06739_ ) );
AOI211_X1 _14722_ ( .A(_06434_ ), .B(_06739_ ), .C1(_03752_ ), .C2(_06446_ ), .ZN(_06740_ ) );
OR2_X1 _14723_ ( .A1(_06738_ ), .A2(_06740_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
INV_X1 _14724_ ( .A(\EX_LS_result_csreg_mem [31] ), .ZN(_06741_ ) );
NAND4_X1 _14725_ ( .A1(_04789_ ), .A2(_06741_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_06742_ ) );
NAND3_X1 _14726_ ( .A1(_04839_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04700_ ), .ZN(_06743_ ) );
NAND4_X1 _14727_ ( .A1(_04738_ ), .A2(_05193_ ), .A3(\mycsreg.CSReg[3][31] ), .A4(_04741_ ), .ZN(_06744_ ) );
NAND4_X1 _14728_ ( .A1(_05372_ ), .A2(_05373_ ), .A3(_06743_ ), .A4(_06744_ ), .ZN(_06745_ ) );
OAI211_X1 _14729_ ( .A(_06742_ ), .B(_06458_ ), .C1(_06542_ ), .C2(_06745_ ), .ZN(_06746_ ) );
AOI21_X1 _14730_ ( .A(\ID_EX_typ [0] ), .B1(_03161_ ), .B2(_03183_ ), .ZN(_06747_ ) );
AND2_X1 _14731_ ( .A1(\ID_EX_typ [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_06748_ ) );
OAI21_X1 _14732_ ( .A(_06746_ ), .B1(_06747_ ), .B2(_06748_ ), .ZN(_06749_ ) );
AND3_X1 _14733_ ( .A1(_04839_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04749_ ), .ZN(_06750_ ) );
NAND4_X1 _14734_ ( .A1(_04836_ ), .A2(_03437_ ), .A3(\mycsreg.CSReg[3][31] ), .A4(_04741_ ), .ZN(_06751_ ) );
NAND4_X1 _14735_ ( .A1(_03429_ ), .A2(_03437_ ), .A3(\mepc [31] ), .A4(_04741_ ), .ZN(_06752_ ) );
NAND2_X1 _14736_ ( .A1(_06751_ ), .A2(_06752_ ), .ZN(_06753_ ) );
NOR2_X1 _14737_ ( .A1(_06750_ ), .A2(_06753_ ), .ZN(_06754_ ) );
AOI22_X1 _14738_ ( .A1(_06754_ ), .A2(_05373_ ), .B1(_04731_ ), .B2(_04732_ ), .ZN(_06755_ ) );
AND3_X1 _14739_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [31] ), .ZN(_06756_ ) );
NOR2_X1 _14740_ ( .A1(_06755_ ), .A2(_06756_ ), .ZN(_06757_ ) );
INV_X1 _14741_ ( .A(_06757_ ), .ZN(_06758_ ) );
OAI211_X1 _14742_ ( .A(_06749_ ), .B(_06457_ ), .C1(_05402_ ), .C2(_06758_ ), .ZN(_06759_ ) );
AND3_X1 _14743_ ( .A1(_06490_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06760_ ) );
AOI21_X1 _14744_ ( .A(_06760_ ), .B1(_03676_ ), .B2(_06580_ ), .ZN(_06761_ ) );
OAI21_X1 _14745_ ( .A(_06759_ ), .B1(_06462_ ), .B2(_06761_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
OR2_X1 _14746_ ( .A1(_05356_ ), .A2(_06432_ ), .ZN(_06762_ ) );
NOR3_X1 _14747_ ( .A1(_04299_ ), .A2(\ID_EX_typ [1] ), .A3(\ID_EX_typ [0] ), .ZN(_06763_ ) );
AND2_X2 _14748_ ( .A1(fanout_net_10 ), .A2(\ID_EX_typ [2] ), .ZN(_06764_ ) );
AND2_X1 _14749_ ( .A1(_06763_ ), .A2(_06764_ ), .ZN(_06765_ ) );
BUF_X4 _14750_ ( .A(_06765_ ), .Z(_06766_ ) );
NAND2_X1 _14751_ ( .A1(_05343_ ), .A2(_06766_ ), .ZN(_06767_ ) );
NOR3_X1 _14752_ ( .A1(_04292_ ), .A2(\ID_EX_typ [0] ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_06768_ ) );
AND2_X2 _14753_ ( .A1(_06768_ ), .A2(_06764_ ), .ZN(_06769_ ) );
INV_X1 _14754_ ( .A(_06769_ ), .ZN(_06770_ ) );
OAI21_X1 _14755_ ( .A(_06767_ ), .B1(_02442_ ), .B2(_06770_ ), .ZN(_06771_ ) );
INV_X1 _14756_ ( .A(_04589_ ), .ZN(_06772_ ) );
NAND2_X1 _14757_ ( .A1(_06772_ ), .A2(_03898_ ), .ZN(_06773_ ) );
AND2_X1 _14758_ ( .A1(_06773_ ), .A2(_04601_ ), .ZN(_06774_ ) );
INV_X1 _14759_ ( .A(_03801_ ), .ZN(_06775_ ) );
OR2_X1 _14760_ ( .A1(_06774_ ), .A2(_06775_ ), .ZN(_06776_ ) );
AND2_X1 _14761_ ( .A1(_06776_ ), .A2(_04607_ ), .ZN(_06777_ ) );
XNOR2_X1 _14762_ ( .A(_06777_ ), .B(_03779_ ), .ZN(_06778_ ) );
AND3_X1 _14763_ ( .A1(_03467_ ), .A2(\ID_EX_typ [3] ), .A3(_04649_ ), .ZN(_06779_ ) );
AND2_X1 _14764_ ( .A1(_06779_ ), .A2(_04299_ ), .ZN(_06780_ ) );
BUF_X4 _14765_ ( .A(_06780_ ), .Z(_06781_ ) );
BUF_X4 _14766_ ( .A(_06781_ ), .Z(_06782_ ) );
AOI21_X1 _14767_ ( .A(_06771_ ), .B1(_06778_ ), .B2(_06782_ ), .ZN(_06783_ ) );
AND2_X1 _14768_ ( .A1(_02263_ ), .A2(_02270_ ), .ZN(_06784_ ) );
INV_X1 _14769_ ( .A(_06784_ ), .ZN(_06785_ ) );
BUF_X4 _14770_ ( .A(_06785_ ), .Z(_06786_ ) );
BUF_X4 _14771_ ( .A(_06786_ ), .Z(_06787_ ) );
OAI21_X1 _14772_ ( .A(_04661_ ), .B1(_06783_ ), .B2(_06787_ ), .ZN(_06788_ ) );
AND2_X2 _14773_ ( .A1(_04338_ ), .A2(_04343_ ), .ZN(_06789_ ) );
AND3_X4 _14774_ ( .A1(_06789_ ), .A2(_04333_ ), .A3(_04326_ ), .ZN(_06790_ ) );
INV_X2 _14775_ ( .A(_06790_ ), .ZN(_06791_ ) );
AND2_X1 _14776_ ( .A1(_04361_ ), .A2(_04427_ ), .ZN(_06792_ ) );
AND3_X1 _14777_ ( .A1(_04351_ ), .A2(_04355_ ), .A3(_06792_ ), .ZN(_06793_ ) );
INV_X1 _14778_ ( .A(_06793_ ), .ZN(_06794_ ) );
INV_X1 _14779_ ( .A(_04373_ ), .ZN(_06795_ ) );
INV_X1 _14780_ ( .A(_04071_ ), .ZN(_06796_ ) );
NOR2_X4 _14781_ ( .A1(_04386_ ), .A2(_06796_ ), .ZN(_06797_ ) );
INV_X1 _14782_ ( .A(_06797_ ), .ZN(_06798_ ) );
NOR3_X2 _14783_ ( .A1(_06798_ ), .A2(_04382_ ), .A3(_04383_ ), .ZN(_06799_ ) );
INV_X1 _14784_ ( .A(_06799_ ), .ZN(_06800_ ) );
INV_X1 _14785_ ( .A(_04382_ ), .ZN(_06801_ ) );
AOI21_X2 _14786_ ( .A(_06795_ ), .B1(_06800_ ), .B2(_06801_ ), .ZN(_06802_ ) );
INV_X1 _14787_ ( .A(_06802_ ), .ZN(_06803_ ) );
BUF_X4 _14788_ ( .A(_04376_ ), .Z(_06804_ ) );
INV_X1 _14789_ ( .A(_06804_ ), .ZN(_06805_ ) );
OAI221_X1 _14790_ ( .A(_06803_ ), .B1(_02833_ ), .B2(_06805_ ), .C1(_04389_ ), .C2(_04372_ ), .ZN(_06806_ ) );
NOR2_X1 _14791_ ( .A1(_06804_ ), .A2(_02829_ ), .ZN(_06807_ ) );
INV_X1 _14792_ ( .A(_06807_ ), .ZN(_06808_ ) );
AND2_X1 _14793_ ( .A1(_04409_ ), .A2(_04414_ ), .ZN(_06809_ ) );
AND3_X1 _14794_ ( .A1(_04399_ ), .A2(_06809_ ), .A3(_04403_ ), .ZN(_06810_ ) );
NAND3_X1 _14795_ ( .A1(_06806_ ), .A2(_06808_ ), .A3(_06810_ ), .ZN(_06811_ ) );
INV_X2 _14796_ ( .A(_04403_ ), .ZN(_06812_ ) );
INV_X1 _14797_ ( .A(_04421_ ), .ZN(_06813_ ) );
INV_X1 _14798_ ( .A(_02677_ ), .ZN(_06814_ ) );
NOR2_X4 _14799_ ( .A1(_04413_ ), .A2(_06814_ ), .ZN(_06815_ ) );
OAI21_X1 _14800_ ( .A(_06813_ ), .B1(_04420_ ), .B2(_06815_ ), .ZN(_06816_ ) );
NOR4_X1 _14801_ ( .A1(_06812_ ), .A2(_06816_ ), .A3(_04397_ ), .A4(_04398_ ), .ZN(_06817_ ) );
NOR2_X1 _14802_ ( .A1(_04402_ ), .A2(_04417_ ), .ZN(_06818_ ) );
AOI211_X1 _14803_ ( .A(_04397_ ), .B(_06817_ ), .C1(_04399_ ), .C2(_06818_ ), .ZN(_06819_ ) );
AOI211_X2 _14804_ ( .A(_06791_ ), .B(_06794_ ), .C1(_06811_ ), .C2(_06819_ ), .ZN(_06820_ ) );
NOR2_X4 _14805_ ( .A1(_04360_ ), .A2(_04428_ ), .ZN(_06821_ ) );
AOI21_X1 _14806_ ( .A(_04367_ ), .B1(_04427_ ), .B2(_06821_ ), .ZN(_06822_ ) );
INV_X1 _14807_ ( .A(_04355_ ), .ZN(_06823_ ) );
OR4_X1 _14808_ ( .A1(_04350_ ), .A2(_06822_ ), .A3(_04349_ ), .A4(_06823_ ), .ZN(_06824_ ) );
NOR2_X1 _14809_ ( .A1(_04354_ ), .A2(_04434_ ), .ZN(_06825_ ) );
AOI21_X1 _14810_ ( .A(_04349_ ), .B1(_04351_ ), .B2(_06825_ ), .ZN(_06826_ ) );
AOI21_X2 _14811_ ( .A(_06791_ ), .B1(_06824_ ), .B2(_06826_ ), .ZN(_06827_ ) );
INV_X1 _14812_ ( .A(_04194_ ), .ZN(_06828_ ) );
NOR2_X1 _14813_ ( .A1(_04337_ ), .A2(_06828_ ), .ZN(_06829_ ) );
AND2_X1 _14814_ ( .A1(_04337_ ), .A2(_06828_ ), .ZN(_06830_ ) );
INV_X1 _14815_ ( .A(_06830_ ), .ZN(_06831_ ) );
AND2_X1 _14816_ ( .A1(_04341_ ), .A2(_02862_ ), .ZN(_06832_ ) );
AOI21_X1 _14817_ ( .A(_06829_ ), .B1(_06831_ ), .B2(_06832_ ), .ZN(_06833_ ) );
INV_X1 _14818_ ( .A(_04326_ ), .ZN(_06834_ ) );
NOR4_X1 _14819_ ( .A1(_06833_ ), .A2(_06834_ ), .A3(_04332_ ), .A4(_04331_ ), .ZN(_06835_ ) );
NOR4_X1 _14820_ ( .A1(_04331_ ), .A2(_04332_ ), .A3(_04442_ ), .A4(_04325_ ), .ZN(_06836_ ) );
OR4_X4 _14821_ ( .A1(_04331_ ), .A2(_06827_ ), .A3(_06835_ ), .A4(_06836_ ), .ZN(_06837_ ) );
NOR2_X4 _14822_ ( .A1(_06820_ ), .A2(_06837_ ), .ZN(_06838_ ) );
INV_X1 _14823_ ( .A(_06838_ ), .ZN(_06839_ ) );
INV_X1 _14824_ ( .A(_04487_ ), .ZN(_06840_ ) );
NOR3_X1 _14825_ ( .A1(_04490_ ), .A2(_06840_ ), .A3(_04491_ ), .ZN(_06841_ ) );
AND4_X4 _14826_ ( .A1(_04496_ ), .A2(_06839_ ), .A3(_04476_ ), .A4(_06841_ ), .ZN(_06842_ ) );
INV_X1 _14827_ ( .A(_02580_ ), .ZN(_06843_ ) );
NOR2_X1 _14828_ ( .A1(_04486_ ), .A2(_06843_ ), .ZN(_06844_ ) );
AOI21_X1 _14829_ ( .A(_04491_ ), .B1(_04472_ ), .B2(_06844_ ), .ZN(_06845_ ) );
NOR3_X1 _14830_ ( .A1(_06845_ ), .A2(_04497_ ), .A3(_04477_ ), .ZN(_06846_ ) );
NOR2_X1 _14831_ ( .A1(_04475_ ), .A2(_06472_ ), .ZN(_06847_ ) );
INV_X1 _14832_ ( .A(_06847_ ), .ZN(_06848_ ) );
NOR2_X1 _14833_ ( .A1(_04482_ ), .A2(_06848_ ), .ZN(_06849_ ) );
NOR3_X1 _14834_ ( .A1(_06846_ ), .A2(_04481_ ), .A3(_06849_ ), .ZN(_06850_ ) );
INV_X1 _14835_ ( .A(_06850_ ), .ZN(_06851_ ) );
NOR2_X4 _14836_ ( .A1(_06842_ ), .A2(_06851_ ), .ZN(_06852_ ) );
NOR2_X1 _14837_ ( .A1(_06852_ ), .A2(_04466_ ), .ZN(_06853_ ) );
INV_X1 _14838_ ( .A(_02485_ ), .ZN(_06854_ ) );
NOR2_X1 _14839_ ( .A1(_04464_ ), .A2(_06854_ ), .ZN(_06855_ ) );
OR3_X1 _14840_ ( .A1(_06853_ ), .A2(_04460_ ), .A3(_06855_ ), .ZN(_06856_ ) );
BUF_X4 _14841_ ( .A(_04290_ ), .Z(_06857_ ) );
NOR2_X1 _14842_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06858_ ) );
INV_X1 _14843_ ( .A(_06858_ ), .ZN(_06859_ ) );
NOR2_X1 _14844_ ( .A1(_06857_ ), .A2(_06859_ ), .ZN(_06860_ ) );
BUF_X4 _14845_ ( .A(_06860_ ), .Z(_06861_ ) );
BUF_X4 _14846_ ( .A(_06861_ ), .Z(_06862_ ) );
OAI21_X1 _14847_ ( .A(_04460_ ), .B1(_06853_ ), .B2(_06855_ ), .ZN(_06863_ ) );
NAND3_X1 _14848_ ( .A1(_06856_ ), .A2(_06862_ ), .A3(_06863_ ), .ZN(_06864_ ) );
AND2_X2 _14849_ ( .A1(_04644_ ), .A2(\ID_EX_typ [2] ), .ZN(_06865_ ) );
BUF_X2 _14850_ ( .A(_06865_ ), .Z(_06866_ ) );
INV_X1 _14851_ ( .A(_03185_ ), .ZN(_06867_ ) );
INV_X1 _14852_ ( .A(_04396_ ), .ZN(_06868_ ) );
NAND2_X1 _14853_ ( .A1(_04300_ ), .A2(_04301_ ), .ZN(_06869_ ) );
OR4_X1 _14854_ ( .A1(_06868_ ), .A2(_04418_ ), .A3(_06869_ ), .A4(_04308_ ), .ZN(_06870_ ) );
NAND2_X1 _14855_ ( .A1(_04511_ ), .A2(_04517_ ), .ZN(_06871_ ) );
NOR4_X1 _14856_ ( .A1(_06870_ ), .A2(_04313_ ), .A3(_04318_ ), .A4(_06871_ ), .ZN(_06872_ ) );
AND4_X1 _14857_ ( .A1(_04448_ ), .A2(_06872_ ), .A3(_04526_ ), .A4(_04530_ ), .ZN(_06873_ ) );
AND4_X1 _14858_ ( .A1(_04360_ ), .A2(_04347_ ), .A3(_04325_ ), .A4(_04486_ ), .ZN(_06874_ ) );
AND3_X1 _14859_ ( .A1(_04469_ ), .A2(_04470_ ), .A3(_04475_ ), .ZN(_06875_ ) );
NAND4_X1 _14860_ ( .A1(_06874_ ), .A2(_04459_ ), .A3(_04480_ ), .A4(_06875_ ), .ZN(_06876_ ) );
INV_X1 _14861_ ( .A(_04337_ ), .ZN(_06877_ ) );
INV_X1 _14862_ ( .A(_04365_ ), .ZN(_06878_ ) );
NOR4_X1 _14863_ ( .A1(_06877_ ), .A2(_06878_ ), .A3(_04438_ ), .A4(_04341_ ), .ZN(_06879_ ) );
NAND3_X1 _14864_ ( .A1(_06879_ ), .A2(_04354_ ), .A3(_04464_ ), .ZN(_06880_ ) );
NOR2_X1 _14865_ ( .A1(_06876_ ), .A2(_06880_ ), .ZN(_06881_ ) );
INV_X1 _14866_ ( .A(_04407_ ), .ZN(_06882_ ) );
AND2_X1 _14867_ ( .A1(_04380_ ), .A2(_04386_ ), .ZN(_06883_ ) );
AND2_X1 _14868_ ( .A1(_06883_ ), .A2(_04372_ ), .ZN(_06884_ ) );
AND2_X1 _14869_ ( .A1(_06884_ ), .A2(_06805_ ), .ZN(_06885_ ) );
AND2_X2 _14870_ ( .A1(_06885_ ), .A2(_04413_ ), .ZN(_06886_ ) );
OAI211_X1 _14871_ ( .A(_06873_ ), .B(_06881_ ), .C1(_06882_ ), .C2(_06886_ ), .ZN(_06887_ ) );
AOI21_X1 _14872_ ( .A(_06867_ ), .B1(_06887_ ), .B2(_04454_ ), .ZN(_06888_ ) );
NAND4_X1 _14873_ ( .A1(_04432_ ), .A2(_06878_ ), .A3(_04429_ ), .A4(_04435_ ), .ZN(_06889_ ) );
AOI21_X1 _14874_ ( .A(_04486_ ), .B1(_04394_ ), .B2(_04395_ ), .ZN(_06890_ ) );
NAND3_X1 _14875_ ( .A1(_06890_ ), .A2(_04418_ ), .A3(_04407_ ), .ZN(_06891_ ) );
NAND4_X1 _14876_ ( .A1(_06877_ ), .A2(_04438_ ), .A3(_04443_ ), .A4(_04341_ ), .ZN(_06892_ ) );
NOR3_X1 _14877_ ( .A1(_06889_ ), .A2(_06891_ ), .A3(_06892_ ), .ZN(_06893_ ) );
NAND4_X1 _14878_ ( .A1(_04311_ ), .A2(_04316_ ), .A3(_04312_ ), .A4(_04317_ ), .ZN(_06894_ ) );
NOR3_X1 _14879_ ( .A1(_04511_ ), .A2(_06894_ ), .A3(_04517_ ), .ZN(_06895_ ) );
AND3_X1 _14880_ ( .A1(_06895_ ), .A2(_06869_ ), .A3(_04308_ ), .ZN(_06896_ ) );
NOR4_X1 _14881_ ( .A1(_04471_ ), .A2(_04480_ ), .A3(_04459_ ), .A4(_04475_ ), .ZN(_06897_ ) );
NOR4_X1 _14882_ ( .A1(_04448_ ), .A2(_04530_ ), .A3(_04464_ ), .A4(_04526_ ), .ZN(_06898_ ) );
NAND4_X1 _14883_ ( .A1(_06893_ ), .A2(_06896_ ), .A3(_06897_ ), .A4(_06898_ ), .ZN(_06899_ ) );
OAI21_X1 _14884_ ( .A(_04501_ ), .B1(_06899_ ), .B2(_06886_ ), .ZN(_06900_ ) );
AND2_X1 _14885_ ( .A1(_06888_ ), .A2(_06900_ ), .ZN(_06901_ ) );
XNOR2_X1 _14886_ ( .A(_06886_ ), .B(_04407_ ), .ZN(_06902_ ) );
AND2_X2 _14887_ ( .A1(_06901_ ), .A2(_06902_ ), .ZN(_06903_ ) );
BUF_X4 _14888_ ( .A(_06903_ ), .Z(_06904_ ) );
BUF_X4 _14889_ ( .A(_04413_ ), .Z(_06905_ ) );
XNOR2_X1 _14890_ ( .A(_06885_ ), .B(_06905_ ), .ZN(_06906_ ) );
NOR2_X1 _14891_ ( .A1(_06906_ ), .A2(_04407_ ), .ZN(_06907_ ) );
BUF_X2 _14892_ ( .A(_06907_ ), .Z(_06908_ ) );
BUF_X2 _14893_ ( .A(_06906_ ), .Z(_06909_ ) );
BUF_X2 _14894_ ( .A(_06901_ ), .Z(_06910_ ) );
BUF_X4 _14895_ ( .A(_04380_ ), .Z(_06911_ ) );
BUF_X4 _14896_ ( .A(_06911_ ), .Z(_06912_ ) );
BUF_X4 _14897_ ( .A(_06912_ ), .Z(_06913_ ) );
BUF_X4 _14898_ ( .A(_06913_ ), .Z(_06914_ ) );
BUF_X4 _14899_ ( .A(_04386_ ), .Z(_06915_ ) );
BUF_X4 _14900_ ( .A(_06915_ ), .Z(_06916_ ) );
BUF_X4 _14901_ ( .A(_06916_ ), .Z(_06917_ ) );
XNOR2_X1 _14902_ ( .A(_06914_ ), .B(_06917_ ), .ZN(_06918_ ) );
BUF_X4 _14903_ ( .A(_04390_ ), .Z(_06919_ ) );
BUF_X4 _14904_ ( .A(_06919_ ), .Z(_06920_ ) );
BUF_X4 _14905_ ( .A(_06920_ ), .Z(_06921_ ) );
NOR2_X1 _14906_ ( .A1(_06918_ ), .A2(_06921_ ), .ZN(_06922_ ) );
INV_X1 _14907_ ( .A(_06922_ ), .ZN(_06923_ ) );
XNOR2_X1 _14908_ ( .A(_06884_ ), .B(_06804_ ), .ZN(_06924_ ) );
INV_X1 _14909_ ( .A(_06924_ ), .ZN(_06925_ ) );
BUF_X2 _14910_ ( .A(_06925_ ), .Z(_06926_ ) );
AND3_X1 _14911_ ( .A1(_06910_ ), .A2(_06923_ ), .A3(_06926_ ), .ZN(_06927_ ) );
OAI221_X1 _14912_ ( .A(_06866_ ), .B1(_06904_ ), .B2(_06908_ ), .C1(_06909_ ), .C2(_06927_ ), .ZN(_06928_ ) );
INV_X1 _14913_ ( .A(_04642_ ), .ZN(_06929_ ) );
BUF_X4 _14914_ ( .A(_04372_ ), .Z(_06930_ ) );
BUF_X4 _14915_ ( .A(_06930_ ), .Z(_06931_ ) );
BUF_X4 _14916_ ( .A(_06931_ ), .Z(_06932_ ) );
INV_X1 _14917_ ( .A(_04380_ ), .ZN(_06933_ ) );
BUF_X4 _14918_ ( .A(_06933_ ), .Z(_06934_ ) );
BUF_X4 _14919_ ( .A(_04386_ ), .Z(_06935_ ) );
BUF_X4 _14920_ ( .A(_06935_ ), .Z(_06936_ ) );
NOR2_X1 _14921_ ( .A1(_06936_ ), .A2(_02580_ ), .ZN(_06937_ ) );
BUF_X4 _14922_ ( .A(_04384_ ), .Z(_06938_ ) );
BUF_X4 _14923_ ( .A(_06938_ ), .Z(_06939_ ) );
BUF_X4 _14924_ ( .A(_04385_ ), .Z(_06940_ ) );
BUF_X4 _14925_ ( .A(_06940_ ), .Z(_06941_ ) );
AOI21_X1 _14926_ ( .A(_02557_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_06942_ ) );
OR3_X1 _14927_ ( .A1(_06934_ ), .A2(_06937_ ), .A3(_06942_ ), .ZN(_06943_ ) );
NOR2_X1 _14928_ ( .A1(_06936_ ), .A2(_02629_ ), .ZN(_06944_ ) );
BUF_X2 _14929_ ( .A(_06911_ ), .Z(_06945_ ) );
AOI21_X1 _14930_ ( .A(_02606_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_06946_ ) );
OR3_X1 _14931_ ( .A1(_06944_ ), .A2(_06945_ ), .A3(_06946_ ), .ZN(_06947_ ) );
AOI21_X1 _14932_ ( .A(_06932_ ), .B1(_06943_ ), .B2(_06947_ ), .ZN(_06948_ ) );
BUF_X4 _14933_ ( .A(_06934_ ), .Z(_06949_ ) );
BUF_X4 _14934_ ( .A(_06949_ ), .Z(_06950_ ) );
NOR2_X1 _14935_ ( .A1(_06936_ ), .A2(_02510_ ), .ZN(_06951_ ) );
AOI21_X1 _14936_ ( .A(_02533_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_06952_ ) );
OAI21_X1 _14937_ ( .A(_06950_ ), .B1(_06951_ ), .B2(_06952_ ), .ZN(_06953_ ) );
BUF_X2 _14938_ ( .A(_06912_ ), .Z(_06954_ ) );
NOR2_X1 _14939_ ( .A1(_06936_ ), .A2(_02485_ ), .ZN(_06955_ ) );
AOI21_X1 _14940_ ( .A(_03777_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_06956_ ) );
OAI21_X1 _14941_ ( .A(_06954_ ), .B1(_06955_ ), .B2(_06956_ ), .ZN(_06957_ ) );
BUF_X4 _14942_ ( .A(_06930_ ), .Z(_06958_ ) );
BUF_X4 _14943_ ( .A(_06958_ ), .Z(_06959_ ) );
AND3_X1 _14944_ ( .A1(_06953_ ), .A2(_06957_ ), .A3(_06959_ ), .ZN(_06960_ ) );
BUF_X4 _14945_ ( .A(_06804_ ), .Z(_06961_ ) );
BUF_X4 _14946_ ( .A(_06961_ ), .Z(_06962_ ) );
BUF_X4 _14947_ ( .A(_06962_ ), .Z(_06963_ ) );
OR3_X1 _14948_ ( .A1(_06948_ ), .A2(_06960_ ), .A3(_06963_ ), .ZN(_06964_ ) );
BUF_X4 _14949_ ( .A(_06905_ ), .Z(_06965_ ) );
BUF_X2 _14950_ ( .A(_06965_ ), .Z(_06966_ ) );
BUF_X2 _14951_ ( .A(_06966_ ), .Z(_06967_ ) );
BUF_X2 _14952_ ( .A(_06962_ ), .Z(_06968_ ) );
NOR2_X1 _14953_ ( .A1(_06936_ ), .A2(_02912_ ), .ZN(_06969_ ) );
INV_X1 _14954_ ( .A(_06969_ ), .ZN(_06970_ ) );
INV_X1 _14955_ ( .A(_06935_ ), .ZN(_06971_ ) );
OAI211_X1 _14956_ ( .A(_06970_ ), .B(_06949_ ), .C1(_02936_ ), .C2(_06971_ ), .ZN(_06972_ ) );
BUF_X2 _14957_ ( .A(_06931_ ), .Z(_06973_ ) );
AOI21_X1 _14958_ ( .A(_04194_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_06974_ ) );
INV_X1 _14959_ ( .A(_06974_ ), .ZN(_06975_ ) );
BUF_X2 _14960_ ( .A(_06911_ ), .Z(_06976_ ) );
OAI211_X1 _14961_ ( .A(_06975_ ), .B(_06976_ ), .C1(_02863_ ), .C2(_06916_ ), .ZN(_06977_ ) );
AND3_X1 _14962_ ( .A1(_06972_ ), .A2(_06973_ ), .A3(_06977_ ), .ZN(_06978_ ) );
NOR2_X1 _14963_ ( .A1(_06935_ ), .A2(_02729_ ), .ZN(_06979_ ) );
AOI21_X1 _14964_ ( .A(_02706_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_06980_ ) );
OAI21_X1 _14965_ ( .A(_06950_ ), .B1(_06979_ ), .B2(_06980_ ), .ZN(_06981_ ) );
NOR2_X1 _14966_ ( .A1(_06936_ ), .A2(_02960_ ), .ZN(_06982_ ) );
AOI21_X1 _14967_ ( .A(_02983_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_06983_ ) );
OAI21_X1 _14968_ ( .A(_06954_ ), .B1(_06982_ ), .B2(_06983_ ), .ZN(_06984_ ) );
AOI21_X1 _14969_ ( .A(_06973_ ), .B1(_06981_ ), .B2(_06984_ ), .ZN(_06985_ ) );
OAI21_X1 _14970_ ( .A(_06968_ ), .B1(_06978_ ), .B2(_06985_ ), .ZN(_06986_ ) );
NAND3_X1 _14971_ ( .A1(_06964_ ), .A2(_06967_ ), .A3(_06986_ ), .ZN(_06987_ ) );
BUF_X4 _14972_ ( .A(_04384_ ), .Z(_06988_ ) );
BUF_X4 _14973_ ( .A(_04385_ ), .Z(_06989_ ) );
AOI21_X1 _14974_ ( .A(_02760_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_06990_ ) );
AOI21_X1 _14975_ ( .A(_06990_ ), .B1(_06971_ ), .B2(_06796_ ), .ZN(_06991_ ) );
BUF_X2 _14976_ ( .A(_06913_ ), .Z(_06992_ ) );
NAND3_X1 _14977_ ( .A1(_06991_ ), .A2(_06920_ ), .A3(_06992_ ), .ZN(_06993_ ) );
NOR2_X1 _14978_ ( .A1(_06915_ ), .A2(_02806_ ), .ZN(_06994_ ) );
AOI21_X1 _14979_ ( .A(_02829_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_06995_ ) );
OAI21_X1 _14980_ ( .A(_06950_ ), .B1(_06994_ ), .B2(_06995_ ), .ZN(_06996_ ) );
NOR2_X1 _14981_ ( .A1(_06935_ ), .A2(_02677_ ), .ZN(_06997_ ) );
AOI21_X1 _14982_ ( .A(_02652_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_06998_ ) );
OAI21_X1 _14983_ ( .A(_06954_ ), .B1(_06997_ ), .B2(_06998_ ), .ZN(_06999_ ) );
NAND2_X1 _14984_ ( .A1(_06996_ ), .A2(_06999_ ), .ZN(_07000_ ) );
BUF_X2 _14985_ ( .A(_06919_ ), .Z(_07001_ ) );
OAI21_X1 _14986_ ( .A(_06993_ ), .B1(_07000_ ), .B2(_07001_ ), .ZN(_07002_ ) );
INV_X1 _14987_ ( .A(_06905_ ), .ZN(_07003_ ) );
BUF_X4 _14988_ ( .A(_07003_ ), .Z(_07004_ ) );
BUF_X4 _14989_ ( .A(_07004_ ), .Z(_07005_ ) );
BUF_X4 _14990_ ( .A(_06805_ ), .Z(_07006_ ) );
BUF_X2 _14991_ ( .A(_07006_ ), .Z(_07007_ ) );
BUF_X2 _14992_ ( .A(_07007_ ), .Z(_07008_ ) );
NAND3_X1 _14993_ ( .A1(_07002_ ), .A2(_07005_ ), .A3(_07008_ ), .ZN(_07009_ ) );
AOI21_X1 _14994_ ( .A(_06929_ ), .B1(_06987_ ), .B2(_07009_ ), .ZN(_07010_ ) );
BUF_X2 _14995_ ( .A(_04645_ ), .Z(_07011_ ) );
AND2_X1 _14996_ ( .A1(_04460_ ), .A2(_07011_ ), .ZN(_07012_ ) );
AND2_X2 _14997_ ( .A1(_04293_ ), .A2(\ID_EX_typ [2] ), .ZN(_07013_ ) );
NOR2_X1 _14998_ ( .A1(_07013_ ), .A2(_06865_ ), .ZN(_07014_ ) );
AND2_X1 _14999_ ( .A1(_06915_ ), .A2(_03185_ ), .ZN(_07015_ ) );
INV_X1 _15000_ ( .A(_07015_ ), .ZN(_07016_ ) );
AND3_X1 _15001_ ( .A1(_02358_ ), .A2(_04384_ ), .A3(_04385_ ), .ZN(_07017_ ) );
AOI21_X1 _15002_ ( .A(_03150_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_07018_ ) );
OR2_X1 _15003_ ( .A1(_07017_ ), .A2(_07018_ ), .ZN(_07019_ ) );
MUX2_X1 _15004_ ( .A(_07016_ ), .B(_07019_ ), .S(_06912_ ), .Z(_07020_ ) );
INV_X1 _15005_ ( .A(_07020_ ), .ZN(_07021_ ) );
BUF_X4 _15006_ ( .A(_06959_ ), .Z(_07022_ ) );
BUF_X4 _15007_ ( .A(_07022_ ), .Z(_07023_ ) );
NAND3_X1 _15008_ ( .A1(_07021_ ), .A2(_06963_ ), .A3(_07023_ ), .ZN(_07024_ ) );
NOR2_X1 _15009_ ( .A1(_06935_ ), .A2(_03047_ ), .ZN(_07025_ ) );
AOI21_X1 _15010_ ( .A(_02438_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_07026_ ) );
OAI21_X1 _15011_ ( .A(_06950_ ), .B1(_07025_ ), .B2(_07026_ ), .ZN(_07027_ ) );
NOR2_X1 _15012_ ( .A1(_06936_ ), .A2(_02411_ ), .ZN(_07028_ ) );
OAI21_X1 _15013_ ( .A(_06913_ ), .B1(_07028_ ), .B2(_06956_ ), .ZN(_07029_ ) );
NAND2_X1 _15014_ ( .A1(_07027_ ), .A2(_07029_ ), .ZN(_07030_ ) );
NAND2_X1 _15015_ ( .A1(_07030_ ), .A2(_06959_ ), .ZN(_07031_ ) );
NOR2_X1 _15016_ ( .A1(_06935_ ), .A2(_02388_ ), .ZN(_07032_ ) );
AOI21_X1 _15017_ ( .A(_03560_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_07033_ ) );
OAI21_X1 _15018_ ( .A(_06949_ ), .B1(_07032_ ), .B2(_07033_ ), .ZN(_07034_ ) );
NOR2_X1 _15019_ ( .A1(_06935_ ), .A2(_03120_ ), .ZN(_07035_ ) );
AOI21_X1 _15020_ ( .A(_03073_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07036_ ) );
OAI21_X1 _15021_ ( .A(_06976_ ), .B1(_07035_ ), .B2(_07036_ ), .ZN(_07037_ ) );
NAND2_X1 _15022_ ( .A1(_07034_ ), .A2(_07037_ ), .ZN(_07038_ ) );
BUF_X2 _15023_ ( .A(_06919_ ), .Z(_07039_ ) );
NAND2_X1 _15024_ ( .A1(_07038_ ), .A2(_07039_ ), .ZN(_07040_ ) );
BUF_X2 _15025_ ( .A(_07006_ ), .Z(_07041_ ) );
BUF_X4 _15026_ ( .A(_07041_ ), .Z(_07042_ ) );
NAND3_X1 _15027_ ( .A1(_07031_ ), .A2(_07040_ ), .A3(_07042_ ), .ZN(_07043_ ) );
AOI211_X1 _15028_ ( .A(_07005_ ), .B(_07014_ ), .C1(_07024_ ), .C2(_07043_ ), .ZN(_07044_ ) );
BUF_X4 _15029_ ( .A(_04291_ ), .Z(_07045_ ) );
NOR3_X1 _15030_ ( .A1(_04459_ ), .A2(_03778_ ), .A3(_07045_ ), .ZN(_07046_ ) );
BUF_X4 _15031_ ( .A(_04295_ ), .Z(_07047_ ) );
AOI21_X1 _15032_ ( .A(_07047_ ), .B1(_04459_ ), .B2(_03778_ ), .ZN(_07048_ ) );
OR2_X1 _15033_ ( .A1(_07046_ ), .A2(_07048_ ), .ZN(_07049_ ) );
NOR4_X1 _15034_ ( .A1(_07010_ ), .A2(_07012_ ), .A3(_07044_ ), .A4(_07049_ ), .ZN(_07050_ ) );
NAND3_X1 _15035_ ( .A1(_06864_ ), .A2(_06928_ ), .A3(_07050_ ), .ZN(_07051_ ) );
OAI21_X1 _15036_ ( .A(_06764_ ), .B1(_06763_ ), .B2(_06768_ ), .ZN(_07052_ ) );
NOR2_X1 _15037_ ( .A1(_03372_ ), .A2(\ID_EX_typ [2] ), .ZN(_07053_ ) );
OAI211_X1 _15038_ ( .A(_07053_ ), .B(_04292_ ), .C1(_04299_ ), .C2(_03250_ ), .ZN(_07054_ ) );
AND2_X1 _15039_ ( .A1(_07052_ ), .A2(_07054_ ), .ZN(_07055_ ) );
NOR2_X1 _15040_ ( .A1(_07055_ ), .A2(_06785_ ), .ZN(_07056_ ) );
INV_X2 _15041_ ( .A(_07056_ ), .ZN(_07057_ ) );
BUF_X4 _15042_ ( .A(_07057_ ), .Z(_07058_ ) );
AOI21_X1 _15043_ ( .A(_06788_ ), .B1(_07051_ ), .B2(_07058_ ), .ZN(_07059_ ) );
NAND2_X1 _15044_ ( .A1(_05347_ ), .A2(_05320_ ), .ZN(_07060_ ) );
NAND2_X1 _15045_ ( .A1(_07060_ ), .A2(_06424_ ), .ZN(_07061_ ) );
OAI21_X1 _15046_ ( .A(_06762_ ), .B1(_07059_ ), .B2(_07061_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
NAND2_X1 _15047_ ( .A1(_04753_ ), .A2(_06435_ ), .ZN(_07062_ ) );
NAND3_X1 _15048_ ( .A1(_06773_ ), .A2(_06775_ ), .A3(_04601_ ), .ZN(_07063_ ) );
NAND3_X1 _15049_ ( .A1(_06776_ ), .A2(_06782_ ), .A3(_07063_ ), .ZN(_07064_ ) );
BUF_X2 _15050_ ( .A(_06766_ ), .Z(_07065_ ) );
BUF_X4 _15051_ ( .A(_06769_ ), .Z(_07066_ ) );
AOI22_X1 _15052_ ( .A1(_04726_ ), .A2(_07065_ ), .B1(\ID_EX_imm [20] ), .B2(_07066_ ), .ZN(_07067_ ) );
AOI21_X1 _15053_ ( .A(_06787_ ), .B1(_07064_ ), .B2(_07067_ ), .ZN(_07068_ ) );
OR2_X1 _15054_ ( .A1(_07068_ ), .A2(_05224_ ), .ZN(_07069_ ) );
BUF_X4 _15055_ ( .A(_07057_ ), .Z(_07070_ ) );
INV_X1 _15056_ ( .A(_06865_ ), .ZN(_07071_ ) );
BUF_X4 _15057_ ( .A(_07071_ ), .Z(_07072_ ) );
INV_X1 _15058_ ( .A(_06901_ ), .ZN(_07073_ ) );
AOI21_X1 _15059_ ( .A(_06920_ ), .B1(_06992_ ), .B2(_06917_ ), .ZN(_07074_ ) );
NOR3_X1 _15060_ ( .A1(_07073_ ), .A2(_06924_ ), .A3(_07074_ ), .ZN(_07075_ ) );
OAI22_X1 _15061_ ( .A1(_07075_ ), .A2(_06909_ ), .B1(_06908_ ), .B2(_06904_ ), .ZN(_07076_ ) );
NOR2_X1 _15062_ ( .A1(_04386_ ), .A2(_03150_ ), .ZN(_07077_ ) );
AOI21_X1 _15063_ ( .A(_02388_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_07078_ ) );
NOR2_X1 _15064_ ( .A1(_07077_ ), .A2(_07078_ ), .ZN(_07079_ ) );
INV_X1 _15065_ ( .A(_02358_ ), .ZN(_07080_ ) );
MUX2_X1 _15066_ ( .A(_03185_ ), .B(_07080_ ), .S(_04386_ ), .Z(_07081_ ) );
MUX2_X1 _15067_ ( .A(_07079_ ), .B(_07081_ ), .S(_06933_ ), .Z(_07082_ ) );
NAND3_X1 _15068_ ( .A1(_07082_ ), .A2(_06962_ ), .A3(_07022_ ), .ZN(_07083_ ) );
BUF_X2 _15069_ ( .A(_06961_ ), .Z(_07084_ ) );
NOR2_X1 _15070_ ( .A1(_04386_ ), .A2(_03560_ ), .ZN(_07085_ ) );
AOI21_X1 _15071_ ( .A(_03120_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_07086_ ) );
OAI21_X1 _15072_ ( .A(_06933_ ), .B1(_07085_ ), .B2(_07086_ ), .ZN(_07087_ ) );
NOR2_X1 _15073_ ( .A1(_04386_ ), .A2(_03073_ ), .ZN(_07088_ ) );
AOI21_X1 _15074_ ( .A(_03047_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_07089_ ) );
OAI21_X1 _15075_ ( .A(_06911_ ), .B1(_07088_ ), .B2(_07089_ ), .ZN(_07090_ ) );
NAND3_X1 _15076_ ( .A1(_07087_ ), .A2(_07090_ ), .A3(_07039_ ), .ZN(_07091_ ) );
NOR2_X1 _15077_ ( .A1(_06915_ ), .A2(_02438_ ), .ZN(_07092_ ) );
AOI21_X1 _15078_ ( .A(_02411_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07093_ ) );
OAI21_X1 _15079_ ( .A(_06934_ ), .B1(_07092_ ), .B2(_07093_ ), .ZN(_07094_ ) );
NOR2_X1 _15080_ ( .A1(_06915_ ), .A2(_03777_ ), .ZN(_07095_ ) );
AOI21_X1 _15081_ ( .A(_02485_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07096_ ) );
OAI21_X1 _15082_ ( .A(_06945_ ), .B1(_07095_ ), .B2(_07096_ ), .ZN(_07097_ ) );
NAND3_X1 _15083_ ( .A1(_07094_ ), .A2(_07097_ ), .A3(_06931_ ), .ZN(_07098_ ) );
AND2_X1 _15084_ ( .A1(_07091_ ), .A2(_07098_ ), .ZN(_07099_ ) );
OAI21_X1 _15085_ ( .A(_07083_ ), .B1(_07084_ ), .B2(_07099_ ), .ZN(_07100_ ) );
BUF_X4 _15086_ ( .A(_06965_ ), .Z(_07101_ ) );
BUF_X2 _15087_ ( .A(_07101_ ), .Z(_07102_ ) );
NAND2_X1 _15088_ ( .A1(_07100_ ), .A2(_07102_ ), .ZN(_07103_ ) );
AOI21_X1 _15089_ ( .A(_07072_ ), .B1(_07076_ ), .B2(_07103_ ), .ZN(_07104_ ) );
NOR2_X1 _15090_ ( .A1(_06935_ ), .A2(_02829_ ), .ZN(_07105_ ) );
AOI21_X1 _15091_ ( .A(_02677_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07106_ ) );
NOR3_X1 _15092_ ( .A1(_06933_ ), .A2(_07105_ ), .A3(_07106_ ), .ZN(_07107_ ) );
NOR2_X1 _15093_ ( .A1(_06935_ ), .A2(_02760_ ), .ZN(_07108_ ) );
AOI21_X1 _15094_ ( .A(_02806_ ), .B1(_06938_ ), .B2(_06940_ ), .ZN(_07109_ ) );
NOR3_X1 _15095_ ( .A1(_07108_ ), .A2(_06911_ ), .A3(_07109_ ), .ZN(_07110_ ) );
OAI21_X1 _15096_ ( .A(_06973_ ), .B1(_07107_ ), .B2(_07110_ ), .ZN(_07111_ ) );
AND2_X1 _15097_ ( .A1(_06935_ ), .A2(_04071_ ), .ZN(_07112_ ) );
NAND3_X1 _15098_ ( .A1(_07112_ ), .A2(_07001_ ), .A3(_06992_ ), .ZN(_07113_ ) );
AND2_X1 _15099_ ( .A1(_07111_ ), .A2(_07113_ ), .ZN(_07114_ ) );
OR3_X1 _15100_ ( .A1(_07114_ ), .A2(_07101_ ), .A3(_06968_ ), .ZN(_07115_ ) );
BUF_X2 _15101_ ( .A(_06934_ ), .Z(_07116_ ) );
BUF_X4 _15102_ ( .A(_07116_ ), .Z(_07117_ ) );
NOR2_X1 _15103_ ( .A1(_06915_ ), .A2(_02557_ ), .ZN(_07118_ ) );
AOI21_X1 _15104_ ( .A(_02510_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07119_ ) );
OAI21_X1 _15105_ ( .A(_07117_ ), .B1(_07118_ ), .B2(_07119_ ), .ZN(_07120_ ) );
NOR2_X1 _15106_ ( .A1(_06915_ ), .A2(_02533_ ), .ZN(_07121_ ) );
OAI21_X1 _15107_ ( .A(_06914_ ), .B1(_07121_ ), .B2(_07096_ ), .ZN(_07122_ ) );
AND3_X1 _15108_ ( .A1(_07120_ ), .A2(_07122_ ), .A3(_06932_ ), .ZN(_07123_ ) );
AOI21_X1 _15109_ ( .A(_02629_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_07124_ ) );
INV_X1 _15110_ ( .A(_07124_ ), .ZN(_07125_ ) );
OAI211_X1 _15111_ ( .A(_07116_ ), .B(_07125_ ), .C1(_04194_ ), .C2(_06916_ ), .ZN(_07126_ ) );
AOI21_X1 _15112_ ( .A(_02580_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07127_ ) );
INV_X1 _15113_ ( .A(_07127_ ), .ZN(_07128_ ) );
OAI211_X1 _15114_ ( .A(_07128_ ), .B(_06913_ ), .C1(_02606_ ), .C2(_06916_ ), .ZN(_07129_ ) );
AOI21_X1 _15115_ ( .A(_06973_ ), .B1(_07126_ ), .B2(_07129_ ), .ZN(_07130_ ) );
OR3_X1 _15116_ ( .A1(_07123_ ), .A2(_07130_ ), .A3(_07084_ ), .ZN(_07131_ ) );
AOI21_X1 _15117_ ( .A(_02912_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_07132_ ) );
INV_X1 _15118_ ( .A(_07132_ ), .ZN(_07133_ ) );
OAI211_X1 _15119_ ( .A(_07116_ ), .B(_07133_ ), .C1(_02983_ ), .C2(_06917_ ), .ZN(_07134_ ) );
AOI21_X1 _15120_ ( .A(_02863_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_07135_ ) );
INV_X1 _15121_ ( .A(_07135_ ), .ZN(_07136_ ) );
OAI211_X1 _15122_ ( .A(_07136_ ), .B(_06913_ ), .C1(_02936_ ), .C2(_06916_ ), .ZN(_07137_ ) );
AND3_X1 _15123_ ( .A1(_07134_ ), .A2(_06959_ ), .A3(_07137_ ), .ZN(_07138_ ) );
NOR2_X1 _15124_ ( .A1(_06915_ ), .A2(_02652_ ), .ZN(_07139_ ) );
AOI21_X1 _15125_ ( .A(_02729_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07140_ ) );
OAI21_X1 _15126_ ( .A(_06933_ ), .B1(_07139_ ), .B2(_07140_ ), .ZN(_07141_ ) );
NOR2_X1 _15127_ ( .A1(_06915_ ), .A2(_02706_ ), .ZN(_07142_ ) );
AOI21_X1 _15128_ ( .A(_02960_ ), .B1(_06988_ ), .B2(_06989_ ), .ZN(_07143_ ) );
OAI21_X1 _15129_ ( .A(_06911_ ), .B1(_07142_ ), .B2(_07143_ ), .ZN(_07144_ ) );
AOI21_X1 _15130_ ( .A(_06959_ ), .B1(_07141_ ), .B2(_07144_ ), .ZN(_07145_ ) );
OAI21_X1 _15131_ ( .A(_06968_ ), .B1(_07138_ ), .B2(_07145_ ), .ZN(_07146_ ) );
NAND3_X1 _15132_ ( .A1(_07131_ ), .A2(_06967_ ), .A3(_07146_ ), .ZN(_07147_ ) );
AOI21_X1 _15133_ ( .A(_06929_ ), .B1(_07115_ ), .B2(_07147_ ), .ZN(_07148_ ) );
BUF_X2 _15134_ ( .A(_07013_ ), .Z(_07149_ ) );
AND3_X1 _15135_ ( .A1(_07100_ ), .A2(_06967_ ), .A3(_07149_ ), .ZN(_07150_ ) );
NOR3_X1 _15136_ ( .A1(_07104_ ), .A2(_07148_ ), .A3(_07150_ ), .ZN(_07151_ ) );
INV_X1 _15137_ ( .A(_06860_ ), .ZN(_07152_ ) );
BUF_X2 _15138_ ( .A(_07152_ ), .Z(_07153_ ) );
INV_X4 _15139_ ( .A(_06852_ ), .ZN(_07154_ ) );
AOI21_X1 _15140_ ( .A(_07153_ ), .B1(_07154_ ), .B2(_04465_ ), .ZN(_07155_ ) );
OAI21_X1 _15141_ ( .A(_07155_ ), .B1(_04465_ ), .B2(_07154_ ), .ZN(_07156_ ) );
AND2_X1 _15142_ ( .A1(_04465_ ), .A2(_07011_ ), .ZN(_07157_ ) );
NOR3_X1 _15143_ ( .A1(_04464_ ), .A2(_06854_ ), .A3(_07045_ ), .ZN(_07158_ ) );
BUF_X2 _15144_ ( .A(_07047_ ), .Z(_07159_ ) );
AOI21_X1 _15145_ ( .A(_07159_ ), .B1(_04464_ ), .B2(_06854_ ), .ZN(_07160_ ) );
NOR3_X1 _15146_ ( .A1(_07157_ ), .A2(_07158_ ), .A3(_07160_ ), .ZN(_07161_ ) );
NAND3_X1 _15147_ ( .A1(_07151_ ), .A2(_07156_ ), .A3(_07161_ ), .ZN(_07162_ ) );
AOI21_X1 _15148_ ( .A(_07069_ ), .B1(_07070_ ), .B2(_07162_ ), .ZN(_07163_ ) );
OAI21_X1 _15149_ ( .A(_06488_ ), .B1(_04723_ ), .B2(_02275_ ), .ZN(_07164_ ) );
OAI21_X1 _15150_ ( .A(_07062_ ), .B1(_07163_ ), .B2(_07164_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
INV_X1 _15151_ ( .A(_06467_ ), .ZN(_07165_ ) );
BUF_X4 _15152_ ( .A(_06786_ ), .Z(_07166_ ) );
AND2_X1 _15153_ ( .A1(_02510_ ), .A2(_03848_ ), .ZN(_07167_ ) );
AND2_X1 _15154_ ( .A1(_02580_ ), .A2(_03871_ ), .ZN(_07168_ ) );
AOI21_X1 _15155_ ( .A(_07168_ ), .B1(_06772_ ), .B2(_03872_ ), .ZN(_07169_ ) );
OAI21_X1 _15156_ ( .A(_04597_ ), .B1(_07169_ ), .B2(_04593_ ), .ZN(_07170_ ) );
AOI21_X1 _15157_ ( .A(_07167_ ), .B1(_07170_ ), .B2(_03849_ ), .ZN(_07171_ ) );
XNOR2_X1 _15158_ ( .A(_07171_ ), .B(_03827_ ), .ZN(_07172_ ) );
NAND2_X1 _15159_ ( .A1(_07172_ ), .A2(_06782_ ), .ZN(_07173_ ) );
AOI22_X1 _15160_ ( .A1(_04769_ ), .A2(_07065_ ), .B1(\ID_EX_imm [19] ), .B2(_07066_ ), .ZN(_07174_ ) );
AOI21_X1 _15161_ ( .A(_07166_ ), .B1(_07173_ ), .B2(_07174_ ), .ZN(_07175_ ) );
OR2_X1 _15162_ ( .A1(_07175_ ), .A2(_05224_ ), .ZN(_07176_ ) );
OR3_X1 _15163_ ( .A1(_07116_ ), .A2(_06955_ ), .A3(_06952_ ), .ZN(_07177_ ) );
OR3_X1 _15164_ ( .A1(_07028_ ), .A2(_06976_ ), .A3(_06956_ ), .ZN(_07178_ ) );
AOI21_X1 _15165_ ( .A(_07039_ ), .B1(_07177_ ), .B2(_07178_ ), .ZN(_07179_ ) );
OAI21_X1 _15166_ ( .A(_06933_ ), .B1(_07035_ ), .B2(_07036_ ), .ZN(_07180_ ) );
OAI21_X1 _15167_ ( .A(_06911_ ), .B1(_07025_ ), .B2(_07026_ ), .ZN(_07181_ ) );
AND3_X1 _15168_ ( .A1(_07180_ ), .A2(_07181_ ), .A3(_07039_ ), .ZN(_07182_ ) );
OAI21_X1 _15169_ ( .A(_07041_ ), .B1(_07179_ ), .B2(_07182_ ), .ZN(_07183_ ) );
AND2_X1 _15170_ ( .A1(_07015_ ), .A2(_06912_ ), .ZN(_07184_ ) );
INV_X1 _15171_ ( .A(_07184_ ), .ZN(_07185_ ) );
NOR3_X1 _15172_ ( .A1(_06933_ ), .A2(_07032_ ), .A3(_07033_ ), .ZN(_07186_ ) );
NOR3_X1 _15173_ ( .A1(_07017_ ), .A2(_06911_ ), .A3(_07018_ ), .ZN(_07187_ ) );
NOR2_X1 _15174_ ( .A1(_07186_ ), .A2(_07187_ ), .ZN(_07188_ ) );
MUX2_X1 _15175_ ( .A(_07185_ ), .B(_07188_ ), .S(_06958_ ), .Z(_07189_ ) );
OAI21_X1 _15176_ ( .A(_07183_ ), .B1(_07189_ ), .B2(_07041_ ), .ZN(_07190_ ) );
AND2_X1 _15177_ ( .A1(_07190_ ), .A2(_06966_ ), .ZN(_07191_ ) );
AOI21_X1 _15178_ ( .A(_07191_ ), .B1(_06904_ ), .B2(_06909_ ), .ZN(_07192_ ) );
XNOR2_X1 _15179_ ( .A(_06883_ ), .B(_06958_ ), .ZN(_07193_ ) );
NAND4_X1 _15180_ ( .A1(_06910_ ), .A2(_06926_ ), .A3(_07193_ ), .A4(_06902_ ), .ZN(_07194_ ) );
AOI21_X1 _15181_ ( .A(_07072_ ), .B1(_07192_ ), .B2(_07194_ ), .ZN(_07195_ ) );
BUF_X2 _15182_ ( .A(_06965_ ), .Z(_07196_ ) );
AND3_X1 _15183_ ( .A1(_07190_ ), .A2(_07196_ ), .A3(_07149_ ), .ZN(_07197_ ) );
BUF_X2 _15184_ ( .A(_04646_ ), .Z(_07198_ ) );
NOR3_X1 _15185_ ( .A1(_04481_ ), .A2(_04482_ ), .A3(_07198_ ), .ZN(_07199_ ) );
NOR3_X1 _15186_ ( .A1(_04480_ ), .A2(_03803_ ), .A3(_07045_ ), .ZN(_07200_ ) );
NOR2_X1 _15187_ ( .A1(_04482_ ), .A2(_07047_ ), .ZN(_07201_ ) );
OR2_X1 _15188_ ( .A1(_07200_ ), .A2(_07201_ ), .ZN(_07202_ ) );
NOR4_X1 _15189_ ( .A1(_07195_ ), .A2(_07197_ ), .A3(_07199_ ), .A4(_07202_ ), .ZN(_07203_ ) );
OAI21_X1 _15190_ ( .A(_06841_ ), .B1(_06820_ ), .B2(_06837_ ), .ZN(_07204_ ) );
AOI21_X1 _15191_ ( .A(_04477_ ), .B1(_07204_ ), .B2(_06845_ ), .ZN(_07205_ ) );
INV_X1 _15192_ ( .A(_07205_ ), .ZN(_07206_ ) );
AOI21_X1 _15193_ ( .A(_04496_ ), .B1(_07206_ ), .B2(_06848_ ), .ZN(_07207_ ) );
NOR3_X1 _15194_ ( .A1(_07205_ ), .A2(_04497_ ), .A3(_06847_ ), .ZN(_07208_ ) );
OAI21_X1 _15195_ ( .A(_06862_ ), .B1(_07207_ ), .B2(_07208_ ), .ZN(_07209_ ) );
OAI21_X1 _15196_ ( .A(_06945_ ), .B1(_06994_ ), .B2(_06995_ ), .ZN(_07210_ ) );
OAI21_X1 _15197_ ( .A(_07210_ ), .B1(_06912_ ), .B2(_06991_ ), .ZN(_07211_ ) );
INV_X1 _15198_ ( .A(_07211_ ), .ZN(_07212_ ) );
NAND3_X1 _15199_ ( .A1(_07212_ ), .A2(_07006_ ), .A3(_06932_ ), .ZN(_07213_ ) );
AOI21_X1 _15200_ ( .A(_06929_ ), .B1(_07213_ ), .B2(_07005_ ), .ZN(_07214_ ) );
OAI21_X1 _15201_ ( .A(_06934_ ), .B1(_06937_ ), .B2(_06942_ ), .ZN(_07215_ ) );
OAI21_X1 _15202_ ( .A(_06912_ ), .B1(_06951_ ), .B2(_06952_ ), .ZN(_07216_ ) );
AOI21_X1 _15203_ ( .A(_07001_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_07217_ ) );
NOR2_X1 _15204_ ( .A1(_06936_ ), .A2(_02863_ ), .ZN(_07218_ ) );
OAI21_X1 _15205_ ( .A(_06949_ ), .B1(_07218_ ), .B2(_06974_ ), .ZN(_07219_ ) );
OAI21_X1 _15206_ ( .A(_06976_ ), .B1(_06944_ ), .B2(_06946_ ), .ZN(_07220_ ) );
AOI21_X1 _15207_ ( .A(_06932_ ), .B1(_07219_ ), .B2(_07220_ ), .ZN(_07221_ ) );
NOR2_X1 _15208_ ( .A1(_07217_ ), .A2(_07221_ ), .ZN(_07222_ ) );
NOR3_X1 _15209_ ( .A1(_06933_ ), .A2(_06979_ ), .A3(_06980_ ), .ZN(_07223_ ) );
NOR3_X1 _15210_ ( .A1(_06997_ ), .A2(_06911_ ), .A3(_06998_ ), .ZN(_07224_ ) );
NOR3_X1 _15211_ ( .A1(_07223_ ), .A2(_07224_ ), .A3(_06932_ ), .ZN(_07225_ ) );
AOI21_X1 _15212_ ( .A(_02936_ ), .B1(_06939_ ), .B2(_06941_ ), .ZN(_07226_ ) );
NOR3_X1 _15213_ ( .A1(_06949_ ), .A2(_06969_ ), .A3(_07226_ ), .ZN(_07227_ ) );
NOR3_X1 _15214_ ( .A1(_06982_ ), .A2(_06912_ ), .A3(_06983_ ), .ZN(_07228_ ) );
NOR3_X1 _15215_ ( .A1(_07227_ ), .A2(_07228_ ), .A3(_06920_ ), .ZN(_07229_ ) );
NOR2_X1 _15216_ ( .A1(_07225_ ), .A2(_07229_ ), .ZN(_07230_ ) );
BUF_X4 _15217_ ( .A(_06963_ ), .Z(_07231_ ) );
MUX2_X1 _15218_ ( .A(_07222_ ), .B(_07230_ ), .S(_07231_ ), .Z(_07232_ ) );
OAI21_X1 _15219_ ( .A(_07214_ ), .B1(_07232_ ), .B2(_07005_ ), .ZN(_07233_ ) );
NAND3_X1 _15220_ ( .A1(_07203_ ), .A2(_07209_ ), .A3(_07233_ ), .ZN(_07234_ ) );
AOI21_X1 _15221_ ( .A(_07176_ ), .B1(_07070_ ), .B2(_07234_ ), .ZN(_07235_ ) );
BUF_X4 _15222_ ( .A(_06422_ ), .Z(_07236_ ) );
OAI21_X1 _15223_ ( .A(_07236_ ), .B1(_04763_ ), .B2(_02275_ ), .ZN(_07237_ ) );
OAI21_X1 _15224_ ( .A(_07165_ ), .B1(_07235_ ), .B2(_07237_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _15225_ ( .A1(_04806_ ), .A2(_04809_ ), .A3(_06559_ ), .ZN(_07238_ ) );
INV_X1 _15226_ ( .A(_06780_ ), .ZN(_07239_ ) );
BUF_X2 _15227_ ( .A(_07239_ ), .Z(_07240_ ) );
AOI21_X1 _15228_ ( .A(_07240_ ), .B1(_07170_ ), .B2(_03849_ ), .ZN(_07241_ ) );
OAI21_X1 _15229_ ( .A(_07241_ ), .B1(_03849_ ), .B2(_07170_ ), .ZN(_07242_ ) );
AOI22_X1 _15230_ ( .A1(_04813_ ), .A2(_07065_ ), .B1(\ID_EX_imm [18] ), .B2(_07066_ ), .ZN(_07243_ ) );
AOI21_X1 _15231_ ( .A(_07166_ ), .B1(_07242_ ), .B2(_07243_ ), .ZN(_07244_ ) );
OR2_X1 _15232_ ( .A1(_07244_ ), .A2(_05224_ ), .ZN(_07245_ ) );
NOR2_X1 _15233_ ( .A1(_06904_ ), .A2(_06908_ ), .ZN(_07246_ ) );
AND2_X1 _15234_ ( .A1(_06901_ ), .A2(_07193_ ), .ZN(_07247_ ) );
INV_X1 _15235_ ( .A(_07247_ ), .ZN(_07248_ ) );
AND2_X1 _15236_ ( .A1(_06971_ ), .A2(_06992_ ), .ZN(_07249_ ) );
OR3_X1 _15237_ ( .A1(_07248_ ), .A2(_07249_ ), .A3(_06924_ ), .ZN(_07250_ ) );
INV_X1 _15238_ ( .A(_06909_ ), .ZN(_07251_ ) );
AOI21_X1 _15239_ ( .A(_07246_ ), .B1(_07250_ ), .B2(_07251_ ), .ZN(_07252_ ) );
NOR3_X1 _15240_ ( .A1(_06950_ ), .A2(_07121_ ), .A3(_07119_ ), .ZN(_07253_ ) );
NOR3_X1 _15241_ ( .A1(_07095_ ), .A2(_06954_ ), .A3(_07096_ ), .ZN(_07254_ ) );
OAI21_X1 _15242_ ( .A(_06932_ ), .B1(_07253_ ), .B2(_07254_ ), .ZN(_07255_ ) );
OAI21_X1 _15243_ ( .A(_06934_ ), .B1(_07088_ ), .B2(_07089_ ), .ZN(_07256_ ) );
OAI21_X1 _15244_ ( .A(_06945_ ), .B1(_07092_ ), .B2(_07093_ ), .ZN(_07257_ ) );
NAND3_X1 _15245_ ( .A1(_07256_ ), .A2(_07257_ ), .A3(_06920_ ), .ZN(_07258_ ) );
AND3_X1 _15246_ ( .A1(_07255_ ), .A2(_07041_ ), .A3(_07258_ ), .ZN(_07259_ ) );
NOR3_X1 _15247_ ( .A1(_06934_ ), .A2(_07085_ ), .A3(_07086_ ), .ZN(_07260_ ) );
NOR3_X1 _15248_ ( .A1(_07077_ ), .A2(_06945_ ), .A3(_07078_ ), .ZN(_07261_ ) );
OR3_X1 _15249_ ( .A1(_07260_ ), .A2(_07261_ ), .A3(_06919_ ), .ZN(_07262_ ) );
AND2_X1 _15250_ ( .A1(_07081_ ), .A2(_06954_ ), .ZN(_07263_ ) );
OAI21_X1 _15251_ ( .A(_07262_ ), .B1(_06932_ ), .B2(_07263_ ), .ZN(_07264_ ) );
AOI21_X1 _15252_ ( .A(_07259_ ), .B1(_07264_ ), .B2(_06963_ ), .ZN(_07265_ ) );
AND2_X1 _15253_ ( .A1(_07265_ ), .A2(_07102_ ), .ZN(_07266_ ) );
OAI21_X1 _15254_ ( .A(_06866_ ), .B1(_07252_ ), .B2(_07266_ ), .ZN(_07267_ ) );
NAND3_X1 _15255_ ( .A1(_07204_ ), .A2(_04477_ ), .A3(_06845_ ), .ZN(_07268_ ) );
NAND3_X1 _15256_ ( .A1(_07206_ ), .A2(_06862_ ), .A3(_07268_ ), .ZN(_07269_ ) );
OAI21_X1 _15257_ ( .A(_06976_ ), .B1(_07108_ ), .B2(_07109_ ), .ZN(_07270_ ) );
OAI211_X1 _15258_ ( .A(_04378_ ), .B(_04379_ ), .C1(_06971_ ), .C2(_06796_ ), .ZN(_07271_ ) );
NAND2_X1 _15259_ ( .A1(_07270_ ), .A2(_07271_ ), .ZN(_07272_ ) );
NOR3_X1 _15260_ ( .A1(_07272_ ), .A2(_06963_ ), .A3(_06921_ ), .ZN(_07273_ ) );
OAI21_X1 _15261_ ( .A(_04642_ ), .B1(_07273_ ), .B2(_07196_ ), .ZN(_07274_ ) );
OR3_X1 _15262_ ( .A1(_06949_ ), .A2(_07118_ ), .A3(_07119_ ), .ZN(_07275_ ) );
OAI211_X1 _15263_ ( .A(_07116_ ), .B(_07128_ ), .C1(_02606_ ), .C2(_06916_ ), .ZN(_07276_ ) );
NAND3_X1 _15264_ ( .A1(_07275_ ), .A2(_07022_ ), .A3(_07276_ ), .ZN(_07277_ ) );
OAI211_X1 _15265_ ( .A(_06950_ ), .B(_07136_ ), .C1(_02936_ ), .C2(_06917_ ), .ZN(_07278_ ) );
OAI211_X1 _15266_ ( .A(_07125_ ), .B(_06913_ ), .C1(_04194_ ), .C2(_06917_ ), .ZN(_07279_ ) );
NAND3_X1 _15267_ ( .A1(_07278_ ), .A2(_06921_ ), .A3(_07279_ ), .ZN(_07280_ ) );
NAND2_X1 _15268_ ( .A1(_07277_ ), .A2(_07280_ ), .ZN(_07281_ ) );
NOR3_X1 _15269_ ( .A1(_06934_ ), .A2(_07139_ ), .A3(_07140_ ), .ZN(_07282_ ) );
NOR3_X1 _15270_ ( .A1(_07105_ ), .A2(_06945_ ), .A3(_07106_ ), .ZN(_07283_ ) );
OR3_X1 _15271_ ( .A1(_07282_ ), .A2(_07283_ ), .A3(_06930_ ), .ZN(_07284_ ) );
OAI21_X1 _15272_ ( .A(_06949_ ), .B1(_07142_ ), .B2(_07143_ ), .ZN(_07285_ ) );
NOR2_X1 _15273_ ( .A1(_06936_ ), .A2(_02983_ ), .ZN(_07286_ ) );
OAI21_X1 _15274_ ( .A(_06976_ ), .B1(_07286_ ), .B2(_07132_ ), .ZN(_07287_ ) );
NAND2_X1 _15275_ ( .A1(_07285_ ), .A2(_07287_ ), .ZN(_07288_ ) );
NAND2_X1 _15276_ ( .A1(_07288_ ), .A2(_06958_ ), .ZN(_07289_ ) );
NAND2_X1 _15277_ ( .A1(_07284_ ), .A2(_07289_ ), .ZN(_07290_ ) );
MUX2_X1 _15278_ ( .A(_07281_ ), .B(_07290_ ), .S(_06963_ ), .Z(_07291_ ) );
AOI21_X1 _15279_ ( .A(_07274_ ), .B1(_07291_ ), .B2(_07102_ ), .ZN(_07292_ ) );
AND3_X1 _15280_ ( .A1(_07265_ ), .A2(_07196_ ), .A3(_07149_ ), .ZN(_07293_ ) );
NOR3_X1 _15281_ ( .A1(_04475_ ), .A2(_06472_ ), .A3(_07045_ ), .ZN(_07294_ ) );
NAND3_X1 _15282_ ( .A1(_06472_ ), .A2(_04474_ ), .A3(_04473_ ), .ZN(_07295_ ) );
BUF_X4 _15283_ ( .A(_04294_ ), .Z(_07296_ ) );
NAND2_X1 _15284_ ( .A1(_07295_ ), .A2(_07296_ ), .ZN(_07297_ ) );
OAI21_X1 _15285_ ( .A(_07297_ ), .B1(_04477_ ), .B2(_07198_ ), .ZN(_07298_ ) );
NOR4_X1 _15286_ ( .A1(_07292_ ), .A2(_07293_ ), .A3(_07294_ ), .A4(_07298_ ), .ZN(_07299_ ) );
NAND3_X1 _15287_ ( .A1(_07267_ ), .A2(_07269_ ), .A3(_07299_ ), .ZN(_07300_ ) );
AOI21_X1 _15288_ ( .A(_07245_ ), .B1(_07070_ ), .B2(_07300_ ), .ZN(_07301_ ) );
NAND2_X1 _15289_ ( .A1(_04816_ ), .A2(_05320_ ), .ZN(_07302_ ) );
NAND2_X1 _15290_ ( .A1(_07302_ ), .A2(_06424_ ), .ZN(_07303_ ) );
OAI21_X1 _15291_ ( .A(_07238_ ), .B1(_07301_ ), .B2(_07303_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
NAND2_X1 _15292_ ( .A1(_06484_ ), .A2(_06435_ ), .ZN(_07304_ ) );
INV_X1 _15293_ ( .A(_06766_ ), .ZN(_07305_ ) );
OAI22_X1 _15294_ ( .A1(_04831_ ), .A2(_07305_ ), .B1(_02558_ ), .B2(_06770_ ), .ZN(_07306_ ) );
XNOR2_X1 _15295_ ( .A(_07169_ ), .B(_03897_ ), .ZN(_07307_ ) );
AOI21_X1 _15296_ ( .A(_07306_ ), .B1(_07307_ ), .B2(_06782_ ), .ZN(_07308_ ) );
OAI21_X1 _15297_ ( .A(_04661_ ), .B1(_07308_ ), .B2(_06787_ ), .ZN(_07309_ ) );
AND3_X1 _15298_ ( .A1(_06910_ ), .A2(_06925_ ), .A3(_07193_ ), .ZN(_07310_ ) );
NAND2_X1 _15299_ ( .A1(_07310_ ), .A2(_06918_ ), .ZN(_07311_ ) );
INV_X1 _15300_ ( .A(_06903_ ), .ZN(_07312_ ) );
INV_X1 _15301_ ( .A(_06908_ ), .ZN(_07313_ ) );
AOI22_X1 _15302_ ( .A1(_07311_ ), .A2(_07251_ ), .B1(_07312_ ), .B2(_07313_ ), .ZN(_07314_ ) );
OR3_X1 _15303_ ( .A1(_07116_ ), .A2(_06951_ ), .A3(_06942_ ), .ZN(_07315_ ) );
OR3_X1 _15304_ ( .A1(_06955_ ), .A2(_06913_ ), .A3(_06952_ ), .ZN(_07316_ ) );
NAND3_X1 _15305_ ( .A1(_07315_ ), .A2(_07316_ ), .A3(_06959_ ), .ZN(_07317_ ) );
NAND2_X1 _15306_ ( .A1(_07030_ ), .A2(_06920_ ), .ZN(_07318_ ) );
AND2_X1 _15307_ ( .A1(_07317_ ), .A2(_07318_ ), .ZN(_07319_ ) );
MUX2_X1 _15308_ ( .A(_07038_ ), .B(_07020_ ), .S(_07039_ ), .Z(_07320_ ) );
INV_X1 _15309_ ( .A(_07320_ ), .ZN(_07321_ ) );
MUX2_X1 _15310_ ( .A(_07319_ ), .B(_07321_ ), .S(_07084_ ), .Z(_07322_ ) );
AND2_X1 _15311_ ( .A1(_07322_ ), .A2(_07102_ ), .ZN(_07323_ ) );
OAI21_X1 _15312_ ( .A(_06866_ ), .B1(_07314_ ), .B2(_07323_ ), .ZN(_07324_ ) );
NOR2_X1 _15313_ ( .A1(_06838_ ), .A2(_06840_ ), .ZN(_07325_ ) );
OR3_X1 _15314_ ( .A1(_07325_ ), .A2(_04472_ ), .A3(_06844_ ), .ZN(_07326_ ) );
OAI21_X1 _15315_ ( .A(_04472_ ), .B1(_07325_ ), .B2(_06844_ ), .ZN(_07327_ ) );
NAND3_X1 _15316_ ( .A1(_07326_ ), .A2(_06862_ ), .A3(_07327_ ), .ZN(_07328_ ) );
AND3_X1 _15317_ ( .A1(_07322_ ), .A2(_06967_ ), .A3(_07149_ ), .ZN(_07329_ ) );
AND3_X1 _15318_ ( .A1(_06991_ ), .A2(_06973_ ), .A3(_06992_ ), .ZN(_07330_ ) );
AND2_X1 _15319_ ( .A1(_07330_ ), .A2(_07007_ ), .ZN(_07331_ ) );
OAI21_X1 _15320_ ( .A(_04642_ ), .B1(_07331_ ), .B2(_07101_ ), .ZN(_07332_ ) );
AOI21_X1 _15321_ ( .A(_06919_ ), .B1(_06943_ ), .B2(_06947_ ), .ZN(_07333_ ) );
AOI21_X1 _15322_ ( .A(_06958_ ), .B1(_06972_ ), .B2(_06977_ ), .ZN(_07334_ ) );
OR2_X1 _15323_ ( .A1(_07333_ ), .A2(_07334_ ), .ZN(_07335_ ) );
AOI21_X1 _15324_ ( .A(_07004_ ), .B1(_07335_ ), .B2(_07008_ ), .ZN(_07336_ ) );
NAND2_X1 _15325_ ( .A1(_06981_ ), .A2(_06984_ ), .ZN(_07337_ ) );
NAND2_X1 _15326_ ( .A1(_07337_ ), .A2(_06959_ ), .ZN(_07338_ ) );
NAND2_X1 _15327_ ( .A1(_07000_ ), .A2(_06920_ ), .ZN(_07339_ ) );
NAND3_X1 _15328_ ( .A1(_07338_ ), .A2(_07339_ ), .A3(_07231_ ), .ZN(_07340_ ) );
AOI21_X1 _15329_ ( .A(_07332_ ), .B1(_07336_ ), .B2(_07340_ ), .ZN(_07341_ ) );
NOR3_X1 _15330_ ( .A1(_04490_ ), .A2(_04491_ ), .A3(_07198_ ), .ZN(_07342_ ) );
OR3_X1 _15331_ ( .A1(_04471_ ), .A2(_03873_ ), .A3(_04291_ ), .ZN(_07343_ ) );
OAI21_X1 _15332_ ( .A(_07343_ ), .B1(_04490_ ), .B2(_07159_ ), .ZN(_07344_ ) );
NOR4_X1 _15333_ ( .A1(_07329_ ), .A2(_07341_ ), .A3(_07342_ ), .A4(_07344_ ), .ZN(_07345_ ) );
NAND3_X1 _15334_ ( .A1(_07324_ ), .A2(_07328_ ), .A3(_07345_ ), .ZN(_07346_ ) );
AOI21_X1 _15335_ ( .A(_07309_ ), .B1(_07070_ ), .B2(_07346_ ), .ZN(_07347_ ) );
OAI21_X1 _15336_ ( .A(_07236_ ), .B1(_04825_ ), .B2(_02275_ ), .ZN(_07348_ ) );
OAI21_X1 _15337_ ( .A(_07304_ ), .B1(_07347_ ), .B2(_07348_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
CLKBUF_X2 _15338_ ( .A(_06422_ ), .Z(_07349_ ) );
OR2_X1 _15339_ ( .A1(_06495_ ), .A2(_07349_ ), .ZN(_07350_ ) );
AOI21_X1 _15340_ ( .A(_07240_ ), .B1(_06772_ ), .B2(_03872_ ), .ZN(_07351_ ) );
OAI21_X1 _15341_ ( .A(_07351_ ), .B1(_03872_ ), .B2(_06772_ ), .ZN(_07352_ ) );
NAND2_X1 _15342_ ( .A1(_04853_ ), .A2(_07065_ ), .ZN(_07353_ ) );
NAND3_X1 _15343_ ( .A1(_06768_ ), .A2(\ID_EX_imm [16] ), .A3(_06764_ ), .ZN(_07354_ ) );
AND3_X1 _15344_ ( .A1(_07352_ ), .A2(_07353_ ), .A3(_07354_ ), .ZN(_07355_ ) );
OAI21_X1 _15345_ ( .A(_04661_ ), .B1(_07355_ ), .B2(_06787_ ), .ZN(_07356_ ) );
OAI211_X1 _15346_ ( .A(_06904_ ), .B(_06866_ ), .C1(_07005_ ), .C2(_06885_ ), .ZN(_07357_ ) );
NAND3_X1 _15347_ ( .A1(_07094_ ), .A2(_07097_ ), .A3(_06919_ ), .ZN(_07358_ ) );
OAI21_X1 _15348_ ( .A(_06934_ ), .B1(_07121_ ), .B2(_07119_ ), .ZN(_07359_ ) );
OAI21_X1 _15349_ ( .A(_06945_ ), .B1(_07118_ ), .B2(_07127_ ), .ZN(_07360_ ) );
NAND3_X1 _15350_ ( .A1(_07359_ ), .A2(_07360_ ), .A3(_06930_ ), .ZN(_07361_ ) );
AND3_X1 _15351_ ( .A1(_07358_ ), .A2(_07361_ ), .A3(_06805_ ), .ZN(_07362_ ) );
AND3_X1 _15352_ ( .A1(_07087_ ), .A2(_07090_ ), .A3(_04372_ ), .ZN(_07363_ ) );
AOI21_X1 _15353_ ( .A(_07363_ ), .B1(_07082_ ), .B2(_06919_ ), .ZN(_07364_ ) );
AOI21_X1 _15354_ ( .A(_07362_ ), .B1(_07364_ ), .B2(_06961_ ), .ZN(_07365_ ) );
NAND2_X1 _15355_ ( .A1(_07365_ ), .A2(_06967_ ), .ZN(_07366_ ) );
AOI21_X1 _15356_ ( .A(_07014_ ), .B1(_07357_ ), .B2(_07366_ ), .ZN(_07367_ ) );
OAI21_X1 _15357_ ( .A(_06861_ ), .B1(_06838_ ), .B2(_06840_ ), .ZN(_07368_ ) );
AOI21_X1 _15358_ ( .A(_07368_ ), .B1(_06840_ ), .B2(_06838_ ), .ZN(_07369_ ) );
AND3_X1 _15359_ ( .A1(_07112_ ), .A2(_04372_ ), .A3(_06911_ ), .ZN(_07370_ ) );
AND2_X1 _15360_ ( .A1(_07006_ ), .A2(_07370_ ), .ZN(_07371_ ) );
OAI21_X1 _15361_ ( .A(_04642_ ), .B1(_07371_ ), .B2(_06965_ ), .ZN(_07372_ ) );
AOI21_X1 _15362_ ( .A(_06931_ ), .B1(_07134_ ), .B2(_07137_ ), .ZN(_07373_ ) );
AOI21_X1 _15363_ ( .A(_07039_ ), .B1(_07126_ ), .B2(_07129_ ), .ZN(_07374_ ) );
NOR2_X1 _15364_ ( .A1(_07373_ ), .A2(_07374_ ), .ZN(_07375_ ) );
NOR3_X1 _15365_ ( .A1(_07107_ ), .A2(_07110_ ), .A3(_04372_ ), .ZN(_07376_ ) );
AOI21_X1 _15366_ ( .A(_04390_ ), .B1(_07141_ ), .B2(_07144_ ), .ZN(_07377_ ) );
OR2_X1 _15367_ ( .A1(_07376_ ), .A2(_07377_ ), .ZN(_07378_ ) );
BUF_X2 _15368_ ( .A(_06961_ ), .Z(_07379_ ) );
MUX2_X1 _15369_ ( .A(_07375_ ), .B(_07378_ ), .S(_07379_ ), .Z(_07380_ ) );
AOI21_X1 _15370_ ( .A(_07372_ ), .B1(_07380_ ), .B2(_06966_ ), .ZN(_07381_ ) );
AND2_X1 _15371_ ( .A1(_04487_ ), .A2(_04645_ ), .ZN(_07382_ ) );
AOI21_X1 _15372_ ( .A(_07047_ ), .B1(_04486_ ), .B2(_06843_ ), .ZN(_07383_ ) );
NOR3_X1 _15373_ ( .A1(_04486_ ), .A2(_06843_ ), .A3(_04291_ ), .ZN(_07384_ ) );
OR4_X1 _15374_ ( .A1(_07381_ ), .A2(_07382_ ), .A3(_07383_ ), .A4(_07384_ ), .ZN(_07385_ ) );
OR3_X1 _15375_ ( .A1(_07367_ ), .A2(_07369_ ), .A3(_07385_ ), .ZN(_07386_ ) );
AOI21_X1 _15376_ ( .A(_07356_ ), .B1(_07070_ ), .B2(_07386_ ), .ZN(_07387_ ) );
OAI21_X1 _15377_ ( .A(_07236_ ), .B1(_04851_ ), .B2(_04720_ ), .ZN(_07388_ ) );
OAI21_X1 _15378_ ( .A(_07350_ ), .B1(_07387_ ), .B2(_07388_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OR2_X1 _15379_ ( .A1(_04896_ ), .A2(_07349_ ), .ZN(_07389_ ) );
INV_X1 _15380_ ( .A(_04216_ ), .ZN(_07390_ ) );
INV_X1 _15381_ ( .A(_04238_ ), .ZN(_07391_ ) );
NAND2_X1 _15382_ ( .A1(_04571_ ), .A2(_04192_ ), .ZN(_07392_ ) );
AOI211_X1 _15383_ ( .A(_07390_ ), .B(_07391_ ), .C1(_07392_ ), .C2(_04585_ ), .ZN(_07393_ ) );
OAI21_X1 _15384_ ( .A(_04283_ ), .B1(_07393_ ), .B2(_04577_ ), .ZN(_07394_ ) );
NAND2_X1 _15385_ ( .A1(_02629_ ), .A2(_04282_ ), .ZN(_07395_ ) );
AND2_X1 _15386_ ( .A1(_07394_ ), .A2(_07395_ ), .ZN(_07396_ ) );
XNOR2_X1 _15387_ ( .A(_07396_ ), .B(_04261_ ), .ZN(_07397_ ) );
NAND2_X1 _15388_ ( .A1(_07397_ ), .A2(_06782_ ), .ZN(_07398_ ) );
AOI22_X1 _15389_ ( .A1(_04881_ ), .A2(_07065_ ), .B1(\ID_EX_imm [15] ), .B2(_07066_ ), .ZN(_07399_ ) );
AOI21_X1 _15390_ ( .A(_07166_ ), .B1(_07398_ ), .B2(_07399_ ), .ZN(_07400_ ) );
OR2_X1 _15391_ ( .A1(_07400_ ), .A2(_05224_ ), .ZN(_07401_ ) );
AND2_X1 _15392_ ( .A1(_06811_ ), .A2(_06819_ ), .ZN(_07402_ ) );
OR2_X1 _15393_ ( .A1(_07402_ ), .A2(_06794_ ), .ZN(_07403_ ) );
AND2_X1 _15394_ ( .A1(_06824_ ), .A2(_06826_ ), .ZN(_07404_ ) );
AND2_X1 _15395_ ( .A1(_07403_ ), .A2(_07404_ ), .ZN(_07405_ ) );
INV_X1 _15396_ ( .A(_07405_ ), .ZN(_07406_ ) );
NAND2_X1 _15397_ ( .A1(_07406_ ), .A2(_06789_ ), .ZN(_07407_ ) );
AOI21_X1 _15398_ ( .A(_06834_ ), .B1(_07407_ ), .B2(_06833_ ), .ZN(_07408_ ) );
NOR2_X1 _15399_ ( .A1(_04325_ ), .A2(_04442_ ), .ZN(_07409_ ) );
OR3_X1 _15400_ ( .A1(_07408_ ), .A2(_04333_ ), .A3(_07409_ ), .ZN(_07410_ ) );
OAI21_X1 _15401_ ( .A(_04333_ ), .B1(_07408_ ), .B2(_07409_ ), .ZN(_07411_ ) );
NAND3_X1 _15402_ ( .A1(_07410_ ), .A2(_06862_ ), .A3(_07411_ ), .ZN(_07412_ ) );
NAND3_X1 _15403_ ( .A1(_06904_ ), .A2(_06909_ ), .A3(_06865_ ), .ZN(_07413_ ) );
NOR3_X1 _15404_ ( .A1(_07186_ ), .A2(_07187_ ), .A3(_04372_ ), .ZN(_07414_ ) );
AOI21_X1 _15405_ ( .A(_04390_ ), .B1(_07180_ ), .B2(_07181_ ), .ZN(_07415_ ) );
OAI21_X1 _15406_ ( .A(_06968_ ), .B1(_07414_ ), .B2(_07415_ ), .ZN(_07416_ ) );
AOI21_X1 _15407_ ( .A(_07022_ ), .B1(_07177_ ), .B2(_07178_ ), .ZN(_07417_ ) );
OR3_X1 _15408_ ( .A1(_06950_ ), .A2(_06937_ ), .A3(_06946_ ), .ZN(_07418_ ) );
OR3_X1 _15409_ ( .A1(_06951_ ), .A2(_06954_ ), .A3(_06942_ ), .ZN(_07419_ ) );
AOI21_X1 _15410_ ( .A(_06921_ ), .B1(_07418_ ), .B2(_07419_ ), .ZN(_07420_ ) );
OR2_X1 _15411_ ( .A1(_07417_ ), .A2(_07420_ ), .ZN(_07421_ ) );
OAI211_X1 _15412_ ( .A(_07196_ ), .B(_07416_ ), .C1(_07421_ ), .C2(_07231_ ), .ZN(_07422_ ) );
NAND4_X1 _15413_ ( .A1(_07008_ ), .A2(_07184_ ), .A3(_07005_ ), .A4(_07023_ ), .ZN(_07423_ ) );
AOI21_X1 _15414_ ( .A(_07014_ ), .B1(_07422_ ), .B2(_07423_ ), .ZN(_07424_ ) );
OR3_X1 _15415_ ( .A1(_07223_ ), .A2(_07224_ ), .A3(_04390_ ), .ZN(_07425_ ) );
OAI21_X1 _15416_ ( .A(_07425_ ), .B1(_07212_ ), .B2(_06958_ ), .ZN(_07426_ ) );
NAND2_X1 _15417_ ( .A1(_07426_ ), .A2(_06961_ ), .ZN(_07427_ ) );
OAI21_X1 _15418_ ( .A(_06919_ ), .B1(_07227_ ), .B2(_07228_ ), .ZN(_07428_ ) );
NAND3_X1 _15419_ ( .A1(_07219_ ), .A2(_07220_ ), .A3(_06930_ ), .ZN(_07429_ ) );
NAND3_X1 _15420_ ( .A1(_07428_ ), .A2(_07006_ ), .A3(_07429_ ), .ZN(_07430_ ) );
AND2_X2 _15421_ ( .A1(_06905_ ), .A2(_04642_ ), .ZN(_07431_ ) );
BUF_X2 _15422_ ( .A(_07431_ ), .Z(_07432_ ) );
AND3_X1 _15423_ ( .A1(_07427_ ), .A2(_07430_ ), .A3(_07432_ ), .ZN(_07433_ ) );
NOR3_X1 _15424_ ( .A1(_04331_ ), .A2(_04332_ ), .A3(_07198_ ), .ZN(_07434_ ) );
NAND3_X1 _15425_ ( .A1(_04438_ ), .A2(_02606_ ), .A3(_06857_ ), .ZN(_07435_ ) );
OAI21_X1 _15426_ ( .A(_07435_ ), .B1(_04332_ ), .B2(_07159_ ), .ZN(_07436_ ) );
NOR4_X1 _15427_ ( .A1(_07424_ ), .A2(_07433_ ), .A3(_07434_ ), .A4(_07436_ ), .ZN(_07437_ ) );
NAND3_X1 _15428_ ( .A1(_07412_ ), .A2(_07413_ ), .A3(_07437_ ), .ZN(_07438_ ) );
AOI21_X1 _15429_ ( .A(_07401_ ), .B1(_07070_ ), .B2(_07438_ ), .ZN(_07439_ ) );
NAND2_X1 _15430_ ( .A1(_04885_ ), .A2(_05320_ ), .ZN(_07440_ ) );
BUF_X4 _15431_ ( .A(_06423_ ), .Z(_07441_ ) );
NAND2_X1 _15432_ ( .A1(_07440_ ), .A2(_07441_ ), .ZN(_07442_ ) );
OAI21_X1 _15433_ ( .A(_07389_ ), .B1(_07439_ ), .B2(_07442_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
OR2_X1 _15434_ ( .A1(_04916_ ), .A2(_07349_ ), .ZN(_07443_ ) );
OR3_X1 _15435_ ( .A1(_07393_ ), .A2(_04283_ ), .A3(_04577_ ), .ZN(_07444_ ) );
NAND3_X1 _15436_ ( .A1(_07444_ ), .A2(_06782_ ), .A3(_07394_ ), .ZN(_07445_ ) );
BUF_X4 _15437_ ( .A(_06766_ ), .Z(_07446_ ) );
AOI22_X1 _15438_ ( .A1(_04901_ ), .A2(_07446_ ), .B1(\ID_EX_imm [14] ), .B2(_07066_ ), .ZN(_07447_ ) );
AOI21_X1 _15439_ ( .A(_07166_ ), .B1(_07445_ ), .B2(_07447_ ), .ZN(_07448_ ) );
OR2_X1 _15440_ ( .A1(_07448_ ), .A2(_05224_ ), .ZN(_07449_ ) );
AND3_X1 _15441_ ( .A1(_07407_ ), .A2(_06834_ ), .A3(_06833_ ), .ZN(_07450_ ) );
OR3_X1 _15442_ ( .A1(_07450_ ), .A2(_07408_ ), .A3(_07153_ ), .ZN(_07451_ ) );
AND2_X2 _15443_ ( .A1(_06902_ ), .A2(_06906_ ), .ZN(_07452_ ) );
AND2_X1 _15444_ ( .A1(_06901_ ), .A2(_06925_ ), .ZN(_07453_ ) );
NAND3_X1 _15445_ ( .A1(_06913_ ), .A2(_06971_ ), .A3(_06930_ ), .ZN(_07454_ ) );
AND3_X1 _15446_ ( .A1(_06888_ ), .A2(_06900_ ), .A3(_07454_ ), .ZN(_07455_ ) );
OAI211_X1 _15447_ ( .A(_06866_ ), .B(_07452_ ), .C1(_07453_ ), .C2(_07455_ ), .ZN(_07456_ ) );
NOR3_X1 _15448_ ( .A1(_07260_ ), .A2(_07261_ ), .A3(_06930_ ), .ZN(_07457_ ) );
AOI21_X1 _15449_ ( .A(_04390_ ), .B1(_07256_ ), .B2(_07257_ ), .ZN(_07458_ ) );
OR3_X1 _15450_ ( .A1(_07457_ ), .A2(_07041_ ), .A3(_07458_ ), .ZN(_07459_ ) );
OAI21_X1 _15451_ ( .A(_06920_ ), .B1(_07253_ ), .B2(_07254_ ), .ZN(_07460_ ) );
NOR2_X1 _15452_ ( .A1(_06916_ ), .A2(_02606_ ), .ZN(_07461_ ) );
NOR3_X1 _15453_ ( .A1(_06950_ ), .A2(_07461_ ), .A3(_07124_ ), .ZN(_07462_ ) );
NOR3_X1 _15454_ ( .A1(_07118_ ), .A2(_06954_ ), .A3(_07127_ ), .ZN(_07463_ ) );
OAI21_X1 _15455_ ( .A(_06959_ ), .B1(_07462_ ), .B2(_07463_ ), .ZN(_07464_ ) );
AND2_X1 _15456_ ( .A1(_07460_ ), .A2(_07464_ ), .ZN(_07465_ ) );
OAI211_X1 _15457_ ( .A(_07459_ ), .B(_07101_ ), .C1(_06968_ ), .C2(_07465_ ), .ZN(_07466_ ) );
INV_X1 _15458_ ( .A(_07014_ ), .ZN(_07467_ ) );
AND3_X1 _15459_ ( .A1(_07081_ ), .A2(_06931_ ), .A3(_06914_ ), .ZN(_07468_ ) );
AND2_X1 _15460_ ( .A1(_07468_ ), .A2(_07041_ ), .ZN(_07469_ ) );
OAI211_X1 _15461_ ( .A(_07466_ ), .B(_07467_ ), .C1(_06967_ ), .C2(_07469_ ), .ZN(_07470_ ) );
NOR2_X1 _15462_ ( .A1(_07282_ ), .A2(_07283_ ), .ZN(_07471_ ) );
MUX2_X1 _15463_ ( .A(_07272_ ), .B(_07471_ ), .S(_06958_ ), .Z(_07472_ ) );
NOR2_X1 _15464_ ( .A1(_07472_ ), .A2(_07041_ ), .ZN(_07473_ ) );
AND3_X1 _15465_ ( .A1(_07278_ ), .A2(_06931_ ), .A3(_07279_ ), .ZN(_07474_ ) );
AOI21_X1 _15466_ ( .A(_06931_ ), .B1(_07285_ ), .B2(_07287_ ), .ZN(_07475_ ) );
NOR3_X1 _15467_ ( .A1(_07474_ ), .A2(_07379_ ), .A3(_07475_ ), .ZN(_07476_ ) );
OAI21_X1 _15468_ ( .A(_07432_ ), .B1(_07473_ ), .B2(_07476_ ), .ZN(_07477_ ) );
BUF_X4 _15469_ ( .A(_06857_ ), .Z(_07478_ ) );
NAND3_X1 _15470_ ( .A1(_04443_ ), .A2(_02629_ ), .A3(_07478_ ), .ZN(_07479_ ) );
AOI21_X1 _15471_ ( .A(_07047_ ), .B1(_04325_ ), .B2(_04442_ ), .ZN(_07480_ ) );
AOI21_X1 _15472_ ( .A(_07480_ ), .B1(_04326_ ), .B2(_04645_ ), .ZN(_07481_ ) );
AND4_X1 _15473_ ( .A1(_07470_ ), .A2(_07477_ ), .A3(_07479_ ), .A4(_07481_ ), .ZN(_07482_ ) );
NAND3_X1 _15474_ ( .A1(_07451_ ), .A2(_07456_ ), .A3(_07482_ ), .ZN(_07483_ ) );
AOI21_X1 _15475_ ( .A(_07449_ ), .B1(_07070_ ), .B2(_07483_ ), .ZN(_07484_ ) );
NAND2_X1 _15476_ ( .A1(_04905_ ), .A2(_05320_ ), .ZN(_07485_ ) );
NAND2_X1 _15477_ ( .A1(_07485_ ), .A2(_07441_ ), .ZN(_07486_ ) );
OAI21_X1 _15478_ ( .A(_07443_ ), .B1(_07484_ ), .B2(_07486_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
INV_X1 _15479_ ( .A(_06514_ ), .ZN(_07487_ ) );
AND2_X1 _15480_ ( .A1(_07392_ ), .A2(_04585_ ), .ZN(_07488_ ) );
OR2_X1 _15481_ ( .A1(_07488_ ), .A2(_07391_ ), .ZN(_07489_ ) );
INV_X1 _15482_ ( .A(_04574_ ), .ZN(_07490_ ) );
AND3_X1 _15483_ ( .A1(_07489_ ), .A2(_07390_ ), .A3(_07490_ ), .ZN(_07491_ ) );
AOI21_X1 _15484_ ( .A(_07390_ ), .B1(_07489_ ), .B2(_07490_ ), .ZN(_07492_ ) );
NOR3_X1 _15485_ ( .A1(_07491_ ), .A2(_07492_ ), .A3(_07240_ ), .ZN(_07493_ ) );
AND2_X1 _15486_ ( .A1(_04921_ ), .A2(_07065_ ), .ZN(_07494_ ) );
AND3_X1 _15487_ ( .A1(_06768_ ), .A2(\ID_EX_imm [13] ), .A3(_06764_ ), .ZN(_07495_ ) );
NOR3_X1 _15488_ ( .A1(_07493_ ), .A2(_07494_ ), .A3(_07495_ ), .ZN(_07496_ ) );
OAI21_X1 _15489_ ( .A(_04661_ ), .B1(_07496_ ), .B2(_06787_ ), .ZN(_07497_ ) );
NAND4_X1 _15490_ ( .A1(_07021_ ), .A2(_07004_ ), .A3(_07042_ ), .A4(_07023_ ), .ZN(_07498_ ) );
AND3_X1 _15491_ ( .A1(_07031_ ), .A2(_07040_ ), .A3(_07379_ ), .ZN(_07499_ ) );
NAND3_X1 _15492_ ( .A1(_07315_ ), .A2(_07316_ ), .A3(_06920_ ), .ZN(_07500_ ) );
OR3_X1 _15493_ ( .A1(_06937_ ), .A2(_06913_ ), .A3(_06946_ ), .ZN(_07501_ ) );
OAI211_X1 _15494_ ( .A(_06975_ ), .B(_06954_ ), .C1(_02629_ ), .C2(_06917_ ), .ZN(_07502_ ) );
NAND3_X1 _15495_ ( .A1(_07501_ ), .A2(_06959_ ), .A3(_07502_ ), .ZN(_07503_ ) );
AND2_X1 _15496_ ( .A1(_07500_ ), .A2(_07503_ ), .ZN(_07504_ ) );
AOI21_X1 _15497_ ( .A(_07499_ ), .B1(_07504_ ), .B2(_07042_ ), .ZN(_07505_ ) );
AND2_X1 _15498_ ( .A1(_06924_ ), .A2(_06922_ ), .ZN(_07506_ ) );
OAI221_X1 _15499_ ( .A(_07498_ ), .B1(_07004_ ), .B2(_07505_ ), .C1(_07413_ ), .C2(_07506_ ), .ZN(_07507_ ) );
AND2_X1 _15500_ ( .A1(_07507_ ), .A2(_07467_ ), .ZN(_07508_ ) );
INV_X1 _15501_ ( .A(_04343_ ), .ZN(_07509_ ) );
AOI21_X1 _15502_ ( .A(_07509_ ), .B1(_07403_ ), .B2(_07404_ ), .ZN(_07510_ ) );
OR4_X1 _15503_ ( .A1(_06829_ ), .A2(_07510_ ), .A3(_06830_ ), .A4(_06832_ ), .ZN(_07511_ ) );
OAI22_X1 _15504_ ( .A1(_07510_ ), .A2(_06832_ ), .B1(_06829_ ), .B2(_06830_ ), .ZN(_07512_ ) );
AOI21_X1 _15505_ ( .A(_07153_ ), .B1(_07511_ ), .B2(_07512_ ), .ZN(_07513_ ) );
NAND3_X1 _15506_ ( .A1(_06877_ ), .A2(_04194_ ), .A3(_07478_ ), .ZN(_07514_ ) );
AOI22_X1 _15507_ ( .A1(_04338_ ), .A2(_04645_ ), .B1(_06831_ ), .B2(_07296_ ), .ZN(_07515_ ) );
NOR3_X1 _15508_ ( .A1(_06978_ ), .A2(_07084_ ), .A3(_06985_ ), .ZN(_07516_ ) );
AND2_X1 _15509_ ( .A1(_07002_ ), .A2(_07084_ ), .ZN(_07517_ ) );
NOR2_X1 _15510_ ( .A1(_07516_ ), .A2(_07517_ ), .ZN(_07518_ ) );
INV_X1 _15511_ ( .A(_07431_ ), .ZN(_07519_ ) );
OAI211_X1 _15512_ ( .A(_07514_ ), .B(_07515_ ), .C1(_07518_ ), .C2(_07519_ ), .ZN(_07520_ ) );
OR3_X1 _15513_ ( .A1(_07508_ ), .A2(_07513_ ), .A3(_07520_ ), .ZN(_07521_ ) );
AOI21_X1 _15514_ ( .A(_07497_ ), .B1(_07070_ ), .B2(_07521_ ), .ZN(_07522_ ) );
NAND2_X1 _15515_ ( .A1(_04924_ ), .A2(_05320_ ), .ZN(_07523_ ) );
NAND2_X1 _15516_ ( .A1(_07523_ ), .A2(_07441_ ), .ZN(_07524_ ) );
OAI21_X1 _15517_ ( .A(_07487_ ), .B1(_07522_ ), .B2(_07524_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
NAND2_X1 _15518_ ( .A1(_04952_ ), .A2(_06435_ ), .ZN(_07525_ ) );
NAND3_X1 _15519_ ( .A1(_07392_ ), .A2(_07391_ ), .A3(_04585_ ), .ZN(_07526_ ) );
NAND3_X1 _15520_ ( .A1(_07489_ ), .A2(_06781_ ), .A3(_07526_ ), .ZN(_07527_ ) );
AOI22_X1 _15521_ ( .A1(_04940_ ), .A2(_07446_ ), .B1(\ID_EX_imm [12] ), .B2(_07066_ ), .ZN(_07528_ ) );
AOI21_X1 _15522_ ( .A(_07166_ ), .B1(_07527_ ), .B2(_07528_ ), .ZN(_07529_ ) );
OR2_X1 _15523_ ( .A1(_07529_ ), .A2(_05224_ ), .ZN(_07530_ ) );
NOR3_X1 _15524_ ( .A1(_07073_ ), .A2(_06925_ ), .A3(_07074_ ), .ZN(_07531_ ) );
OAI211_X1 _15525_ ( .A(_06866_ ), .B(_07452_ ), .C1(_07531_ ), .C2(_07453_ ), .ZN(_07532_ ) );
NOR2_X1 _15526_ ( .A1(_07510_ ), .A2(_07153_ ), .ZN(_07533_ ) );
OAI21_X1 _15527_ ( .A(_07533_ ), .B1(_04343_ ), .B2(_07406_ ), .ZN(_07534_ ) );
AOI21_X1 _15528_ ( .A(_07007_ ), .B1(_07091_ ), .B2(_07098_ ), .ZN(_07535_ ) );
NAND3_X1 _15529_ ( .A1(_07359_ ), .A2(_07360_ ), .A3(_07039_ ), .ZN(_07536_ ) );
OAI21_X1 _15530_ ( .A(_06949_ ), .B1(_07461_ ), .B2(_07124_ ), .ZN(_07537_ ) );
NOR2_X1 _15531_ ( .A1(_06936_ ), .A2(_04194_ ), .ZN(_07538_ ) );
OAI21_X1 _15532_ ( .A(_06912_ ), .B1(_07538_ ), .B2(_07135_ ), .ZN(_07539_ ) );
NAND3_X1 _15533_ ( .A1(_07537_ ), .A2(_07539_ ), .A3(_06931_ ), .ZN(_07540_ ) );
NAND2_X1 _15534_ ( .A1(_07536_ ), .A2(_07540_ ), .ZN(_07541_ ) );
AOI211_X1 _15535_ ( .A(_07004_ ), .B(_07535_ ), .C1(_07008_ ), .C2(_07541_ ), .ZN(_07542_ ) );
NAND3_X1 _15536_ ( .A1(_07082_ ), .A2(_07006_ ), .A3(_06973_ ), .ZN(_07543_ ) );
AOI211_X1 _15537_ ( .A(_07014_ ), .B(_07542_ ), .C1(_07005_ ), .C2(_07543_ ), .ZN(_07544_ ) );
OR3_X1 _15538_ ( .A1(_07138_ ), .A2(_06962_ ), .A3(_07145_ ), .ZN(_07545_ ) );
OAI21_X1 _15539_ ( .A(_07545_ ), .B1(_07114_ ), .B2(_07008_ ), .ZN(_07546_ ) );
AND2_X1 _15540_ ( .A1(_07546_ ), .A2(_07432_ ), .ZN(_07547_ ) );
AND3_X1 _15541_ ( .A1(_04341_ ), .A2(_02863_ ), .A3(_06857_ ), .ZN(_07548_ ) );
OAI21_X1 _15542_ ( .A(_07296_ ), .B1(_04341_ ), .B2(_02863_ ), .ZN(_07549_ ) );
OAI21_X1 _15543_ ( .A(_07549_ ), .B1(_07509_ ), .B2(_07198_ ), .ZN(_07550_ ) );
NOR4_X1 _15544_ ( .A1(_07544_ ), .A2(_07547_ ), .A3(_07548_ ), .A4(_07550_ ), .ZN(_07551_ ) );
NAND3_X1 _15545_ ( .A1(_07532_ ), .A2(_07534_ ), .A3(_07551_ ), .ZN(_07552_ ) );
AOI21_X1 _15546_ ( .A(_07530_ ), .B1(_07070_ ), .B2(_07552_ ), .ZN(_07553_ ) );
OAI21_X1 _15547_ ( .A(_07236_ ), .B1(_04939_ ), .B2(_04720_ ), .ZN(_07554_ ) );
OAI21_X1 _15548_ ( .A(_07525_ ), .B1(_07553_ ), .B2(_07554_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
OAI211_X1 _15549_ ( .A(_06541_ ), .B(_06457_ ), .C1(_06543_ ), .C2(\EX_LS_result_csreg_mem [30] ), .ZN(_07555_ ) );
AND2_X1 _15550_ ( .A1(_04460_ ), .A2(_04465_ ), .ZN(_07556_ ) );
NAND4_X2 _15551_ ( .A1(_07154_ ), .A2(_04451_ ), .A3(_04455_ ), .A4(_07556_ ), .ZN(_07557_ ) );
INV_X1 _15552_ ( .A(_04451_ ), .ZN(_07558_ ) );
NOR2_X1 _15553_ ( .A1(_04459_ ), .A2(_03778_ ), .ZN(_07559_ ) );
AOI21_X1 _15554_ ( .A(_07559_ ), .B1(_04460_ ), .B2(_06855_ ), .ZN(_07560_ ) );
INV_X1 _15555_ ( .A(_04455_ ), .ZN(_07561_ ) );
NOR3_X1 _15556_ ( .A1(_07558_ ), .A2(_07560_ ), .A3(_07561_ ), .ZN(_07562_ ) );
OR2_X1 _15557_ ( .A1(_04454_ ), .A2(_04500_ ), .ZN(_07563_ ) );
NOR3_X1 _15558_ ( .A1(_04449_ ), .A2(_04450_ ), .A3(_07563_ ), .ZN(_07564_ ) );
NOR3_X1 _15559_ ( .A1(_07562_ ), .A2(_04449_ ), .A3(_07564_ ), .ZN(_07565_ ) );
AND2_X4 _15560_ ( .A1(_07557_ ), .A2(_07565_ ), .ZN(_07566_ ) );
NAND4_X1 _15561_ ( .A1(_04514_ ), .A2(_04534_ ), .A3(_04521_ ), .A4(_04527_ ), .ZN(_07567_ ) );
OR2_X4 _15562_ ( .A1(_07566_ ), .A2(_07567_ ), .ZN(_07568_ ) );
INV_X1 _15563_ ( .A(_04514_ ), .ZN(_07569_ ) );
INV_X1 _15564_ ( .A(_04538_ ), .ZN(_07570_ ) );
AOI21_X1 _15565_ ( .A(_04539_ ), .B1(_07570_ ), .B2(_04532_ ), .ZN(_07571_ ) );
NOR3_X1 _15566_ ( .A1(_07569_ ), .A2(_07571_ ), .A3(_04542_ ), .ZN(_07572_ ) );
AOI211_X1 _15567_ ( .A(_04519_ ), .B(_07572_ ), .C1(_04521_ ), .C2(_04512_ ), .ZN(_07573_ ) );
AND2_X4 _15568_ ( .A1(_07568_ ), .A2(_07573_ ), .ZN(_07574_ ) );
INV_X4 _15569_ ( .A(_07574_ ), .ZN(_07575_ ) );
NAND3_X4 _15570_ ( .A1(_07575_ ), .A2(_04314_ ), .A3(_04320_ ), .ZN(_07576_ ) );
INV_X1 _15571_ ( .A(_04309_ ), .ZN(_07577_ ) );
AND2_X1 _15572_ ( .A1(_04318_ ), .A2(_02388_ ), .ZN(_07578_ ) );
AND2_X1 _15573_ ( .A1(_04314_ ), .A2(_07578_ ), .ZN(_07579_ ) );
AOI21_X1 _15574_ ( .A(_07579_ ), .B1(_03150_ ), .B2(_04313_ ), .ZN(_07580_ ) );
AND3_X1 _15575_ ( .A1(_07576_ ), .A2(_07577_ ), .A3(_07580_ ), .ZN(_07581_ ) );
AOI21_X2 _15576_ ( .A(_07577_ ), .B1(_07576_ ), .B2(_07580_ ), .ZN(_07582_ ) );
OR3_X1 _15577_ ( .A1(_07581_ ), .A2(_07582_ ), .A3(_07153_ ), .ZN(_07583_ ) );
NAND2_X1 _15578_ ( .A1(_04309_ ), .A2(_07011_ ), .ZN(_07584_ ) );
INV_X1 _15579_ ( .A(_07455_ ), .ZN(_07585_ ) );
AOI21_X1 _15580_ ( .A(_07585_ ), .B1(_07312_ ), .B2(_07313_ ), .ZN(_07586_ ) );
AOI21_X1 _15581_ ( .A(_07586_ ), .B1(_06966_ ), .B2(_07469_ ), .ZN(_07587_ ) );
AND2_X1 _15582_ ( .A1(_06903_ ), .A2(_06909_ ), .ZN(_07588_ ) );
AND4_X1 _15583_ ( .A1(_06925_ ), .A2(_06888_ ), .A3(_06900_ ), .A4(_06907_ ), .ZN(_07589_ ) );
NOR2_X1 _15584_ ( .A1(_07588_ ), .A2(_07589_ ), .ZN(_07590_ ) );
AOI21_X1 _15585_ ( .A(_07071_ ), .B1(_07587_ ), .B2(_07590_ ), .ZN(_07591_ ) );
AND2_X1 _15586_ ( .A1(_06916_ ), .A2(_02358_ ), .ZN(_07592_ ) );
OR3_X1 _15587_ ( .A1(_07592_ ), .A2(_07116_ ), .A3(_07077_ ), .ZN(_07593_ ) );
NOR2_X1 _15588_ ( .A1(_07085_ ), .A2(_07078_ ), .ZN(_07594_ ) );
INV_X1 _15589_ ( .A(_07594_ ), .ZN(_07595_ ) );
OAI211_X1 _15590_ ( .A(_07593_ ), .B(_06959_ ), .C1(_06992_ ), .C2(_07595_ ), .ZN(_07596_ ) );
OR3_X1 _15591_ ( .A1(_07116_ ), .A2(_07088_ ), .A3(_07086_ ), .ZN(_07597_ ) );
OR3_X1 _15592_ ( .A1(_07092_ ), .A2(_06976_ ), .A3(_07089_ ), .ZN(_07598_ ) );
NAND3_X1 _15593_ ( .A1(_07597_ ), .A2(_07598_ ), .A3(_07039_ ), .ZN(_07599_ ) );
AOI21_X1 _15594_ ( .A(_06961_ ), .B1(_07596_ ), .B2(_07599_ ), .ZN(_07600_ ) );
NAND3_X1 _15595_ ( .A1(_07275_ ), .A2(_07039_ ), .A3(_07276_ ), .ZN(_07601_ ) );
OAI21_X1 _15596_ ( .A(_07116_ ), .B1(_07121_ ), .B2(_07096_ ), .ZN(_07602_ ) );
OAI21_X1 _15597_ ( .A(_06913_ ), .B1(_07095_ ), .B2(_07093_ ), .ZN(_07603_ ) );
NAND2_X1 _15598_ ( .A1(_07602_ ), .A2(_07603_ ), .ZN(_07604_ ) );
NAND2_X1 _15599_ ( .A1(_07604_ ), .A2(_06931_ ), .ZN(_07605_ ) );
AOI21_X1 _15600_ ( .A(_07006_ ), .B1(_07601_ ), .B2(_07605_ ), .ZN(_07606_ ) );
OR3_X1 _15601_ ( .A1(_07600_ ), .A2(_07003_ ), .A3(_07606_ ), .ZN(_07607_ ) );
OAI21_X1 _15602_ ( .A(_07003_ ), .B1(_07473_ ), .B2(_07476_ ), .ZN(_07608_ ) );
AOI21_X1 _15603_ ( .A(_06929_ ), .B1(_07607_ ), .B2(_07608_ ), .ZN(_07609_ ) );
AND3_X1 _15604_ ( .A1(_07469_ ), .A2(_06966_ ), .A3(_07013_ ), .ZN(_07610_ ) );
NOR3_X1 _15605_ ( .A1(_07591_ ), .A2(_07609_ ), .A3(_07610_ ), .ZN(_07611_ ) );
NAND3_X1 _15606_ ( .A1(_04308_ ), .A2(_07080_ ), .A3(_07478_ ), .ZN(_07612_ ) );
OAI21_X1 _15607_ ( .A(_07296_ ), .B1(_04308_ ), .B2(_07080_ ), .ZN(_07613_ ) );
AND4_X1 _15608_ ( .A1(_07584_ ), .A2(_07611_ ), .A3(_07612_ ), .A4(_07613_ ), .ZN(_07614_ ) );
AOI21_X1 _15609_ ( .A(_07056_ ), .B1(_07583_ ), .B2(_07614_ ), .ZN(_07615_ ) );
NAND2_X1 _15610_ ( .A1(_06772_ ), .A2(_03899_ ), .ZN(_07616_ ) );
AND2_X1 _15611_ ( .A1(_07616_ ), .A2(_04615_ ), .ZN(_07617_ ) );
INV_X1 _15612_ ( .A(_03611_ ), .ZN(_07618_ ) );
OAI21_X1 _15613_ ( .A(_04626_ ), .B1(_07617_ ), .B2(_07618_ ), .ZN(_07619_ ) );
NAND2_X1 _15614_ ( .A1(_07619_ ), .A2(_03655_ ), .ZN(_07620_ ) );
AND3_X1 _15615_ ( .A1(_07620_ ), .A2(_04633_ ), .A3(_04632_ ), .ZN(_07621_ ) );
AOI21_X1 _15616_ ( .A(_04633_ ), .B1(_07620_ ), .B2(_04632_ ), .ZN(_07622_ ) );
OR3_X1 _15617_ ( .A1(_07621_ ), .A2(_07622_ ), .A3(_07240_ ), .ZN(_07623_ ) );
AND3_X1 _15618_ ( .A1(_06768_ ), .A2(\ID_EX_imm [30] ), .A3(_06764_ ), .ZN(_07624_ ) );
AOI21_X1 _15619_ ( .A(_07624_ ), .B1(_03370_ ), .B2(_07065_ ), .ZN(_07625_ ) );
AOI21_X1 _15620_ ( .A(_06787_ ), .B1(_07623_ ), .B2(_07625_ ), .ZN(_07626_ ) );
NOR3_X1 _15621_ ( .A1(_07615_ ), .A2(_07626_ ), .A3(_05320_ ), .ZN(_07627_ ) );
OAI21_X1 _15622_ ( .A(_07236_ ), .B1(_03466_ ), .B2(_04720_ ), .ZN(_07628_ ) );
OAI21_X1 _15623_ ( .A(_07555_ ), .B1(_07627_ ), .B2(_07628_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
INV_X1 _15624_ ( .A(_04167_ ), .ZN(_07629_ ) );
NOR4_X1 _15625_ ( .A1(_04570_ ), .A2(_07629_ ), .A3(_04189_ ), .A4(_04190_ ), .ZN(_07630_ ) );
OR3_X1 _15626_ ( .A1(_07630_ ), .A2(_04189_ ), .A3(_04580_ ), .ZN(_07631_ ) );
XOR2_X1 _15627_ ( .A(_02912_ ), .B(_04142_ ), .Z(_07632_ ) );
AND2_X1 _15628_ ( .A1(_07631_ ), .A2(_07632_ ), .ZN(_07633_ ) );
OR3_X1 _15629_ ( .A1(_07633_ ), .A2(_04121_ ), .A3(_04143_ ), .ZN(_07634_ ) );
OAI21_X1 _15630_ ( .A(_04121_ ), .B1(_07633_ ), .B2(_04143_ ), .ZN(_07635_ ) );
AOI21_X1 _15631_ ( .A(_07240_ ), .B1(_07634_ ), .B2(_07635_ ), .ZN(_07636_ ) );
OAI22_X1 _15632_ ( .A1(_04966_ ), .A2(_07305_ ), .B1(_02937_ ), .B2(_06770_ ), .ZN(_07637_ ) );
OAI21_X1 _15633_ ( .A(_06784_ ), .B1(_07636_ ), .B2(_07637_ ), .ZN(_07638_ ) );
NAND2_X1 _15634_ ( .A1(_07638_ ), .A2(_04720_ ), .ZN(_07639_ ) );
OAI211_X1 _15635_ ( .A(_06910_ ), .B(_07452_ ), .C1(_06926_ ), .C2(_07193_ ), .ZN(_07640_ ) );
NOR2_X1 _15636_ ( .A1(_07640_ ), .A2(_07072_ ), .ZN(_07641_ ) );
OR3_X1 _15637_ ( .A1(_07179_ ), .A2(_07182_ ), .A3(_07041_ ), .ZN(_07642_ ) );
NAND3_X1 _15638_ ( .A1(_07418_ ), .A2(_07419_ ), .A3(_07001_ ), .ZN(_07643_ ) );
OAI21_X1 _15639_ ( .A(_07117_ ), .B1(_06944_ ), .B2(_06974_ ), .ZN(_07644_ ) );
OAI21_X1 _15640_ ( .A(_06914_ ), .B1(_07218_ ), .B2(_07226_ ), .ZN(_07645_ ) );
NAND2_X1 _15641_ ( .A1(_07644_ ), .A2(_07645_ ), .ZN(_07646_ ) );
NAND2_X1 _15642_ ( .A1(_07646_ ), .A2(_07022_ ), .ZN(_07647_ ) );
AND2_X1 _15643_ ( .A1(_07643_ ), .A2(_07647_ ), .ZN(_07648_ ) );
OAI211_X1 _15644_ ( .A(_07642_ ), .B(_07101_ ), .C1(_06968_ ), .C2(_07648_ ), .ZN(_07649_ ) );
OR3_X1 _15645_ ( .A1(_07189_ ), .A2(_06966_ ), .A3(_06963_ ), .ZN(_07650_ ) );
AOI21_X1 _15646_ ( .A(_07014_ ), .B1(_07649_ ), .B2(_07650_ ), .ZN(_07651_ ) );
OR3_X1 _15647_ ( .A1(_04349_ ), .A2(_04350_ ), .A3(_04646_ ), .ZN(_07652_ ) );
NAND3_X1 _15648_ ( .A1(_04432_ ), .A2(_02936_ ), .A3(_06857_ ), .ZN(_07653_ ) );
OR2_X1 _15649_ ( .A1(_04350_ ), .A2(_07047_ ), .ZN(_07654_ ) );
NAND3_X1 _15650_ ( .A1(_07652_ ), .A2(_07653_ ), .A3(_07654_ ), .ZN(_07655_ ) );
NAND2_X1 _15651_ ( .A1(_07230_ ), .A2(_07042_ ), .ZN(_07656_ ) );
NAND3_X1 _15652_ ( .A1(_07212_ ), .A2(_07084_ ), .A3(_07022_ ), .ZN(_07657_ ) );
AOI21_X1 _15653_ ( .A(_07519_ ), .B1(_07656_ ), .B2(_07657_ ), .ZN(_07658_ ) );
NOR4_X1 _15654_ ( .A1(_07641_ ), .A2(_07651_ ), .A3(_07655_ ), .A4(_07658_ ), .ZN(_07659_ ) );
INV_X1 _15655_ ( .A(_07402_ ), .ZN(_07660_ ) );
NAND2_X1 _15656_ ( .A1(_07660_ ), .A2(_06792_ ), .ZN(_07661_ ) );
AOI21_X1 _15657_ ( .A(_06823_ ), .B1(_07661_ ), .B2(_06822_ ), .ZN(_07662_ ) );
OR3_X1 _15658_ ( .A1(_07662_ ), .A2(_04351_ ), .A3(_06825_ ), .ZN(_07663_ ) );
OAI21_X1 _15659_ ( .A(_04351_ ), .B1(_07662_ ), .B2(_06825_ ), .ZN(_07664_ ) );
NAND3_X1 _15660_ ( .A1(_07663_ ), .A2(_06861_ ), .A3(_07664_ ), .ZN(_07665_ ) );
AOI21_X1 _15661_ ( .A(_07056_ ), .B1(_07659_ ), .B2(_07665_ ), .ZN(_07666_ ) );
OAI221_X1 _15662_ ( .A(_06488_ ), .B1(_04720_ ), .B2(_04959_ ), .C1(_07639_ ), .C2(_07666_ ), .ZN(_07667_ ) );
INV_X1 _15663_ ( .A(_06550_ ), .ZN(_07668_ ) );
NAND2_X1 _15664_ ( .A1(_07667_ ), .A2(_07668_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
OR2_X1 _15665_ ( .A1(_06554_ ), .A2(_07349_ ), .ZN(_07669_ ) );
AOI21_X1 _15666_ ( .A(_07240_ ), .B1(_07631_ ), .B2(_07632_ ), .ZN(_07670_ ) );
OAI21_X1 _15667_ ( .A(_07670_ ), .B1(_07632_ ), .B2(_07631_ ), .ZN(_07671_ ) );
AOI22_X1 _15668_ ( .A1(_05007_ ), .A2(_07446_ ), .B1(\ID_EX_imm [10] ), .B2(_07066_ ), .ZN(_07672_ ) );
AOI21_X1 _15669_ ( .A(_07166_ ), .B1(_07671_ ), .B2(_07672_ ), .ZN(_07673_ ) );
OR2_X1 _15670_ ( .A1(_07673_ ), .A2(_05224_ ), .ZN(_07674_ ) );
INV_X1 _15671_ ( .A(_07453_ ), .ZN(_07675_ ) );
OAI21_X1 _15672_ ( .A(_07675_ ), .B1(_07248_ ), .B2(_07249_ ), .ZN(_07676_ ) );
NAND2_X1 _15673_ ( .A1(_07676_ ), .A2(_07452_ ), .ZN(_07677_ ) );
OR3_X1 _15674_ ( .A1(_07264_ ), .A2(_06965_ ), .A3(_06962_ ), .ZN(_07678_ ) );
NOR3_X1 _15675_ ( .A1(_07462_ ), .A2(_07463_ ), .A3(_06932_ ), .ZN(_07679_ ) );
OAI21_X1 _15676_ ( .A(_07117_ ), .B1(_07538_ ), .B2(_07135_ ), .ZN(_07680_ ) );
NOR2_X1 _15677_ ( .A1(_06916_ ), .A2(_02936_ ), .ZN(_07681_ ) );
OAI21_X1 _15678_ ( .A(_06914_ ), .B1(_07681_ ), .B2(_07132_ ), .ZN(_07682_ ) );
AOI21_X1 _15679_ ( .A(_07001_ ), .B1(_07680_ ), .B2(_07682_ ), .ZN(_07683_ ) );
OAI21_X1 _15680_ ( .A(_07007_ ), .B1(_07679_ ), .B2(_07683_ ), .ZN(_07684_ ) );
NAND3_X1 _15681_ ( .A1(_07255_ ), .A2(_06962_ ), .A3(_07258_ ), .ZN(_07685_ ) );
NAND3_X1 _15682_ ( .A1(_07684_ ), .A2(_06966_ ), .A3(_07685_ ), .ZN(_07686_ ) );
AND2_X1 _15683_ ( .A1(_07678_ ), .A2(_07686_ ), .ZN(_07687_ ) );
AOI21_X1 _15684_ ( .A(_07072_ ), .B1(_07677_ ), .B2(_07687_ ), .ZN(_07688_ ) );
AND3_X1 _15685_ ( .A1(_07661_ ), .A2(_06823_ ), .A3(_06822_ ), .ZN(_07689_ ) );
NOR3_X1 _15686_ ( .A1(_07689_ ), .A2(_07662_ ), .A3(_07152_ ), .ZN(_07690_ ) );
NAND3_X1 _15687_ ( .A1(_07284_ ), .A2(_07006_ ), .A3(_07289_ ), .ZN(_07691_ ) );
NAND4_X1 _15688_ ( .A1(_07270_ ), .A2(_06961_ ), .A3(_07271_ ), .A4(_06931_ ), .ZN(_07692_ ) );
AOI21_X1 _15689_ ( .A(_07519_ ), .B1(_07691_ ), .B2(_07692_ ), .ZN(_07693_ ) );
AOI221_X4 _15690_ ( .A(_07693_ ), .B1(_06825_ ), .B2(_06857_ ), .C1(_04355_ ), .C2(_04645_ ), .ZN(_07694_ ) );
OAI21_X1 _15691_ ( .A(_07296_ ), .B1(_04435_ ), .B2(_02912_ ), .ZN(_07695_ ) );
INV_X1 _15692_ ( .A(_07013_ ), .ZN(_07696_ ) );
OAI211_X1 _15693_ ( .A(_07694_ ), .B(_07695_ ), .C1(_07696_ ), .C2(_07687_ ), .ZN(_07697_ ) );
OR3_X1 _15694_ ( .A1(_07688_ ), .A2(_07690_ ), .A3(_07697_ ), .ZN(_07698_ ) );
AOI21_X1 _15695_ ( .A(_07674_ ), .B1(_07070_ ), .B2(_07698_ ), .ZN(_07699_ ) );
NAND2_X1 _15696_ ( .A1(_05005_ ), .A2(_05320_ ), .ZN(_07700_ ) );
NAND2_X1 _15697_ ( .A1(_07700_ ), .A2(_07441_ ), .ZN(_07701_ ) );
OAI21_X1 _15698_ ( .A(_07669_ ), .B1(_07699_ ), .B2(_07701_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
OR2_X1 _15699_ ( .A1(_05037_ ), .A2(_07349_ ), .ZN(_07702_ ) );
NOR2_X1 _15700_ ( .A1(_04570_ ), .A2(_07629_ ), .ZN(_07703_ ) );
AOI21_X1 _15701_ ( .A(_07703_ ), .B1(_02960_ ), .B2(_04166_ ), .ZN(_07704_ ) );
XNOR2_X1 _15702_ ( .A(_07704_ ), .B(_04191_ ), .ZN(_07705_ ) );
NAND2_X1 _15703_ ( .A1(_07705_ ), .A2(_06782_ ), .ZN(_07706_ ) );
AOI22_X1 _15704_ ( .A1(_05026_ ), .A2(_07446_ ), .B1(\ID_EX_imm [9] ), .B2(_07066_ ), .ZN(_07707_ ) );
AOI21_X1 _15705_ ( .A(_07166_ ), .B1(_07706_ ), .B2(_07707_ ), .ZN(_07708_ ) );
OR2_X1 _15706_ ( .A1(_07708_ ), .A2(_05224_ ), .ZN(_07709_ ) );
NAND3_X1 _15707_ ( .A1(_07317_ ), .A2(_07318_ ), .A3(_07084_ ), .ZN(_07710_ ) );
OAI21_X1 _15708_ ( .A(_06950_ ), .B1(_07218_ ), .B2(_07226_ ), .ZN(_07711_ ) );
OAI21_X1 _15709_ ( .A(_06914_ ), .B1(_06969_ ), .B2(_06983_ ), .ZN(_07712_ ) );
NAND2_X1 _15710_ ( .A1(_07711_ ), .A2(_07712_ ), .ZN(_07713_ ) );
NAND2_X1 _15711_ ( .A1(_07713_ ), .A2(_06973_ ), .ZN(_07714_ ) );
NAND3_X1 _15712_ ( .A1(_07501_ ), .A2(_07001_ ), .A3(_07502_ ), .ZN(_07715_ ) );
NAND3_X1 _15713_ ( .A1(_07714_ ), .A2(_07715_ ), .A3(_07007_ ), .ZN(_07716_ ) );
AOI21_X1 _15714_ ( .A(_07004_ ), .B1(_07710_ ), .B2(_07716_ ), .ZN(_07717_ ) );
NOR3_X1 _15715_ ( .A1(_07320_ ), .A2(_06966_ ), .A3(_06963_ ), .ZN(_07718_ ) );
AOI211_X1 _15716_ ( .A(_07717_ ), .B(_07718_ ), .C1(_07453_ ), .C2(_07452_ ), .ZN(_07719_ ) );
NAND4_X1 _15717_ ( .A1(_07247_ ), .A2(_06918_ ), .A3(_06924_ ), .A4(_07452_ ), .ZN(_07720_ ) );
AOI21_X1 _15718_ ( .A(_07072_ ), .B1(_07719_ ), .B2(_07720_ ), .ZN(_07721_ ) );
AOI21_X1 _15719_ ( .A(_04362_ ), .B1(_06811_ ), .B2(_06819_ ), .ZN(_07722_ ) );
OR3_X1 _15720_ ( .A1(_07722_ ), .A2(_04427_ ), .A3(_06821_ ), .ZN(_07723_ ) );
OAI21_X1 _15721_ ( .A(_04427_ ), .B1(_07722_ ), .B2(_06821_ ), .ZN(_07724_ ) );
AND3_X1 _15722_ ( .A1(_07723_ ), .A2(_06861_ ), .A3(_07724_ ), .ZN(_07725_ ) );
OAI21_X1 _15723_ ( .A(_07149_ ), .B1(_07718_ ), .B2(_07717_ ), .ZN(_07726_ ) );
NAND3_X1 _15724_ ( .A1(_07338_ ), .A2(_07339_ ), .A3(_07041_ ), .ZN(_07727_ ) );
NAND4_X1 _15725_ ( .A1(_07379_ ), .A2(_06973_ ), .A3(_06992_ ), .A4(_06991_ ), .ZN(_07728_ ) );
NAND2_X1 _15726_ ( .A1(_07727_ ), .A2(_07728_ ), .ZN(_07729_ ) );
NAND2_X1 _15727_ ( .A1(_07729_ ), .A2(_07432_ ), .ZN(_07730_ ) );
NOR3_X1 _15728_ ( .A1(_04367_ ), .A2(_04368_ ), .A3(_04646_ ), .ZN(_07731_ ) );
NOR3_X1 _15729_ ( .A1(_04365_ ), .A2(_04366_ ), .A3(_07045_ ), .ZN(_07732_ ) );
AOI21_X1 _15730_ ( .A(_07047_ ), .B1(_04365_ ), .B2(_04366_ ), .ZN(_07733_ ) );
NOR3_X1 _15731_ ( .A1(_07731_ ), .A2(_07732_ ), .A3(_07733_ ), .ZN(_07734_ ) );
NAND3_X1 _15732_ ( .A1(_07726_ ), .A2(_07730_ ), .A3(_07734_ ), .ZN(_07735_ ) );
OR3_X1 _15733_ ( .A1(_07721_ ), .A2(_07725_ ), .A3(_07735_ ), .ZN(_07736_ ) );
AOI21_X1 _15734_ ( .A(_07709_ ), .B1(_07058_ ), .B2(_07736_ ), .ZN(_07737_ ) );
NAND2_X1 _15735_ ( .A1(_05028_ ), .A2(_05320_ ), .ZN(_07738_ ) );
NAND2_X1 _15736_ ( .A1(_07738_ ), .A2(_07441_ ), .ZN(_07739_ ) );
OAI21_X1 _15737_ ( .A(_07702_ ), .B1(_07737_ ), .B2(_07739_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _15738_ ( .A(_07239_ ), .B1(_04571_ ), .B2(_04167_ ), .ZN(_07740_ ) );
OAI21_X1 _15739_ ( .A(_07740_ ), .B1(_04167_ ), .B2(_04571_ ), .ZN(_07741_ ) );
AND3_X1 _15740_ ( .A1(_06768_ ), .A2(\ID_EX_imm [8] ), .A3(_06764_ ), .ZN(_07742_ ) );
AOI21_X1 _15741_ ( .A(_07742_ ), .B1(_05046_ ), .B2(_06766_ ), .ZN(_07743_ ) );
AOI21_X1 _15742_ ( .A(_06785_ ), .B1(_07741_ ), .B2(_07743_ ), .ZN(_07744_ ) );
NOR2_X1 _15743_ ( .A1(_07744_ ), .A2(_02272_ ), .ZN(_07745_ ) );
NOR2_X1 _15744_ ( .A1(_06884_ ), .A2(_07379_ ), .ZN(_07746_ ) );
INV_X1 _15745_ ( .A(_07746_ ), .ZN(_07747_ ) );
NAND4_X1 _15746_ ( .A1(_06910_ ), .A2(_06909_ ), .A3(_07747_ ), .A4(_06902_ ), .ZN(_07748_ ) );
OR3_X1 _15747_ ( .A1(_07364_ ), .A2(_06905_ ), .A3(_06804_ ), .ZN(_07749_ ) );
NAND3_X1 _15748_ ( .A1(_07358_ ), .A2(_07361_ ), .A3(_06804_ ), .ZN(_07750_ ) );
NAND3_X1 _15749_ ( .A1(_07537_ ), .A2(_07539_ ), .A3(_06919_ ), .ZN(_07751_ ) );
OAI21_X1 _15750_ ( .A(_06949_ ), .B1(_07681_ ), .B2(_07132_ ), .ZN(_07752_ ) );
OAI21_X1 _15751_ ( .A(_06976_ ), .B1(_07286_ ), .B2(_07143_ ), .ZN(_07753_ ) );
NAND3_X1 _15752_ ( .A1(_07752_ ), .A2(_07753_ ), .A3(_06930_ ), .ZN(_07754_ ) );
NAND2_X1 _15753_ ( .A1(_07751_ ), .A2(_07754_ ), .ZN(_07755_ ) );
OAI211_X1 _15754_ ( .A(_07750_ ), .B(_06905_ ), .C1(_07755_ ), .C2(_06961_ ), .ZN(_07756_ ) );
AND2_X1 _15755_ ( .A1(_07749_ ), .A2(_07756_ ), .ZN(_07757_ ) );
AOI21_X1 _15756_ ( .A(_07072_ ), .B1(_07748_ ), .B2(_07757_ ), .ZN(_07758_ ) );
NOR2_X1 _15757_ ( .A1(_07722_ ), .A2(_07152_ ), .ZN(_07759_ ) );
OAI21_X1 _15758_ ( .A(_07759_ ), .B1(_04361_ ), .B2(_07660_ ), .ZN(_07760_ ) );
OR2_X1 _15759_ ( .A1(_07757_ ), .A2(_07696_ ), .ZN(_07761_ ) );
OAI21_X1 _15760_ ( .A(_07296_ ), .B1(_04429_ ), .B2(_02960_ ), .ZN(_07762_ ) );
OAI21_X1 _15761_ ( .A(_06805_ ), .B1(_07376_ ), .B2(_07377_ ), .ZN(_07763_ ) );
OR2_X1 _15762_ ( .A1(_06805_ ), .A2(_07370_ ), .ZN(_07764_ ) );
AND3_X1 _15763_ ( .A1(_07763_ ), .A2(_07431_ ), .A3(_07764_ ), .ZN(_07765_ ) );
AOI221_X4 _15764_ ( .A(_07765_ ), .B1(_06821_ ), .B2(_06857_ ), .C1(_04361_ ), .C2(_04645_ ), .ZN(_07766_ ) );
NAND4_X1 _15765_ ( .A1(_07760_ ), .A2(_07761_ ), .A3(_07762_ ), .A4(_07766_ ), .ZN(_07767_ ) );
OAI21_X1 _15766_ ( .A(_07057_ ), .B1(_07758_ ), .B2(_07767_ ), .ZN(_07768_ ) );
AOI221_X4 _15767_ ( .A(_06421_ ), .B1(_02272_ ), .B2(_05048_ ), .C1(_07745_ ), .C2(_07768_ ), .ZN(_07769_ ) );
AOI21_X1 _15768_ ( .A(_07349_ ), .B1(_05057_ ), .B2(_05058_ ), .ZN(_07770_ ) );
OR2_X1 _15769_ ( .A1(_07769_ ), .A2(_07770_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
OR2_X1 _15770_ ( .A1(_05078_ ), .A2(_07349_ ), .ZN(_07771_ ) );
AOI21_X1 _15771_ ( .A(_07240_ ), .B1(_04567_ ), .B2(_03924_ ), .ZN(_07772_ ) );
OAI21_X1 _15772_ ( .A(_07772_ ), .B1(_03924_ ), .B2(_04567_ ), .ZN(_07773_ ) );
BUF_X4 _15773_ ( .A(_06769_ ), .Z(_07774_ ) );
AOI22_X1 _15774_ ( .A1(_05067_ ), .A2(_07446_ ), .B1(\ID_EX_imm [7] ), .B2(_07774_ ), .ZN(_07775_ ) );
AOI21_X1 _15775_ ( .A(_07166_ ), .B1(_07773_ ), .B2(_07775_ ), .ZN(_07776_ ) );
OR2_X1 _15776_ ( .A1(_07776_ ), .A2(_05224_ ), .ZN(_07777_ ) );
AND4_X1 _15777_ ( .A1(_06926_ ), .A2(_06910_ ), .A3(_06866_ ), .A4(_07452_ ), .ZN(_07778_ ) );
OR3_X1 _15778_ ( .A1(_07414_ ), .A2(_06804_ ), .A3(_07415_ ), .ZN(_07779_ ) );
NAND4_X1 _15779_ ( .A1(_06804_ ), .A2(_03185_ ), .A3(_06883_ ), .A4(_06958_ ), .ZN(_07780_ ) );
NAND2_X1 _15780_ ( .A1(_07779_ ), .A2(_07780_ ), .ZN(_07781_ ) );
NAND2_X1 _15781_ ( .A1(_07781_ ), .A2(_07005_ ), .ZN(_07782_ ) );
OAI21_X1 _15782_ ( .A(_06914_ ), .B1(_06982_ ), .B2(_06980_ ), .ZN(_07783_ ) );
OAI21_X1 _15783_ ( .A(_06950_ ), .B1(_06969_ ), .B2(_06983_ ), .ZN(_07784_ ) );
NAND3_X1 _15784_ ( .A1(_07783_ ), .A2(_07784_ ), .A3(_07023_ ), .ZN(_07785_ ) );
OAI211_X1 _15785_ ( .A(_07785_ ), .B(_07008_ ), .C1(_07023_ ), .C2(_07646_ ), .ZN(_07786_ ) );
OAI211_X1 _15786_ ( .A(_06967_ ), .B(_07786_ ), .C1(_07421_ ), .C2(_07008_ ), .ZN(_07787_ ) );
NAND2_X1 _15787_ ( .A1(_07782_ ), .A2(_07787_ ), .ZN(_07788_ ) );
OAI21_X1 _15788_ ( .A(_07467_ ), .B1(_07778_ ), .B2(_07788_ ), .ZN(_07789_ ) );
NAND3_X1 _15789_ ( .A1(_06806_ ), .A2(_06808_ ), .A3(_06809_ ), .ZN(_07790_ ) );
AOI21_X1 _15790_ ( .A(_06812_ ), .B1(_07790_ ), .B2(_06816_ ), .ZN(_07791_ ) );
OR3_X1 _15791_ ( .A1(_07791_ ), .A2(_04399_ ), .A3(_06818_ ), .ZN(_07792_ ) );
OAI21_X1 _15792_ ( .A(_04399_ ), .B1(_07791_ ), .B2(_06818_ ), .ZN(_07793_ ) );
NAND3_X1 _15793_ ( .A1(_07792_ ), .A2(_06862_ ), .A3(_07793_ ), .ZN(_07794_ ) );
NAND3_X1 _15794_ ( .A1(_06868_ ), .A2(_02706_ ), .A3(_06857_ ), .ZN(_07795_ ) );
OAI21_X1 _15795_ ( .A(_07795_ ), .B1(_04398_ ), .B2(_07159_ ), .ZN(_07796_ ) );
NOR3_X1 _15796_ ( .A1(_07426_ ), .A2(_07231_ ), .A3(_07519_ ), .ZN(_07797_ ) );
AOI211_X1 _15797_ ( .A(_07796_ ), .B(_07797_ ), .C1(_04399_ ), .C2(_07011_ ), .ZN(_07798_ ) );
NAND3_X1 _15798_ ( .A1(_07789_ ), .A2(_07794_ ), .A3(_07798_ ), .ZN(_07799_ ) );
AOI21_X1 _15799_ ( .A(_07777_ ), .B1(_07799_ ), .B2(_07057_ ), .ZN(_07800_ ) );
NAND2_X1 _15800_ ( .A1(_05069_ ), .A2(_04755_ ), .ZN(_07801_ ) );
NAND2_X1 _15801_ ( .A1(_07801_ ), .A2(_07441_ ), .ZN(_07802_ ) );
OAI21_X1 _15802_ ( .A(_07771_ ), .B1(_07800_ ), .B2(_07802_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
AOI21_X1 _15803_ ( .A(_05093_ ), .B1(_04776_ ), .B2(_04789_ ), .ZN(_07803_ ) );
NAND2_X1 _15804_ ( .A1(_04781_ ), .A2(\mepc [6] ), .ZN(_07804_ ) );
NAND3_X1 _15805_ ( .A1(_04839_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_04700_ ), .ZN(_07805_ ) );
NAND2_X1 _15806_ ( .A1(_07804_ ), .A2(_07805_ ), .ZN(_07806_ ) );
AND4_X1 _15807_ ( .A1(\mycsreg.CSReg[3][6] ), .A2(_04738_ ), .A3(_05193_ ), .A4(_04701_ ), .ZN(_07807_ ) );
NOR3_X1 _15808_ ( .A1(_07806_ ), .A2(_05136_ ), .A3(_07807_ ), .ZN(_07808_ ) );
NAND2_X1 _15809_ ( .A1(_07803_ ), .A2(_07808_ ), .ZN(_07809_ ) );
NAND4_X1 _15810_ ( .A1(_04789_ ), .A2(_06318_ ), .A3(_04791_ ), .A4(_04792_ ), .ZN(_07810_ ) );
NAND3_X1 _15811_ ( .A1(_07809_ ), .A2(_07810_ ), .A3(_06559_ ), .ZN(_07811_ ) );
NAND2_X1 _15812_ ( .A1(_04563_ ), .A2(_04564_ ), .ZN(_07812_ ) );
NAND3_X1 _15813_ ( .A1(_04565_ ), .A2(_06781_ ), .A3(_07812_ ), .ZN(_07813_ ) );
AOI22_X1 _15814_ ( .A1(_05089_ ), .A2(_07446_ ), .B1(\ID_EX_imm [6] ), .B2(_07774_ ), .ZN(_07814_ ) );
AOI21_X1 _15815_ ( .A(_07166_ ), .B1(_07813_ ), .B2(_07814_ ), .ZN(_07815_ ) );
OR2_X1 _15816_ ( .A1(_07815_ ), .A2(_05319_ ), .ZN(_07816_ ) );
AND3_X1 _15817_ ( .A1(_07455_ ), .A2(_06926_ ), .A3(_07452_ ), .ZN(_07817_ ) );
OR2_X1 _15818_ ( .A1(_07465_ ), .A2(_07007_ ), .ZN(_07818_ ) );
OR3_X1 _15819_ ( .A1(_07117_ ), .A2(_07142_ ), .A3(_07140_ ), .ZN(_07819_ ) );
OR3_X1 _15820_ ( .A1(_07286_ ), .A2(_06914_ ), .A3(_07143_ ), .ZN(_07820_ ) );
AOI21_X1 _15821_ ( .A(_06921_ ), .B1(_07819_ ), .B2(_07820_ ), .ZN(_07821_ ) );
AND3_X1 _15822_ ( .A1(_07680_ ), .A2(_07682_ ), .A3(_07001_ ), .ZN(_07822_ ) );
OAI21_X1 _15823_ ( .A(_07042_ ), .B1(_07821_ ), .B2(_07822_ ), .ZN(_07823_ ) );
AOI21_X1 _15824_ ( .A(_07004_ ), .B1(_07818_ ), .B2(_07823_ ), .ZN(_07824_ ) );
OR3_X1 _15825_ ( .A1(_07457_ ), .A2(_06804_ ), .A3(_07458_ ), .ZN(_07825_ ) );
NAND4_X1 _15826_ ( .A1(_07081_ ), .A2(_06804_ ), .A3(_06958_ ), .A4(_06954_ ), .ZN(_07826_ ) );
AOI21_X1 _15827_ ( .A(_07101_ ), .B1(_07825_ ), .B2(_07826_ ), .ZN(_07827_ ) );
OR2_X1 _15828_ ( .A1(_07824_ ), .A2(_07827_ ), .ZN(_07828_ ) );
OAI21_X1 _15829_ ( .A(_06866_ ), .B1(_07817_ ), .B2(_07828_ ), .ZN(_07829_ ) );
AND3_X1 _15830_ ( .A1(_07790_ ), .A2(_06812_ ), .A3(_06816_ ), .ZN(_07830_ ) );
OR3_X1 _15831_ ( .A1(_07830_ ), .A2(_07791_ ), .A3(_07153_ ), .ZN(_07831_ ) );
OAI21_X1 _15832_ ( .A(_07149_ ), .B1(_07824_ ), .B2(_07827_ ), .ZN(_07832_ ) );
OR3_X1 _15833_ ( .A1(_07472_ ), .A2(_06968_ ), .A3(_07519_ ), .ZN(_07833_ ) );
NAND3_X1 _15834_ ( .A1(_04418_ ), .A2(_02729_ ), .A3(_07478_ ), .ZN(_07834_ ) );
AOI21_X1 _15835_ ( .A(_07159_ ), .B1(_04402_ ), .B2(_04417_ ), .ZN(_07835_ ) );
AOI21_X1 _15836_ ( .A(_07835_ ), .B1(_04403_ ), .B2(_07011_ ), .ZN(_07836_ ) );
AND4_X1 _15837_ ( .A1(_07832_ ), .A2(_07833_ ), .A3(_07834_ ), .A4(_07836_ ), .ZN(_07837_ ) );
NAND3_X1 _15838_ ( .A1(_07829_ ), .A2(_07831_ ), .A3(_07837_ ), .ZN(_07838_ ) );
AOI21_X1 _15839_ ( .A(_07816_ ), .B1(_07838_ ), .B2(_07057_ ), .ZN(_07839_ ) );
NAND2_X1 _15840_ ( .A1(_05091_ ), .A2(_04755_ ), .ZN(_07840_ ) );
NAND2_X1 _15841_ ( .A1(_07840_ ), .A2(_07441_ ), .ZN(_07841_ ) );
OAI21_X1 _15842_ ( .A(_07811_ ), .B1(_07839_ ), .B2(_07841_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
OR2_X1 _15843_ ( .A1(_05120_ ), .A2(_07349_ ), .ZN(_07842_ ) );
NAND3_X1 _15844_ ( .A1(_04560_ ), .A2(_03973_ ), .A3(_04561_ ), .ZN(_07843_ ) );
NAND2_X1 _15845_ ( .A1(_03972_ ), .A2(_02677_ ), .ZN(_07844_ ) );
AND2_X1 _15846_ ( .A1(_07843_ ), .A2(_07844_ ), .ZN(_07845_ ) );
XNOR2_X1 _15847_ ( .A(_07845_ ), .B(_03996_ ), .ZN(_07846_ ) );
NAND2_X1 _15848_ ( .A1(_07846_ ), .A2(_06782_ ), .ZN(_07847_ ) );
AOI22_X1 _15849_ ( .A1(_05109_ ), .A2(_07446_ ), .B1(\ID_EX_imm [5] ), .B2(_07774_ ), .ZN(_07848_ ) );
AOI21_X1 _15850_ ( .A(_07166_ ), .B1(_07847_ ), .B2(_07848_ ), .ZN(_07849_ ) );
OR2_X1 _15851_ ( .A1(_07849_ ), .A2(_05319_ ), .ZN(_07850_ ) );
AND2_X1 _15852_ ( .A1(_07452_ ), .A2(_06865_ ), .ZN(_07851_ ) );
NAND4_X1 _15853_ ( .A1(_06910_ ), .A2(_06923_ ), .A3(_06926_ ), .A4(_07851_ ), .ZN(_07852_ ) );
NAND2_X1 _15854_ ( .A1(_06806_ ), .A2(_06808_ ), .ZN(_07853_ ) );
NOR2_X1 _15855_ ( .A1(_07853_ ), .A2(_04415_ ), .ZN(_07854_ ) );
OAI21_X1 _15856_ ( .A(_04409_ ), .B1(_07854_ ), .B2(_06815_ ), .ZN(_07855_ ) );
INV_X1 _15857_ ( .A(_06815_ ), .ZN(_07856_ ) );
OAI211_X1 _15858_ ( .A(_04410_ ), .B(_07856_ ), .C1(_07853_ ), .C2(_04415_ ), .ZN(_07857_ ) );
NAND3_X1 _15859_ ( .A1(_07855_ ), .A2(_06862_ ), .A3(_07857_ ), .ZN(_07858_ ) );
AOI21_X1 _15860_ ( .A(_07007_ ), .B1(_07500_ ), .B2(_07503_ ), .ZN(_07859_ ) );
OAI21_X1 _15861_ ( .A(_07117_ ), .B1(_06982_ ), .B2(_06980_ ), .ZN(_07860_ ) );
OAI21_X1 _15862_ ( .A(_06992_ ), .B1(_06979_ ), .B2(_06998_ ), .ZN(_07861_ ) );
NAND2_X1 _15863_ ( .A1(_07860_ ), .A2(_07861_ ), .ZN(_07862_ ) );
MUX2_X1 _15864_ ( .A(_07862_ ), .B(_07713_ ), .S(_07001_ ), .Z(_07863_ ) );
AOI211_X1 _15865_ ( .A(_07004_ ), .B(_07859_ ), .C1(_07008_ ), .C2(_07863_ ), .ZN(_07864_ ) );
AOI21_X1 _15866_ ( .A(_07101_ ), .B1(_07024_ ), .B2(_07043_ ), .ZN(_07865_ ) );
OAI21_X1 _15867_ ( .A(_07467_ ), .B1(_07864_ ), .B2(_07865_ ), .ZN(_07866_ ) );
NAND3_X1 _15868_ ( .A1(_07002_ ), .A2(_07008_ ), .A3(_07432_ ), .ZN(_07867_ ) );
NAND3_X1 _15869_ ( .A1(_04407_ ), .A2(_02652_ ), .A3(_07478_ ), .ZN(_07868_ ) );
AOI22_X1 _15870_ ( .A1(_04409_ ), .A2(_07011_ ), .B1(_06813_ ), .B2(_07296_ ), .ZN(_07869_ ) );
AND4_X1 _15871_ ( .A1(_07866_ ), .A2(_07867_ ), .A3(_07868_ ), .A4(_07869_ ), .ZN(_07870_ ) );
NAND3_X1 _15872_ ( .A1(_07852_ ), .A2(_07858_ ), .A3(_07870_ ), .ZN(_07871_ ) );
AOI21_X1 _15873_ ( .A(_07850_ ), .B1(_07871_ ), .B2(_07057_ ), .ZN(_07872_ ) );
NAND2_X1 _15874_ ( .A1(_05111_ ), .A2(_04755_ ), .ZN(_07873_ ) );
NAND2_X1 _15875_ ( .A1(_07873_ ), .A2(_07441_ ), .ZN(_07874_ ) );
OAI21_X1 _15876_ ( .A(_07842_ ), .B1(_07872_ ), .B2(_07874_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
AND3_X1 _15877_ ( .A1(_06602_ ), .A2(_06603_ ), .A3(_06434_ ), .ZN(_07875_ ) );
INV_X1 _15878_ ( .A(_07875_ ), .ZN(_07876_ ) );
OAI211_X1 _15879_ ( .A(_07453_ ), .B(_07851_ ), .C1(_06921_ ), .C2(_06883_ ), .ZN(_07877_ ) );
AND3_X1 _15880_ ( .A1(_07752_ ), .A2(_07753_ ), .A3(_07039_ ), .ZN(_07878_ ) );
NOR2_X1 _15881_ ( .A1(_07139_ ), .A2(_07106_ ), .ZN(_07879_ ) );
NAND2_X1 _15882_ ( .A1(_07879_ ), .A2(_06976_ ), .ZN(_07880_ ) );
OR3_X1 _15883_ ( .A1(_07142_ ), .A2(_06945_ ), .A3(_07140_ ), .ZN(_07881_ ) );
NAND2_X1 _15884_ ( .A1(_07880_ ), .A2(_07881_ ), .ZN(_07882_ ) );
AOI211_X1 _15885_ ( .A(_07379_ ), .B(_07878_ ), .C1(_06973_ ), .C2(_07882_ ), .ZN(_07883_ ) );
AND3_X1 _15886_ ( .A1(_07536_ ), .A2(_07540_ ), .A3(_06961_ ), .ZN(_07884_ ) );
OR3_X1 _15887_ ( .A1(_07883_ ), .A2(_07003_ ), .A3(_07884_ ), .ZN(_07885_ ) );
NAND2_X1 _15888_ ( .A1(_07100_ ), .A2(_07004_ ), .ZN(_07886_ ) );
NAND3_X1 _15889_ ( .A1(_07877_ ), .A2(_07885_ ), .A3(_07886_ ), .ZN(_07887_ ) );
AND2_X1 _15890_ ( .A1(_07887_ ), .A2(_07467_ ), .ZN(_07888_ ) );
NOR3_X1 _15891_ ( .A1(_07102_ ), .A2(_06814_ ), .A3(_07045_ ), .ZN(_07889_ ) );
OAI21_X1 _15892_ ( .A(_07296_ ), .B1(_07005_ ), .B2(_02677_ ), .ZN(_07890_ ) );
OAI21_X1 _15893_ ( .A(_07890_ ), .B1(_04415_ ), .B2(_07198_ ), .ZN(_07891_ ) );
NOR3_X1 _15894_ ( .A1(_07114_ ), .A2(_07231_ ), .A3(_07519_ ), .ZN(_07892_ ) );
NOR4_X1 _15895_ ( .A1(_07888_ ), .A2(_07889_ ), .A3(_07891_ ), .A4(_07892_ ), .ZN(_07893_ ) );
AOI21_X1 _15896_ ( .A(_07153_ ), .B1(_07853_ ), .B2(_04415_ ), .ZN(_07894_ ) );
OAI21_X1 _15897_ ( .A(_07894_ ), .B1(_04415_ ), .B2(_07853_ ), .ZN(_07895_ ) );
AOI21_X1 _15898_ ( .A(_07056_ ), .B1(_07893_ ), .B2(_07895_ ), .ZN(_07896_ ) );
OR2_X1 _15899_ ( .A1(_04562_ ), .A2(_03973_ ), .ZN(_07897_ ) );
NAND3_X1 _15900_ ( .A1(_07897_ ), .A2(_07843_ ), .A3(_06782_ ), .ZN(_07898_ ) );
AOI22_X1 _15901_ ( .A1(_05130_ ), .A2(_07065_ ), .B1(\ID_EX_imm [4] ), .B2(_07066_ ), .ZN(_07899_ ) );
AOI21_X1 _15902_ ( .A(_06787_ ), .B1(_07898_ ), .B2(_07899_ ), .ZN(_07900_ ) );
NOR3_X1 _15903_ ( .A1(_07896_ ), .A2(_04756_ ), .A3(_07900_ ), .ZN(_07901_ ) );
OAI21_X1 _15904_ ( .A(_07236_ ), .B1(_05004_ ), .B2(_05129_ ), .ZN(_07902_ ) );
OAI21_X1 _15905_ ( .A(_07876_ ), .B1(_07901_ ), .B2(_07902_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
AND3_X1 _15906_ ( .A1(_06610_ ), .A2(_06611_ ), .A3(_06434_ ), .ZN(_07903_ ) );
INV_X1 _15907_ ( .A(_07903_ ), .ZN(_07904_ ) );
NAND4_X1 _15908_ ( .A1(_06910_ ), .A2(_06926_ ), .A3(_07193_ ), .A4(_07851_ ), .ZN(_07905_ ) );
AND3_X1 _15909_ ( .A1(_07783_ ), .A2(_07784_ ), .A3(_07001_ ), .ZN(_07906_ ) );
NOR2_X1 _15910_ ( .A1(_06997_ ), .A2(_06995_ ), .ZN(_07907_ ) );
NOR2_X1 _15911_ ( .A1(_06979_ ), .A2(_06998_ ), .ZN(_07908_ ) );
MUX2_X1 _15912_ ( .A(_07907_ ), .B(_07908_ ), .S(_07117_ ), .Z(_07909_ ) );
AOI211_X1 _15913_ ( .A(_07084_ ), .B(_07906_ ), .C1(_07023_ ), .C2(_07909_ ), .ZN(_07910_ ) );
AOI21_X1 _15914_ ( .A(_07007_ ), .B1(_07643_ ), .B2(_07647_ ), .ZN(_07911_ ) );
OAI21_X1 _15915_ ( .A(_07196_ ), .B1(_07910_ ), .B2(_07911_ ), .ZN(_07912_ ) );
OAI211_X1 _15916_ ( .A(_07912_ ), .B(_07467_ ), .C1(_06967_ ), .C2(_07190_ ), .ZN(_07913_ ) );
NOR2_X1 _15917_ ( .A1(_07022_ ), .A2(_04389_ ), .ZN(_07914_ ) );
OR3_X1 _15918_ ( .A1(_06802_ ), .A2(_04377_ ), .A3(_07914_ ), .ZN(_07915_ ) );
OAI21_X1 _15919_ ( .A(_04377_ ), .B1(_06802_ ), .B2(_07914_ ), .ZN(_07916_ ) );
NAND3_X1 _15920_ ( .A1(_07915_ ), .A2(_06861_ ), .A3(_07916_ ), .ZN(_07917_ ) );
NAND3_X1 _15921_ ( .A1(_07231_ ), .A2(_02829_ ), .A3(_07478_ ), .ZN(_07918_ ) );
NOR2_X1 _15922_ ( .A1(_07213_ ), .A2(_07519_ ), .ZN(_07919_ ) );
AOI221_X4 _15923_ ( .A(_07919_ ), .B1(_06808_ ), .B2(_04294_ ), .C1(_04377_ ), .C2(_04645_ ), .ZN(_07920_ ) );
AND4_X1 _15924_ ( .A1(_07913_ ), .A2(_07917_ ), .A3(_07918_ ), .A4(_07920_ ), .ZN(_07921_ ) );
AOI21_X1 _15925_ ( .A(_07056_ ), .B1(_07905_ ), .B2(_07921_ ), .ZN(_07922_ ) );
OR2_X1 _15926_ ( .A1(_04559_ ), .A2(_04021_ ), .ZN(_07923_ ) );
AND3_X1 _15927_ ( .A1(_07923_ ), .A2(_04557_ ), .A3(_04045_ ), .ZN(_07924_ ) );
AOI21_X1 _15928_ ( .A(_04045_ ), .B1(_07923_ ), .B2(_04557_ ), .ZN(_07925_ ) );
OR3_X1 _15929_ ( .A1(_07924_ ), .A2(_07925_ ), .A3(_07240_ ), .ZN(_07926_ ) );
AOI22_X1 _15930_ ( .A1(_05160_ ), .A2(_07065_ ), .B1(\ID_EX_imm [3] ), .B2(_07066_ ), .ZN(_07927_ ) );
AOI21_X1 _15931_ ( .A(_06787_ ), .B1(_07926_ ), .B2(_07927_ ), .ZN(_07928_ ) );
NOR3_X1 _15932_ ( .A1(_07922_ ), .A2(_04756_ ), .A3(_07928_ ), .ZN(_07929_ ) );
OAI21_X1 _15933_ ( .A(_07236_ ), .B1(_05004_ ), .B2(_05158_ ), .ZN(_07930_ ) );
OAI21_X1 _15934_ ( .A(_07904_ ), .B1(_07929_ ), .B2(_07930_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
NAND3_X1 _15935_ ( .A1(_05178_ ), .A2(_05180_ ), .A3(_06559_ ), .ZN(_07931_ ) );
NAND3_X1 _15936_ ( .A1(_04558_ ), .A2(_04021_ ), .A3(_04067_ ), .ZN(_07932_ ) );
NAND3_X1 _15937_ ( .A1(_07923_ ), .A2(_06781_ ), .A3(_07932_ ), .ZN(_07933_ ) );
AOI22_X1 _15938_ ( .A1(_05168_ ), .A2(_07446_ ), .B1(\ID_EX_imm [2] ), .B2(_07774_ ), .ZN(_07934_ ) );
AOI21_X1 _15939_ ( .A(_06786_ ), .B1(_07933_ ), .B2(_07934_ ), .ZN(_07935_ ) );
OR2_X1 _15940_ ( .A1(_07935_ ), .A2(_05319_ ), .ZN(_07936_ ) );
NOR2_X1 _15941_ ( .A1(_07248_ ), .A2(_07249_ ), .ZN(_07937_ ) );
NAND3_X1 _15942_ ( .A1(_07937_ ), .A2(_06926_ ), .A3(_07851_ ), .ZN(_07938_ ) );
NAND3_X1 _15943_ ( .A1(_06800_ ), .A2(_06801_ ), .A3(_06795_ ), .ZN(_07939_ ) );
NAND3_X1 _15944_ ( .A1(_06803_ ), .A2(_06861_ ), .A3(_07939_ ), .ZN(_07940_ ) );
NAND2_X1 _15945_ ( .A1(_07273_ ), .A2(_07432_ ), .ZN(_07941_ ) );
NAND3_X1 _15946_ ( .A1(_06921_ ), .A2(_02806_ ), .A3(_07478_ ), .ZN(_07942_ ) );
NAND3_X1 _15947_ ( .A1(_07940_ ), .A2(_07941_ ), .A3(_07942_ ), .ZN(_07943_ ) );
AND2_X1 _15948_ ( .A1(_04373_ ), .A2(_07011_ ), .ZN(_07944_ ) );
AOI21_X1 _15949_ ( .A(_07159_ ), .B1(_07023_ ), .B2(_04389_ ), .ZN(_07945_ ) );
NOR3_X1 _15950_ ( .A1(_07943_ ), .A2(_07944_ ), .A3(_07945_ ), .ZN(_07946_ ) );
OR3_X1 _15951_ ( .A1(_07679_ ), .A2(_07042_ ), .A3(_07683_ ), .ZN(_07947_ ) );
AOI21_X1 _15952_ ( .A(_07023_ ), .B1(_07819_ ), .B2(_07820_ ), .ZN(_07948_ ) );
NOR2_X1 _15953_ ( .A1(_07105_ ), .A2(_07109_ ), .ZN(_07949_ ) );
MUX2_X1 _15954_ ( .A(_07949_ ), .B(_07879_ ), .S(_07117_ ), .Z(_07950_ ) );
AOI21_X1 _15955_ ( .A(_07948_ ), .B1(_07023_ ), .B2(_07950_ ), .ZN(_07951_ ) );
OAI211_X1 _15956_ ( .A(_07947_ ), .B(_07102_ ), .C1(_07951_ ), .C2(_07231_ ), .ZN(_07952_ ) );
OAI211_X1 _15957_ ( .A(_07952_ ), .B(_07467_ ), .C1(_07102_ ), .C2(_07265_ ), .ZN(_07953_ ) );
NAND3_X1 _15958_ ( .A1(_07938_ ), .A2(_07946_ ), .A3(_07953_ ), .ZN(_07954_ ) );
AOI21_X1 _15959_ ( .A(_07936_ ), .B1(_07954_ ), .B2(_07057_ ), .ZN(_07955_ ) );
OAI21_X1 _15960_ ( .A(_07236_ ), .B1(_05004_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07956_ ) );
OAI21_X1 _15961_ ( .A(_07931_ ), .B1(_07955_ ), .B2(_07956_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
AND4_X1 _15962_ ( .A1(\mycsreg.CSReg[3][29] ), .A2(_04738_ ), .A3(_05193_ ), .A4(_04701_ ), .ZN(_07957_ ) );
AND4_X1 _15963_ ( .A1(\mepc [29] ), .A2(_03429_ ), .A3(_05193_ ), .A4(_04741_ ), .ZN(_07958_ ) );
NOR3_X1 _15964_ ( .A1(_04734_ ), .A2(_07957_ ), .A3(_07958_ ), .ZN(_07959_ ) );
AND3_X1 _15965_ ( .A1(_04839_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_04700_ ), .ZN(_07960_ ) );
NOR2_X1 _15966_ ( .A1(_04692_ ), .A2(_07960_ ), .ZN(_07961_ ) );
AOI22_X1 _15967_ ( .A1(_07959_ ), .A2(_07961_ ), .B1(_04731_ ), .B2(_04732_ ), .ZN(_07962_ ) );
AND3_X1 _15968_ ( .A1(_04731_ ), .A2(_04732_ ), .A3(\EX_LS_result_csreg_mem [29] ), .ZN(_07963_ ) );
OAI21_X1 _15969_ ( .A(_06559_ ), .B1(_07962_ ), .B2(_07963_ ), .ZN(_07964_ ) );
AND2_X1 _15970_ ( .A1(_07619_ ), .A2(_03632_ ), .ZN(_07965_ ) );
OR3_X1 _15971_ ( .A1(_07965_ ), .A2(_03654_ ), .A3(_04631_ ), .ZN(_07966_ ) );
OAI21_X1 _15972_ ( .A(_03654_ ), .B1(_07965_ ), .B2(_04631_ ), .ZN(_07967_ ) );
AND3_X1 _15973_ ( .A1(_07966_ ), .A2(_06781_ ), .A3(_07967_ ), .ZN(_07968_ ) );
OAI22_X1 _15974_ ( .A1(_04681_ ), .A2(_07305_ ), .B1(_03151_ ), .B2(_06770_ ), .ZN(_07969_ ) );
OAI21_X1 _15975_ ( .A(_06784_ ), .B1(_07968_ ), .B2(_07969_ ), .ZN(_07970_ ) );
NAND2_X1 _15976_ ( .A1(_07970_ ), .A2(_04661_ ), .ZN(_07971_ ) );
AOI21_X1 _15977_ ( .A(_04321_ ), .B1(_07568_ ), .B2(_07573_ ), .ZN(_07972_ ) );
OR3_X1 _15978_ ( .A1(_07972_ ), .A2(_04314_ ), .A3(_07578_ ), .ZN(_07973_ ) );
OAI21_X1 _15979_ ( .A(_04314_ ), .B1(_07972_ ), .B2(_07578_ ), .ZN(_07974_ ) );
NAND3_X1 _15980_ ( .A1(_07973_ ), .A2(_06862_ ), .A3(_07974_ ), .ZN(_07975_ ) );
NAND2_X1 _15981_ ( .A1(_04314_ ), .A2(_07011_ ), .ZN(_07976_ ) );
OAI21_X1 _15982_ ( .A(_07296_ ), .B1(_04313_ ), .B2(_03150_ ), .ZN(_07977_ ) );
NAND3_X1 _15983_ ( .A1(_04313_ ), .A2(_03150_ ), .A3(_07478_ ), .ZN(_07978_ ) );
AND3_X1 _15984_ ( .A1(_07976_ ), .A2(_07977_ ), .A3(_07978_ ), .ZN(_07979_ ) );
OR3_X1 _15985_ ( .A1(_06948_ ), .A2(_06960_ ), .A3(_07041_ ), .ZN(_07980_ ) );
OR3_X1 _15986_ ( .A1(_07116_ ), .A2(_07025_ ), .A3(_07036_ ), .ZN(_07981_ ) );
OR3_X1 _15987_ ( .A1(_07028_ ), .A2(_06976_ ), .A3(_07026_ ), .ZN(_07982_ ) );
NAND2_X1 _15988_ ( .A1(_07981_ ), .A2(_07982_ ), .ZN(_07983_ ) );
NOR2_X1 _15989_ ( .A1(_07035_ ), .A2(_07033_ ), .ZN(_07984_ ) );
NOR2_X1 _15990_ ( .A1(_07032_ ), .A2(_07018_ ), .ZN(_07985_ ) );
MUX2_X1 _15991_ ( .A(_07984_ ), .B(_07985_ ), .S(_06914_ ), .Z(_07986_ ) );
MUX2_X1 _15992_ ( .A(_07983_ ), .B(_07986_ ), .S(_07022_ ), .Z(_07987_ ) );
OAI211_X1 _15993_ ( .A(_07101_ ), .B(_07980_ ), .C1(_07987_ ), .C2(_06968_ ), .ZN(_07988_ ) );
OAI21_X1 _15994_ ( .A(_07005_ ), .B1(_07516_ ), .B2(_07517_ ), .ZN(_07989_ ) );
AOI21_X1 _15995_ ( .A(_06929_ ), .B1(_07988_ ), .B2(_07989_ ), .ZN(_07990_ ) );
NOR3_X1 _15996_ ( .A1(_07020_ ), .A2(_06963_ ), .A3(_06921_ ), .ZN(_07991_ ) );
AND3_X1 _15997_ ( .A1(_07991_ ), .A2(_07196_ ), .A3(_07013_ ), .ZN(_07992_ ) );
OAI211_X1 _15998_ ( .A(_06910_ ), .B(_06902_ ), .C1(_06923_ ), .C2(_06926_ ), .ZN(_07993_ ) );
NAND2_X1 _15999_ ( .A1(_07991_ ), .A2(_07196_ ), .ZN(_07994_ ) );
OAI211_X1 _16000_ ( .A(_07993_ ), .B(_07994_ ), .C1(_07312_ ), .C2(_07251_ ), .ZN(_07995_ ) );
AOI211_X1 _16001_ ( .A(_07990_ ), .B(_07992_ ), .C1(_07995_ ), .C2(_06866_ ), .ZN(_07996_ ) );
NAND3_X1 _16002_ ( .A1(_07975_ ), .A2(_07979_ ), .A3(_07996_ ), .ZN(_07997_ ) );
AOI21_X1 _16003_ ( .A(_07971_ ), .B1(_07058_ ), .B2(_07997_ ), .ZN(_07998_ ) );
OAI21_X1 _16004_ ( .A(_07236_ ), .B1(_04676_ ), .B2(_04720_ ), .ZN(_07999_ ) );
OAI21_X1 _16005_ ( .A(_07964_ ), .B1(_07998_ ), .B2(_07999_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
OAI21_X1 _16006_ ( .A(_06559_ ), .B1(_06642_ ), .B2(_06643_ ), .ZN(_08000_ ) );
NAND2_X1 _16007_ ( .A1(_04070_ ), .A2(_04094_ ), .ZN(_08001_ ) );
NAND3_X1 _16008_ ( .A1(_04558_ ), .A2(_06781_ ), .A3(_08001_ ), .ZN(_08002_ ) );
AOI22_X1 _16009_ ( .A1(_05187_ ), .A2(_07446_ ), .B1(\ID_EX_imm [1] ), .B2(_07774_ ), .ZN(_08003_ ) );
AOI21_X1 _16010_ ( .A(_06786_ ), .B1(_08002_ ), .B2(_08003_ ), .ZN(_08004_ ) );
OR2_X1 _16011_ ( .A1(_08004_ ), .A2(_05319_ ), .ZN(_08005_ ) );
NAND4_X1 _16012_ ( .A1(_07247_ ), .A2(_06918_ ), .A3(_06926_ ), .A4(_07851_ ), .ZN(_08006_ ) );
NAND3_X1 _16013_ ( .A1(_07714_ ), .A2(_07715_ ), .A3(_07231_ ), .ZN(_08007_ ) );
OAI21_X1 _16014_ ( .A(_06992_ ), .B1(_06994_ ), .B2(_06990_ ), .ZN(_08008_ ) );
OAI21_X1 _16015_ ( .A(_08008_ ), .B1(_07907_ ), .B2(_06992_ ), .ZN(_08009_ ) );
MUX2_X1 _16016_ ( .A(_07862_ ), .B(_08009_ ), .S(_07023_ ), .Z(_08010_ ) );
OAI211_X1 _16017_ ( .A(_07102_ ), .B(_08007_ ), .C1(_08010_ ), .C2(_07231_ ), .ZN(_08011_ ) );
OAI211_X1 _16018_ ( .A(_07467_ ), .B(_08011_ ), .C1(_07322_ ), .C2(_07102_ ), .ZN(_08012_ ) );
AND3_X1 _16019_ ( .A1(_07330_ ), .A2(_07008_ ), .A3(_07432_ ), .ZN(_08013_ ) );
NOR2_X1 _16020_ ( .A1(_04382_ ), .A2(_04383_ ), .ZN(_08014_ ) );
OAI21_X1 _16021_ ( .A(_06861_ ), .B1(_08014_ ), .B2(_06797_ ), .ZN(_08015_ ) );
NOR2_X1 _16022_ ( .A1(_08015_ ), .A2(_06799_ ), .ZN(_08016_ ) );
NOR3_X1 _16023_ ( .A1(_04382_ ), .A2(_04383_ ), .A3(_07198_ ), .ZN(_08017_ ) );
OAI22_X1 _16024_ ( .A1(_06801_ ), .A2(_07045_ ), .B1(_04383_ ), .B2(_07159_ ), .ZN(_08018_ ) );
NOR4_X1 _16025_ ( .A1(_08013_ ), .A2(_08016_ ), .A3(_08017_ ), .A4(_08018_ ), .ZN(_08019_ ) );
NAND3_X1 _16026_ ( .A1(_08006_ ), .A2(_08012_ ), .A3(_08019_ ), .ZN(_08020_ ) );
AOI21_X1 _16027_ ( .A(_08005_ ), .B1(_08020_ ), .B2(_07057_ ), .ZN(_08021_ ) );
OAI21_X1 _16028_ ( .A(_07236_ ), .B1(_04729_ ), .B2(\ID_EX_pc [1] ), .ZN(_08022_ ) );
OAI21_X1 _16029_ ( .A(_08000_ ), .B1(_08021_ ), .B2(_08022_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
AND3_X1 _16030_ ( .A1(_04289_ ), .A2(_07053_ ), .A3(_04299_ ), .ZN(_08023_ ) );
AND4_X1 _16031_ ( .A1(\ID_EX_typ [4] ), .A2(_03467_ ), .A3(\ID_EX_typ [3] ), .A4(_04649_ ), .ZN(_08024_ ) );
OR2_X1 _16032_ ( .A1(_08023_ ), .A2(_08024_ ), .ZN(_08025_ ) );
AND3_X1 _16033_ ( .A1(_04546_ ), .A2(_04552_ ), .A3(_08025_ ), .ZN(_08026_ ) );
OAI21_X1 _16034_ ( .A(_06780_ ), .B1(_04096_ ), .B2(_04094_ ), .ZN(_08027_ ) );
NAND3_X1 _16035_ ( .A1(_05225_ ), .A2(_06764_ ), .A3(_06763_ ), .ZN(_08028_ ) );
OAI211_X1 _16036_ ( .A(_08027_ ), .B(_08028_ ), .C1(_02763_ ), .C2(_06770_ ), .ZN(_08029_ ) );
OAI21_X1 _16037_ ( .A(_06784_ ), .B1(_08026_ ), .B2(_08029_ ), .ZN(_08030_ ) );
OAI21_X1 _16038_ ( .A(_04650_ ), .B1(_06869_ ), .B2(_06867_ ), .ZN(_08031_ ) );
AOI211_X1 _16039_ ( .A(_04548_ ), .B(_08031_ ), .C1(_04551_ ), .C2(_04310_ ), .ZN(_08032_ ) );
AND2_X1 _16040_ ( .A1(_04546_ ), .A2(_08032_ ), .ZN(_08033_ ) );
NAND4_X1 _16041_ ( .A1(_06888_ ), .A2(_04407_ ), .A3(_06886_ ), .A4(_06900_ ), .ZN(_08034_ ) );
OR2_X1 _16042_ ( .A1(_07365_ ), .A2(_06905_ ), .ZN(_08035_ ) );
AOI21_X1 _16043_ ( .A(_07108_ ), .B1(_06796_ ), .B2(_06916_ ), .ZN(_08036_ ) );
MUX2_X1 _16044_ ( .A(_07949_ ), .B(_08036_ ), .S(_06912_ ), .Z(_08037_ ) );
MUX2_X1 _16045_ ( .A(_07882_ ), .B(_08037_ ), .S(_06958_ ), .Z(_08038_ ) );
NAND2_X1 _16046_ ( .A1(_08038_ ), .A2(_07006_ ), .ZN(_08039_ ) );
NAND2_X1 _16047_ ( .A1(_07755_ ), .A2(_06961_ ), .ZN(_08040_ ) );
NAND3_X1 _16048_ ( .A1(_08039_ ), .A2(_06965_ ), .A3(_08040_ ), .ZN(_08041_ ) );
NAND2_X1 _16049_ ( .A1(_08035_ ), .A2(_08041_ ), .ZN(_00340_ ) );
AOI21_X1 _16050_ ( .A(_07071_ ), .B1(_08034_ ), .B2(_00340_ ), .ZN(_00341_ ) );
NAND3_X1 _16051_ ( .A1(_08035_ ), .A2(_07013_ ), .A3(_08041_ ), .ZN(_00342_ ) );
NAND3_X1 _16052_ ( .A1(_07042_ ), .A2(_07370_ ), .A3(_07431_ ), .ZN(_00343_ ) );
AND2_X1 _16053_ ( .A1(_06917_ ), .A2(_06796_ ), .ZN(_00344_ ) );
NOR3_X1 _16054_ ( .A1(_00344_ ), .A2(_06797_ ), .A3(_04646_ ), .ZN(_00345_ ) );
NOR3_X1 _16055_ ( .A1(_00344_ ), .A2(_06797_ ), .A3(_07152_ ), .ZN(_00346_ ) );
NOR3_X1 _16056_ ( .A1(_06917_ ), .A2(_06796_ ), .A3(_04291_ ), .ZN(_00347_ ) );
AOI21_X1 _16057_ ( .A(_07047_ ), .B1(_06917_ ), .B2(_06796_ ), .ZN(_00348_ ) );
NOR4_X1 _16058_ ( .A1(_00345_ ), .A2(_00346_ ), .A3(_00347_ ), .A4(_00348_ ), .ZN(_00349_ ) );
NAND3_X1 _16059_ ( .A1(_00342_ ), .A2(_00343_ ), .A3(_00349_ ), .ZN(_00350_ ) );
NOR3_X1 _16060_ ( .A1(_08033_ ), .A2(_00341_ ), .A3(_00350_ ), .ZN(_00351_ ) );
OAI21_X1 _16061_ ( .A(_08030_ ), .B1(_00351_ ), .B2(_07056_ ), .ZN(_00352_ ) );
MUX2_X1 _16062_ ( .A(\ID_EX_pc [0] ), .B(_00352_ ), .S(_02273_ ), .Z(_00353_ ) );
MUX2_X1 _16063_ ( .A(_06662_ ), .B(_00353_ ), .S(_06432_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
OAI21_X1 _16064_ ( .A(_06559_ ), .B1(_06669_ ), .B2(_06670_ ), .ZN(_00354_ ) );
NOR2_X1 _16065_ ( .A1(_07619_ ), .A2(_03632_ ), .ZN(_00355_ ) );
NOR3_X1 _16066_ ( .A1(_07965_ ), .A2(_00355_ ), .A3(_07240_ ), .ZN(_00356_ ) );
NOR2_X1 _16067_ ( .A1(_04989_ ), .A2(_07305_ ), .ZN(_00357_ ) );
AND3_X1 _16068_ ( .A1(_06768_ ), .A2(\ID_EX_imm [28] ), .A3(_06764_ ), .ZN(_00358_ ) );
NOR3_X1 _16069_ ( .A1(_00356_ ), .A2(_00357_ ), .A3(_00358_ ), .ZN(_00359_ ) );
OAI21_X1 _16070_ ( .A(_04661_ ), .B1(_00359_ ), .B2(_06787_ ), .ZN(_00360_ ) );
NOR2_X1 _16071_ ( .A1(_07972_ ), .A2(_07153_ ), .ZN(_00361_ ) );
OAI21_X1 _16072_ ( .A(_00361_ ), .B1(_04320_ ), .B2(_07575_ ), .ZN(_00362_ ) );
NAND2_X1 _16073_ ( .A1(_04320_ ), .A2(_07011_ ), .ZN(_00363_ ) );
OAI21_X1 _16074_ ( .A(_07296_ ), .B1(_04318_ ), .B2(_02388_ ), .ZN(_00364_ ) );
NAND3_X1 _16075_ ( .A1(_04318_ ), .A2(_02388_ ), .A3(_07478_ ), .ZN(_00365_ ) );
AND3_X1 _16076_ ( .A1(_00363_ ), .A2(_00364_ ), .A3(_00365_ ), .ZN(_00366_ ) );
NOR2_X1 _16077_ ( .A1(_07543_ ), .A2(_07003_ ), .ZN(_00367_ ) );
NOR3_X1 _16078_ ( .A1(_07588_ ), .A2(_07589_ ), .A3(_00367_ ), .ZN(_00368_ ) );
OAI21_X1 _16079_ ( .A(_07531_ ), .B1(_06908_ ), .B2(_06904_ ), .ZN(_00369_ ) );
AOI21_X1 _16080_ ( .A(_07072_ ), .B1(_00368_ ), .B2(_00369_ ), .ZN(_00370_ ) );
AOI21_X1 _16081_ ( .A(_00370_ ), .B1(_07149_ ), .B2(_00367_ ), .ZN(_00371_ ) );
OR3_X1 _16082_ ( .A1(_07088_ ), .A2(_06954_ ), .A3(_07086_ ), .ZN(_00372_ ) );
OAI211_X1 _16083_ ( .A(_00372_ ), .B(_06973_ ), .C1(_07595_ ), .C2(_07117_ ), .ZN(_00373_ ) );
OAI21_X1 _16084_ ( .A(_07117_ ), .B1(_07095_ ), .B2(_07093_ ), .ZN(_00374_ ) );
OAI21_X1 _16085_ ( .A(_06914_ ), .B1(_07092_ ), .B2(_07089_ ), .ZN(_00375_ ) );
AND2_X1 _16086_ ( .A1(_00374_ ), .A2(_00375_ ), .ZN(_00376_ ) );
OAI211_X1 _16087_ ( .A(_00373_ ), .B(_07007_ ), .C1(_07022_ ), .C2(_00376_ ), .ZN(_00377_ ) );
OAI21_X1 _16088_ ( .A(_07084_ ), .B1(_07123_ ), .B2(_07130_ ), .ZN(_00378_ ) );
NAND3_X1 _16089_ ( .A1(_00377_ ), .A2(_07101_ ), .A3(_00378_ ), .ZN(_00379_ ) );
AND2_X1 _16090_ ( .A1(_00379_ ), .A2(_04642_ ), .ZN(_00380_ ) );
OAI21_X1 _16091_ ( .A(_00380_ ), .B1(_07102_ ), .B2(_07546_ ), .ZN(_00381_ ) );
AND2_X1 _16092_ ( .A1(_00371_ ), .A2(_00381_ ), .ZN(_00382_ ) );
NAND3_X1 _16093_ ( .A1(_00362_ ), .A2(_00366_ ), .A3(_00382_ ), .ZN(_00383_ ) );
AOI21_X1 _16094_ ( .A(_00360_ ), .B1(_07058_ ), .B2(_00383_ ), .ZN(_00384_ ) );
OAI21_X1 _16095_ ( .A(_06432_ ), .B1(_04987_ ), .B2(_04720_ ), .ZN(_00385_ ) );
OAI21_X1 _16096_ ( .A(_00354_ ), .B1(_00384_ ), .B2(_00385_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
OR2_X1 _16097_ ( .A1(_06680_ ), .A2(_07349_ ), .ZN(_00386_ ) );
INV_X1 _16098_ ( .A(_03587_ ), .ZN(_00387_ ) );
NOR2_X1 _16099_ ( .A1(_07617_ ), .A2(_00387_ ), .ZN(_00388_ ) );
NOR3_X1 _16100_ ( .A1(_00388_ ), .A2(_04619_ ), .A3(_04621_ ), .ZN(_00389_ ) );
AOI21_X1 _16101_ ( .A(_00389_ ), .B1(_04537_ ), .B2(_03609_ ), .ZN(_00390_ ) );
AND2_X1 _16102_ ( .A1(_00390_ ), .A2(_03538_ ), .ZN(_00391_ ) );
OR3_X1 _16103_ ( .A1(_00391_ ), .A2(_03561_ ), .A3(_04624_ ), .ZN(_00392_ ) );
OAI21_X1 _16104_ ( .A(_03561_ ), .B1(_00391_ ), .B2(_04624_ ), .ZN(_00393_ ) );
NAND3_X1 _16105_ ( .A1(_00392_ ), .A2(_06781_ ), .A3(_00393_ ), .ZN(_00394_ ) );
AOI22_X1 _16106_ ( .A1(_05208_ ), .A2(_07446_ ), .B1(\ID_EX_imm [27] ), .B2(_07774_ ), .ZN(_00395_ ) );
AOI21_X1 _16107_ ( .A(_06786_ ), .B1(_00394_ ), .B2(_00395_ ), .ZN(_00396_ ) );
OR2_X1 _16108_ ( .A1(_00396_ ), .A2(_05319_ ), .ZN(_00397_ ) );
INV_X1 _16109_ ( .A(_04527_ ), .ZN(_00398_ ) );
INV_X1 _16110_ ( .A(_04534_ ), .ZN(_00399_ ) );
OR3_X1 _16111_ ( .A1(_07566_ ), .A2(_00398_ ), .A3(_00399_ ), .ZN(_00400_ ) );
AOI21_X1 _16112_ ( .A(_07569_ ), .B1(_00400_ ), .B2(_07571_ ), .ZN(_00401_ ) );
INV_X1 _16113_ ( .A(_00401_ ), .ZN(_00402_ ) );
INV_X1 _16114_ ( .A(_04512_ ), .ZN(_00403_ ) );
AOI21_X1 _16115_ ( .A(_04521_ ), .B1(_00402_ ), .B2(_00403_ ), .ZN(_00404_ ) );
NOR3_X1 _16116_ ( .A1(_00401_ ), .A2(_04542_ ), .A3(_04512_ ), .ZN(_00405_ ) );
OAI21_X1 _16117_ ( .A(_06862_ ), .B1(_00404_ ), .B2(_00405_ ), .ZN(_00406_ ) );
AOI21_X1 _16118_ ( .A(_07047_ ), .B1(_04517_ ), .B2(_04518_ ), .ZN(_00407_ ) );
NAND2_X1 _16119_ ( .A1(_07656_ ), .A2(_07657_ ), .ZN(_00408_ ) );
NOR2_X1 _16120_ ( .A1(_06905_ ), .A2(_06929_ ), .ZN(_00409_ ) );
OAI21_X1 _16121_ ( .A(_06949_ ), .B1(_06955_ ), .B2(_06956_ ), .ZN(_00410_ ) );
OAI21_X1 _16122_ ( .A(_06912_ ), .B1(_07028_ ), .B2(_07026_ ), .ZN(_00411_ ) );
AND2_X1 _16123_ ( .A1(_00410_ ), .A2(_00411_ ), .ZN(_00412_ ) );
OAI21_X1 _16124_ ( .A(_06934_ ), .B1(_07025_ ), .B2(_07036_ ), .ZN(_00413_ ) );
OAI21_X1 _16125_ ( .A(_06945_ ), .B1(_07035_ ), .B2(_07033_ ), .ZN(_00414_ ) );
AND2_X1 _16126_ ( .A1(_00413_ ), .A2(_00414_ ), .ZN(_00415_ ) );
MUX2_X1 _16127_ ( .A(_00412_ ), .B(_00415_ ), .S(_06932_ ), .Z(_00416_ ) );
MUX2_X1 _16128_ ( .A(_07222_ ), .B(_00416_ ), .S(_07042_ ), .Z(_00417_ ) );
AOI221_X4 _16129_ ( .A(_00407_ ), .B1(_00408_ ), .B2(_00409_ ), .C1(_00417_ ), .C2(_07432_ ), .ZN(_00418_ ) );
NOR2_X1 _16130_ ( .A1(_07189_ ), .A2(_07379_ ), .ZN(_00419_ ) );
AOI221_X4 _16131_ ( .A(_07589_ ), .B1(_06965_ ), .B2(_00419_ ), .C1(_06903_ ), .C2(_06909_ ), .ZN(_00420_ ) );
OAI211_X1 _16132_ ( .A(_06910_ ), .B(_07193_ ), .C1(_06902_ ), .C2(_06908_ ), .ZN(_00421_ ) );
AOI21_X1 _16133_ ( .A(_07072_ ), .B1(_00420_ ), .B2(_00421_ ), .ZN(_00422_ ) );
NOR3_X1 _16134_ ( .A1(_04519_ ), .A2(_04520_ ), .A3(_07198_ ), .ZN(_00423_ ) );
NOR3_X1 _16135_ ( .A1(_04517_ ), .A2(_04518_ ), .A3(_07045_ ), .ZN(_00424_ ) );
AND3_X1 _16136_ ( .A1(_00419_ ), .A2(_07196_ ), .A3(_07013_ ), .ZN(_00425_ ) );
NOR4_X1 _16137_ ( .A1(_00422_ ), .A2(_00423_ ), .A3(_00424_ ), .A4(_00425_ ), .ZN(_00426_ ) );
NAND3_X1 _16138_ ( .A1(_00406_ ), .A2(_00418_ ), .A3(_00426_ ), .ZN(_00427_ ) );
AOI21_X1 _16139_ ( .A(_00397_ ), .B1(_07058_ ), .B2(_00427_ ), .ZN(_00428_ ) );
NAND2_X1 _16140_ ( .A1(_05211_ ), .A2(_04755_ ), .ZN(_00429_ ) );
NAND2_X1 _16141_ ( .A1(_00429_ ), .A2(_07441_ ), .ZN(_00430_ ) );
OAI21_X1 _16142_ ( .A(_00386_ ), .B1(_00428_ ), .B2(_00430_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
OAI21_X1 _16143_ ( .A(_06559_ ), .B1(_06692_ ), .B2(_06693_ ), .ZN(_00431_ ) );
AOI21_X1 _16144_ ( .A(_07240_ ), .B1(_00390_ ), .B2(_03538_ ), .ZN(_00432_ ) );
OAI21_X1 _16145_ ( .A(_00432_ ), .B1(_03538_ ), .B2(_00390_ ), .ZN(_00433_ ) );
AOI22_X1 _16146_ ( .A1(_05242_ ), .A2(_06766_ ), .B1(\ID_EX_imm [26] ), .B2(_07774_ ), .ZN(_00434_ ) );
AOI21_X1 _16147_ ( .A(_06786_ ), .B1(_00433_ ), .B2(_00434_ ), .ZN(_00435_ ) );
OR2_X1 _16148_ ( .A1(_00435_ ), .A2(_05319_ ), .ZN(_00436_ ) );
NAND3_X1 _16149_ ( .A1(_00400_ ), .A2(_07569_ ), .A3(_07571_ ), .ZN(_00437_ ) );
NAND3_X1 _16150_ ( .A1(_00402_ ), .A2(_06862_ ), .A3(_00437_ ), .ZN(_00438_ ) );
NOR2_X1 _16151_ ( .A1(_07264_ ), .A2(_06962_ ), .ZN(_00439_ ) );
AND3_X1 _16152_ ( .A1(_00439_ ), .A2(_06967_ ), .A3(_07149_ ), .ZN(_00440_ ) );
NOR3_X1 _16153_ ( .A1(_04512_ ), .A2(_04513_ ), .A3(_07198_ ), .ZN(_00441_ ) );
NOR3_X1 _16154_ ( .A1(_04511_ ), .A2(_03126_ ), .A3(_07045_ ), .ZN(_00442_ ) );
AOI21_X1 _16155_ ( .A(_07159_ ), .B1(_04511_ ), .B2(_03126_ ), .ZN(_00443_ ) );
NOR4_X1 _16156_ ( .A1(_00440_ ), .A2(_00441_ ), .A3(_00442_ ), .A4(_00443_ ), .ZN(_00444_ ) );
AND2_X1 _16157_ ( .A1(_00439_ ), .A2(_06966_ ), .ZN(_00445_ ) );
AOI211_X1 _16158_ ( .A(_07589_ ), .B(_00445_ ), .C1(_06904_ ), .C2(_06909_ ), .ZN(_00446_ ) );
OAI221_X1 _16159_ ( .A(_07247_ ), .B1(_07117_ ), .B2(_06917_ ), .C1(_06904_ ), .C2(_06908_ ), .ZN(_00447_ ) );
AOI21_X1 _16160_ ( .A(_07072_ ), .B1(_00446_ ), .B2(_00447_ ), .ZN(_00448_ ) );
NAND2_X1 _16161_ ( .A1(_07691_ ), .A2(_07692_ ), .ZN(_00449_ ) );
AND2_X1 _16162_ ( .A1(_00449_ ), .A2(_00409_ ), .ZN(_00450_ ) );
AOI21_X1 _16163_ ( .A(_06921_ ), .B1(_07597_ ), .B2(_07598_ ), .ZN(_00451_ ) );
AND3_X1 _16164_ ( .A1(_07602_ ), .A2(_07603_ ), .A3(_07001_ ), .ZN(_00452_ ) );
OR3_X1 _16165_ ( .A1(_00451_ ), .A2(_00452_ ), .A3(_06963_ ), .ZN(_00453_ ) );
NAND2_X1 _16166_ ( .A1(_07281_ ), .A2(_07231_ ), .ZN(_00454_ ) );
AND3_X1 _16167_ ( .A1(_00453_ ), .A2(_07432_ ), .A3(_00454_ ), .ZN(_00455_ ) );
NOR3_X1 _16168_ ( .A1(_00448_ ), .A2(_00450_ ), .A3(_00455_ ), .ZN(_00456_ ) );
NAND3_X1 _16169_ ( .A1(_00438_ ), .A2(_00444_ ), .A3(_00456_ ), .ZN(_00457_ ) );
AOI21_X1 _16170_ ( .A(_00436_ ), .B1(_07058_ ), .B2(_00457_ ), .ZN(_00458_ ) );
OAI21_X1 _16171_ ( .A(_06432_ ), .B1(_05240_ ), .B2(_04720_ ), .ZN(_00459_ ) );
OAI21_X1 _16172_ ( .A(_00431_ ), .B1(_00458_ ), .B2(_00459_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
INV_X1 _16173_ ( .A(_05275_ ), .ZN(_00460_ ) );
OAI211_X1 _16174_ ( .A(_00460_ ), .B(_06457_ ), .C1(_06542_ ), .C2(_05272_ ), .ZN(_00461_ ) );
OR3_X1 _16175_ ( .A1(_00388_ ), .A2(_04619_ ), .A3(_03610_ ), .ZN(_00462_ ) );
OAI21_X1 _16176_ ( .A(_03610_ ), .B1(_00388_ ), .B2(_04619_ ), .ZN(_00463_ ) );
NAND3_X1 _16177_ ( .A1(_00462_ ), .A2(_06781_ ), .A3(_00463_ ), .ZN(_00464_ ) );
AOI22_X1 _16178_ ( .A1(_05258_ ), .A2(_06766_ ), .B1(\ID_EX_imm [25] ), .B2(_07774_ ), .ZN(_00465_ ) );
AOI21_X1 _16179_ ( .A(_06786_ ), .B1(_00464_ ), .B2(_00465_ ), .ZN(_00466_ ) );
OR2_X1 _16180_ ( .A1(_00466_ ), .A2(_05319_ ), .ZN(_00467_ ) );
AOI21_X1 _16181_ ( .A(_00399_ ), .B1(_07557_ ), .B2(_07565_ ), .ZN(_00468_ ) );
OR3_X1 _16182_ ( .A1(_00468_ ), .A2(_04527_ ), .A3(_04532_ ), .ZN(_00469_ ) );
OAI21_X1 _16183_ ( .A(_04527_ ), .B1(_00468_ ), .B2(_04532_ ), .ZN(_00470_ ) );
AND3_X1 _16184_ ( .A1(_00469_ ), .A2(_06861_ ), .A3(_00470_ ), .ZN(_00471_ ) );
INV_X1 _16185_ ( .A(_07590_ ), .ZN(_00472_ ) );
NOR2_X1 _16186_ ( .A1(_07320_ ), .A2(_06962_ ), .ZN(_00473_ ) );
AOI21_X1 _16187_ ( .A(_00472_ ), .B1(_06967_ ), .B2(_00473_ ), .ZN(_00474_ ) );
AND3_X1 _16188_ ( .A1(_07247_ ), .A2(_06918_ ), .A3(_06924_ ), .ZN(_00475_ ) );
OAI21_X1 _16189_ ( .A(_00475_ ), .B1(_06908_ ), .B2(_06904_ ), .ZN(_00476_ ) );
AOI21_X1 _16190_ ( .A(_07072_ ), .B1(_00474_ ), .B2(_00476_ ), .ZN(_00477_ ) );
AND2_X1 _16191_ ( .A1(_07335_ ), .A2(_07379_ ), .ZN(_00478_ ) );
NAND2_X1 _16192_ ( .A1(_07983_ ), .A2(_06932_ ), .ZN(_00479_ ) );
NAND3_X1 _16193_ ( .A1(_06953_ ), .A2(_06957_ ), .A3(_06920_ ), .ZN(_00480_ ) );
AOI21_X1 _16194_ ( .A(_07379_ ), .B1(_00479_ ), .B2(_00480_ ), .ZN(_00481_ ) );
OAI21_X1 _16195_ ( .A(_07431_ ), .B1(_00478_ ), .B2(_00481_ ), .ZN(_00482_ ) );
AOI22_X1 _16196_ ( .A1(_07570_ ), .A2(_04294_ ), .B1(_04539_ ), .B2(_06857_ ), .ZN(_00483_ ) );
OAI211_X1 _16197_ ( .A(_00482_ ), .B(_00483_ ), .C1(_00398_ ), .C2(_04646_ ), .ZN(_00484_ ) );
AND2_X1 _16198_ ( .A1(_07729_ ), .A2(_00409_ ), .ZN(_00485_ ) );
AND3_X1 _16199_ ( .A1(_00473_ ), .A2(_06965_ ), .A3(_07013_ ), .ZN(_00486_ ) );
OR3_X1 _16200_ ( .A1(_00484_ ), .A2(_00485_ ), .A3(_00486_ ), .ZN(_00487_ ) );
OR3_X1 _16201_ ( .A1(_00471_ ), .A2(_00477_ ), .A3(_00487_ ), .ZN(_00488_ ) );
AOI21_X1 _16202_ ( .A(_00467_ ), .B1(_07058_ ), .B2(_00488_ ), .ZN(_00489_ ) );
NAND2_X1 _16203_ ( .A1(_05265_ ), .A2(_04755_ ), .ZN(_00490_ ) );
NAND2_X1 _16204_ ( .A1(_00490_ ), .A2(_07441_ ), .ZN(_00491_ ) );
OAI21_X1 _16205_ ( .A(_00461_ ), .B1(_00489_ ), .B2(_00491_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _16206_ ( .A1(_05289_ ), .A2(_06435_ ), .ZN(_00492_ ) );
OAI21_X1 _16207_ ( .A(_06781_ ), .B1(_07617_ ), .B2(_00387_ ), .ZN(_00493_ ) );
AOI21_X1 _16208_ ( .A(_00493_ ), .B1(_00387_ ), .B2(_07617_ ), .ZN(_00494_ ) );
AND2_X1 _16209_ ( .A1(_05291_ ), .A2(_07065_ ), .ZN(_00495_ ) );
AND3_X1 _16210_ ( .A1(_06768_ ), .A2(\ID_EX_imm [24] ), .A3(_06764_ ), .ZN(_00496_ ) );
NOR3_X1 _16211_ ( .A1(_00494_ ), .A2(_00495_ ), .A3(_00496_ ), .ZN(_00497_ ) );
OAI21_X1 _16212_ ( .A(_04661_ ), .B1(_00497_ ), .B2(_06787_ ), .ZN(_00498_ ) );
OAI21_X1 _16213_ ( .A(_06861_ ), .B1(_07566_ ), .B2(_00399_ ), .ZN(_00499_ ) );
AOI21_X1 _16214_ ( .A(_00499_ ), .B1(_00399_ ), .B2(_07566_ ), .ZN(_00500_ ) );
OR3_X1 _16215_ ( .A1(_04532_ ), .A2(_04533_ ), .A3(_07198_ ), .ZN(_00501_ ) );
OR3_X1 _16216_ ( .A1(_04530_ ), .A2(_04531_ ), .A3(_07045_ ), .ZN(_00502_ ) );
OR2_X1 _16217_ ( .A1(_04533_ ), .A2(_07159_ ), .ZN(_00503_ ) );
NAND3_X1 _16218_ ( .A1(_00501_ ), .A2(_00502_ ), .A3(_00503_ ), .ZN(_00504_ ) );
NAND4_X1 _16219_ ( .A1(_06888_ ), .A2(_07747_ ), .A3(_06900_ ), .A4(_06908_ ), .ZN(_00505_ ) );
NOR2_X1 _16220_ ( .A1(_07364_ ), .A2(_06962_ ), .ZN(_00506_ ) );
NAND2_X1 _16221_ ( .A1(_00506_ ), .A2(_06966_ ), .ZN(_00507_ ) );
NAND2_X1 _16222_ ( .A1(_00505_ ), .A2(_00507_ ), .ZN(_00508_ ) );
OAI21_X1 _16223_ ( .A(_06865_ ), .B1(_07588_ ), .B2(_00508_ ), .ZN(_00509_ ) );
NAND3_X1 _16224_ ( .A1(_07763_ ), .A2(_07764_ ), .A3(_00409_ ), .ZN(_00510_ ) );
NAND2_X1 _16225_ ( .A1(_07375_ ), .A2(_06968_ ), .ZN(_00511_ ) );
AOI21_X1 _16226_ ( .A(_07022_ ), .B1(_07120_ ), .B2(_07122_ ), .ZN(_00512_ ) );
AOI21_X1 _16227_ ( .A(_06921_ ), .B1(_00374_ ), .B2(_00375_ ), .ZN(_00513_ ) );
OAI21_X1 _16228_ ( .A(_07042_ ), .B1(_00512_ ), .B2(_00513_ ), .ZN(_00514_ ) );
NAND3_X1 _16229_ ( .A1(_00511_ ), .A2(_07432_ ), .A3(_00514_ ), .ZN(_00515_ ) );
NAND3_X1 _16230_ ( .A1(_00506_ ), .A2(_07196_ ), .A3(_07013_ ), .ZN(_00516_ ) );
NAND4_X1 _16231_ ( .A1(_00509_ ), .A2(_00510_ ), .A3(_00515_ ), .A4(_00516_ ), .ZN(_00517_ ) );
OR3_X1 _16232_ ( .A1(_00500_ ), .A2(_00504_ ), .A3(_00517_ ), .ZN(_00518_ ) );
AOI21_X1 _16233_ ( .A(_00498_ ), .B1(_07058_ ), .B2(_00518_ ), .ZN(_00519_ ) );
OAI21_X1 _16234_ ( .A(_06432_ ), .B1(_05290_ ), .B2(_04720_ ), .ZN(_00520_ ) );
OAI21_X1 _16235_ ( .A(_00492_ ), .B1(_00519_ ), .B2(_00520_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
OR3_X1 _16236_ ( .A1(_05313_ ), .A2(_05315_ ), .A3(_06422_ ), .ZN(_00521_ ) );
NOR4_X1 _16237_ ( .A1(_06774_ ), .A2(_04605_ ), .A3(_04606_ ), .A4(_06775_ ), .ZN(_00522_ ) );
OAI21_X1 _16238_ ( .A(_03753_ ), .B1(_00522_ ), .B2(_04609_ ), .ZN(_00523_ ) );
INV_X1 _16239_ ( .A(_04612_ ), .ZN(_00524_ ) );
AND2_X1 _16240_ ( .A1(_00523_ ), .A2(_00524_ ), .ZN(_00525_ ) );
XNOR2_X1 _16241_ ( .A(_00525_ ), .B(_03731_ ), .ZN(_00526_ ) );
NAND2_X1 _16242_ ( .A1(_00526_ ), .A2(_06782_ ), .ZN(_00527_ ) );
AOI22_X1 _16243_ ( .A1(_05302_ ), .A2(_06766_ ), .B1(\ID_EX_imm [23] ), .B2(_07774_ ), .ZN(_00528_ ) );
AOI21_X1 _16244_ ( .A(_06786_ ), .B1(_00527_ ), .B2(_00528_ ), .ZN(_00529_ ) );
OR2_X1 _16245_ ( .A1(_00529_ ), .A2(_05319_ ), .ZN(_00530_ ) );
OAI21_X1 _16246_ ( .A(_07556_ ), .B1(_06842_ ), .B2(_06851_ ), .ZN(_00531_ ) );
AND2_X1 _16247_ ( .A1(_00531_ ), .A2(_07560_ ), .ZN(_00532_ ) );
OR2_X1 _16248_ ( .A1(_00532_ ), .A2(_07561_ ), .ZN(_00533_ ) );
AND3_X1 _16249_ ( .A1(_00533_ ), .A2(_07558_ ), .A3(_07563_ ), .ZN(_00534_ ) );
AOI21_X1 _16250_ ( .A(_07558_ ), .B1(_00533_ ), .B2(_07563_ ), .ZN(_00535_ ) );
NOR3_X1 _16251_ ( .A1(_00534_ ), .A2(_00535_ ), .A3(_07153_ ), .ZN(_00536_ ) );
NAND3_X1 _16252_ ( .A1(_07781_ ), .A2(_07196_ ), .A3(_07149_ ), .ZN(_00537_ ) );
OAI21_X1 _16253_ ( .A(_00537_ ), .B1(_04450_ ), .B2(_07159_ ), .ZN(_00538_ ) );
AND2_X1 _16254_ ( .A1(_07781_ ), .A2(_06905_ ), .ZN(_00539_ ) );
AOI211_X1 _16255_ ( .A(_07589_ ), .B(_00539_ ), .C1(_06903_ ), .C2(_06909_ ), .ZN(_00540_ ) );
NOR2_X1 _16256_ ( .A1(_00540_ ), .A2(_07071_ ), .ZN(_00541_ ) );
OR3_X1 _16257_ ( .A1(_07426_ ), .A2(_06965_ ), .A3(_07379_ ), .ZN(_00542_ ) );
NAND3_X1 _16258_ ( .A1(_07428_ ), .A2(_06962_ ), .A3(_07429_ ), .ZN(_00543_ ) );
AOI21_X1 _16259_ ( .A(_06919_ ), .B1(_00410_ ), .B2(_00411_ ), .ZN(_00544_ ) );
AOI21_X1 _16260_ ( .A(_06930_ ), .B1(_07215_ ), .B2(_07216_ ), .ZN(_00545_ ) );
NOR2_X1 _16261_ ( .A1(_00544_ ), .A2(_00545_ ), .ZN(_00546_ ) );
OAI211_X1 _16262_ ( .A(_00543_ ), .B(_06965_ ), .C1(_00546_ ), .C2(_07084_ ), .ZN(_00547_ ) );
AOI21_X1 _16263_ ( .A(_06929_ ), .B1(_00542_ ), .B2(_00547_ ), .ZN(_00548_ ) );
OR3_X1 _16264_ ( .A1(_04448_ ), .A2(_03703_ ), .A3(_04291_ ), .ZN(_00549_ ) );
OAI21_X1 _16265_ ( .A(_00549_ ), .B1(_07558_ ), .B2(_04646_ ), .ZN(_00550_ ) );
OR3_X1 _16266_ ( .A1(_00541_ ), .A2(_00548_ ), .A3(_00550_ ), .ZN(_00551_ ) );
OR3_X1 _16267_ ( .A1(_00536_ ), .A2(_00538_ ), .A3(_00551_ ), .ZN(_00552_ ) );
AOI21_X1 _16268_ ( .A(_00530_ ), .B1(_07058_ ), .B2(_00552_ ), .ZN(_00553_ ) );
NAND2_X1 _16269_ ( .A1(_05305_ ), .A2(_04755_ ), .ZN(_00554_ ) );
NAND2_X1 _16270_ ( .A1(_00554_ ), .A2(_06488_ ), .ZN(_00555_ ) );
OAI21_X1 _16271_ ( .A(_00521_ ), .B1(_00553_ ), .B2(_00555_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
OR2_X1 _16272_ ( .A1(_06733_ ), .A2(_07349_ ), .ZN(_00556_ ) );
OR3_X1 _16273_ ( .A1(_00522_ ), .A2(_03753_ ), .A3(_04609_ ), .ZN(_00557_ ) );
NAND3_X1 _16274_ ( .A1(_00557_ ), .A2(_06781_ ), .A3(_00523_ ), .ZN(_00558_ ) );
AOI22_X1 _16275_ ( .A1(_05324_ ), .A2(_06766_ ), .B1(\ID_EX_imm [22] ), .B2(_07774_ ), .ZN(_00559_ ) );
AOI21_X1 _16276_ ( .A(_06786_ ), .B1(_00558_ ), .B2(_00559_ ), .ZN(_00560_ ) );
OR2_X1 _16277_ ( .A1(_00560_ ), .A2(_05319_ ), .ZN(_00561_ ) );
OR3_X1 _16278_ ( .A1(_07474_ ), .A2(_07007_ ), .A3(_07475_ ), .ZN(_00562_ ) );
NAND3_X1 _16279_ ( .A1(_07601_ ), .A2(_07605_ ), .A3(_07042_ ), .ZN(_00563_ ) );
AOI21_X1 _16280_ ( .A(_07004_ ), .B1(_00562_ ), .B2(_00563_ ), .ZN(_00564_ ) );
NOR3_X1 _16281_ ( .A1(_07472_ ), .A2(_07101_ ), .A3(_06968_ ), .ZN(_00565_ ) );
OAI21_X1 _16282_ ( .A(_04642_ ), .B1(_00564_ ), .B2(_00565_ ), .ZN(_00566_ ) );
AND3_X1 _16283_ ( .A1(_07455_ ), .A2(_06925_ ), .A3(_06908_ ), .ZN(_00567_ ) );
NAND2_X1 _16284_ ( .A1(_07825_ ), .A2(_07826_ ), .ZN(_00568_ ) );
AND2_X1 _16285_ ( .A1(_00568_ ), .A2(_06905_ ), .ZN(_00569_ ) );
OR3_X1 _16286_ ( .A1(_07588_ ), .A2(_00567_ ), .A3(_00569_ ), .ZN(_00570_ ) );
AOI22_X1 _16287_ ( .A1(_00570_ ), .A2(_06866_ ), .B1(_07149_ ), .B2(_00569_ ), .ZN(_00571_ ) );
NAND3_X1 _16288_ ( .A1(_04501_ ), .A2(_02411_ ), .A3(_07478_ ), .ZN(_00572_ ) );
AOI21_X1 _16289_ ( .A(_07047_ ), .B1(_04454_ ), .B2(_04500_ ), .ZN(_00573_ ) );
AOI21_X1 _16290_ ( .A(_00573_ ), .B1(_04455_ ), .B2(_07011_ ), .ZN(_00574_ ) );
AND4_X1 _16291_ ( .A1(_00566_ ), .A2(_00571_ ), .A3(_00572_ ), .A4(_00574_ ), .ZN(_00575_ ) );
XNOR2_X1 _16292_ ( .A(_00532_ ), .B(_07561_ ), .ZN(_00576_ ) );
OAI21_X1 _16293_ ( .A(_00575_ ), .B1(_07153_ ), .B2(_00576_ ), .ZN(_00577_ ) );
AOI21_X1 _16294_ ( .A(_00561_ ), .B1(_07058_ ), .B2(_00577_ ), .ZN(_00578_ ) );
NAND2_X1 _16295_ ( .A1(_05322_ ), .A2(_04755_ ), .ZN(_00579_ ) );
NAND2_X1 _16296_ ( .A1(_00579_ ), .A2(_06488_ ), .ZN(_00580_ ) );
OAI21_X1 _16297_ ( .A(_00556_ ), .B1(_00578_ ), .B2(_00580_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NOR2_X1 _16298_ ( .A1(_07622_ ), .A2(_04637_ ), .ZN(_00581_ ) );
AOI21_X1 _16299_ ( .A(_07239_ ), .B1(_00581_ ), .B2(_04634_ ), .ZN(_00582_ ) );
OAI21_X1 _16300_ ( .A(_00582_ ), .B1(_04634_ ), .B2(_00581_ ), .ZN(_00583_ ) );
AOI22_X1 _16301_ ( .A1(_05369_ ), .A2(_06766_ ), .B1(\ID_EX_imm [31] ), .B2(_06769_ ), .ZN(_00584_ ) );
AOI21_X1 _16302_ ( .A(_06786_ ), .B1(_00583_ ), .B2(_00584_ ), .ZN(_00585_ ) );
AND3_X1 _16303_ ( .A1(_07080_ ), .A2(_04307_ ), .A3(_04306_ ), .ZN(_00586_ ) );
OR3_X2 _16304_ ( .A1(_07582_ ), .A2(_04305_ ), .A3(_00586_ ), .ZN(_00587_ ) );
OAI21_X1 _16305_ ( .A(_04305_ ), .B1(_07582_ ), .B2(_00586_ ), .ZN(_00588_ ) );
NAND3_X1 _16306_ ( .A1(_00587_ ), .A2(_06861_ ), .A3(_00588_ ), .ZN(_00589_ ) );
NAND3_X1 _16307_ ( .A1(_07427_ ), .A2(_07430_ ), .A3(_00409_ ), .ZN(_00590_ ) );
OAI21_X1 _16308_ ( .A(_04294_ ), .B1(_06869_ ), .B2(_03185_ ), .ZN(_00591_ ) );
NAND3_X1 _16309_ ( .A1(_06886_ ), .A2(_03185_ ), .A3(_07013_ ), .ZN(_00592_ ) );
AND3_X1 _16310_ ( .A1(_06869_ ), .A2(_03185_ ), .A3(_06857_ ), .ZN(_00593_ ) );
AOI21_X1 _16311_ ( .A(_00593_ ), .B1(_04305_ ), .B2(_04645_ ), .ZN(_00594_ ) );
NAND4_X1 _16312_ ( .A1(_00590_ ), .A2(_00591_ ), .A3(_00592_ ), .A4(_00594_ ), .ZN(_00595_ ) );
AOI21_X1 _16313_ ( .A(_07017_ ), .B1(_06867_ ), .B2(_06915_ ), .ZN(_00596_ ) );
MUX2_X1 _16314_ ( .A(_07985_ ), .B(_00596_ ), .S(_06945_ ), .Z(_00597_ ) );
MUX2_X1 _16315_ ( .A(_00415_ ), .B(_00597_ ), .S(_06930_ ), .Z(_00598_ ) );
MUX2_X1 _16316_ ( .A(_00546_ ), .B(_00598_ ), .S(_07006_ ), .Z(_00599_ ) );
AND2_X1 _16317_ ( .A1(_06886_ ), .A2(_03185_ ), .ZN(_00600_ ) );
OR2_X1 _16318_ ( .A1(_06903_ ), .A2(_00600_ ), .ZN(_00601_ ) );
AOI221_X4 _16319_ ( .A(_00595_ ), .B1(_07431_ ), .B2(_00599_ ), .C1(_00601_ ), .C2(_06865_ ), .ZN(_00602_ ) );
AOI21_X1 _16320_ ( .A(_07056_ ), .B1(_00589_ ), .B2(_00602_ ), .ZN(_00603_ ) );
OAI21_X1 _16321_ ( .A(_02273_ ), .B1(_00585_ ), .B2(_00603_ ), .ZN(_00604_ ) );
OAI21_X1 _16322_ ( .A(_00604_ ), .B1(_04661_ ), .B2(_05363_ ), .ZN(_00605_ ) );
MUX2_X2 _16323_ ( .A(_06758_ ), .B(_00605_ ), .S(_06432_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_D ) );
NAND2_X1 _16324_ ( .A1(_05671_ ), .A2(IDU_valid_EXU ), .ZN(_00606_ ) );
OAI21_X1 _16325_ ( .A(_00606_ ), .B1(_05584_ ), .B2(_05637_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16326_ ( .A1(_05583_ ), .A2(_05637_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16327_ ( .A1(_05583_ ), .A2(_05637_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16328_ ( .A(_05632_ ), .ZN(_00607_ ) );
NOR4_X1 _16329_ ( .A1(_05583_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_05431_ ), .A4(_00607_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_NOR__A_Y ) );
AOI21_X1 _16330_ ( .A(_06159_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16331_ ( .A(_00606_ ), .B1(_00607_ ), .B2(_05671_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16332_ ( .A1(_05632_ ), .A2(_05671_ ), .B1(_02186_ ), .B2(_02260_ ), .ZN(_00608_ ) );
INV_X1 _16333_ ( .A(loaduse_clear ), .ZN(_00609_ ) );
AOI221_X4 _16334_ ( .A(_00608_ ), .B1(\myidu.state [2] ), .B2(_00609_ ), .C1(_05583_ ), .C2(_06159_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _16335_ ( .A1(_05572_ ), .A2(_05578_ ), .ZN(_00610_ ) );
NOR3_X1 _16336_ ( .A1(_00610_ ), .A2(_05573_ ), .A3(_05551_ ), .ZN(_00611_ ) );
NAND2_X1 _16337_ ( .A1(_05698_ ), .A2(_05699_ ), .ZN(_00612_ ) );
NOR2_X1 _16338_ ( .A1(_05530_ ), .A2(_00612_ ), .ZN(_00613_ ) );
BUF_X2 _16339_ ( .A(_00613_ ), .Z(_00614_ ) );
AND3_X1 _16340_ ( .A1(_00611_ ), .A2(_05657_ ), .A3(_00614_ ), .ZN(_00615_ ) );
OAI211_X1 _16341_ ( .A(_05580_ ), .B(_05696_ ), .C1(_05692_ ), .C2(_00615_ ), .ZN(_00616_ ) );
AND2_X1 _16342_ ( .A1(_05634_ ), .A2(_05417_ ), .ZN(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ) );
AOI22_X1 _16343_ ( .A1(_00616_ ), .A2(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .B1(loaduse_clear ), .B2(_00244_ ), .ZN(_00617_ ) );
NAND3_X1 _16344_ ( .A1(_05493_ ), .A2(IDU_valid_EXU ), .A3(_06203_ ), .ZN(_00618_ ) );
NAND2_X1 _16345_ ( .A1(_00617_ ), .A2(_00618_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16346_ ( .A(_02261_ ), .B(_05493_ ), .C1(_05632_ ), .C2(_05671_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
NAND4_X1 _16347_ ( .A1(_05632_ ), .A2(IDU_ready_IFU ), .A3(_05417_ ), .A4(_05692_ ), .ZN(_00619_ ) );
NAND3_X1 _16348_ ( .A1(_05680_ ), .A2(_05682_ ), .A3(_05683_ ), .ZN(_00620_ ) );
OR2_X1 _16349_ ( .A1(_05674_ ), .A2(_00620_ ), .ZN(_00621_ ) );
AOI21_X1 _16350_ ( .A(_00619_ ), .B1(_00615_ ), .B2(_00621_ ), .ZN(_00622_ ) );
AND3_X1 _16351_ ( .A1(_05493_ ), .A2(\myidu.state [2] ), .A3(_00609_ ), .ZN(_00623_ ) );
OR2_X1 _16352_ ( .A1(_00622_ ), .A2(_00623_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
AND4_X1 _16353_ ( .A1(\ID_EX_typ [7] ), .A2(_02267_ ), .A3(_06218_ ), .A4(IDU_valid_EXU ), .ZN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16354_ ( .A1(_05629_ ), .A2(IDU_ready_IFU ), .ZN(_00624_ ) );
OAI21_X1 _16355_ ( .A(_01634_ ), .B1(_05629_ ), .B2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00625_ ) );
INV_X1 _16356_ ( .A(\myifu.state [0] ), .ZN(_00626_ ) );
AOI211_X1 _16357_ ( .A(_00624_ ), .B(_00625_ ), .C1(_00626_ ), .C2(_05629_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
OR3_X1 _16358_ ( .A1(_02101_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06277_ ), .ZN(_00627_ ) );
OAI21_X1 _16359_ ( .A(_00627_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06278_ ), .ZN(_00628_ ) );
MUX2_X1 _16360_ ( .A(\io_master_rdata [31] ), .B(_00628_ ), .S(_02207_ ), .Z(_00629_ ) );
AND2_X1 _16361_ ( .A1(_00629_ ), .A2(_06231_ ), .ZN(\myifu.data_in [31] ) );
OR4_X1 _16362_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [22] ), .A3(\io_master_araddr [20] ), .A4(\io_master_araddr [23] ), .ZN(_00630_ ) );
OR2_X1 _16363_ ( .A1(\io_master_araddr [18] ), .A2(\io_master_araddr [17] ), .ZN(_00631_ ) );
OR4_X4 _16364_ ( .A1(\io_master_araddr [19] ), .A2(_00630_ ), .A3(\io_master_araddr [16] ), .A4(_00631_ ), .ZN(_00632_ ) );
OR4_X2 _16365_ ( .A1(\io_master_araddr [28] ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [29] ), .A4(\io_master_araddr [31] ), .ZN(_00633_ ) );
NAND2_X1 _16366_ ( .A1(_02178_ ), .A2(\io_master_araddr [25] ), .ZN(_00634_ ) );
OR4_X4 _16367_ ( .A1(\io_master_araddr [27] ), .A2(_00633_ ), .A3(\io_master_araddr [26] ), .A4(_00634_ ), .ZN(_00635_ ) );
NOR2_X4 _16368_ ( .A1(_00632_ ), .A2(_00635_ ), .ZN(_00636_ ) );
BUF_X4 _16369_ ( .A(_00636_ ), .Z(_00637_ ) );
CLKBUF_X2 _16370_ ( .A(_06277_ ), .Z(_00638_ ) );
OR3_X1 _16371_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00639_ ) );
OAI211_X1 _16372_ ( .A(_00637_ ), .B(_00639_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00640_ ) );
OAI21_X1 _16373_ ( .A(_00640_ ), .B1(\io_master_rdata [30] ), .B2(_00637_ ), .ZN(_00641_ ) );
NOR2_X1 _16374_ ( .A1(_00641_ ), .A2(_06249_ ), .ZN(\myifu.data_in [30] ) );
BUF_X2 _16375_ ( .A(_00637_ ), .Z(_00642_ ) );
CLKBUF_X2 _16376_ ( .A(_00642_ ), .Z(_00643_ ) );
OR2_X1 _16377_ ( .A1(_00643_ ), .A2(\io_master_rdata [21] ), .ZN(_00644_ ) );
BUF_X4 _16378_ ( .A(_00637_ ), .Z(_00645_ ) );
BUF_X4 _16379_ ( .A(_00645_ ), .Z(_00646_ ) );
BUF_X4 _16380_ ( .A(_00646_ ), .Z(_00647_ ) );
CLKBUF_X2 _16381_ ( .A(_00638_ ), .Z(_00648_ ) );
OR3_X1 _16382_ ( .A1(_02104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00649_ ) );
OAI211_X1 _16383_ ( .A(_00647_ ), .B(_00649_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00650_ ) );
AND3_X1 _16384_ ( .A1(_00644_ ), .A2(_00650_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [21] ) );
OR2_X1 _16385_ ( .A1(_00645_ ), .A2(\io_master_rdata [20] ), .ZN(_00651_ ) );
CLKBUF_X2 _16386_ ( .A(_00638_ ), .Z(_00652_ ) );
OR3_X1 _16387_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00653_ ) );
OAI211_X1 _16388_ ( .A(_00642_ ), .B(_00653_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00654_ ) );
AND3_X1 _16389_ ( .A1(_00651_ ), .A2(_00654_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [20] ) );
OR2_X1 _16390_ ( .A1(_00643_ ), .A2(\io_master_rdata [19] ), .ZN(_00655_ ) );
OR3_X1 _16391_ ( .A1(_02104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00656_ ) );
OAI211_X1 _16392_ ( .A(_00647_ ), .B(_00656_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00657_ ) );
AND3_X1 _16393_ ( .A1(_00655_ ), .A2(_00657_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [19] ) );
OR2_X1 _16394_ ( .A1(_00642_ ), .A2(\io_master_rdata [18] ), .ZN(_00658_ ) );
OR3_X1 _16395_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00659_ ) );
OAI211_X1 _16396_ ( .A(_00646_ ), .B(_00659_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06280_ ), .ZN(_00660_ ) );
CLKBUF_X2 _16397_ ( .A(_06231_ ), .Z(_00661_ ) );
AND3_X1 _16398_ ( .A1(_00658_ ), .A2(_00660_ ), .A3(_00661_ ), .ZN(\myifu.data_in [18] ) );
OR2_X1 _16399_ ( .A1(_00645_ ), .A2(\io_master_rdata [17] ), .ZN(_00662_ ) );
OR3_X1 _16400_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00663_ ) );
OAI211_X1 _16401_ ( .A(_00642_ ), .B(_00663_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00664_ ) );
AND3_X1 _16402_ ( .A1(_00662_ ), .A2(_00664_ ), .A3(_00661_ ), .ZN(\myifu.data_in [17] ) );
OR2_X1 _16403_ ( .A1(_00645_ ), .A2(\io_master_rdata [16] ), .ZN(_00665_ ) );
OR3_X1 _16404_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00666_ ) );
OAI211_X1 _16405_ ( .A(_00645_ ), .B(_00666_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00667_ ) );
AND3_X1 _16406_ ( .A1(_00665_ ), .A2(_00667_ ), .A3(_00661_ ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16407_ ( .A1(_02101_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06277_ ), .ZN(_00668_ ) );
OAI211_X1 _16408_ ( .A(_00636_ ), .B(_00668_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06278_ ), .ZN(_00669_ ) );
OAI21_X2 _16409_ ( .A(_00669_ ), .B1(\io_master_rdata [15] ), .B2(_00636_ ), .ZN(_00670_ ) );
BUF_X4 _16410_ ( .A(_06282_ ), .Z(_00671_ ) );
NOR2_X1 _16411_ ( .A1(_00670_ ), .A2(_00671_ ), .ZN(\myifu.data_in [15] ) );
OR2_X1 _16412_ ( .A1(_00637_ ), .A2(\io_master_rdata [14] ), .ZN(_00672_ ) );
OR3_X1 _16413_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00673_ ) );
OAI211_X1 _16414_ ( .A(_00645_ ), .B(_00673_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00674_ ) );
AND3_X1 _16415_ ( .A1(_00672_ ), .A2(_00674_ ), .A3(_06231_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16416_ ( .A1(_00642_ ), .A2(\io_master_rdata [13] ), .ZN(_00675_ ) );
OR3_X1 _16417_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00676_ ) );
OAI211_X1 _16418_ ( .A(_00646_ ), .B(_00676_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06280_ ), .ZN(_00677_ ) );
AND3_X1 _16419_ ( .A1(_00675_ ), .A2(_00677_ ), .A3(_00661_ ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _16420_ ( .A1(_00643_ ), .A2(\io_master_rdata [12] ), .ZN(_00678_ ) );
OR3_X1 _16421_ ( .A1(_02104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00679_ ) );
OAI211_X1 _16422_ ( .A(_00643_ ), .B(_00679_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00680_ ) );
AND3_X1 _16423_ ( .A1(_00678_ ), .A2(_00680_ ), .A3(_00661_ ), .ZN(\myifu.data_in [12] ) );
OR2_X1 _16424_ ( .A1(_00645_ ), .A2(\io_master_rdata [29] ), .ZN(_00681_ ) );
OR3_X1 _16425_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00682_ ) );
OAI211_X1 _16426_ ( .A(_00642_ ), .B(_00682_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06280_ ), .ZN(_00683_ ) );
AND3_X1 _16427_ ( .A1(_00681_ ), .A2(_00683_ ), .A3(_06231_ ), .ZN(\myifu.data_in [29] ) );
MUX2_X1 _16428_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06280_ ), .Z(_00684_ ) );
NAND2_X1 _16429_ ( .A1(_00647_ ), .A2(_00684_ ), .ZN(_00685_ ) );
INV_X1 _16430_ ( .A(\io_master_rdata [11] ), .ZN(_00686_ ) );
OAI21_X1 _16431_ ( .A(_00686_ ), .B1(_00632_ ), .B2(_00635_ ), .ZN(_00687_ ) );
AND3_X1 _16432_ ( .A1(_00685_ ), .A2(_06231_ ), .A3(_00687_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16433_ ( .A1(_00643_ ), .A2(\io_master_rdata [10] ), .ZN(_00688_ ) );
OR3_X1 _16434_ ( .A1(_02104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00689_ ) );
OAI211_X1 _16435_ ( .A(_00643_ ), .B(_00689_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00690_ ) );
AND3_X1 _16436_ ( .A1(_00688_ ), .A2(_00690_ ), .A3(_06231_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16437_ ( .A1(_00646_ ), .A2(\io_master_rdata [9] ), .ZN(_00691_ ) );
OR3_X1 _16438_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00692_ ) );
OAI211_X1 _16439_ ( .A(_00646_ ), .B(_00692_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06280_ ), .ZN(_00693_ ) );
AND3_X1 _16440_ ( .A1(_00691_ ), .A2(_00693_ ), .A3(_00661_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16441_ ( .A1(_00643_ ), .A2(\io_master_rdata [8] ), .ZN(_00694_ ) );
OR3_X1 _16442_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00695_ ) );
OAI211_X1 _16443_ ( .A(_00643_ ), .B(_00695_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00696_ ) );
AND3_X1 _16444_ ( .A1(_00694_ ), .A2(_00696_ ), .A3(_00661_ ), .ZN(\myifu.data_in [8] ) );
OR3_X1 _16445_ ( .A1(_02101_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00697_ ) );
OAI211_X1 _16446_ ( .A(_00636_ ), .B(_00697_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06278_ ), .ZN(_00698_ ) );
OAI21_X1 _16447_ ( .A(_00698_ ), .B1(\io_master_rdata [7] ), .B2(_00637_ ), .ZN(_00699_ ) );
NOR2_X1 _16448_ ( .A1(_00699_ ), .A2(_00671_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16449_ ( .A1(_02101_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00700_ ) );
OAI211_X1 _16450_ ( .A(_00636_ ), .B(_00700_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06278_ ), .ZN(_00701_ ) );
OAI21_X1 _16451_ ( .A(_00701_ ), .B1(\io_master_rdata [6] ), .B2(_00637_ ), .ZN(_00702_ ) );
NOR2_X1 _16452_ ( .A1(_00702_ ), .A2(_00671_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16453_ ( .A1(_02104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00703_ ) );
OAI211_X1 _16454_ ( .A(_00647_ ), .B(_00703_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00704_ ) );
OAI21_X1 _16455_ ( .A(_00704_ ), .B1(\io_master_rdata [5] ), .B2(_00647_ ), .ZN(_00705_ ) );
NOR2_X1 _16456_ ( .A1(_00705_ ), .A2(_00671_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16457_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00706_ ) );
OAI211_X1 _16458_ ( .A(_00646_ ), .B(_00706_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06280_ ), .ZN(_00707_ ) );
OAI21_X1 _16459_ ( .A(_00707_ ), .B1(\io_master_rdata [4] ), .B2(_00646_ ), .ZN(_00708_ ) );
NOR2_X1 _16460_ ( .A1(_00708_ ), .A2(_00671_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16461_ ( .A1(_02104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00709_ ) );
OAI211_X1 _16462_ ( .A(_00647_ ), .B(_00709_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00710_ ) );
OAI21_X1 _16463_ ( .A(_00710_ ), .B1(\io_master_rdata [3] ), .B2(_00647_ ), .ZN(_00711_ ) );
NOR2_X1 _16464_ ( .A1(_00711_ ), .A2(_00671_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16465_ ( .A1(_02104_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00712_ ) );
OAI211_X1 _16466_ ( .A(_00647_ ), .B(_00712_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00713_ ) );
OAI21_X1 _16467_ ( .A(_00713_ ), .B1(\io_master_rdata [2] ), .B2(_00647_ ), .ZN(_00714_ ) );
NOR2_X1 _16468_ ( .A1(_00714_ ), .A2(_00671_ ), .ZN(\myifu.data_in [2] ) );
OR2_X1 _16469_ ( .A1(_00645_ ), .A2(\io_master_rdata [28] ), .ZN(_00715_ ) );
OR3_X1 _16470_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00716_ ) );
OAI211_X1 _16471_ ( .A(_00642_ ), .B(_00716_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00717_ ) );
AND3_X1 _16472_ ( .A1(_00715_ ), .A2(_00717_ ), .A3(_00661_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16473_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00718_ ) );
OAI211_X1 _16474_ ( .A(_00646_ ), .B(_00718_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06280_ ), .ZN(_00719_ ) );
OAI21_X1 _16475_ ( .A(_00719_ ), .B1(\io_master_rdata [1] ), .B2(_00646_ ), .ZN(_00720_ ) );
NOR2_X1 _16476_ ( .A1(_00720_ ), .A2(_00671_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16477_ ( .A1(_02103_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00652_ ), .ZN(_00721_ ) );
OAI211_X1 _16478_ ( .A(_00642_ ), .B(_00721_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(_06280_ ), .ZN(_00722_ ) );
OAI21_X1 _16479_ ( .A(_00722_ ), .B1(\io_master_rdata [0] ), .B2(_00646_ ), .ZN(_00723_ ) );
NOR2_X1 _16480_ ( .A1(_00723_ ), .A2(_00671_ ), .ZN(\myifu.data_in [0] ) );
MUX2_X1 _16481_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_06280_ ), .Z(_00724_ ) );
NAND2_X1 _16482_ ( .A1(_00647_ ), .A2(_00724_ ), .ZN(_00725_ ) );
INV_X1 _16483_ ( .A(\io_master_rdata [27] ), .ZN(_00726_ ) );
OAI21_X1 _16484_ ( .A(_00726_ ), .B1(_00632_ ), .B2(_00635_ ), .ZN(_00727_ ) );
AND3_X1 _16485_ ( .A1(_00725_ ), .A2(\io_master_arburst [0] ), .A3(_00727_ ), .ZN(\myifu.data_in [27] ) );
OR2_X1 _16486_ ( .A1(_00645_ ), .A2(\io_master_rdata [26] ), .ZN(_00728_ ) );
OR3_X1 _16487_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00729_ ) );
OAI211_X1 _16488_ ( .A(_00642_ ), .B(_00729_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00730_ ) );
AND3_X1 _16489_ ( .A1(_00728_ ), .A2(_00730_ ), .A3(_00661_ ), .ZN(\myifu.data_in [26] ) );
OR2_X1 _16490_ ( .A1(_00643_ ), .A2(\io_master_rdata [25] ), .ZN(_00731_ ) );
OR3_X1 _16491_ ( .A1(_02103_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00648_ ), .ZN(_00732_ ) );
OAI211_X1 _16492_ ( .A(_00643_ ), .B(_00732_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00733_ ) );
AND3_X1 _16493_ ( .A1(_00731_ ), .A2(_00733_ ), .A3(_00661_ ), .ZN(\myifu.data_in [25] ) );
OR2_X1 _16494_ ( .A1(_00645_ ), .A2(\io_master_rdata [24] ), .ZN(_00734_ ) );
OR3_X1 _16495_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00652_ ), .ZN(_00735_ ) );
OAI211_X1 _16496_ ( .A(_00642_ ), .B(_00735_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00736_ ) );
AND3_X1 _16497_ ( .A1(_00734_ ), .A2(_00736_ ), .A3(_06231_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16498_ ( .A1(_02101_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00737_ ) );
OAI211_X2 _16499_ ( .A(_00636_ ), .B(_00737_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06278_ ), .ZN(_00738_ ) );
OAI21_X2 _16500_ ( .A(_00738_ ), .B1(\io_master_rdata [23] ), .B2(_00637_ ), .ZN(_00739_ ) );
NOR2_X1 _16501_ ( .A1(_00739_ ), .A2(_00671_ ), .ZN(\myifu.data_in [23] ) );
OR3_X1 _16502_ ( .A1(_02102_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00638_ ), .ZN(_00740_ ) );
OAI211_X1 _16503_ ( .A(_00637_ ), .B(_00740_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06279_ ), .ZN(_00741_ ) );
OAI21_X2 _16504_ ( .A(_00741_ ), .B1(\io_master_rdata [22] ), .B2(_00637_ ), .ZN(_00742_ ) );
NOR2_X1 _16505_ ( .A1(_00742_ ), .A2(_06250_ ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16506_ ( .A(_00278_ ), .ZN(_00743_ ) );
NAND2_X1 _16507_ ( .A1(_00743_ ), .A2(_02144_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16508_ ( .A1(_06078_ ), .A2(fanout_net_12 ), .ZN(_00744_ ) );
INV_X1 _16509_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00745_ ) );
OAI21_X1 _16510_ ( .A(_02144_ ), .B1(_00744_ ), .B2(_00745_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16511_ ( .A1(_06087_ ), .A2(fanout_net_16 ), .ZN(_00746_ ) );
OAI21_X1 _16512_ ( .A(_02144_ ), .B1(_00746_ ), .B2(_00745_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16513_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .ZN(_00747_ ) );
OAI21_X1 _16514_ ( .A(_02144_ ), .B1(_00747_ ), .B2(_00745_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
OAI21_X1 _16515_ ( .A(\IF_ID_inst [8] ), .B1(_05530_ ), .B2(_00612_ ), .ZN(_00748_ ) );
AND2_X1 _16516_ ( .A1(_00613_ ), .A2(_05727_ ), .ZN(_00749_ ) );
NAND2_X1 _16517_ ( .A1(_05570_ ), .A2(_05717_ ), .ZN(_00750_ ) );
AND4_X1 _16518_ ( .A1(_05414_ ), .A2(_05460_ ), .A3(_05675_ ), .A4(_00750_ ), .ZN(_00751_ ) );
OAI211_X1 _16519_ ( .A(_05709_ ), .B(_05710_ ), .C1(_05575_ ), .C2(_05576_ ), .ZN(_00752_ ) );
INV_X1 _16520_ ( .A(_00752_ ), .ZN(_00753_ ) );
AND4_X1 _16521_ ( .A1(_05505_ ), .A2(_00753_ ), .A3(_05574_ ), .A4(_05712_ ), .ZN(_00754_ ) );
NAND3_X1 _16522_ ( .A1(_00749_ ), .A2(_00751_ ), .A3(_00754_ ), .ZN(_00755_ ) );
AND2_X1 _16523_ ( .A1(_00755_ ), .A2(_05505_ ), .ZN(_00756_ ) );
OAI221_X1 _16524_ ( .A(_00748_ ), .B1(_05639_ ), .B2(_05415_ ), .C1(_00756_ ), .C2(_05422_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
NOR2_X1 _16525_ ( .A1(_05673_ ), .A2(_05562_ ), .ZN(_00757_ ) );
NOR2_X1 _16526_ ( .A1(_00757_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_00758_ ) );
AND3_X1 _16527_ ( .A1(_05762_ ), .A2(_05478_ ), .A3(\IF_ID_inst [31] ), .ZN(_00759_ ) );
NOR2_X1 _16528_ ( .A1(_00758_ ), .A2(_00759_ ), .ZN(_00760_ ) );
BUF_X4 _16529_ ( .A(_00760_ ), .Z(_00761_ ) );
OAI21_X1 _16530_ ( .A(_00761_ ), .B1(_00749_ ), .B2(_05416_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
OR2_X1 _16531_ ( .A1(_00613_ ), .A2(_05416_ ), .ZN(_00762_ ) );
BUF_X4 _16532_ ( .A(_00762_ ), .Z(_00763_ ) );
BUF_X4 _16533_ ( .A(_00763_ ), .Z(_00764_ ) );
BUF_X4 _16534_ ( .A(_05727_ ), .Z(_00765_ ) );
OAI211_X1 _16535_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05421_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16536_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05422_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16537_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05425_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
BUF_X4 _16538_ ( .A(_00757_ ), .Z(_00766_ ) );
OAI221_X1 _16539_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00766_ ), .C1(_05518_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI221_X1 _16540_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00766_ ), .C1(_05519_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI221_X1 _16541_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00766_ ), .C1(_05520_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16542_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00757_ ), .C1(_05639_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _16543_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00757_ ), .C1(_05437_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16544_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00757_ ), .C1(_05534_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16545_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00757_ ), .C1(_05470_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16546_ ( .A(_00763_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B2(_00757_ ), .C1(_05435_ ), .C2(_05693_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16547_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05426_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
AOI22_X1 _16548_ ( .A1(_05530_ ), .A2(\IF_ID_inst [31] ), .B1(_00612_ ), .B2(\IF_ID_inst [7] ), .ZN(_00767_ ) );
OAI221_X1 _16549_ ( .A(_00767_ ), .B1(_05425_ ), .B2(_05505_ ), .C1(_00766_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16550_ ( .A(_05857_ ), .ZN(_00768_ ) );
OAI221_X1 _16551_ ( .A(_00768_ ), .B1(_05421_ ), .B2(_00614_ ), .C1(_00766_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
INV_X1 _16552_ ( .A(_05853_ ), .ZN(_00769_ ) );
OAI221_X1 _16553_ ( .A(_00769_ ), .B1(_05426_ ), .B2(_00614_ ), .C1(_00766_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16554_ ( .A(_05820_ ), .ZN(_00770_ ) );
OAI221_X1 _16555_ ( .A(_00770_ ), .B1(_05427_ ), .B2(_00614_ ), .C1(_00766_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
OAI221_X1 _16556_ ( .A(_05767_ ), .B1(_05428_ ), .B2(_00614_ ), .C1(_00766_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16557_ ( .A(_05807_ ), .ZN(_00771_ ) );
OAI221_X1 _16558_ ( .A(_00771_ ), .B1(_05429_ ), .B2(_00614_ ), .C1(_00766_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16559_ ( .A(_05804_ ), .ZN(_00772_ ) );
OAI221_X1 _16560_ ( .A(_00772_ ), .B1(_05430_ ), .B2(_00614_ ), .C1(_00766_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16561_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05427_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16562_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05428_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16563_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05429_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16564_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05430_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16565_ ( .A(_00761_ ), .B(_00764_ ), .C1(_05432_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16566_ ( .A(_00760_ ), .B(_00764_ ), .C1(_05433_ ), .C2(_00765_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16567_ ( .A(_00760_ ), .B(_00763_ ), .C1(_05434_ ), .C2(_05727_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16568_ ( .A(\IF_ID_inst [19] ), .B1(_05409_ ), .B2(_05413_ ), .ZN(_00773_ ) );
OAI221_X1 _16569_ ( .A(_00773_ ), .B1(_05442_ ), .B2(_00614_ ), .C1(_00756_ ), .C2(_05432_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16570_ ( .A(\IF_ID_inst [18] ), .B1(_05409_ ), .B2(_05413_ ), .ZN(_00774_ ) );
OAI221_X1 _16571_ ( .A(_00774_ ), .B1(_05443_ ), .B2(_00614_ ), .C1(_00756_ ), .C2(_05433_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16572_ ( .A(\IF_ID_inst [17] ), .B1(_05409_ ), .B2(_05413_ ), .ZN(_00775_ ) );
OAI221_X1 _16573_ ( .A(_00775_ ), .B1(_05444_ ), .B2(_00614_ ), .C1(_00756_ ), .C2(_05434_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16574_ ( .A1(_05474_ ), .A2(_05436_ ), .ZN(_00776_ ) );
OAI221_X1 _16575_ ( .A(_00776_ ), .B1(_05437_ ), .B2(_05414_ ), .C1(_00755_ ), .C2(_05425_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
BUF_X4 _16576_ ( .A(_06153_ ), .Z(_00777_ ) );
AOI21_X1 _16577_ ( .A(\IF_ID_pc [1] ), .B1(_06156_ ), .B2(\IF_ID_pc [2] ), .ZN(_00778_ ) );
INV_X1 _16578_ ( .A(_00778_ ), .ZN(_00779_ ) );
OAI21_X1 _16579_ ( .A(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .B1(_06156_ ), .B2(\IF_ID_pc [2] ), .ZN(_00780_ ) );
NOR2_X2 _16580_ ( .A1(_00779_ ), .A2(_00780_ ), .ZN(_00781_ ) );
BUF_X4 _16581_ ( .A(_00781_ ), .Z(_00782_ ) );
NAND2_X1 _16582_ ( .A1(_00694_ ), .A2(_00696_ ), .ZN(_00783_ ) );
OAI211_X1 _16583_ ( .A(_00777_ ), .B(_00782_ ), .C1(_06249_ ), .C2(_00783_ ), .ZN(_00784_ ) );
AND2_X4 _16584_ ( .A1(_06153_ ), .A2(_00781_ ), .ZN(_00785_ ) );
BUF_X4 _16585_ ( .A(_00785_ ), .Z(_00786_ ) );
BUF_X4 _16586_ ( .A(_00786_ ), .Z(_00787_ ) );
OAI211_X1 _16587_ ( .A(_00784_ ), .B(\myifu.state [2] ), .C1(_00787_ ), .C2(_05777_ ), .ZN(_00788_ ) );
AND3_X1 _16588_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00789_ ) );
AND3_X1 _16589_ ( .A1(_06077_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00790_ ) );
AOI211_X1 _16590_ ( .A(_00789_ ), .B(_00790_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_06230_ ), .ZN(_00791_ ) );
NAND2_X2 _16591_ ( .A1(_00745_ ), .A2(\IF_ID_pc [2] ), .ZN(_00792_ ) );
BUF_X2 _16592_ ( .A(_00792_ ), .Z(_00793_ ) );
NAND2_X2 _16593_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00794_ ) );
BUF_X4 _16594_ ( .A(_00794_ ), .Z(_00795_ ) );
NAND3_X1 _16595_ ( .A1(_06087_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00796_ ) );
NAND4_X1 _16596_ ( .A1(_00791_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00796_ ), .ZN(_00797_ ) );
NOR2_X1 _16597_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00798_ ) );
BUF_X4 _16598_ ( .A(_00798_ ), .Z(_00799_ ) );
BUF_X4 _16599_ ( .A(_00799_ ), .Z(_00800_ ) );
BUF_X2 _16600_ ( .A(_05793_ ), .Z(_00801_ ) );
BUF_X4 _16601_ ( .A(_00801_ ), .Z(_00802_ ) );
NAND3_X1 _16602_ ( .A1(_00802_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00803_ ) );
NAND3_X1 _16603_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00804_ ) );
AND2_X1 _16604_ ( .A1(_00803_ ), .A2(_00804_ ), .ZN(_00805_ ) );
NAND2_X1 _16605_ ( .A1(_00792_ ), .A2(_00794_ ), .ZN(_00806_ ) );
BUF_X2 _16606_ ( .A(_00806_ ), .Z(_00807_ ) );
BUF_X4 _16607_ ( .A(_06085_ ), .Z(_00808_ ) );
BUF_X4 _16608_ ( .A(_00808_ ), .Z(_00809_ ) );
NAND3_X1 _16609_ ( .A1(_00809_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00810_ ) );
BUF_X4 _16610_ ( .A(_06086_ ), .Z(_00811_ ) );
NAND3_X1 _16611_ ( .A1(_06078_ ), .A2(_00811_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00812_ ) );
NAND4_X1 _16612_ ( .A1(_00805_ ), .A2(_00807_ ), .A3(_00810_ ), .A4(_00812_ ), .ZN(_00813_ ) );
NAND3_X1 _16613_ ( .A1(_00797_ ), .A2(_00800_ ), .A3(_00813_ ), .ZN(_00814_ ) );
NAND2_X1 _16614_ ( .A1(_00788_ ), .A2(_00814_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16615_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00815_ ) );
AND3_X1 _16616_ ( .A1(_00801_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00816_ ) );
BUF_X4 _16617_ ( .A(_06229_ ), .Z(_00817_ ) );
AOI211_X1 _16618_ ( .A(_00815_ ), .B(_00816_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00817_ ), .ZN(_00818_ ) );
BUF_X4 _16619_ ( .A(_00792_ ), .Z(_00819_ ) );
BUF_X4 _16620_ ( .A(_00794_ ), .Z(_00820_ ) );
NAND3_X1 _16621_ ( .A1(_00811_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00821_ ) );
NAND4_X1 _16622_ ( .A1(_00818_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_00821_ ), .ZN(_00822_ ) );
BUF_X4 _16623_ ( .A(_06076_ ), .Z(_00823_ ) );
NAND3_X1 _16624_ ( .A1(_00823_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00824_ ) );
NAND3_X1 _16625_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00825_ ) );
AND2_X1 _16626_ ( .A1(_00824_ ), .A2(_00825_ ), .ZN(_00826_ ) );
BUF_X4 _16627_ ( .A(_00806_ ), .Z(_00827_ ) );
BUF_X4 _16628_ ( .A(_06086_ ), .Z(_00828_ ) );
NAND3_X1 _16629_ ( .A1(_00828_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00829_ ) );
BUF_X4 _16630_ ( .A(_06077_ ), .Z(_00830_ ) );
NAND3_X1 _16631_ ( .A1(_00830_ ), .A2(_00828_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00831_ ) );
NAND4_X1 _16632_ ( .A1(_00826_ ), .A2(_00827_ ), .A3(_00829_ ), .A4(_00831_ ), .ZN(_00832_ ) );
NAND3_X1 _16633_ ( .A1(_00822_ ), .A2(_00799_ ), .A3(_00832_ ), .ZN(_00833_ ) );
INV_X2 _16634_ ( .A(_00785_ ), .ZN(_00834_ ) );
BUF_X4 _16635_ ( .A(_00834_ ), .Z(_00835_ ) );
NOR2_X1 _16636_ ( .A1(_00835_ ), .A2(\myifu.data_in [31] ), .ZN(_00836_ ) );
OAI21_X1 _16637_ ( .A(\myifu.state [2] ), .B1(_00787_ ), .B2(_05833_ ), .ZN(_00837_ ) );
OAI21_X1 _16638_ ( .A(_00833_ ), .B1(_00836_ ), .B2(_00837_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
AND3_X1 _16639_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00838_ ) );
AND3_X1 _16640_ ( .A1(_00801_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00839_ ) );
AOI211_X1 _16641_ ( .A(_00838_ ), .B(_00839_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_00817_ ), .ZN(_00840_ ) );
NAND3_X1 _16642_ ( .A1(_00811_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00841_ ) );
NAND4_X1 _16643_ ( .A1(_00840_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_00841_ ), .ZN(_00842_ ) );
NAND3_X1 _16644_ ( .A1(_00823_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00843_ ) );
NAND3_X1 _16645_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00844_ ) );
AND2_X1 _16646_ ( .A1(_00843_ ), .A2(_00844_ ), .ZN(_00845_ ) );
NAND3_X1 _16647_ ( .A1(_00828_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00846_ ) );
NAND3_X1 _16648_ ( .A1(_00830_ ), .A2(_00828_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00847_ ) );
NAND4_X1 _16649_ ( .A1(_00845_ ), .A2(_00827_ ), .A3(_00846_ ), .A4(_00847_ ), .ZN(_00848_ ) );
NAND3_X1 _16650_ ( .A1(_00842_ ), .A2(_00799_ ), .A3(_00848_ ), .ZN(_00849_ ) );
NOR2_X1 _16651_ ( .A1(_00835_ ), .A2(\myifu.data_in [30] ), .ZN(_00850_ ) );
OAI21_X1 _16652_ ( .A(\myifu.state [2] ), .B1(_00787_ ), .B2(_05858_ ), .ZN(_00851_ ) );
OAI21_X1 _16653_ ( .A(_00849_ ), .B1(_00850_ ), .B2(_00851_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
INV_X2 _16654_ ( .A(\myifu.state [2] ), .ZN(_00852_ ) );
BUF_X4 _16655_ ( .A(_00852_ ), .Z(_00853_ ) );
AOI21_X1 _16656_ ( .A(_00853_ ), .B1(_00835_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00854_ ) );
BUF_X4 _16657_ ( .A(_06249_ ), .Z(_00855_ ) );
NAND2_X1 _16658_ ( .A1(_00644_ ), .A2(_00650_ ), .ZN(_00856_ ) );
OAI211_X1 _16659_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_00856_ ), .ZN(_00857_ ) );
NAND2_X1 _16660_ ( .A1(_00854_ ), .A2(_00857_ ), .ZN(_00858_ ) );
AND3_X1 _16661_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00859_ ) );
CLKBUF_X2 _16662_ ( .A(_06076_ ), .Z(_00860_ ) );
AND3_X1 _16663_ ( .A1(_00860_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00861_ ) );
AOI211_X1 _16664_ ( .A(_00859_ ), .B(_00861_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_06230_ ), .ZN(_00862_ ) );
NAND3_X1 _16665_ ( .A1(_06087_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00863_ ) );
NAND4_X1 _16666_ ( .A1(_00862_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00863_ ), .ZN(_00864_ ) );
NAND3_X1 _16667_ ( .A1(_00802_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00865_ ) );
NAND3_X1 _16668_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00866_ ) );
AND2_X1 _16669_ ( .A1(_00865_ ), .A2(_00866_ ), .ZN(_00867_ ) );
BUF_X4 _16670_ ( .A(_00808_ ), .Z(_00868_ ) );
NAND3_X1 _16671_ ( .A1(_00868_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00869_ ) );
NAND3_X1 _16672_ ( .A1(_06078_ ), .A2(_00811_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00870_ ) );
NAND4_X1 _16673_ ( .A1(_00867_ ), .A2(_00807_ ), .A3(_00869_ ), .A4(_00870_ ), .ZN(_00871_ ) );
NAND3_X1 _16674_ ( .A1(_00864_ ), .A2(_00800_ ), .A3(_00871_ ), .ZN(_00872_ ) );
NAND2_X1 _16675_ ( .A1(_00858_ ), .A2(_00872_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
AOI21_X1 _16676_ ( .A(_00853_ ), .B1(_00835_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00873_ ) );
NAND2_X1 _16677_ ( .A1(_00651_ ), .A2(_00654_ ), .ZN(_00874_ ) );
OAI21_X1 _16678_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00874_ ), .ZN(_00875_ ) );
NAND2_X1 _16679_ ( .A1(_00873_ ), .A2(_00875_ ), .ZN(_00876_ ) );
AND3_X1 _16680_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00877_ ) );
AND3_X1 _16681_ ( .A1(_00860_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00878_ ) );
AOI211_X1 _16682_ ( .A(_00877_ ), .B(_00878_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_06230_ ), .ZN(_00879_ ) );
NAND3_X1 _16683_ ( .A1(_06087_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00880_ ) );
NAND4_X1 _16684_ ( .A1(_00879_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00880_ ), .ZN(_00881_ ) );
NAND3_X1 _16685_ ( .A1(_00802_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00882_ ) );
NAND3_X1 _16686_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00883_ ) );
AND2_X1 _16687_ ( .A1(_00882_ ), .A2(_00883_ ), .ZN(_00884_ ) );
NAND3_X1 _16688_ ( .A1(_00868_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00885_ ) );
BUF_X4 _16689_ ( .A(_06086_ ), .Z(_00886_ ) );
NAND3_X1 _16690_ ( .A1(_06078_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00887_ ) );
NAND4_X1 _16691_ ( .A1(_00884_ ), .A2(_00807_ ), .A3(_00885_ ), .A4(_00887_ ), .ZN(_00888_ ) );
NAND3_X1 _16692_ ( .A1(_00881_ ), .A2(_00800_ ), .A3(_00888_ ), .ZN(_00889_ ) );
NAND2_X1 _16693_ ( .A1(_00876_ ), .A2(_00889_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
AOI21_X1 _16694_ ( .A(_00853_ ), .B1(_00835_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00890_ ) );
NAND2_X1 _16695_ ( .A1(_00655_ ), .A2(_00657_ ), .ZN(_00891_ ) );
OAI211_X1 _16696_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_00891_ ), .ZN(_00892_ ) );
NAND2_X1 _16697_ ( .A1(_00890_ ), .A2(_00892_ ), .ZN(_00893_ ) );
AND3_X1 _16698_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00894_ ) );
AND3_X1 _16699_ ( .A1(_00860_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00895_ ) );
AOI211_X1 _16700_ ( .A(_00894_ ), .B(_00895_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_06230_ ), .ZN(_00896_ ) );
NAND3_X1 _16701_ ( .A1(_06087_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00897_ ) );
NAND4_X1 _16702_ ( .A1(_00896_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00897_ ), .ZN(_00898_ ) );
NAND3_X1 _16703_ ( .A1(_00802_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00899_ ) );
NAND3_X1 _16704_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00900_ ) );
AND2_X1 _16705_ ( .A1(_00899_ ), .A2(_00900_ ), .ZN(_00901_ ) );
BUF_X4 _16706_ ( .A(_00827_ ), .Z(_00902_ ) );
NAND3_X1 _16707_ ( .A1(_00868_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00903_ ) );
NAND3_X1 _16708_ ( .A1(_06078_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00904_ ) );
NAND4_X1 _16709_ ( .A1(_00901_ ), .A2(_00902_ ), .A3(_00903_ ), .A4(_00904_ ), .ZN(_00905_ ) );
NAND3_X1 _16710_ ( .A1(_00898_ ), .A2(_00800_ ), .A3(_00905_ ), .ZN(_00906_ ) );
NAND2_X1 _16711_ ( .A1(_00893_ ), .A2(_00906_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
BUF_X4 _16712_ ( .A(_00834_ ), .Z(_00907_ ) );
AOI21_X1 _16713_ ( .A(_00853_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00908_ ) );
NAND2_X1 _16714_ ( .A1(_00658_ ), .A2(_00660_ ), .ZN(_00909_ ) );
OAI21_X1 _16715_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00909_ ), .ZN(_00910_ ) );
NAND2_X1 _16716_ ( .A1(_00908_ ), .A2(_00910_ ), .ZN(_00911_ ) );
AND3_X1 _16717_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00912_ ) );
AND3_X1 _16718_ ( .A1(_00860_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00913_ ) );
AOI211_X1 _16719_ ( .A(_00912_ ), .B(_00913_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_06230_ ), .ZN(_00914_ ) );
BUF_X4 _16720_ ( .A(_00808_ ), .Z(_00915_ ) );
NAND3_X1 _16721_ ( .A1(_00915_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00916_ ) );
NAND4_X1 _16722_ ( .A1(_00914_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00916_ ), .ZN(_00917_ ) );
NAND3_X1 _16723_ ( .A1(_00802_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00918_ ) );
NAND3_X1 _16724_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00919_ ) );
AND2_X1 _16725_ ( .A1(_00918_ ), .A2(_00919_ ), .ZN(_00920_ ) );
NAND3_X1 _16726_ ( .A1(_00868_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00921_ ) );
NAND3_X1 _16727_ ( .A1(_06078_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00922_ ) );
NAND4_X1 _16728_ ( .A1(_00920_ ), .A2(_00902_ ), .A3(_00921_ ), .A4(_00922_ ), .ZN(_00923_ ) );
NAND3_X1 _16729_ ( .A1(_00917_ ), .A2(_00800_ ), .A3(_00923_ ), .ZN(_00924_ ) );
NAND2_X1 _16730_ ( .A1(_00911_ ), .A2(_00924_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
AOI21_X1 _16731_ ( .A(_00853_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00925_ ) );
NAND2_X1 _16732_ ( .A1(_00662_ ), .A2(_00664_ ), .ZN(_00926_ ) );
OAI21_X1 _16733_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00926_ ), .ZN(_00927_ ) );
NAND2_X1 _16734_ ( .A1(_00925_ ), .A2(_00927_ ), .ZN(_00928_ ) );
AND3_X1 _16735_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00929_ ) );
AND3_X1 _16736_ ( .A1(_00860_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00930_ ) );
AOI211_X1 _16737_ ( .A(_00929_ ), .B(_00930_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_06230_ ), .ZN(_00931_ ) );
NAND3_X1 _16738_ ( .A1(_00915_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00932_ ) );
NAND4_X1 _16739_ ( .A1(_00931_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00932_ ), .ZN(_00933_ ) );
NAND3_X1 _16740_ ( .A1(_00802_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00934_ ) );
NAND3_X1 _16741_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00935_ ) );
AND2_X1 _16742_ ( .A1(_00934_ ), .A2(_00935_ ), .ZN(_00936_ ) );
NAND3_X1 _16743_ ( .A1(_00868_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00937_ ) );
BUF_X4 _16744_ ( .A(_06077_ ), .Z(_00938_ ) );
NAND3_X1 _16745_ ( .A1(_00938_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00939_ ) );
NAND4_X1 _16746_ ( .A1(_00936_ ), .A2(_00902_ ), .A3(_00937_ ), .A4(_00939_ ), .ZN(_00940_ ) );
NAND3_X1 _16747_ ( .A1(_00933_ ), .A2(_00800_ ), .A3(_00940_ ), .ZN(_00941_ ) );
NAND2_X1 _16748_ ( .A1(_00928_ ), .A2(_00941_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
NAND2_X1 _16749_ ( .A1(_00665_ ), .A2(_00667_ ), .ZN(_00942_ ) );
OAI211_X1 _16750_ ( .A(_06153_ ), .B(_00781_ ), .C1(_06249_ ), .C2(_00942_ ), .ZN(_00943_ ) );
NAND2_X1 _16751_ ( .A1(_00943_ ), .A2(\myifu.state [2] ), .ZN(_00944_ ) );
AOI21_X1 _16752_ ( .A(_00944_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00834_ ), .ZN(_00945_ ) );
AND3_X1 _16753_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00946_ ) );
AND3_X1 _16754_ ( .A1(_06076_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00947_ ) );
AOI211_X1 _16755_ ( .A(_00946_ ), .B(_00947_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_06229_ ), .ZN(_00948_ ) );
NAND3_X1 _16756_ ( .A1(_00808_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00949_ ) );
NAND4_X1 _16757_ ( .A1(_00948_ ), .A2(_00792_ ), .A3(_00794_ ), .A4(_00949_ ), .ZN(_00950_ ) );
NAND3_X1 _16758_ ( .A1(_06076_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00951_ ) );
NAND3_X1 _16759_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00952_ ) );
AND2_X1 _16760_ ( .A1(_00951_ ), .A2(_00952_ ), .ZN(_00953_ ) );
NAND3_X1 _16761_ ( .A1(_06086_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00954_ ) );
NAND3_X1 _16762_ ( .A1(_06077_ ), .A2(_06086_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00955_ ) );
NAND4_X1 _16763_ ( .A1(_00953_ ), .A2(_00827_ ), .A3(_00954_ ), .A4(_00955_ ), .ZN(_00956_ ) );
AND3_X1 _16764_ ( .A1(_00950_ ), .A2(_00798_ ), .A3(_00956_ ), .ZN(_00957_ ) );
OR2_X1 _16765_ ( .A1(_00945_ ), .A2(_00957_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
AOI21_X1 _16766_ ( .A(_00853_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00958_ ) );
OAI21_X1 _16767_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00670_ ), .ZN(_00959_ ) );
NAND2_X1 _16768_ ( .A1(_00958_ ), .A2(_00959_ ), .ZN(_00960_ ) );
AND3_X1 _16769_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00961_ ) );
AND3_X1 _16770_ ( .A1(_00860_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00962_ ) );
BUF_X4 _16771_ ( .A(_06229_ ), .Z(_00963_ ) );
AOI211_X1 _16772_ ( .A(_00961_ ), .B(_00962_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_00963_ ), .ZN(_00964_ ) );
NAND3_X1 _16773_ ( .A1(_00915_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00965_ ) );
NAND4_X1 _16774_ ( .A1(_00964_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00965_ ), .ZN(_00966_ ) );
BUF_X4 _16775_ ( .A(_00801_ ), .Z(_00967_ ) );
NAND3_X1 _16776_ ( .A1(_00967_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00968_ ) );
NAND3_X1 _16777_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00969_ ) );
AND2_X1 _16778_ ( .A1(_00968_ ), .A2(_00969_ ), .ZN(_00970_ ) );
NAND3_X1 _16779_ ( .A1(_00868_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00971_ ) );
NAND3_X1 _16780_ ( .A1(_00938_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00972_ ) );
NAND4_X1 _16781_ ( .A1(_00970_ ), .A2(_00902_ ), .A3(_00971_ ), .A4(_00972_ ), .ZN(_00973_ ) );
NAND3_X1 _16782_ ( .A1(_00966_ ), .A2(_00800_ ), .A3(_00973_ ), .ZN(_00974_ ) );
NAND2_X1 _16783_ ( .A1(_00960_ ), .A2(_00974_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
AND3_X1 _16784_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00975_ ) );
AND3_X1 _16785_ ( .A1(_00801_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00976_ ) );
AOI211_X1 _16786_ ( .A(_00975_ ), .B(_00976_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_00817_ ), .ZN(_00977_ ) );
NAND3_X1 _16787_ ( .A1(_00811_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00978_ ) );
NAND4_X1 _16788_ ( .A1(_00977_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_00978_ ), .ZN(_00979_ ) );
NAND3_X1 _16789_ ( .A1(_00823_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00980_ ) );
NAND3_X1 _16790_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00981_ ) );
AND2_X1 _16791_ ( .A1(_00980_ ), .A2(_00981_ ), .ZN(_00982_ ) );
NAND3_X1 _16792_ ( .A1(_00828_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00983_ ) );
NAND3_X1 _16793_ ( .A1(_00802_ ), .A2(_00828_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00984_ ) );
NAND4_X1 _16794_ ( .A1(_00982_ ), .A2(_00827_ ), .A3(_00983_ ), .A4(_00984_ ), .ZN(_00985_ ) );
NAND3_X1 _16795_ ( .A1(_00979_ ), .A2(_00799_ ), .A3(_00985_ ), .ZN(_00986_ ) );
AND2_X1 _16796_ ( .A1(_00835_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00987_ ) );
OAI21_X1 _16797_ ( .A(\myifu.state [2] ), .B1(_00835_ ), .B2(\myifu.data_in [14] ), .ZN(_00988_ ) );
OAI21_X1 _16798_ ( .A(_00986_ ), .B1(_00987_ ), .B2(_00988_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
AOI21_X1 _16799_ ( .A(_00853_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00989_ ) );
NAND2_X1 _16800_ ( .A1(_00675_ ), .A2(_00677_ ), .ZN(_00990_ ) );
OAI21_X1 _16801_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00990_ ), .ZN(_00991_ ) );
NAND2_X1 _16802_ ( .A1(_00989_ ), .A2(_00991_ ), .ZN(_00992_ ) );
AND3_X1 _16803_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00993_ ) );
AND3_X1 _16804_ ( .A1(_00860_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00994_ ) );
AOI211_X1 _16805_ ( .A(_00993_ ), .B(_00994_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_00963_ ), .ZN(_00995_ ) );
NAND3_X1 _16806_ ( .A1(_00915_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00996_ ) );
NAND4_X1 _16807_ ( .A1(_00995_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_00996_ ), .ZN(_00997_ ) );
NAND3_X1 _16808_ ( .A1(_00967_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00998_ ) );
NAND3_X1 _16809_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00999_ ) );
AND2_X1 _16810_ ( .A1(_00998_ ), .A2(_00999_ ), .ZN(_01000_ ) );
NAND3_X1 _16811_ ( .A1(_00868_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_01001_ ) );
NAND3_X1 _16812_ ( .A1(_00938_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_01002_ ) );
NAND4_X1 _16813_ ( .A1(_01000_ ), .A2(_00902_ ), .A3(_01001_ ), .A4(_01002_ ), .ZN(_01003_ ) );
NAND3_X1 _16814_ ( .A1(_00997_ ), .A2(_00800_ ), .A3(_01003_ ), .ZN(_01004_ ) );
NAND2_X1 _16815_ ( .A1(_00992_ ), .A2(_01004_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
AOI21_X1 _16816_ ( .A(_00853_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01005_ ) );
NAND2_X1 _16817_ ( .A1(_00678_ ), .A2(_00680_ ), .ZN(_01006_ ) );
OAI211_X1 _16818_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_01006_ ), .ZN(_01007_ ) );
NAND2_X1 _16819_ ( .A1(_01005_ ), .A2(_01007_ ), .ZN(_01008_ ) );
AND3_X1 _16820_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_01009_ ) );
AND3_X1 _16821_ ( .A1(_00860_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_01010_ ) );
AOI211_X1 _16822_ ( .A(_01009_ ), .B(_01010_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_00963_ ), .ZN(_01011_ ) );
NAND3_X1 _16823_ ( .A1(_00915_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_01012_ ) );
NAND4_X1 _16824_ ( .A1(_01011_ ), .A2(_00793_ ), .A3(_00795_ ), .A4(_01012_ ), .ZN(_01013_ ) );
NAND3_X1 _16825_ ( .A1(_00967_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_01014_ ) );
NAND3_X1 _16826_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_01015_ ) );
AND2_X1 _16827_ ( .A1(_01014_ ), .A2(_01015_ ), .ZN(_01016_ ) );
NAND3_X1 _16828_ ( .A1(_00868_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_01017_ ) );
NAND3_X1 _16829_ ( .A1(_00938_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_01018_ ) );
NAND4_X1 _16830_ ( .A1(_01016_ ), .A2(_00902_ ), .A3(_01017_ ), .A4(_01018_ ), .ZN(_01019_ ) );
NAND3_X1 _16831_ ( .A1(_01013_ ), .A2(_00800_ ), .A3(_01019_ ), .ZN(_01020_ ) );
NAND2_X1 _16832_ ( .A1(_01008_ ), .A2(_01020_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
AND3_X1 _16833_ ( .A1(fanout_net_18 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_01021_ ) );
AND3_X1 _16834_ ( .A1(_00801_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_01022_ ) );
AOI211_X1 _16835_ ( .A(_01021_ ), .B(_01022_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_06229_ ), .ZN(_01023_ ) );
NAND3_X1 _16836_ ( .A1(_00811_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_01024_ ) );
NAND4_X1 _16837_ ( .A1(_01023_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_01024_ ), .ZN(_01025_ ) );
NAND3_X1 _16838_ ( .A1(_06077_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_01026_ ) );
NAND3_X1 _16839_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_01027_ ) );
AND2_X1 _16840_ ( .A1(_01026_ ), .A2(_01027_ ), .ZN(_01028_ ) );
NAND3_X1 _16841_ ( .A1(_00828_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_01029_ ) );
NAND3_X1 _16842_ ( .A1(_00802_ ), .A2(_00808_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_01030_ ) );
NAND4_X1 _16843_ ( .A1(_01028_ ), .A2(_00827_ ), .A3(_01029_ ), .A4(_01030_ ), .ZN(_01031_ ) );
NAND3_X1 _16844_ ( .A1(_01025_ ), .A2(_00799_ ), .A3(_01031_ ), .ZN(_01032_ ) );
NOR2_X1 _16845_ ( .A1(_00835_ ), .A2(\myifu.data_in [29] ), .ZN(_01033_ ) );
OAI21_X1 _16846_ ( .A(\myifu.state [2] ), .B1(_00787_ ), .B2(_05854_ ), .ZN(_01034_ ) );
OAI21_X1 _16847_ ( .A(_01032_ ), .B1(_01033_ ), .B2(_01034_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16848_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_01035_ ) );
AND3_X1 _16849_ ( .A1(_00801_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_01036_ ) );
AOI211_X1 _16850_ ( .A(_01035_ ), .B(_01036_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_06229_ ), .ZN(_01037_ ) );
NAND3_X1 _16851_ ( .A1(_00811_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_01038_ ) );
NAND4_X1 _16852_ ( .A1(_01037_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_01038_ ), .ZN(_01039_ ) );
NAND3_X1 _16853_ ( .A1(_06077_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_01040_ ) );
NAND3_X1 _16854_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_01041_ ) );
AND2_X1 _16855_ ( .A1(_01040_ ), .A2(_01041_ ), .ZN(_01042_ ) );
NAND3_X1 _16856_ ( .A1(_00828_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_01043_ ) );
NAND3_X1 _16857_ ( .A1(_00802_ ), .A2(_00808_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_01044_ ) );
NAND4_X1 _16858_ ( .A1(_01042_ ), .A2(_00827_ ), .A3(_01043_ ), .A4(_01044_ ), .ZN(_01045_ ) );
NAND3_X1 _16859_ ( .A1(_01039_ ), .A2(_00799_ ), .A3(_01045_ ), .ZN(_01046_ ) );
NOR2_X1 _16860_ ( .A1(_00835_ ), .A2(\myifu.data_in [11] ), .ZN(_01047_ ) );
OAI21_X1 _16861_ ( .A(\myifu.state [2] ), .B1(_00787_ ), .B2(_05789_ ), .ZN(_01048_ ) );
OAI21_X1 _16862_ ( .A(_01046_ ), .B1(_01047_ ), .B2(_01048_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
AND3_X1 _16863_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_01049_ ) );
AND3_X1 _16864_ ( .A1(_00801_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_01050_ ) );
AOI211_X1 _16865_ ( .A(_01049_ ), .B(_01050_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_06229_ ), .ZN(_01051_ ) );
NAND3_X1 _16866_ ( .A1(_00811_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_01052_ ) );
NAND4_X1 _16867_ ( .A1(_01051_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_01052_ ), .ZN(_01053_ ) );
NAND3_X1 _16868_ ( .A1(_06077_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_01054_ ) );
NAND3_X1 _16869_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_01055_ ) );
AND2_X1 _16870_ ( .A1(_01054_ ), .A2(_01055_ ), .ZN(_01056_ ) );
NAND3_X1 _16871_ ( .A1(_00828_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_01057_ ) );
NAND3_X1 _16872_ ( .A1(_00802_ ), .A2(_00808_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_01058_ ) );
NAND4_X1 _16873_ ( .A1(_01056_ ), .A2(_00827_ ), .A3(_01057_ ), .A4(_01058_ ), .ZN(_01059_ ) );
NAND3_X1 _16874_ ( .A1(_01053_ ), .A2(_00799_ ), .A3(_01059_ ), .ZN(_01060_ ) );
NOR2_X1 _16875_ ( .A1(_00835_ ), .A2(\myifu.data_in [10] ), .ZN(_01061_ ) );
OAI21_X1 _16876_ ( .A(\myifu.state [2] ), .B1(_00787_ ), .B2(_05784_ ), .ZN(_01062_ ) );
OAI21_X1 _16877_ ( .A(_01060_ ), .B1(_01061_ ), .B2(_01062_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
NAND2_X1 _16878_ ( .A1(_00691_ ), .A2(_00693_ ), .ZN(_01063_ ) );
OAI211_X1 _16879_ ( .A(_06153_ ), .B(_00781_ ), .C1(_02156_ ), .C2(_01063_ ), .ZN(_01064_ ) );
NAND2_X1 _16880_ ( .A1(_01064_ ), .A2(\myifu.state [2] ), .ZN(_01065_ ) );
AOI21_X1 _16881_ ( .A(_01065_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .B2(_00834_ ), .ZN(_01066_ ) );
AND3_X1 _16882_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_01067_ ) );
AND3_X1 _16883_ ( .A1(_06076_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_01068_ ) );
AOI211_X1 _16884_ ( .A(_01067_ ), .B(_01068_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_06229_ ), .ZN(_01069_ ) );
NAND3_X1 _16885_ ( .A1(_00808_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_01070_ ) );
NAND4_X1 _16886_ ( .A1(_01069_ ), .A2(_00792_ ), .A3(_00794_ ), .A4(_01070_ ), .ZN(_01071_ ) );
NAND3_X1 _16887_ ( .A1(_06076_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_01072_ ) );
NAND3_X1 _16888_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_01073_ ) );
AND2_X1 _16889_ ( .A1(_01072_ ), .A2(_01073_ ), .ZN(_01074_ ) );
NAND3_X1 _16890_ ( .A1(_06086_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_01075_ ) );
NAND3_X1 _16891_ ( .A1(_06077_ ), .A2(_06086_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_01076_ ) );
NAND4_X1 _16892_ ( .A1(_01074_ ), .A2(_00827_ ), .A3(_01075_ ), .A4(_01076_ ), .ZN(_01077_ ) );
AND3_X1 _16893_ ( .A1(_01071_ ), .A2(_00798_ ), .A3(_01077_ ), .ZN(_01078_ ) );
OR2_X1 _16894_ ( .A1(_01066_ ), .A2(_01078_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
OAI211_X1 _16895_ ( .A(_06153_ ), .B(_00781_ ), .C1(_06249_ ), .C2(_00699_ ), .ZN(_01079_ ) );
OAI211_X1 _16896_ ( .A(_01079_ ), .B(\myifu.state [2] ), .C1(_00787_ ), .C2(_05848_ ), .ZN(_01080_ ) );
AND3_X1 _16897_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_01081_ ) );
AND3_X1 _16898_ ( .A1(_00860_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_01082_ ) );
AOI211_X1 _16899_ ( .A(_01081_ ), .B(_01082_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_00963_ ), .ZN(_01083_ ) );
BUF_X4 _16900_ ( .A(_00792_ ), .Z(_01084_ ) );
BUF_X4 _16901_ ( .A(_00794_ ), .Z(_01085_ ) );
NAND3_X1 _16902_ ( .A1(_00915_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_01086_ ) );
NAND4_X1 _16903_ ( .A1(_01083_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01086_ ), .ZN(_01087_ ) );
NAND3_X1 _16904_ ( .A1(_00967_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_01088_ ) );
NAND3_X1 _16905_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_01089_ ) );
AND2_X1 _16906_ ( .A1(_01088_ ), .A2(_01089_ ), .ZN(_01090_ ) );
NAND3_X1 _16907_ ( .A1(_00868_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_01091_ ) );
NAND3_X1 _16908_ ( .A1(_00938_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_01092_ ) );
NAND4_X1 _16909_ ( .A1(_01090_ ), .A2(_00902_ ), .A3(_01091_ ), .A4(_01092_ ), .ZN(_01093_ ) );
NAND3_X1 _16910_ ( .A1(_01087_ ), .A2(_00800_ ), .A3(_01093_ ), .ZN(_01094_ ) );
NAND2_X1 _16911_ ( .A1(_01080_ ), .A2(_01094_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
OAI211_X1 _16912_ ( .A(_06153_ ), .B(_00781_ ), .C1(_06249_ ), .C2(_00702_ ), .ZN(_01095_ ) );
OAI211_X1 _16913_ ( .A(_01095_ ), .B(\myifu.state [2] ), .C1(_00787_ ), .C2(_05502_ ), .ZN(_01096_ ) );
AND3_X1 _16914_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_01097_ ) );
AND3_X1 _16915_ ( .A1(_00860_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_01098_ ) );
AOI211_X1 _16916_ ( .A(_01097_ ), .B(_01098_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00963_ ), .ZN(_01099_ ) );
NAND3_X1 _16917_ ( .A1(_00915_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_01100_ ) );
NAND4_X1 _16918_ ( .A1(_01099_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01100_ ), .ZN(_01101_ ) );
BUF_X4 _16919_ ( .A(_00798_ ), .Z(_01102_ ) );
NAND3_X1 _16920_ ( .A1(_00967_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_01103_ ) );
NAND3_X1 _16921_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_01104_ ) );
AND2_X1 _16922_ ( .A1(_01103_ ), .A2(_01104_ ), .ZN(_01105_ ) );
NAND3_X1 _16923_ ( .A1(_00868_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_01106_ ) );
NAND3_X1 _16924_ ( .A1(_00938_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_01107_ ) );
NAND4_X1 _16925_ ( .A1(_01105_ ), .A2(_00902_ ), .A3(_01106_ ), .A4(_01107_ ), .ZN(_01108_ ) );
NAND3_X1 _16926_ ( .A1(_01101_ ), .A2(_01102_ ), .A3(_01108_ ), .ZN(_01109_ ) );
NAND2_X1 _16927_ ( .A1(_01096_ ), .A2(_01109_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
AOI21_X1 _16928_ ( .A(_00853_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01110_ ) );
OAI211_X1 _16929_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_00705_ ), .ZN(_01111_ ) );
NAND2_X1 _16930_ ( .A1(_01110_ ), .A2(_01111_ ), .ZN(_01112_ ) );
AND3_X1 _16931_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_01113_ ) );
CLKBUF_X2 _16932_ ( .A(_06076_ ), .Z(_01114_ ) );
AND3_X1 _16933_ ( .A1(_01114_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_01115_ ) );
AOI211_X1 _16934_ ( .A(_01113_ ), .B(_01115_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00963_ ), .ZN(_01116_ ) );
NAND3_X1 _16935_ ( .A1(_00915_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_01117_ ) );
NAND4_X1 _16936_ ( .A1(_01116_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01117_ ), .ZN(_01118_ ) );
NAND3_X1 _16937_ ( .A1(_00967_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_01119_ ) );
NAND3_X1 _16938_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_01120_ ) );
AND2_X1 _16939_ ( .A1(_01119_ ), .A2(_01120_ ), .ZN(_01121_ ) );
BUF_X4 _16940_ ( .A(_00808_ ), .Z(_01122_ ) );
NAND3_X1 _16941_ ( .A1(_01122_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_01123_ ) );
NAND3_X1 _16942_ ( .A1(_00938_ ), .A2(_00886_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_01124_ ) );
NAND4_X1 _16943_ ( .A1(_01121_ ), .A2(_00902_ ), .A3(_01123_ ), .A4(_01124_ ), .ZN(_01125_ ) );
NAND3_X1 _16944_ ( .A1(_01118_ ), .A2(_01102_ ), .A3(_01125_ ), .ZN(_01126_ ) );
NAND2_X1 _16945_ ( .A1(_01112_ ), .A2(_01126_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
AOI21_X1 _16946_ ( .A(_00853_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01127_ ) );
OAI21_X1 _16947_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00708_ ), .ZN(_01128_ ) );
NAND2_X1 _16948_ ( .A1(_01127_ ), .A2(_01128_ ), .ZN(_01129_ ) );
AND3_X1 _16949_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_01130_ ) );
AND3_X1 _16950_ ( .A1(_01114_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_01131_ ) );
AOI211_X1 _16951_ ( .A(_01130_ ), .B(_01131_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00963_ ), .ZN(_01132_ ) );
NAND3_X1 _16952_ ( .A1(_00915_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_01133_ ) );
NAND4_X1 _16953_ ( .A1(_01132_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01133_ ), .ZN(_01134_ ) );
NAND3_X1 _16954_ ( .A1(_00967_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_01135_ ) );
NAND3_X1 _16955_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_01136_ ) );
AND2_X1 _16956_ ( .A1(_01135_ ), .A2(_01136_ ), .ZN(_01137_ ) );
NAND3_X1 _16957_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_01138_ ) );
BUF_X4 _16958_ ( .A(_06086_ ), .Z(_01139_ ) );
NAND3_X1 _16959_ ( .A1(_00938_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_01140_ ) );
NAND4_X1 _16960_ ( .A1(_01137_ ), .A2(_00902_ ), .A3(_01138_ ), .A4(_01140_ ), .ZN(_01141_ ) );
NAND3_X1 _16961_ ( .A1(_01134_ ), .A2(_01102_ ), .A3(_01141_ ), .ZN(_01142_ ) );
NAND2_X1 _16962_ ( .A1(_01129_ ), .A2(_01142_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _16963_ ( .A(_00852_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01143_ ) );
OAI211_X1 _16964_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_00711_ ), .ZN(_01144_ ) );
NAND2_X1 _16965_ ( .A1(_01143_ ), .A2(_01144_ ), .ZN(_01145_ ) );
AND3_X1 _16966_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_01146_ ) );
AND3_X1 _16967_ ( .A1(_01114_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_01147_ ) );
AOI211_X1 _16968_ ( .A(_01146_ ), .B(_01147_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00963_ ), .ZN(_01148_ ) );
NAND3_X1 _16969_ ( .A1(_00915_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_01149_ ) );
NAND4_X1 _16970_ ( .A1(_01148_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01149_ ), .ZN(_01150_ ) );
NAND3_X1 _16971_ ( .A1(_00967_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_01151_ ) );
NAND3_X1 _16972_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_01152_ ) );
AND2_X1 _16973_ ( .A1(_01151_ ), .A2(_01152_ ), .ZN(_01153_ ) );
BUF_X4 _16974_ ( .A(_00827_ ), .Z(_01154_ ) );
NAND3_X1 _16975_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_01155_ ) );
NAND3_X1 _16976_ ( .A1(_00938_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_01156_ ) );
NAND4_X1 _16977_ ( .A1(_01153_ ), .A2(_01154_ ), .A3(_01155_ ), .A4(_01156_ ), .ZN(_01157_ ) );
NAND3_X1 _16978_ ( .A1(_01150_ ), .A2(_01102_ ), .A3(_01157_ ), .ZN(_01158_ ) );
NAND2_X1 _16979_ ( .A1(_01145_ ), .A2(_01158_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
AOI21_X1 _16980_ ( .A(_00852_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01159_ ) );
OAI211_X1 _16981_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_00714_ ), .ZN(_01160_ ) );
NAND2_X1 _16982_ ( .A1(_01159_ ), .A2(_01160_ ), .ZN(_01161_ ) );
AND3_X1 _16983_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_01162_ ) );
AND3_X1 _16984_ ( .A1(_01114_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_01163_ ) );
AOI211_X1 _16985_ ( .A(_01162_ ), .B(_01163_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_00963_ ), .ZN(_01164_ ) );
NAND3_X1 _16986_ ( .A1(_00809_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_01165_ ) );
NAND4_X1 _16987_ ( .A1(_01164_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01165_ ), .ZN(_01166_ ) );
NAND3_X1 _16988_ ( .A1(_00967_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_01167_ ) );
NAND3_X1 _16989_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_01168_ ) );
AND2_X1 _16990_ ( .A1(_01167_ ), .A2(_01168_ ), .ZN(_01169_ ) );
NAND3_X1 _16991_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_01170_ ) );
NAND3_X1 _16992_ ( .A1(_00938_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_01171_ ) );
NAND4_X1 _16993_ ( .A1(_01169_ ), .A2(_01154_ ), .A3(_01170_ ), .A4(_01171_ ), .ZN(_01172_ ) );
NAND3_X1 _16994_ ( .A1(_01166_ ), .A2(_01102_ ), .A3(_01172_ ), .ZN(_01173_ ) );
NAND2_X1 _16995_ ( .A1(_01161_ ), .A2(_01173_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
AOI21_X1 _16996_ ( .A(_00852_ ), .B1(_00907_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01174_ ) );
OAI21_X1 _16997_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00720_ ), .ZN(_01175_ ) );
NAND2_X1 _16998_ ( .A1(_01174_ ), .A2(_01175_ ), .ZN(_01176_ ) );
AND3_X1 _16999_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01177_ ) );
AND3_X1 _17000_ ( .A1(_01114_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01178_ ) );
AOI211_X1 _17001_ ( .A(_01177_ ), .B(_01178_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_00963_ ), .ZN(_01179_ ) );
NAND3_X1 _17002_ ( .A1(_00809_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01180_ ) );
NAND4_X1 _17003_ ( .A1(_01179_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01180_ ), .ZN(_01181_ ) );
NAND3_X1 _17004_ ( .A1(_00967_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01182_ ) );
NAND3_X1 _17005_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01183_ ) );
AND2_X1 _17006_ ( .A1(_01182_ ), .A2(_01183_ ), .ZN(_01184_ ) );
NAND3_X1 _17007_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01185_ ) );
NAND3_X1 _17008_ ( .A1(_00830_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01186_ ) );
NAND4_X1 _17009_ ( .A1(_01184_ ), .A2(_01154_ ), .A3(_01185_ ), .A4(_01186_ ), .ZN(_01187_ ) );
NAND3_X1 _17010_ ( .A1(_01181_ ), .A2(_01102_ ), .A3(_01187_ ), .ZN(_01188_ ) );
NAND2_X1 _17011_ ( .A1(_01176_ ), .A2(_01188_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
NAND2_X1 _17012_ ( .A1(_00715_ ), .A2(_00717_ ), .ZN(_01189_ ) );
OAI211_X1 _17013_ ( .A(_06153_ ), .B(_00781_ ), .C1(_06249_ ), .C2(_01189_ ), .ZN(_01190_ ) );
OAI211_X1 _17014_ ( .A(_01190_ ), .B(\myifu.state [2] ), .C1(_00787_ ), .C2(_05821_ ), .ZN(_01191_ ) );
AND3_X1 _17015_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01192_ ) );
AND3_X1 _17016_ ( .A1(_01114_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01193_ ) );
AOI211_X1 _17017_ ( .A(_01192_ ), .B(_01193_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00817_ ), .ZN(_01194_ ) );
NAND3_X1 _17018_ ( .A1(_00809_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01195_ ) );
NAND4_X1 _17019_ ( .A1(_01194_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01195_ ), .ZN(_01196_ ) );
NAND3_X1 _17020_ ( .A1(_00823_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01197_ ) );
NAND3_X1 _17021_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01198_ ) );
AND2_X1 _17022_ ( .A1(_01197_ ), .A2(_01198_ ), .ZN(_01199_ ) );
NAND3_X1 _17023_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01200_ ) );
NAND3_X1 _17024_ ( .A1(_00830_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01201_ ) );
NAND4_X1 _17025_ ( .A1(_01199_ ), .A2(_01154_ ), .A3(_01200_ ), .A4(_01201_ ), .ZN(_01202_ ) );
NAND3_X1 _17026_ ( .A1(_01196_ ), .A2(_01102_ ), .A3(_01202_ ), .ZN(_01203_ ) );
NAND2_X1 _17027_ ( .A1(_01191_ ), .A2(_01203_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
AOI21_X1 _17028_ ( .A(_00852_ ), .B1(_00834_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01204_ ) );
OAI21_X1 _17029_ ( .A(_00786_ ), .B1(_06282_ ), .B2(_00723_ ), .ZN(_01205_ ) );
NAND2_X1 _17030_ ( .A1(_01204_ ), .A2(_01205_ ), .ZN(_01206_ ) );
AND3_X1 _17031_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01207_ ) );
AND3_X1 _17032_ ( .A1(_01114_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01208_ ) );
AOI211_X1 _17033_ ( .A(_01207_ ), .B(_01208_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_00817_ ), .ZN(_01209_ ) );
NAND3_X1 _17034_ ( .A1(_00809_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01210_ ) );
NAND4_X1 _17035_ ( .A1(_01209_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01210_ ), .ZN(_01211_ ) );
NAND3_X1 _17036_ ( .A1(_00823_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01212_ ) );
NAND3_X1 _17037_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01213_ ) );
AND2_X1 _17038_ ( .A1(_01212_ ), .A2(_01213_ ), .ZN(_01214_ ) );
NAND3_X1 _17039_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01215_ ) );
NAND3_X1 _17040_ ( .A1(_00830_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01216_ ) );
NAND4_X1 _17041_ ( .A1(_01214_ ), .A2(_01154_ ), .A3(_01215_ ), .A4(_01216_ ), .ZN(_01217_ ) );
NAND3_X1 _17042_ ( .A1(_01211_ ), .A2(_01102_ ), .A3(_01217_ ), .ZN(_01218_ ) );
NAND2_X1 _17043_ ( .A1(_01206_ ), .A2(_01218_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
AOI21_X1 _17044_ ( .A(_00852_ ), .B1(_00834_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_01219_ ) );
NAND2_X1 _17045_ ( .A1(_00725_ ), .A2(_00727_ ), .ZN(_01220_ ) );
OAI211_X1 _17046_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_01220_ ), .ZN(_01221_ ) );
NAND2_X1 _17047_ ( .A1(_01219_ ), .A2(_01221_ ), .ZN(_01222_ ) );
AND3_X1 _17048_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01223_ ) );
AND3_X1 _17049_ ( .A1(_01114_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01224_ ) );
AOI211_X1 _17050_ ( .A(_01223_ ), .B(_01224_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00817_ ), .ZN(_01225_ ) );
NAND3_X1 _17051_ ( .A1(_00809_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01226_ ) );
NAND4_X1 _17052_ ( .A1(_01225_ ), .A2(_01084_ ), .A3(_01085_ ), .A4(_01226_ ), .ZN(_01227_ ) );
NAND3_X1 _17053_ ( .A1(_00823_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01228_ ) );
NAND3_X1 _17054_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01229_ ) );
AND2_X1 _17055_ ( .A1(_01228_ ), .A2(_01229_ ), .ZN(_01230_ ) );
NAND3_X1 _17056_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01231_ ) );
NAND3_X1 _17057_ ( .A1(_00830_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01232_ ) );
NAND4_X1 _17058_ ( .A1(_01230_ ), .A2(_01154_ ), .A3(_01231_ ), .A4(_01232_ ), .ZN(_01233_ ) );
NAND3_X1 _17059_ ( .A1(_01227_ ), .A2(_01102_ ), .A3(_01233_ ), .ZN(_01234_ ) );
NAND2_X1 _17060_ ( .A1(_01222_ ), .A2(_01234_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
NAND2_X1 _17061_ ( .A1(_00728_ ), .A2(_00730_ ), .ZN(_01235_ ) );
OAI211_X1 _17062_ ( .A(_06153_ ), .B(_00781_ ), .C1(_06249_ ), .C2(_01235_ ), .ZN(_01236_ ) );
OAI211_X1 _17063_ ( .A(_01236_ ), .B(\myifu.state [2] ), .C1(_00787_ ), .C2(_05808_ ), .ZN(_01237_ ) );
AND3_X1 _17064_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01238_ ) );
AND3_X1 _17065_ ( .A1(_01114_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01239_ ) );
AOI211_X1 _17066_ ( .A(_01238_ ), .B(_01239_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_00817_ ), .ZN(_01240_ ) );
NAND3_X1 _17067_ ( .A1(_00809_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01241_ ) );
NAND4_X1 _17068_ ( .A1(_01240_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_01241_ ), .ZN(_01242_ ) );
NAND3_X1 _17069_ ( .A1(_00823_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01243_ ) );
NAND3_X1 _17070_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01244_ ) );
AND2_X1 _17071_ ( .A1(_01243_ ), .A2(_01244_ ), .ZN(_01245_ ) );
NAND3_X1 _17072_ ( .A1(_01122_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01246_ ) );
NAND3_X1 _17073_ ( .A1(_00830_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01247_ ) );
NAND4_X1 _17074_ ( .A1(_01245_ ), .A2(_01154_ ), .A3(_01246_ ), .A4(_01247_ ), .ZN(_01248_ ) );
NAND3_X1 _17075_ ( .A1(_01242_ ), .A2(_01102_ ), .A3(_01248_ ), .ZN(_01249_ ) );
NAND2_X1 _17076_ ( .A1(_01237_ ), .A2(_01249_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
AOI21_X1 _17077_ ( .A(_00852_ ), .B1(_00834_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_01250_ ) );
NAND2_X1 _17078_ ( .A1(_00731_ ), .A2(_00733_ ), .ZN(_01251_ ) );
OAI211_X1 _17079_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_01251_ ), .ZN(_01252_ ) );
NAND2_X1 _17080_ ( .A1(_01250_ ), .A2(_01252_ ), .ZN(_01253_ ) );
AND3_X1 _17081_ ( .A1(\IF_ID_pc [4] ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01254_ ) );
AND3_X1 _17082_ ( .A1(_01114_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01255_ ) );
AOI211_X1 _17083_ ( .A(_01254_ ), .B(_01255_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00817_ ), .ZN(_01256_ ) );
NAND3_X1 _17084_ ( .A1(_00809_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01257_ ) );
NAND4_X1 _17085_ ( .A1(_01256_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_01257_ ), .ZN(_01258_ ) );
NAND3_X1 _17086_ ( .A1(_00823_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01259_ ) );
NAND3_X1 _17087_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01260_ ) );
AND2_X1 _17088_ ( .A1(_01259_ ), .A2(_01260_ ), .ZN(_01261_ ) );
NAND3_X1 _17089_ ( .A1(_01122_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01262_ ) );
NAND3_X1 _17090_ ( .A1(_00830_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01263_ ) );
NAND4_X1 _17091_ ( .A1(_01261_ ), .A2(_01154_ ), .A3(_01262_ ), .A4(_01263_ ), .ZN(_01264_ ) );
NAND3_X1 _17092_ ( .A1(_01258_ ), .A2(_00799_ ), .A3(_01264_ ), .ZN(_01265_ ) );
NAND2_X1 _17093_ ( .A1(_01253_ ), .A2(_01265_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
NAND2_X1 _17094_ ( .A1(_00734_ ), .A2(_00736_ ), .ZN(_01266_ ) );
OAI211_X1 _17095_ ( .A(_06153_ ), .B(_00781_ ), .C1(_02156_ ), .C2(_01266_ ), .ZN(_01267_ ) );
NAND2_X1 _17096_ ( .A1(_01267_ ), .A2(\myifu.state [2] ), .ZN(_01268_ ) );
AOI21_X1 _17097_ ( .A(_01268_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00834_ ), .ZN(_01269_ ) );
AND3_X1 _17098_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01270_ ) );
AND3_X1 _17099_ ( .A1(_06076_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01271_ ) );
AOI211_X1 _17100_ ( .A(_01270_ ), .B(_01271_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_06229_ ), .ZN(_01272_ ) );
NAND3_X1 _17101_ ( .A1(_00808_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01273_ ) );
NAND4_X1 _17102_ ( .A1(_01272_ ), .A2(_00792_ ), .A3(_00794_ ), .A4(_01273_ ), .ZN(_01274_ ) );
NAND3_X1 _17103_ ( .A1(_06076_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01275_ ) );
NAND3_X1 _17104_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01276_ ) );
AND2_X1 _17105_ ( .A1(_01275_ ), .A2(_01276_ ), .ZN(_01277_ ) );
NAND3_X1 _17106_ ( .A1(_06086_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01278_ ) );
NAND3_X1 _17107_ ( .A1(_06077_ ), .A2(_06085_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01279_ ) );
NAND4_X1 _17108_ ( .A1(_01277_ ), .A2(_00806_ ), .A3(_01278_ ), .A4(_01279_ ), .ZN(_01280_ ) );
AND3_X1 _17109_ ( .A1(_01274_ ), .A2(_00798_ ), .A3(_01280_ ), .ZN(_01281_ ) );
OR2_X1 _17110_ ( .A1(_01269_ ), .A2(_01281_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
AOI21_X1 _17111_ ( .A(_00852_ ), .B1(_00834_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01282_ ) );
OAI211_X1 _17112_ ( .A(_00777_ ), .B(_00782_ ), .C1(_00855_ ), .C2(_00739_ ), .ZN(_01283_ ) );
NAND2_X1 _17113_ ( .A1(_01282_ ), .A2(_01283_ ), .ZN(_01284_ ) );
AND3_X1 _17114_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01285_ ) );
AND3_X1 _17115_ ( .A1(_00801_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01286_ ) );
AOI211_X1 _17116_ ( .A(_01285_ ), .B(_01286_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_00817_ ), .ZN(_01287_ ) );
NAND3_X1 _17117_ ( .A1(_00809_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01288_ ) );
NAND4_X1 _17118_ ( .A1(_01287_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_01288_ ), .ZN(_01289_ ) );
NAND3_X1 _17119_ ( .A1(_00823_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01290_ ) );
NAND3_X1 _17120_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01291_ ) );
AND2_X1 _17121_ ( .A1(_01290_ ), .A2(_01291_ ), .ZN(_01292_ ) );
NAND3_X1 _17122_ ( .A1(_00811_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01293_ ) );
NAND3_X1 _17123_ ( .A1(_00830_ ), .A2(_01139_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01294_ ) );
NAND4_X1 _17124_ ( .A1(_01292_ ), .A2(_01154_ ), .A3(_01293_ ), .A4(_01294_ ), .ZN(_01295_ ) );
NAND3_X1 _17125_ ( .A1(_01289_ ), .A2(_00799_ ), .A3(_01295_ ), .ZN(_01296_ ) );
NAND2_X1 _17126_ ( .A1(_01284_ ), .A2(_01296_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
AOI21_X1 _17127_ ( .A(_00852_ ), .B1(_00834_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_01297_ ) );
OAI21_X1 _17128_ ( .A(_00786_ ), .B1(_00855_ ), .B2(_00742_ ), .ZN(_01298_ ) );
NAND2_X1 _17129_ ( .A1(_01297_ ), .A2(_01298_ ), .ZN(_01299_ ) );
AND3_X1 _17130_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01300_ ) );
AND3_X1 _17131_ ( .A1(_00801_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01301_ ) );
AOI211_X1 _17132_ ( .A(_01300_ ), .B(_01301_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_00817_ ), .ZN(_01302_ ) );
NAND3_X1 _17133_ ( .A1(_00809_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01303_ ) );
NAND4_X1 _17134_ ( .A1(_01302_ ), .A2(_00819_ ), .A3(_00820_ ), .A4(_01303_ ), .ZN(_01304_ ) );
NAND3_X1 _17135_ ( .A1(_00823_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01305_ ) );
NAND3_X1 _17136_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01306_ ) );
AND2_X1 _17137_ ( .A1(_01305_ ), .A2(_01306_ ), .ZN(_01307_ ) );
NAND3_X1 _17138_ ( .A1(_00811_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01308_ ) );
NAND3_X1 _17139_ ( .A1(_00830_ ), .A2(_00828_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01309_ ) );
NAND4_X1 _17140_ ( .A1(_01307_ ), .A2(_01154_ ), .A3(_01308_ ), .A4(_01309_ ), .ZN(_01310_ ) );
NAND3_X1 _17141_ ( .A1(_01304_ ), .A2(_00799_ ), .A3(_01310_ ), .ZN(_01311_ ) );
NAND2_X1 _17142_ ( .A1(_01299_ ), .A2(_01311_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI21_X1 _17143_ ( .A(_06079_ ), .B1(_05972_ ), .B2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _17144_ ( .A1(_06146_ ), .A2(\myifu.state [2] ), .A3(_06154_ ), .A4(_06151_ ), .ZN(_01312_ ) );
NOR2_X1 _17145_ ( .A1(_02096_ ), .A2(_00626_ ), .ZN(_01313_ ) );
INV_X1 _17146_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01314_ ) );
AOI21_X1 _17147_ ( .A(_00624_ ), .B1(_01313_ ), .B2(_01314_ ), .ZN(_01315_ ) );
AOI21_X1 _17148_ ( .A(fanout_net_6 ), .B1(_01312_ ), .B2(_01315_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17149_ ( .A1(_05390_ ), .A2(_06231_ ), .ZN(_01316_ ) );
NAND3_X1 _17150_ ( .A1(_01316_ ), .A2(_01314_ ), .A3(_02097_ ), .ZN(_01317_ ) );
OAI211_X1 _17151_ ( .A(_01317_ ), .B(_06074_ ), .C1(_01314_ ), .C2(_00626_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _17152_ ( .A1(_06155_ ), .A2(_01794_ ), .A3(\myifu.state [2] ), .ZN(_01318_ ) );
NAND3_X1 _17153_ ( .A1(_05390_ ), .A2(\io_master_arburst [0] ), .A3(_02145_ ), .ZN(_01319_ ) );
NAND2_X1 _17154_ ( .A1(_01318_ ), .A2(_01319_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _17155_ ( .A1(_06146_ ), .A2(\myifu.state [2] ), .A3(_06151_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17156_ ( .A1(_06369_ ), .A2(exception_quest_IDU ), .A3(_02256_ ), .ZN(_01320_ ) );
NOR3_X1 _17157_ ( .A1(_01320_ ), .A2(fanout_net_6 ), .A3(_02259_ ), .ZN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_B_$_MUX__Y_A_$_NOR__B_Y ) );
INV_X1 _17158_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01321_ ) );
NOR3_X1 _17159_ ( .A1(_01321_ ), .A2(_00746_ ), .A3(_00807_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
NOR3_X1 _17160_ ( .A1(_01321_ ), .A2(_00747_ ), .A3(_00807_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _17161_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00807_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17162_ ( .A1(\IF_ID_pc [4] ), .A2(_06228_ ), .A3(_06087_ ), .A4(_00807_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
NOR3_X1 _17163_ ( .A1(_01321_ ), .A2(_00744_ ), .A3(_00807_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17164_ ( .A1(_06078_ ), .A2(_06228_ ), .A3(\IF_ID_pc [3] ), .A4(_00807_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
AND3_X1 _17165_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06230_ ), .A3(_00807_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17166_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06230_ ), .A3(_00793_ ), .A4(_00795_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
AND3_X1 _17167_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06078_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
AND3_X1 _17168_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_06087_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
AND3_X1 _17169_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
AND3_X1 _17170_ ( .A1(_02144_ ), .A2(_06230_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
AOI21_X1 _17171_ ( .A(_00624_ ), .B1(\myidu.stall_quest_fencei ), .B2(\myifu.state [0] ), .ZN(_01322_ ) );
NAND3_X1 _17172_ ( .A1(_00626_ ), .A2(_05629_ ), .A3(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01323_ ) );
NAND3_X1 _17173_ ( .A1(_01322_ ), .A2(_05631_ ), .A3(_01323_ ), .ZN(_01324_ ) );
OR2_X1 _17174_ ( .A1(_01313_ ), .A2(_01324_ ), .ZN(_01325_ ) );
AOI221_X4 _17175_ ( .A(_01325_ ), .B1(\myifu.state [0] ), .B2(_01316_ ), .C1(_06155_ ), .C2(_02098_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17176_ ( .A1(_05953_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_05631_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
AOI211_X1 _17177_ ( .A(_05671_ ), .B(_00607_ ), .C1(_05415_ ), .C2(_05501_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
AOI211_X1 _17178_ ( .A(fanout_net_6 ), .B(_01324_ ), .C1(_02096_ ), .C2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _17179_ ( .A(_06162_ ), .B(_06218_ ), .S(\mylsu.state [0] ), .Z(_01326_ ) );
NOR2_X1 _17180_ ( .A1(_06297_ ), .A2(_01326_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17181_ ( .A1(_06297_ ), .A2(_04663_ ), .A3(_01326_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
AND2_X1 _17182_ ( .A1(_02129_ ), .A2(_06217_ ), .ZN(_01327_ ) );
AND2_X1 _17183_ ( .A1(_05393_ ), .A2(_06203_ ), .ZN(_01328_ ) );
NAND4_X1 _17184_ ( .A1(_05392_ ), .A2(\mylsu.state [0] ), .A3(_01327_ ), .A4(_01328_ ), .ZN(_01329_ ) );
AND2_X1 _17185_ ( .A1(_06146_ ), .A2(_06296_ ), .ZN(_01330_ ) );
OAI21_X1 _17186_ ( .A(_01329_ ), .B1(_06225_ ), .B2(_01330_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND2_X1 _17187_ ( .A1(_02277_ ), .A2(\mylsu.state [0] ), .ZN(_01331_ ) );
AND2_X1 _17188_ ( .A1(_01331_ ), .A2(_06203_ ), .ZN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
BUF_X2 _17189_ ( .A(_02132_ ), .Z(_01332_ ) );
OAI211_X1 _17190_ ( .A(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .B(_01332_ ), .C1(io_master_wready ), .C2(io_master_awready ), .ZN(_01333_ ) );
NOR3_X1 _17191_ ( .A1(_02133_ ), .A2(_02140_ ), .A3(_01333_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _17192_ ( .A1(_06169_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01334_ ) );
AND2_X1 _17193_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01335_ ) );
NOR3_X1 _17194_ ( .A1(_01335_ ), .A2(fanout_net_6 ), .A3(excp_written ), .ZN(_01336_ ) );
AND4_X1 _17195_ ( .A1(io_master_awready ), .A2(_01334_ ), .A3(_01332_ ), .A4(_01336_ ), .ZN(_01337_ ) );
NAND3_X1 _17196_ ( .A1(_02141_ ), .A2(\mylsu.state [0] ), .A3(_01337_ ), .ZN(_01338_ ) );
INV_X1 _17197_ ( .A(io_master_wready ), .ZN(_01339_ ) );
NAND3_X1 _17198_ ( .A1(_02279_ ), .A2(\mylsu.state [2] ), .A3(_01339_ ), .ZN(_01340_ ) );
NAND2_X1 _17199_ ( .A1(_01338_ ), .A2(_01340_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _17200_ ( .A1(_02132_ ), .A2(EXU_valid_LSU ), .A3(_01335_ ), .ZN(_01341_ ) );
NOR4_X1 _17201_ ( .A1(_02133_ ), .A2(_02140_ ), .A3(_03248_ ), .A4(_01341_ ), .ZN(_01342_ ) );
NAND2_X1 _17202_ ( .A1(_01342_ ), .A2(\mylsu.state [0] ), .ZN(_01343_ ) );
NAND3_X1 _17203_ ( .A1(_02279_ ), .A2(\mylsu.state [4] ), .A3(io_master_awready ), .ZN(_01344_ ) );
NAND3_X1 _17204_ ( .A1(_02278_ ), .A2(\mylsu.state [2] ), .A3(io_master_wready ), .ZN(_01345_ ) );
NAND3_X1 _17205_ ( .A1(_06303_ ), .A2(\mylsu.state [1] ), .A3(_02278_ ), .ZN(_01346_ ) );
NAND4_X1 _17206_ ( .A1(_01343_ ), .A2(_01344_ ), .A3(_01345_ ), .A4(_01346_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
AND2_X1 _17207_ ( .A1(_05395_ ), .A2(_01327_ ), .ZN(_01347_ ) );
AND4_X1 _17208_ ( .A1(_01339_ ), .A2(_01334_ ), .A3(_05398_ ), .A4(_02277_ ), .ZN(_01348_ ) );
AND3_X1 _17209_ ( .A1(_02141_ ), .A2(_01332_ ), .A3(_01348_ ), .ZN(_01349_ ) );
OAI21_X1 _17210_ ( .A(\mylsu.state [0] ), .B1(_01347_ ), .B2(_01349_ ), .ZN(_01350_ ) );
NAND4_X1 _17211_ ( .A1(_02125_ ), .A2(_05393_ ), .A3(_02126_ ), .A4(_06203_ ), .ZN(_01351_ ) );
AOI21_X1 _17212_ ( .A(_01351_ ), .B1(_02118_ ), .B2(_02122_ ), .ZN(_01352_ ) );
AND3_X1 _17213_ ( .A1(_06164_ ), .A2(_01334_ ), .A3(_05394_ ), .ZN(_01353_ ) );
OAI21_X1 _17214_ ( .A(_01331_ ), .B1(_01352_ ), .B2(_01353_ ), .ZN(_01354_ ) );
NAND4_X1 _17215_ ( .A1(_06146_ ), .A2(\mylsu.state [3] ), .A3(_02278_ ), .A4(_06296_ ), .ZN(_01355_ ) );
AND4_X1 _17216_ ( .A1(_02122_ ), .A2(_02118_ ), .A3(_02277_ ), .A4(_01328_ ), .ZN(_01356_ ) );
AND2_X1 _17217_ ( .A1(_02132_ ), .A2(EXU_valid_LSU ), .ZN(_01357_ ) );
NAND3_X1 _17218_ ( .A1(_01357_ ), .A2(_02127_ ), .A3(_06217_ ), .ZN(_01358_ ) );
NOR2_X1 _17219_ ( .A1(_01358_ ), .A2(_02140_ ), .ZN(_01359_ ) );
OAI21_X1 _17220_ ( .A(\mylsu.state [0] ), .B1(_01356_ ), .B2(_01359_ ), .ZN(_01360_ ) );
NAND4_X1 _17221_ ( .A1(_06299_ ), .A2(_06301_ ), .A3(\mylsu.state [1] ), .A4(_02277_ ), .ZN(_01361_ ) );
AND3_X1 _17222_ ( .A1(_01355_ ), .A2(_01360_ ), .A3(_01361_ ), .ZN(_01362_ ) );
NAND4_X1 _17223_ ( .A1(_02140_ ), .A2(\mylsu.state [0] ), .A3(_02278_ ), .A4(_01357_ ), .ZN(_01363_ ) );
OAI211_X1 _17224_ ( .A(\mylsu.state [0] ), .B(_02278_ ), .C1(_06169_ ), .C2(_06218_ ), .ZN(_01364_ ) );
AND3_X1 _17225_ ( .A1(_01363_ ), .A2(_02278_ ), .A3(_01364_ ), .ZN(_01365_ ) );
NAND4_X1 _17226_ ( .A1(_01350_ ), .A2(_01354_ ), .A3(_01362_ ), .A4(_01365_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
AND3_X1 _17227_ ( .A1(_01357_ ), .A2(io_master_wready ), .A3(_05398_ ), .ZN(_01366_ ) );
NAND3_X1 _17228_ ( .A1(_02141_ ), .A2(_01331_ ), .A3(_01366_ ), .ZN(_01367_ ) );
NAND2_X1 _17229_ ( .A1(_02279_ ), .A2(\mylsu.state [4] ), .ZN(_01368_ ) );
AOI21_X1 _17230_ ( .A(io_master_awready ), .B1(_01367_ ), .B2(_01368_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
BUF_X4 _17231_ ( .A(_06170_ ), .Z(_01369_ ) );
BUF_X4 _17232_ ( .A(_01369_ ), .Z(_01370_ ) );
AOI21_X1 _17233_ ( .A(\EX_LS_pc [21] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01371_ ) );
MUX2_X1 _17234_ ( .A(\LS_WB_wdata_csreg [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_02331_ ), .Z(_01372_ ) );
NOR3_X1 _17235_ ( .A1(_06165_ ), .A2(_06171_ ), .A3(_01372_ ), .ZN(_01373_ ) );
NOR2_X1 _17236_ ( .A1(_01371_ ), .A2(_01373_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
AOI21_X1 _17237_ ( .A(\EX_LS_pc [20] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01374_ ) );
OAI21_X1 _17238_ ( .A(_01369_ ), .B1(_04712_ ), .B2(_06325_ ), .ZN(_01375_ ) );
AOI221_X4 _17239_ ( .A(_01375_ ), .B1(\LS_WB_wdata_csreg [20] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_01332_ ), .ZN(_01376_ ) );
NOR2_X1 _17240_ ( .A1(_01374_ ), .A2(_01376_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _17241_ ( .A(\LS_WB_wdata_csreg [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_04715_ ), .Z(_01377_ ) );
MUX2_X1 _17242_ ( .A(_01377_ ), .B(\EX_LS_pc [19] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
BUF_X4 _17243_ ( .A(_02331_ ), .Z(_01378_ ) );
MUX2_X1 _17244_ ( .A(\LS_WB_wdata_csreg [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_01378_ ), .Z(_01379_ ) );
MUX2_X1 _17245_ ( .A(_01379_ ), .B(\EX_LS_pc [18] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
AOI21_X1 _17246_ ( .A(\EX_LS_pc [17] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01380_ ) );
OAI21_X1 _17247_ ( .A(_01369_ ), .B1(_04712_ ), .B2(_06477_ ), .ZN(_01381_ ) );
AOI221_X4 _17248_ ( .A(_01381_ ), .B1(\LS_WB_wdata_csreg [17] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_01332_ ), .ZN(_01382_ ) );
NOR2_X1 _17249_ ( .A1(_01380_ ), .A2(_01382_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
AOI21_X1 _17250_ ( .A(\EX_LS_pc [16] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01383_ ) );
MUX2_X1 _17251_ ( .A(\LS_WB_wdata_csreg [16] ), .B(\EX_LS_result_csreg_mem [16] ), .S(_02331_ ), .Z(_01384_ ) );
NOR3_X1 _17252_ ( .A1(_06165_ ), .A2(_06171_ ), .A3(_01384_ ), .ZN(_01385_ ) );
NOR2_X1 _17253_ ( .A1(_01383_ ), .A2(_01385_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
AOI21_X1 _17254_ ( .A(\EX_LS_pc [15] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01386_ ) );
OAI21_X1 _17255_ ( .A(_01369_ ), .B1(_04712_ ), .B2(_06342_ ), .ZN(_01387_ ) );
AOI221_X4 _17256_ ( .A(_01387_ ), .B1(\LS_WB_wdata_csreg [15] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_01332_ ), .ZN(_01388_ ) );
NOR2_X1 _17257_ ( .A1(_01386_ ), .A2(_01388_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _17258_ ( .A(\LS_WB_wdata_csreg [14] ), .B(\EX_LS_result_csreg_mem [14] ), .S(_01378_ ), .Z(_01389_ ) );
MUX2_X1 _17259_ ( .A(_01389_ ), .B(\EX_LS_pc [14] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _17260_ ( .A(\LS_WB_wdata_csreg [13] ), .B(\EX_LS_result_csreg_mem [13] ), .S(_01378_ ), .Z(_01390_ ) );
MUX2_X1 _17261_ ( .A(_01390_ ), .B(\EX_LS_pc [13] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
AOI21_X1 _17262_ ( .A(\EX_LS_pc [12] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01391_ ) );
OAI21_X1 _17263_ ( .A(_01369_ ), .B1(_04712_ ), .B2(_06326_ ), .ZN(_01392_ ) );
AOI221_X4 _17264_ ( .A(_01392_ ), .B1(\LS_WB_wdata_csreg [12] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_01332_ ), .ZN(_01393_ ) );
NOR2_X1 _17265_ ( .A1(_01391_ ), .A2(_01393_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
MUX2_X1 _17266_ ( .A(\LS_WB_wdata_csreg [30] ), .B(\EX_LS_result_csreg_mem [30] ), .S(_01378_ ), .Z(_01394_ ) );
MUX2_X1 _17267_ ( .A(_01394_ ), .B(\EX_LS_pc [30] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _17268_ ( .A(\LS_WB_wdata_csreg [11] ), .B(\EX_LS_result_csreg_mem [11] ), .S(_01378_ ), .Z(_01395_ ) );
MUX2_X1 _17269_ ( .A(_01395_ ), .B(\EX_LS_pc [11] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _17270_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_01378_ ), .Z(_01396_ ) );
MUX2_X1 _17271_ ( .A(_01396_ ), .B(\EX_LS_pc [10] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _17272_ ( .A(\LS_WB_wdata_csreg [9] ), .B(\EX_LS_result_csreg_mem [9] ), .S(_01378_ ), .Z(_01397_ ) );
MUX2_X1 _17273_ ( .A(_01397_ ), .B(\EX_LS_pc [9] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _17274_ ( .A(\LS_WB_wdata_csreg [8] ), .B(\EX_LS_result_csreg_mem [8] ), .S(_01378_ ), .Z(_01398_ ) );
MUX2_X1 _17275_ ( .A(_01398_ ), .B(\EX_LS_pc [8] ), .S(_06173_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _17276_ ( .A(\LS_WB_wdata_csreg [7] ), .B(\EX_LS_result_csreg_mem [7] ), .S(_01378_ ), .Z(_01399_ ) );
BUF_X4 _17277_ ( .A(_06172_ ), .Z(_01400_ ) );
MUX2_X1 _17278_ ( .A(_01399_ ), .B(\EX_LS_pc [7] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
AOI21_X1 _17279_ ( .A(\EX_LS_pc [6] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01401_ ) );
OAI21_X1 _17280_ ( .A(_01369_ ), .B1(_04712_ ), .B2(_06318_ ), .ZN(_01402_ ) );
AOI221_X4 _17281_ ( .A(_01402_ ), .B1(\LS_WB_wdata_csreg [6] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_01332_ ), .ZN(_01403_ ) );
NOR2_X1 _17282_ ( .A1(_01401_ ), .A2(_01403_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
AOI21_X1 _17283_ ( .A(\EX_LS_pc [5] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01404_ ) );
OAI21_X1 _17284_ ( .A(_01369_ ), .B1(_04712_ ), .B2(_06308_ ), .ZN(_01405_ ) );
AOI221_X4 _17285_ ( .A(_01405_ ), .B1(\LS_WB_wdata_csreg [5] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_01332_ ), .ZN(_01406_ ) );
NOR2_X1 _17286_ ( .A1(_01404_ ), .A2(_01406_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
OAI22_X1 _17287_ ( .A1(_04713_ ), .A2(_05133_ ), .B1(_02232_ ), .B2(\EX_LS_flag [2] ), .ZN(_01407_ ) );
MUX2_X1 _17288_ ( .A(_01407_ ), .B(\EX_LS_pc [4] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _17289_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\EX_LS_result_csreg_mem [3] ), .S(_01378_ ), .Z(_01408_ ) );
MUX2_X1 _17290_ ( .A(_01408_ ), .B(\EX_LS_pc [3] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
MUX2_X1 _17291_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\EX_LS_result_csreg_mem [2] ), .S(_02331_ ), .Z(_01409_ ) );
MUX2_X1 _17292_ ( .A(_01409_ ), .B(\EX_LS_pc [2] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
OAI22_X1 _17293_ ( .A1(_04713_ ), .A2(_06629_ ), .B1(_02224_ ), .B2(\EX_LS_flag [2] ), .ZN(_01410_ ) );
MUX2_X1 _17294_ ( .A(_01410_ ), .B(\EX_LS_pc [29] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
OAI22_X1 _17295_ ( .A1(_04713_ ), .A2(_06309_ ), .B1(_02236_ ), .B2(\EX_LS_flag [2] ), .ZN(_01411_ ) );
MUX2_X1 _17296_ ( .A(_01411_ ), .B(\EX_LS_pc [1] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI21_X1 _17297_ ( .A(\EX_LS_pc [0] ), .B1(_06215_ ), .B2(_01370_ ), .ZN(_01412_ ) );
OAI21_X1 _17298_ ( .A(_01369_ ), .B1(_04712_ ), .B2(_06310_ ), .ZN(_01413_ ) );
AOI221_X4 _17299_ ( .A(_01413_ ), .B1(\LS_WB_wdata_csreg [0] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_01332_ ), .ZN(_01414_ ) );
NOR2_X1 _17300_ ( .A1(_01412_ ), .A2(_01414_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
NAND3_X1 _17301_ ( .A1(_05397_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_result_csreg_mem [28] ), .ZN(_01415_ ) );
OAI21_X1 _17302_ ( .A(_01415_ ), .B1(_02235_ ), .B2(\EX_LS_flag [2] ), .ZN(_01416_ ) );
MUX2_X1 _17303_ ( .A(_01416_ ), .B(\EX_LS_pc [28] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _17304_ ( .A(\LS_WB_wdata_csreg [27] ), .B(\EX_LS_result_csreg_mem [27] ), .S(_02331_ ), .Z(_01417_ ) );
MUX2_X1 _17305_ ( .A(_01417_ ), .B(\EX_LS_pc [27] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI221_X4 _17306_ ( .A(_06172_ ), .B1(\LS_WB_wdata_csreg [26] ), .B2(_05377_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [26] ), .ZN(_01418_ ) );
AOI21_X1 _17307_ ( .A(\EX_LS_pc [26] ), .B1(_06214_ ), .B2(_01369_ ), .ZN(_01419_ ) );
NOR2_X1 _17308_ ( .A1(_01418_ ), .A2(_01419_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
OAI22_X1 _17309_ ( .A1(_04713_ ), .A2(_05274_ ), .B1(_02240_ ), .B2(\EX_LS_flag [2] ), .ZN(_01420_ ) );
MUX2_X1 _17310_ ( .A(_01420_ ), .B(\EX_LS_pc [25] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _17311_ ( .A(\EX_LS_pc [24] ), .B1(_06214_ ), .B2(_01370_ ), .ZN(_01421_ ) );
OAI21_X1 _17312_ ( .A(_06170_ ), .B1(_04712_ ), .B2(_06719_ ), .ZN(_01422_ ) );
AOI221_X4 _17313_ ( .A(_01422_ ), .B1(\LS_WB_wdata_csreg [24] ), .B2(_05377_ ), .C1(_02258_ ), .C2(_02132_ ), .ZN(_01423_ ) );
NOR2_X1 _17314_ ( .A1(_01421_ ), .A2(_01423_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _17315_ ( .A(\LS_WB_wdata_csreg [23] ), .B(\EX_LS_result_csreg_mem [23] ), .S(_02331_ ), .Z(_01424_ ) );
MUX2_X1 _17316_ ( .A(_01424_ ), .B(\EX_LS_pc [23] ), .S(_01400_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
AOI21_X1 _17317_ ( .A(\EX_LS_pc [22] ), .B1(_06214_ ), .B2(_01369_ ), .ZN(_01425_ ) );
MUX2_X1 _17318_ ( .A(\LS_WB_wdata_csreg [22] ), .B(\EX_LS_result_csreg_mem [22] ), .S(_02331_ ), .Z(_01426_ ) );
NOR3_X1 _17319_ ( .A1(_06165_ ), .A2(_06171_ ), .A3(_01426_ ), .ZN(_01427_ ) );
NOR2_X1 _17320_ ( .A1(_01425_ ), .A2(_01427_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
OAI22_X1 _17321_ ( .A1(_04713_ ), .A2(_06741_ ), .B1(_01633_ ), .B2(\EX_LS_flag [2] ), .ZN(_01428_ ) );
MUX2_X1 _17322_ ( .A(_01428_ ), .B(\EX_LS_pc [31] ), .S(_06172_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X2 _17323_ ( .A1(_00670_ ), .A2(_06235_ ), .ZN(_01429_ ) );
NOR2_X1 _17324_ ( .A1(_06241_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01430_ ) );
NOR2_X2 _17325_ ( .A1(_00739_ ), .A2(_06235_ ), .ZN(_01431_ ) );
NOR2_X1 _17326_ ( .A1(_06238_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01432_ ) );
AOI22_X4 _17327_ ( .A1(_01429_ ), .A2(_01430_ ), .B1(_01431_ ), .B2(_01432_ ), .ZN(_01433_ ) );
NOR2_X1 _17328_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01434_ ) );
INV_X1 _17329_ ( .A(_01434_ ), .ZN(_01435_ ) );
OR3_X1 _17330_ ( .A1(_00699_ ), .A2(_06235_ ), .A3(_01435_ ), .ZN(_01436_ ) );
NAND4_X1 _17331_ ( .A1(_00629_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_05391_ ), .ZN(_01437_ ) );
AND3_X4 _17332_ ( .A1(_01433_ ), .A2(_01436_ ), .A3(_01437_ ), .ZN(_01438_ ) );
INV_X1 _17333_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01439_ ) );
AND2_X1 _17334_ ( .A1(_01439_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01440_ ) );
INV_X1 _17335_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_01441_ ) );
AND2_X2 _17336_ ( .A1(_01440_ ), .A2(_01441_ ), .ZN(_01442_ ) );
INV_X2 _17337_ ( .A(_01442_ ), .ZN(_01443_ ) );
NOR2_X4 _17338_ ( .A1(_01438_ ), .A2(_01443_ ), .ZN(_01444_ ) );
NOR2_X1 _17339_ ( .A1(_01444_ ), .A2(_06162_ ), .ZN(_01445_ ) );
OR3_X1 _17340_ ( .A1(_00670_ ), .A2(_06234_ ), .A3(_01435_ ), .ZN(_01446_ ) );
NAND3_X1 _17341_ ( .A1(_00629_ ), .A2(_05391_ ), .A3(_01435_ ), .ZN(_01447_ ) );
NAND2_X2 _17342_ ( .A1(_01446_ ), .A2(_01447_ ), .ZN(_01448_ ) );
AND2_X2 _17343_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01449_ ) );
AND2_X1 _17344_ ( .A1(_01449_ ), .A2(_01439_ ), .ZN(_01450_ ) );
BUF_X4 _17345_ ( .A(_01450_ ), .Z(_01451_ ) );
INV_X1 _17346_ ( .A(_01451_ ), .ZN(_01452_ ) );
NOR2_X2 _17347_ ( .A1(_01448_ ), .A2(_01452_ ), .ZN(_01453_ ) );
NAND2_X1 _17348_ ( .A1(_01441_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01454_ ) );
NOR2_X1 _17349_ ( .A1(_01454_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01455_ ) );
OR2_X1 _17350_ ( .A1(_01442_ ), .A2(_01455_ ), .ZN(_01456_ ) );
NOR2_X4 _17351_ ( .A1(_01453_ ), .A2(_01456_ ), .ZN(_01457_ ) );
BUF_X8 _17352_ ( .A(_01457_ ), .Z(_01458_ ) );
NAND3_X1 _17353_ ( .A1(_00644_ ), .A2(_00650_ ), .A3(\io_master_arid [1] ), .ZN(_01459_ ) );
AND2_X2 _17354_ ( .A1(_01449_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01460_ ) );
NOR2_X1 _17355_ ( .A1(_01459_ ), .A2(_01460_ ), .ZN(_01461_ ) );
BUF_X4 _17356_ ( .A(_01451_ ), .Z(_01462_ ) );
OAI21_X1 _17357_ ( .A(_01458_ ), .B1(_01461_ ), .B2(_01462_ ), .ZN(_01463_ ) );
BUF_X4 _17358_ ( .A(_06162_ ), .Z(_01464_ ) );
AOI22_X1 _17359_ ( .A1(_01445_ ), .A2(_01463_ ), .B1(_01464_ ), .B2(_03774_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
NAND3_X1 _17360_ ( .A1(_00651_ ), .A2(_00654_ ), .A3(_06281_ ), .ZN(_01465_ ) );
NOR2_X1 _17361_ ( .A1(_01465_ ), .A2(_01460_ ), .ZN(_01466_ ) );
OAI21_X1 _17362_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01466_ ), .ZN(_01467_ ) );
BUF_X4 _17363_ ( .A(_01443_ ), .Z(_01468_ ) );
BUF_X4 _17364_ ( .A(_01438_ ), .Z(_01469_ ) );
OAI21_X1 _17365_ ( .A(_01467_ ), .B1(_01468_ ), .B2(_01469_ ), .ZN(_01470_ ) );
MUX2_X1 _17366_ ( .A(\EX_LS_result_reg [20] ), .B(_01470_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _17367_ ( .A1(_00655_ ), .A2(_00657_ ), .A3(\io_master_arid [1] ), .ZN(_01471_ ) );
NOR2_X1 _17368_ ( .A1(_01471_ ), .A2(_01460_ ), .ZN(_01472_ ) );
OAI21_X1 _17369_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01472_ ), .ZN(_01473_ ) );
AOI22_X1 _17370_ ( .A1(_01445_ ), .A2(_01473_ ), .B1(_01464_ ), .B2(_03804_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _17371_ ( .A1(_00658_ ), .A2(_00660_ ), .A3(_06281_ ), .ZN(_01474_ ) );
NOR2_X1 _17372_ ( .A1(_01474_ ), .A2(_01460_ ), .ZN(_01475_ ) );
OAI21_X1 _17373_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01475_ ), .ZN(_01476_ ) );
OAI21_X1 _17374_ ( .A(_01476_ ), .B1(_01468_ ), .B2(_01469_ ), .ZN(_01477_ ) );
MUX2_X1 _17375_ ( .A(\EX_LS_result_reg [18] ), .B(_01477_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _17376_ ( .A1(_00662_ ), .A2(_00664_ ), .A3(\io_master_arid [1] ), .ZN(_01478_ ) );
NOR2_X1 _17377_ ( .A1(_01478_ ), .A2(_01460_ ), .ZN(_01479_ ) );
OAI21_X1 _17378_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01479_ ), .ZN(_01480_ ) );
AOI22_X1 _17379_ ( .A1(_01445_ ), .A2(_01480_ ), .B1(_01464_ ), .B2(_03874_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _17380_ ( .A1(_00665_ ), .A2(_00667_ ), .A3(_06281_ ), .ZN(_01481_ ) );
NOR2_X1 _17381_ ( .A1(_01481_ ), .A2(_01460_ ), .ZN(_01482_ ) );
OAI21_X1 _17382_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01482_ ), .ZN(_01483_ ) );
OAI21_X1 _17383_ ( .A(_01483_ ), .B1(_01468_ ), .B2(_01469_ ), .ZN(_01484_ ) );
MUX2_X1 _17384_ ( .A(\EX_LS_result_reg [16] ), .B(_01484_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
NOR3_X1 _17385_ ( .A1(_01442_ ), .A2(_01449_ ), .A3(_01455_ ), .ZN(_01485_ ) );
NAND2_X1 _17386_ ( .A1(_01429_ ), .A2(_01485_ ), .ZN(_01486_ ) );
NAND2_X1 _17387_ ( .A1(_01448_ ), .A2(_01449_ ), .ZN(_01487_ ) );
OAI211_X1 _17388_ ( .A(_01486_ ), .B(_01487_ ), .C1(_01469_ ), .C2(_01443_ ), .ZN(_01488_ ) );
MUX2_X1 _17389_ ( .A(\EX_LS_result_reg [15] ), .B(_01488_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
NAND2_X1 _17390_ ( .A1(_01435_ ), .A2(_01449_ ), .ZN(_01489_ ) );
OR3_X1 _17391_ ( .A1(_00641_ ), .A2(_06236_ ), .A3(_01489_ ), .ZN(_01490_ ) );
INV_X1 _17392_ ( .A(_01455_ ), .ZN(_01491_ ) );
NAND3_X1 _17393_ ( .A1(_01443_ ), .A2(_01491_ ), .A3(_01489_ ), .ZN(_01492_ ) );
NOR2_X1 _17394_ ( .A1(_06235_ ), .A2(_01492_ ), .ZN(_01493_ ) );
NAND3_X1 _17395_ ( .A1(_00672_ ), .A2(_00674_ ), .A3(_01493_ ), .ZN(_01494_ ) );
OAI211_X1 _17396_ ( .A(_01490_ ), .B(_01494_ ), .C1(_01469_ ), .C2(_01443_ ), .ZN(_01495_ ) );
MUX2_X1 _17397_ ( .A(\EX_LS_result_reg [14] ), .B(_01495_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17398_ ( .A1(_00675_ ), .A2(_00677_ ), .A3(_01493_ ), .ZN(_01496_ ) );
INV_X1 _17399_ ( .A(_01449_ ), .ZN(_01497_ ) );
NOR2_X1 _17400_ ( .A1(_01497_ ), .A2(_01434_ ), .ZN(_01498_ ) );
AND4_X1 _17401_ ( .A1(_05391_ ), .A2(_00683_ ), .A3(_00681_ ), .A4(_01498_ ), .ZN(_01499_ ) );
OR3_X4 _17402_ ( .A1(_01444_ ), .A2(_01496_ ), .A3(_01499_ ), .ZN(_01500_ ) );
MUX2_X2 _17403_ ( .A(\EX_LS_result_reg [13] ), .B(_01500_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _17404_ ( .A1(_00678_ ), .A2(_00680_ ), .A3(_01493_ ), .ZN(_01501_ ) );
NAND4_X1 _17405_ ( .A1(_00715_ ), .A2(_00717_ ), .A3(_06281_ ), .A4(_01498_ ), .ZN(_01502_ ) );
OAI211_X1 _17406_ ( .A(_01501_ ), .B(_01502_ ), .C1(_01469_ ), .C2(_01443_ ), .ZN(_01503_ ) );
MUX2_X1 _17407_ ( .A(\EX_LS_result_reg [12] ), .B(_01503_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
NOR3_X1 _17408_ ( .A1(_00641_ ), .A2(_06236_ ), .A3(_01449_ ), .ZN(_01504_ ) );
OAI21_X1 _17409_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01504_ ), .ZN(_01505_ ) );
OAI21_X1 _17410_ ( .A(_01505_ ), .B1(_01468_ ), .B2(_01469_ ), .ZN(_01506_ ) );
MUX2_X1 _17411_ ( .A(\EX_LS_result_reg [30] ), .B(_01506_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NAND4_X1 _17412_ ( .A1(_00725_ ), .A2(\io_master_arid [1] ), .A3(_00727_ ), .A4(_01498_ ), .ZN(_01507_ ) );
NAND3_X1 _17413_ ( .A1(_00685_ ), .A2(_00687_ ), .A3(_01493_ ), .ZN(_01508_ ) );
AND2_X1 _17414_ ( .A1(_01507_ ), .A2(_01508_ ), .ZN(_01509_ ) );
AOI22_X1 _17415_ ( .A1(_01445_ ), .A2(_01509_ ), .B1(_01464_ ), .B2(_04098_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
NAND3_X1 _17416_ ( .A1(_00688_ ), .A2(_00690_ ), .A3(_01493_ ), .ZN(_01510_ ) );
NAND4_X1 _17417_ ( .A1(_00728_ ), .A2(_00730_ ), .A3(_06281_ ), .A4(_01498_ ), .ZN(_01511_ ) );
OAI211_X1 _17418_ ( .A(_01510_ ), .B(_01511_ ), .C1(_01469_ ), .C2(_01443_ ), .ZN(_01512_ ) );
MUX2_X1 _17419_ ( .A(\EX_LS_result_reg [10] ), .B(_01512_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
NAND3_X1 _17420_ ( .A1(_00691_ ), .A2(_00693_ ), .A3(_01493_ ), .ZN(_01513_ ) );
NAND4_X1 _17421_ ( .A1(_00731_ ), .A2(_00733_ ), .A3(_06281_ ), .A4(_01498_ ), .ZN(_01514_ ) );
OAI211_X1 _17422_ ( .A(_01513_ ), .B(_01514_ ), .C1(_01469_ ), .C2(_01443_ ), .ZN(_01515_ ) );
MUX2_X1 _17423_ ( .A(\EX_LS_result_reg [9] ), .B(_01515_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _17424_ ( .A1(_00694_ ), .A2(_00696_ ), .A3(_01493_ ), .ZN(_01516_ ) );
NAND4_X1 _17425_ ( .A1(_00734_ ), .A2(_00736_ ), .A3(_06281_ ), .A4(_01498_ ), .ZN(_01517_ ) );
OAI211_X1 _17426_ ( .A(_01516_ ), .B(_01517_ ), .C1(_01469_ ), .C2(_01443_ ), .ZN(_01518_ ) );
MUX2_X1 _17427_ ( .A(\EX_LS_result_reg [8] ), .B(_01518_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
AND4_X1 _17428_ ( .A1(_01456_ ), .A2(_01433_ ), .A3(_01436_ ), .A4(_01437_ ), .ZN(_01519_ ) );
NOR2_X1 _17429_ ( .A1(_00699_ ), .A2(_06236_ ), .ZN(_01520_ ) );
OAI221_X1 _17430_ ( .A(\mylsu.state [3] ), .B1(_01520_ ), .B2(_01492_ ), .C1(_01431_ ), .C2(_01489_ ), .ZN(_01521_ ) );
OAI22_X1 _17431_ ( .A1(_01519_ ), .A2(_01521_ ), .B1(\mylsu.state [3] ), .B2(_03900_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
NOR4_X1 _17432_ ( .A1(_00742_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(_06238_ ), .A4(_06235_ ), .ZN(_01522_ ) );
NOR3_X1 _17433_ ( .A1(_00641_ ), .A2(_06235_ ), .A3(_01432_ ), .ZN(_01523_ ) );
OAI22_X1 _17434_ ( .A1(_01522_ ), .A2(_01523_ ), .B1(_06241_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01524_ ) );
NAND4_X1 _17435_ ( .A1(_00672_ ), .A2(_00674_ ), .A3(_05391_ ), .A4(_01430_ ), .ZN(_01525_ ) );
AOI21_X1 _17436_ ( .A(_01434_ ), .B1(_01524_ ), .B2(_01525_ ), .ZN(_01526_ ) );
NOR3_X2 _17437_ ( .A1(_00702_ ), .A2(_06235_ ), .A3(_01435_ ), .ZN(_01527_ ) );
OAI21_X1 _17438_ ( .A(_01442_ ), .B1(_01526_ ), .B2(_01527_ ), .ZN(_01528_ ) );
OAI21_X1 _17439_ ( .A(_01455_ ), .B1(_01526_ ), .B2(_01527_ ), .ZN(_01529_ ) );
NOR3_X1 _17440_ ( .A1(_00742_ ), .A2(_06235_ ), .A3(_01434_ ), .ZN(_01530_ ) );
OAI21_X1 _17441_ ( .A(_01460_ ), .B1(_01530_ ), .B2(_01527_ ), .ZN(_01531_ ) );
OR3_X1 _17442_ ( .A1(_00702_ ), .A2(_06235_ ), .A3(_01460_ ), .ZN(_01532_ ) );
AOI21_X1 _17443_ ( .A(_01451_ ), .B1(_01531_ ), .B2(_01532_ ), .ZN(_01533_ ) );
INV_X1 _17444_ ( .A(_01530_ ), .ZN(_01534_ ) );
INV_X1 _17445_ ( .A(_01527_ ), .ZN(_01535_ ) );
AOI21_X1 _17446_ ( .A(_01452_ ), .B1(_01534_ ), .B2(_01535_ ), .ZN(_01536_ ) );
OAI21_X1 _17447_ ( .A(_01491_ ), .B1(_01533_ ), .B2(_01536_ ), .ZN(_01537_ ) );
AND2_X1 _17448_ ( .A1(_01529_ ), .A2(_01537_ ), .ZN(_01538_ ) );
OAI21_X1 _17449_ ( .A(_01528_ ), .B1(_01538_ ), .B2(_01442_ ), .ZN(_01539_ ) );
MUX2_X1 _17450_ ( .A(\EX_LS_result_reg [6] ), .B(_01539_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NOR2_X1 _17451_ ( .A1(_01485_ ), .A2(_01434_ ), .ZN(_01540_ ) );
INV_X1 _17452_ ( .A(_01540_ ), .ZN(_01541_ ) );
AOI211_X1 _17453_ ( .A(_06162_ ), .B(_06236_ ), .C1(_00705_ ), .C2(_01541_ ), .ZN(_01542_ ) );
AND2_X2 _17454_ ( .A1(_01456_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01543_ ) );
NOR2_X1 _17455_ ( .A1(_01541_ ), .A2(_01543_ ), .ZN(_01544_ ) );
NAND2_X1 _17456_ ( .A1(_00856_ ), .A2(_01544_ ), .ZN(_01545_ ) );
AND3_X1 _17457_ ( .A1(_00681_ ), .A2(_00683_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01546_ ) );
OAI21_X1 _17458_ ( .A(_01543_ ), .B1(_00990_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01547_ ) );
OAI211_X1 _17459_ ( .A(_01542_ ), .B(_01545_ ), .C1(_01546_ ), .C2(_01547_ ), .ZN(_01548_ ) );
NAND2_X1 _17460_ ( .A1(_01464_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_01549_ ) );
NAND2_X1 _17461_ ( .A1(_01548_ ), .A2(_01549_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
AOI221_X4 _17462_ ( .A(_06161_ ), .B1(_00874_ ), .B2(_01544_ ), .C1(_00708_ ), .C2(_01541_ ), .ZN(_01550_ ) );
AND3_X1 _17463_ ( .A1(_00715_ ), .A2(_00717_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01551_ ) );
OAI21_X1 _17464_ ( .A(_01543_ ), .B1(_01006_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01552_ ) );
OAI211_X1 _17465_ ( .A(_01550_ ), .B(\io_master_arid [1] ), .C1(_01551_ ), .C2(_01552_ ), .ZN(_01553_ ) );
NAND2_X1 _17466_ ( .A1(_01464_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_01554_ ) );
NAND2_X1 _17467_ ( .A1(_01553_ ), .A2(_01554_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _17468_ ( .A1(_06162_ ), .A2(\EX_LS_result_reg [3] ), .ZN(_01555_ ) );
AOI211_X1 _17469_ ( .A(_06162_ ), .B(_06236_ ), .C1(_00891_ ), .C2(_01544_ ), .ZN(_01556_ ) );
NAND2_X1 _17470_ ( .A1(_00711_ ), .A2(_01541_ ), .ZN(_01557_ ) );
NAND2_X1 _17471_ ( .A1(_01556_ ), .A2(_01557_ ), .ZN(_01558_ ) );
NAND3_X1 _17472_ ( .A1(_00725_ ), .A2(\mylsu.araddr_tmp [1] ), .A3(_00727_ ), .ZN(_01559_ ) );
NAND3_X1 _17473_ ( .A1(_00685_ ), .A2(_06238_ ), .A3(_00687_ ), .ZN(_01560_ ) );
AND3_X1 _17474_ ( .A1(_01559_ ), .A2(_01560_ ), .A3(_01543_ ), .ZN(_01561_ ) );
OAI21_X1 _17475_ ( .A(_01555_ ), .B1(_01558_ ), .B2(_01561_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
NAND2_X1 _17476_ ( .A1(_06162_ ), .A2(\EX_LS_result_reg [2] ), .ZN(_01562_ ) );
AOI211_X1 _17477_ ( .A(_06162_ ), .B(_06236_ ), .C1(_00909_ ), .C2(_01544_ ), .ZN(_01563_ ) );
NAND2_X1 _17478_ ( .A1(_00714_ ), .A2(_01541_ ), .ZN(_01564_ ) );
NAND2_X1 _17479_ ( .A1(_01563_ ), .A2(_01564_ ), .ZN(_01565_ ) );
NAND3_X1 _17480_ ( .A1(_00728_ ), .A2(_00730_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01566_ ) );
NAND3_X1 _17481_ ( .A1(_00688_ ), .A2(_00690_ ), .A3(_06238_ ), .ZN(_01567_ ) );
AND3_X1 _17482_ ( .A1(_01566_ ), .A2(_01567_ ), .A3(_01543_ ), .ZN(_01568_ ) );
OAI21_X1 _17483_ ( .A(_01562_ ), .B1(_01565_ ), .B2(_01568_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
AND4_X1 _17484_ ( .A1(_06281_ ), .A2(_00681_ ), .A3(_00683_ ), .A4(_01497_ ), .ZN(_01569_ ) );
OAI21_X1 _17485_ ( .A(_01457_ ), .B1(_01451_ ), .B2(_01569_ ), .ZN(_01570_ ) );
OAI21_X1 _17486_ ( .A(_01570_ ), .B1(_01468_ ), .B2(_01438_ ), .ZN(_01571_ ) );
MUX2_X1 _17487_ ( .A(\EX_LS_result_reg [29] ), .B(_01571_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
AOI221_X4 _17488_ ( .A(_06161_ ), .B1(_00926_ ), .B2(_01544_ ), .C1(_00720_ ), .C2(_01541_ ), .ZN(_01572_ ) );
AND3_X1 _17489_ ( .A1(_00731_ ), .A2(_00733_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01573_ ) );
OAI21_X1 _17490_ ( .A(_01543_ ), .B1(_01063_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01574_ ) );
OAI211_X1 _17491_ ( .A(_01572_ ), .B(\io_master_arid [1] ), .C1(_01573_ ), .C2(_01574_ ), .ZN(_01575_ ) );
NAND2_X1 _17492_ ( .A1(_01464_ ), .A2(\EX_LS_result_reg [1] ), .ZN(_01576_ ) );
NAND2_X1 _17493_ ( .A1(_01575_ ), .A2(_01576_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
AOI221_X4 _17494_ ( .A(_06161_ ), .B1(_00942_ ), .B2(_01544_ ), .C1(_00723_ ), .C2(_01541_ ), .ZN(_01577_ ) );
AND3_X1 _17495_ ( .A1(_00734_ ), .A2(_00736_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01578_ ) );
OAI21_X1 _17496_ ( .A(_01543_ ), .B1(_00783_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01579_ ) );
OAI211_X1 _17497_ ( .A(_01577_ ), .B(\io_master_arid [1] ), .C1(_01578_ ), .C2(_01579_ ), .ZN(_01580_ ) );
OAI21_X1 _17498_ ( .A(_01580_ ), .B1(\mylsu.state [3] ), .B2(_04092_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
AND4_X1 _17499_ ( .A1(_05391_ ), .A2(_00715_ ), .A3(_00717_ ), .A4(_01497_ ), .ZN(_01581_ ) );
OAI21_X1 _17500_ ( .A(_01457_ ), .B1(_01451_ ), .B2(_01581_ ), .ZN(_01582_ ) );
OAI21_X1 _17501_ ( .A(_01582_ ), .B1(_01468_ ), .B2(_01438_ ), .ZN(_01583_ ) );
MUX2_X1 _17502_ ( .A(\EX_LS_result_reg [28] ), .B(_01583_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
AND4_X1 _17503_ ( .A1(\io_master_arid [1] ), .A2(_00725_ ), .A3(_00727_ ), .A4(_01497_ ), .ZN(_01584_ ) );
OAI21_X1 _17504_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01584_ ), .ZN(_01585_ ) );
AOI22_X1 _17505_ ( .A1(_01445_ ), .A2(_01585_ ), .B1(_01464_ ), .B2(_03557_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
AND4_X1 _17506_ ( .A1(_05391_ ), .A2(_00728_ ), .A3(_00730_ ), .A4(_01497_ ), .ZN(_01586_ ) );
OAI21_X1 _17507_ ( .A(_01457_ ), .B1(_01451_ ), .B2(_01586_ ), .ZN(_01587_ ) );
OAI21_X1 _17508_ ( .A(_01587_ ), .B1(_01468_ ), .B2(_01438_ ), .ZN(_01588_ ) );
MUX2_X1 _17509_ ( .A(\EX_LS_result_reg [26] ), .B(_01588_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
AND4_X1 _17510_ ( .A1(\io_master_arid [1] ), .A2(_00731_ ), .A3(_00733_ ), .A4(_01497_ ), .ZN(_01589_ ) );
OAI21_X1 _17511_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01589_ ), .ZN(_01590_ ) );
AOI22_X1 _17512_ ( .A1(_01445_ ), .A2(_01590_ ), .B1(_01464_ ), .B2(_03588_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
AND4_X1 _17513_ ( .A1(_05391_ ), .A2(_00734_ ), .A3(_00736_ ), .A4(_01497_ ), .ZN(_01591_ ) );
OAI21_X1 _17514_ ( .A(_01457_ ), .B1(_01451_ ), .B2(_01591_ ), .ZN(_01592_ ) );
OAI21_X1 _17515_ ( .A(_01592_ ), .B1(_01468_ ), .B2(_01438_ ), .ZN(_01593_ ) );
MUX2_X1 _17516_ ( .A(\EX_LS_result_reg [24] ), .B(_01593_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _17517_ ( .A1(_00739_ ), .A2(_06236_ ), .A3(_01449_ ), .ZN(_01594_ ) );
OAI21_X1 _17518_ ( .A(_01458_ ), .B1(_01462_ ), .B2(_01594_ ), .ZN(_01595_ ) );
AOI22_X1 _17519_ ( .A1(_01445_ ), .A2(_01595_ ), .B1(_01464_ ), .B2(_03704_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _17520_ ( .A1(_00742_ ), .A2(_06236_ ), .A3(_01449_ ), .ZN(_01596_ ) );
OAI21_X1 _17521_ ( .A(_01457_ ), .B1(_01451_ ), .B2(_01596_ ), .ZN(_01597_ ) );
OAI21_X1 _17522_ ( .A(_01597_ ), .B1(_01468_ ), .B2(_01438_ ), .ZN(_01598_ ) );
MUX2_X1 _17523_ ( .A(\EX_LS_result_reg [22] ), .B(_01598_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17524_ ( .A1(_00629_ ), .A2(_06281_ ), .A3(_01497_ ), .ZN(_01599_ ) );
OAI21_X1 _17525_ ( .A(_01457_ ), .B1(_01451_ ), .B2(_01599_ ), .ZN(_01600_ ) );
OAI21_X1 _17526_ ( .A(_01600_ ), .B1(_01468_ ), .B2(_01438_ ), .ZN(_01601_ ) );
MUX2_X1 _17527_ ( .A(\EX_LS_result_reg [31] ), .B(_01601_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17528_ ( .A1(\LS_WB_waddr_reg [1] ), .A2(\LS_WB_waddr_reg [0] ), .ZN(_01602_ ) );
INV_X1 _17529_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01603_ ) );
INV_X1 _17530_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01604_ ) );
NAND3_X1 _17531_ ( .A1(_01602_ ), .A2(_01603_ ), .A3(_01604_ ), .ZN(_01605_ ) );
AND2_X1 _17532_ ( .A1(_01634_ ), .A2(LS_WB_wen_reg ), .ZN(_01606_ ) );
NAND2_X1 _17533_ ( .A1(_01605_ ), .A2(_01606_ ), .ZN(_01607_ ) );
BUF_X4 _17534_ ( .A(_01607_ ), .Z(_01608_ ) );
INV_X1 _17535_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01609_ ) );
INV_X1 _17536_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01610_ ) );
AOI21_X1 _17537_ ( .A(_01608_ ), .B1(_01609_ ), .B2(_01610_ ), .ZN(_01611_ ) );
NOR2_X1 _17538_ ( .A1(_01608_ ), .A2(_01604_ ), .ZN(_01612_ ) );
NOR4_X1 _17539_ ( .A1(_01611_ ), .A2(_01612_ ), .A3(_01603_ ), .A4(_01608_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
NOR2_X1 _17540_ ( .A1(_01607_ ), .A2(_01603_ ), .ZN(_01613_ ) );
NOR2_X1 _17541_ ( .A1(_01608_ ), .A2(_01610_ ), .ZN(_01614_ ) );
AND4_X1 _17542_ ( .A1(_01604_ ), .A2(_01613_ ), .A3(_01614_ ), .A4(_01609_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
AOI21_X1 _17543_ ( .A(_01608_ ), .B1(_01603_ ), .B2(_01604_ ), .ZN(_01615_ ) );
NOR4_X1 _17544_ ( .A1(_01615_ ), .A2(_01614_ ), .A3(_01609_ ), .A4(_01608_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR4_X1 _17545_ ( .A1(_01615_ ), .A2(_01609_ ), .A3(_01610_ ), .A4(_01608_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
NOR4_X1 _17546_ ( .A1(_01611_ ), .A2(_01613_ ), .A3(_01604_ ), .A4(_01608_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
AND4_X1 _17547_ ( .A1(_01603_ ), .A2(_01612_ ), .A3(_01614_ ), .A4(_01609_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR2_X1 _17548_ ( .A1(_01607_ ), .A2(_01609_ ), .ZN(_01616_ ) );
AND4_X1 _17549_ ( .A1(_01603_ ), .A2(_01612_ ), .A3(_01616_ ), .A4(_01610_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17550_ ( .A1(_01604_ ), .A2(_01613_ ), .A3(_01616_ ), .A4(_01610_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17551_ ( .A1(_01604_ ), .A2(_01613_ ), .A3(_01616_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _17552_ ( .A1(_01611_ ), .A2(_01603_ ), .A3(_01604_ ), .A4(_01608_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17553_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01613_ ), .A3(_01614_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17554_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01613_ ), .A3(_01614_ ), .A4(_01609_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17555_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01613_ ), .A3(_01616_ ), .A4(_01610_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
CLKBUF_X1 _17556_ ( .A(fanout_net_6 ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
NOR4_X1 _17557_ ( .A1(_01615_ ), .A2(_01616_ ), .A3(_01610_ ), .A4(_01608_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
AND4_X1 _17558_ ( .A1(_01603_ ), .A2(_01612_ ), .A3(_01616_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17559_ ( .A1(_02099_ ), .A2(_01794_ ), .A3(_02148_ ), .ZN(_01617_ ) );
NAND2_X1 _17560_ ( .A1(_01617_ ), .A2(_01794_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17561_ ( .A(fanout_net_6 ), .B(_02099_ ), .C1(_02100_ ), .C2(_06243_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17562_ ( .A(_01605_ ), .Z(_01618_ ) );
CLKBUF_X2 _17563_ ( .A(_01606_ ), .Z(_01619_ ) );
AND3_X1 _17564_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17565_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17566_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17567_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17568_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17569_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17570_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17571_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17572_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17573_ ( .A1(_01618_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01619_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17574_ ( .A(_01605_ ), .Z(_01620_ ) );
CLKBUF_X2 _17575_ ( .A(_01606_ ), .Z(_01621_ ) );
AND3_X1 _17576_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17577_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17578_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17579_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17580_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17581_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17582_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17583_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17584_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17585_ ( .A1(_01620_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01621_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17586_ ( .A(_01605_ ), .Z(_01622_ ) );
CLKBUF_X2 _17587_ ( .A(_01606_ ), .Z(_01623_ ) );
AND3_X1 _17588_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17589_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17590_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17591_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17592_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17593_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17594_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17595_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17596_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17597_ ( .A1(_01622_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01623_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17598_ ( .A1(_01605_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01606_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17599_ ( .A1(_01605_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01606_ ), .ZN(\myreg.Reg[5]_$_DFFE_PP__Q_D ) );
AND3_X1 _17600_ ( .A1(_01794_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17601_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01624_ ) );
AND2_X1 _17602_ ( .A1(_01624_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01625_ ) );
INV_X1 _17603_ ( .A(_01625_ ), .ZN(_01626_ ) );
NOR2_X1 _17604_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01627_ ) );
OAI211_X1 _17605_ ( .A(_01634_ ), .B(\mysc.state [0] ), .C1(_01626_ ), .C2(_01627_ ), .ZN(_01628_ ) );
INV_X1 _17606_ ( .A(_01628_ ), .ZN(_01629_ ) );
OR3_X1 _17607_ ( .A1(_01629_ ), .A2(fanout_net_6 ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17608_ ( .A1(_01626_ ), .A2(fanout_net_6 ), .A3(_01627_ ), .ZN(_01630_ ) );
NAND2_X1 _17609_ ( .A1(_01630_ ), .A2(\mysc.state [0] ), .ZN(_01631_ ) );
OR3_X1 _17610_ ( .A1(_06227_ ), .A2(fanout_net_6 ), .A3(\mylsu.previous_load_done ), .ZN(_01632_ ) );
NAND2_X1 _17611_ ( .A1(_01631_ ), .A2(_01632_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17612_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_08042_ ) );
CLKGATE_X1 _17613_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08043_ ) );
CLKGATE_X1 _17614_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_08044_ ) );
CLKGATE_X1 _17615_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_08045_ ) );
CLKGATE_X1 _17616_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_08046_ ) );
CLKGATE_X1 _17617_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_08047_ ) );
CLKGATE_X1 _17618_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_08048_ ) );
CLKGATE_X1 _17619_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_08049_ ) );
CLKGATE_X1 _17620_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_08050_ ) );
CLKGATE_X1 _17621_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_08051_ ) );
CLKGATE_X1 _17622_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08052_ ) );
CLKGATE_X1 _17623_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08053_ ) );
CLKGATE_X1 _17624_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08054_ ) );
CLKGATE_X1 _17625_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08055_ ) );
CLKGATE_X1 _17626_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08056_ ) );
CLKGATE_X1 _17627_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08057_ ) );
CLKGATE_X1 _17628_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_08058_ ) );
CLKGATE_X1 _17629_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08059_ ) );
CLKGATE_X1 _17630_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_08060_ ) );
CLKGATE_X1 _17631_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ), .GCK(_08061_ ) );
CLKGATE_X1 _17632_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .GCK(_08062_ ) );
CLKGATE_X1 _17633_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08063_ ) );
CLKGATE_X1 _17634_ ( .CK(clock ), .E(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_08064_ ) );
CLKGATE_X1 _17635_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_08065_ ) );
CLKGATE_X1 _17636_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_08066_ ) );
CLKGATE_X1 _17637_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_08067_ ) );
CLKGATE_X1 _17638_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_08068_ ) );
CLKGATE_X1 _17639_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_08069_ ) );
CLKGATE_X1 _17640_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_08070_ ) );
CLKGATE_X1 _17641_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_08071_ ) );
CLKGATE_X1 _17642_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_08072_ ) );
CLKGATE_X1 _17643_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_08073_ ) );
CLKGATE_X1 _17644_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_08074_ ) );
CLKGATE_X1 _17645_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_08075_ ) );
CLKGATE_X1 _17646_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_08076_ ) );
CLKGATE_X1 _17647_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08077_ ) );
CLKGATE_X1 _17648_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08078_ ) );
CLKGATE_X1 _17649_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08079_ ) );
CLKGATE_X1 _17650_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08080_ ) );
CLKGATE_X1 _17651_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08081_ ) );
CLKGATE_X1 _17652_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_08082_ ) );
CLKGATE_X1 _17653_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08083_ ) );
CLKGATE_X1 _17654_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08084_ ) );
CLKGATE_X1 _17655_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08085_ ) );
CLKGATE_X1 _17656_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08086_ ) );
CLKGATE_X1 _17657_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_08087_ ) );
CLKGATE_X1 _17658_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08088_ ) );
CLKGATE_X1 _17659_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08089_ ) );
CLKGATE_X1 _17660_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_08090_ ) );
CLKGATE_X1 _17661_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08091_ ) );
CLKGATE_X1 _17662_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08092_ ) );
CLKGATE_X1 _17663_ ( .CK(clock ), .E(\myidu.state_$_DFF_P__Q_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__B_Y ), .GCK(_08093_ ) );
CLKGATE_X1 _17664_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_NOR__A_Y ), .GCK(_08094_ ) );
CLKGATE_X1 _17665_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08095_ ) );
CLKGATE_X1 _17666_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08096_ ) );
CLKGATE_X1 _17667_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08097_ ) );
CLKGATE_X1 _17668_ ( .CK(clock ), .E(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08098_ ) );
CLKGATE_X1 _17669_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_08099_ ) );
CLKGATE_X1 _17670_ ( .CK(clock ), .E(\mycsreg.excp_written_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08100_ ) );
CLKGATE_X1 _17671_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08101_ ) );
CLKGATE_X1 _17672_ ( .CK(clock ), .E(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_B_$_MUX__Y_A_$_NOR__B_Y ), .GCK(_08102_ ) );
CLKGATE_X1 _17673_ ( .CK(clock ), .E(\mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ), .GCK(_08103_ ) );
CLKGATE_X1 _17674_ ( .CK(clock ), .E(\mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ), .GCK(_08104_ ) );
CLKGATE_X1 _17675_ ( .CK(clock ), .E(\mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ), .GCK(_08105_ ) );
CLKGATE_X1 _17676_ ( .CK(clock ), .E(\mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ), .GCK(_08106_ ) );
LOGIC1_X1 _17677_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17678_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00064_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00065_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08435_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08434_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08433_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08432_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08431_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08430_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08429_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08428_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08427_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08426_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08425_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08424_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08423_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08422_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08421_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08420_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08419_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08418_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08417_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08416_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08415_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08414_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08413_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08412_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08411_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08410_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08409_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08408_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08407_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08406_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08405_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08106_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08404_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08105_ ), .Q(\mtvec [31] ), .QN(_08403_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08105_ ), .Q(\mtvec [30] ), .QN(_08402_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08105_ ), .Q(\mtvec [21] ), .QN(_08401_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08105_ ), .Q(\mtvec [20] ), .QN(_08400_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08105_ ), .Q(\mtvec [19] ), .QN(_08399_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08105_ ), .Q(\mtvec [18] ), .QN(_08398_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08105_ ), .Q(\mtvec [17] ), .QN(_08397_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08105_ ), .Q(\mtvec [16] ), .QN(_08396_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08105_ ), .Q(\mtvec [15] ), .QN(_08395_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08105_ ), .Q(\mtvec [14] ), .QN(_08394_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08105_ ), .Q(\mtvec [13] ), .QN(_08393_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08105_ ), .Q(\mtvec [12] ), .QN(_08392_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08105_ ), .Q(\mtvec [29] ), .QN(_08391_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08105_ ), .Q(\mtvec [11] ), .QN(_08390_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08105_ ), .Q(\mtvec [10] ), .QN(_08389_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08105_ ), .Q(\mtvec [9] ), .QN(_08388_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08105_ ), .Q(\mtvec [8] ), .QN(_08387_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08105_ ), .Q(\mtvec [7] ), .QN(_08386_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08105_ ), .Q(\mtvec [6] ), .QN(_08385_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08105_ ), .Q(\mtvec [5] ), .QN(_08384_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08105_ ), .Q(\mtvec [4] ), .QN(_08383_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08105_ ), .Q(\mtvec [3] ), .QN(_08382_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08105_ ), .Q(\mtvec [2] ), .QN(_08381_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08105_ ), .Q(\mtvec [28] ), .QN(_08380_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08105_ ), .Q(\mtvec [1] ), .QN(_08379_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08105_ ), .Q(\mtvec [0] ), .QN(_08378_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08105_ ), .Q(\mtvec [27] ), .QN(_08377_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08105_ ), .Q(\mtvec [26] ), .QN(_08376_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08105_ ), .Q(\mtvec [25] ), .QN(_08375_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08105_ ), .Q(\mtvec [24] ), .QN(_08374_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08105_ ), .Q(\mtvec [23] ), .QN(_08373_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08105_ ), .Q(\mtvec [22] ), .QN(_08372_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08104_ ), .Q(\mepc [31] ), .QN(_08371_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08104_ ), .Q(\mepc [30] ), .QN(_08370_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08104_ ), .Q(\mepc [21] ), .QN(_08369_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08104_ ), .Q(\mepc [20] ), .QN(_08368_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08104_ ), .Q(\mepc [19] ), .QN(_08367_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08104_ ), .Q(\mepc [18] ), .QN(_08366_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08104_ ), .Q(\mepc [17] ), .QN(_08365_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08104_ ), .Q(\mepc [16] ), .QN(_08364_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08104_ ), .Q(\mepc [15] ), .QN(_08363_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08104_ ), .Q(\mepc [14] ), .QN(_08362_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08104_ ), .Q(\mepc [13] ), .QN(_08361_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08104_ ), .Q(\mepc [12] ), .QN(_08360_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08104_ ), .Q(\mepc [29] ), .QN(_08359_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08104_ ), .Q(\mepc [11] ), .QN(_08358_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08104_ ), .Q(\mepc [10] ), .QN(_08357_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08104_ ), .Q(\mepc [9] ), .QN(_08356_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08104_ ), .Q(\mepc [8] ), .QN(_08355_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08104_ ), .Q(\mepc [7] ), .QN(_08354_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08104_ ), .Q(\mepc [6] ), .QN(_08353_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08104_ ), .Q(\mepc [5] ), .QN(_08352_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08104_ ), .Q(\mepc [4] ), .QN(_08351_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08104_ ), .Q(\mepc [3] ), .QN(_08350_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08104_ ), .Q(\mepc [2] ), .QN(_08349_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08104_ ), .Q(\mepc [28] ), .QN(_08348_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08104_ ), .Q(\mepc [1] ), .QN(_08347_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08104_ ), .Q(\mepc [0] ), .QN(_08346_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08104_ ), .Q(\mepc [27] ), .QN(_08345_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08104_ ), .Q(\mepc [26] ), .QN(_08344_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08104_ ), .Q(\mepc [25] ), .QN(_08343_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08104_ ), .Q(\mepc [24] ), .QN(_08342_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08104_ ), .Q(\mepc [23] ), .QN(_08341_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08104_ ), .Q(\mepc [22] ), .QN(_08340_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q ( .D(_00097_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08339_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_1 ( .D(_00098_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08338_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_10 ( .D(_00099_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08337_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_11 ( .D(_00100_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08336_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_12 ( .D(_00101_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08335_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_13 ( .D(_00102_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08334_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_14 ( .D(_00103_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08333_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_15 ( .D(_00104_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08332_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_16 ( .D(_00105_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08331_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_17 ( .D(_00106_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08330_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_18 ( .D(_00107_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08329_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_19 ( .D(_00108_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08328_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_2 ( .D(_00109_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08327_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_20 ( .D(_00110_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08326_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_21 ( .D(_00111_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08325_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_22 ( .D(_00112_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08324_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_23 ( .D(_00113_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08323_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_24 ( .D(_00114_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08322_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_25 ( .D(_00115_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08321_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_26 ( .D(_00116_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08320_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_27 ( .D(_00117_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08319_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_28 ( .D(_00118_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08318_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_29 ( .D(_00119_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08317_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_3 ( .D(_00120_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08316_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_30 ( .D(_00121_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08315_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_31 ( .D(_00122_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08314_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_4 ( .D(_00123_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08313_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_5 ( .D(_00124_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08312_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_6 ( .D(_00125_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08311_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_7 ( .D(_00126_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08310_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_8 ( .D(_00127_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08309_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_9 ( .D(_00128_ ), .CK(_08103_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08436_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PP0__Q ( .D(_00129_ ), .CK(clock ), .Q(excp_written ), .QN(_08437_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08308_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08438_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08439_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08440_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08441_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08442_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08443_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08444_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08445_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08446_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08447_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08448_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08449_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08450_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08451_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08452_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08453_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08454_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08455_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08456_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08457_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08458_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08459_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08460_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08461_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08462_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08463_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08464_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08465_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08466_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08467_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08102_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08307_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00130_ ), .CK(_08101_ ), .Q(\myec.state [1] ), .QN(_08306_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00131_ ), .CK(_08101_ ), .Q(\myec.state [0] ), .QN(_08468_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PP0__Q ( .D(_00132_ ), .CK(clock ), .Q(check_quest ), .QN(_08469_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08305_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08470_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08471_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08472_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08473_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08474_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08475_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08476_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08477_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08478_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08479_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08304_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00133_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08303_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00134_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08302_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00135_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08301_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00136_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08300_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00137_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08299_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00138_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08298_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00139_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08297_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00140_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08296_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00141_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08295_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00142_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08294_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00143_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08293_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00144_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08292_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00145_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08291_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00146_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08290_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00147_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08289_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00148_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08288_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00149_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08287_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00150_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08286_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00151_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08285_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00152_ ), .CK(_08100_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08284_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q ( .D(_00153_ ), .CK(_08099_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08283_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_1 ( .D(_00154_ ), .CK(_08099_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08282_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_2 ( .D(_00155_ ), .CK(_08099_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08281_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_3 ( .D(_00156_ ), .CK(_08099_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08280_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_4 ( .D(_00157_ ), .CK(_08099_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08279_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q ( .D(_00158_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [30] ), .QN(_08278_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_1 ( .D(_00159_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [29] ), .QN(_08277_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_10 ( .D(_00160_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [20] ), .QN(_08276_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_11 ( .D(_00161_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [19] ), .QN(_08275_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_12 ( .D(_00162_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [18] ), .QN(_08274_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_13 ( .D(_00163_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [17] ), .QN(_08273_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_14 ( .D(_00164_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [16] ), .QN(_08272_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_15 ( .D(_00165_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [15] ), .QN(_08271_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_16 ( .D(_00166_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [14] ), .QN(_08270_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_17 ( .D(_00167_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [13] ), .QN(_08269_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_18 ( .D(_00168_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [12] ), .QN(_08268_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_19 ( .D(_00169_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [11] ), .QN(_08267_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_2 ( .D(_00170_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [28] ), .QN(_08266_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_20 ( .D(_00171_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [10] ), .QN(_08265_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_21 ( .D(_00172_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [9] ), .QN(_08264_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_22 ( .D(_00173_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [8] ), .QN(_08263_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_23 ( .D(_00174_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [7] ), .QN(_08262_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_24 ( .D(_00175_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [6] ), .QN(_08261_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_25 ( .D(_00176_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [5] ), .QN(_08260_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_26 ( .D(_00177_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [4] ), .QN(_08259_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_27 ( .D(_00178_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [3] ), .QN(_08258_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_28 ( .D(_00179_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [2] ), .QN(_08257_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_29 ( .D(_00180_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [1] ), .QN(_08256_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_3 ( .D(_00181_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [27] ), .QN(_08255_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_30 ( .D(_00182_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [0] ), .QN(_08254_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_4 ( .D(_00183_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [26] ), .QN(_08253_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_5 ( .D(_00184_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [25] ), .QN(_08252_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_6 ( .D(_00185_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [24] ), .QN(_08251_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_7 ( .D(_00186_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [23] ), .QN(_08250_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_8 ( .D(_00187_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [22] ), .QN(_08249_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP0P__Q_9 ( .D(_00188_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [21] ), .QN(_08248_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PP1P__Q ( .D(_00189_ ), .CK(_08098_ ), .Q(\myexu.pc_jump [31] ), .QN(_08247_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q ( .D(_00190_ ), .CK(_08099_ ), .Q(\EX_LS_pc [31] ), .QN(_08246_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_1 ( .D(_00191_ ), .CK(_08099_ ), .Q(\EX_LS_pc [30] ), .QN(_08245_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_10 ( .D(_00192_ ), .CK(_08099_ ), .Q(\EX_LS_pc [21] ), .QN(_08244_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_11 ( .D(_00193_ ), .CK(_08099_ ), .Q(\EX_LS_pc [20] ), .QN(_08243_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_12 ( .D(_00194_ ), .CK(_08099_ ), .Q(\EX_LS_pc [19] ), .QN(_08242_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_13 ( .D(_00195_ ), .CK(_08099_ ), .Q(\EX_LS_pc [18] ), .QN(_08241_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_14 ( .D(_00196_ ), .CK(_08099_ ), .Q(\EX_LS_pc [17] ), .QN(_08240_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_15 ( .D(_00197_ ), .CK(_08099_ ), .Q(\EX_LS_pc [16] ), .QN(_08239_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_16 ( .D(_00198_ ), .CK(_08099_ ), .Q(\EX_LS_pc [15] ), .QN(_08238_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_17 ( .D(_00199_ ), .CK(_08099_ ), .Q(\EX_LS_pc [14] ), .QN(_08237_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_18 ( .D(_00200_ ), .CK(_08099_ ), .Q(\EX_LS_pc [13] ), .QN(_08236_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_19 ( .D(_00201_ ), .CK(_08099_ ), .Q(\EX_LS_pc [12] ), .QN(_08235_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_2 ( .D(_00202_ ), .CK(_08099_ ), .Q(\EX_LS_pc [29] ), .QN(_08234_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_20 ( .D(_00203_ ), .CK(_08099_ ), .Q(\EX_LS_pc [11] ), .QN(_08233_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_21 ( .D(_00204_ ), .CK(_08099_ ), .Q(\EX_LS_pc [10] ), .QN(_08232_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_22 ( .D(_00205_ ), .CK(_08099_ ), .Q(\EX_LS_pc [9] ), .QN(_08231_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_23 ( .D(_00206_ ), .CK(_08099_ ), .Q(\EX_LS_pc [8] ), .QN(_08230_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_24 ( .D(_00207_ ), .CK(_08099_ ), .Q(\EX_LS_pc [7] ), .QN(_08229_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_25 ( .D(_00208_ ), .CK(_08099_ ), .Q(\EX_LS_pc [6] ), .QN(_08228_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_26 ( .D(_00209_ ), .CK(_08099_ ), .Q(\EX_LS_pc [5] ), .QN(_08227_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_27 ( .D(_00210_ ), .CK(_08099_ ), .Q(\EX_LS_pc [4] ), .QN(_08226_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_28 ( .D(_00211_ ), .CK(_08099_ ), .Q(\EX_LS_pc [3] ), .QN(_08225_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_29 ( .D(_00212_ ), .CK(_08099_ ), .Q(\EX_LS_pc [2] ), .QN(_08224_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_3 ( .D(_00213_ ), .CK(_08099_ ), .Q(\EX_LS_pc [28] ), .QN(_08223_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_30 ( .D(_00214_ ), .CK(_08099_ ), .Q(\EX_LS_pc [1] ), .QN(_08222_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_31 ( .D(_00215_ ), .CK(_08099_ ), .Q(\EX_LS_pc [0] ), .QN(_08221_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_4 ( .D(_00216_ ), .CK(_08099_ ), .Q(\EX_LS_pc [27] ), .QN(_08220_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_5 ( .D(_00217_ ), .CK(_08099_ ), .Q(\EX_LS_pc [26] ), .QN(_08219_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_6 ( .D(_00218_ ), .CK(_08099_ ), .Q(\EX_LS_pc [25] ), .QN(_08218_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_7 ( .D(_00219_ ), .CK(_08099_ ), .Q(\EX_LS_pc [24] ), .QN(_08217_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_8 ( .D(_00220_ ), .CK(_08099_ ), .Q(\EX_LS_pc [23] ), .QN(_08216_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_9 ( .D(_00221_ ), .CK(_08099_ ), .Q(\EX_LS_pc [22] ), .QN(_08480_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08481_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08482_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08483_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08484_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08485_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08486_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08487_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08488_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08489_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08490_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08491_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08492_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08493_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08494_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08495_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08496_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08497_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08498_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08499_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08500_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08501_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08502_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08503_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08504_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08505_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08506_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08507_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08508_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08509_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08510_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08511_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08100_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08512_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08100_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PP0__Q ( .D(_00223_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q ( .D(_00222_ ), .CK(_08099_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_1 ( .D(_00224_ ), .CK(_08099_ ), .Q(\EX_LS_flag [1] ), .QN(_08215_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_2 ( .D(_00225_ ), .CK(_08099_ ), .Q(\EX_LS_flag [0] ), .QN(_08214_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_3 ( .D(_00226_ ), .CK(_08099_ ), .Q(\EX_LS_typ [4] ), .QN(_08213_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_4 ( .D(_00227_ ), .CK(_08099_ ), .Q(\EX_LS_typ [3] ), .QN(_08212_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_5 ( .D(_00228_ ), .CK(_08099_ ), .Q(\EX_LS_typ [2] ), .QN(_08211_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_6 ( .D(_00229_ ), .CK(_08099_ ), .Q(\EX_LS_typ [1] ), .QN(_08210_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_7 ( .D(_00230_ ), .CK(_08099_ ), .Q(\EX_LS_typ [0] ), .QN(_08209_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_08097_ ), .Q(\ID_EX_csr [11] ), .QN(_08208_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00232_ ), .CK(_08097_ ), .Q(\ID_EX_csr [10] ), .QN(_08207_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00233_ ), .CK(_08097_ ), .Q(\ID_EX_csr [1] ), .QN(_08206_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00234_ ), .CK(_08097_ ), .Q(\ID_EX_csr [0] ), .QN(_08205_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00235_ ), .CK(_08097_ ), .Q(\ID_EX_csr [9] ), .QN(_08204_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00236_ ), .CK(_08097_ ), .Q(\ID_EX_csr [8] ), .QN(_08203_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00237_ ), .CK(_08097_ ), .Q(\ID_EX_csr [7] ), .QN(_08202_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00238_ ), .CK(_08097_ ), .Q(\ID_EX_csr [6] ), .QN(_08201_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00239_ ), .CK(_08097_ ), .Q(\ID_EX_csr [5] ), .QN(_08200_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00240_ ), .CK(_08097_ ), .Q(\ID_EX_csr [4] ), .QN(_08199_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00241_ ), .CK(_08097_ ), .Q(\ID_EX_csr [3] ), .QN(_08198_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00242_ ), .CK(_08097_ ), .Q(\ID_EX_csr [2] ), .QN(_08197_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00243_ ), .CK(_08096_ ), .Q(exception_quest_IDU ), .QN(_08196_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00244_ ), .CK(_08095_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08094_ ), .Q(\ID_EX_imm [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08094_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08094_ ), .Q(\ID_EX_imm [21] ), .QN(_08513_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08094_ ), .Q(\ID_EX_imm [20] ), .QN(_08514_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08094_ ), .Q(\ID_EX_imm [19] ), .QN(_08515_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08094_ ), .Q(\ID_EX_imm [18] ), .QN(_08516_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08094_ ), .Q(\ID_EX_imm [17] ), .QN(_08517_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08094_ ), .Q(\ID_EX_imm [16] ), .QN(_08518_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08094_ ), .Q(\ID_EX_imm [15] ), .QN(_08519_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08094_ ), .Q(\ID_EX_imm [14] ), .QN(_08520_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08094_ ), .Q(\ID_EX_imm [13] ), .QN(_08521_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08094_ ), .Q(\ID_EX_imm [12] ), .QN(_08522_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08094_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08094_ ), .Q(\ID_EX_imm [11] ), .QN(_08523_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08094_ ), .Q(\ID_EX_imm [10] ), .QN(_08524_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08094_ ), .Q(\ID_EX_imm [9] ), .QN(_08525_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08094_ ), .Q(\ID_EX_imm [8] ), .QN(_08526_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08094_ ), .Q(\ID_EX_imm [7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08094_ ), .Q(\ID_EX_imm [6] ), .QN(_08527_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08094_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08094_ ), .Q(\ID_EX_imm [4] ), .QN(_08528_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08094_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08094_ ), .Q(\ID_EX_imm [2] ), .QN(_08529_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08094_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08094_ ), .Q(\ID_EX_imm [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08094_ ), .Q(\ID_EX_imm [0] ), .QN(_08530_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08094_ ), .Q(\ID_EX_imm [27] ), .QN(_08531_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08094_ ), .Q(\ID_EX_imm [26] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_4_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08094_ ), .Q(\ID_EX_imm [25] ), .QN(_08532_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08094_ ), .Q(\ID_EX_imm [24] ), .QN(_08533_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08094_ ), .Q(\ID_EX_imm [23] ), .QN(_08534_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08094_ ), .Q(\ID_EX_imm [22] ), .QN(_08535_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08093_ ), .Q(\ID_EX_pc [31] ), .QN(_08536_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08093_ ), .Q(\ID_EX_pc [30] ), .QN(_08537_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08093_ ), .Q(\ID_EX_pc [21] ), .QN(_08538_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08093_ ), .Q(\ID_EX_pc [20] ), .QN(_08539_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08093_ ), .Q(\ID_EX_pc [19] ), .QN(_08540_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08093_ ), .Q(\ID_EX_pc [18] ), .QN(_08541_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08093_ ), .Q(\ID_EX_pc [17] ), .QN(_08542_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08093_ ), .Q(\ID_EX_pc [16] ), .QN(_08543_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08093_ ), .Q(\ID_EX_pc [15] ), .QN(_08544_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08093_ ), .Q(\ID_EX_pc [14] ), .QN(_08545_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08093_ ), .Q(\ID_EX_pc [13] ), .QN(_08546_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08093_ ), .Q(\ID_EX_pc [12] ), .QN(_08547_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08093_ ), .Q(\ID_EX_pc [29] ), .QN(_08548_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08093_ ), .Q(\ID_EX_pc [11] ), .QN(_08549_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08093_ ), .Q(\ID_EX_pc [10] ), .QN(_08550_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08093_ ), .Q(\ID_EX_pc [9] ), .QN(_08551_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08093_ ), .Q(\ID_EX_pc [8] ), .QN(_08552_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08093_ ), .Q(\ID_EX_pc [7] ), .QN(_08553_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08093_ ), .Q(\ID_EX_pc [6] ), .QN(_08554_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08093_ ), .Q(\ID_EX_pc [5] ), .QN(_08555_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08093_ ), .Q(\ID_EX_pc [4] ), .QN(_08556_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08093_ ), .Q(\ID_EX_pc [3] ), .QN(_08557_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08093_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08093_ ), .Q(\ID_EX_pc [28] ), .QN(_08558_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08093_ ), .Q(\ID_EX_pc [1] ), .QN(_08559_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08093_ ), .Q(\ID_EX_pc [0] ), .QN(_08560_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08093_ ), .Q(\ID_EX_pc [27] ), .QN(_08561_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08093_ ), .Q(\ID_EX_pc [26] ), .QN(_08562_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08093_ ), .Q(\ID_EX_pc [25] ), .QN(_08563_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08093_ ), .Q(\ID_EX_pc [24] ), .QN(_08564_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08093_ ), .Q(\ID_EX_pc [23] ), .QN(_08565_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08093_ ), .Q(\ID_EX_pc [22] ), .QN(_08195_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_08092_ ), .Q(\ID_EX_rd [4] ), .QN(_08194_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_08092_ ), .Q(\ID_EX_rd [3] ), .QN(_08193_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00247_ ), .CK(_08092_ ), .Q(\ID_EX_rd [2] ), .QN(_08192_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00248_ ), .CK(_08092_ ), .Q(\ID_EX_rd [1] ), .QN(_08191_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00249_ ), .CK(_08092_ ), .Q(\ID_EX_rd [0] ), .QN(_08190_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00250_ ), .CK(_08091_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08189_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00251_ ), .CK(_08091_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08188_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00253_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08186_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00252_ ), .CK(_08091_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08187_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00255_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08184_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00254_ ), .CK(_08091_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08185_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00257_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08182_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00256_ ), .CK(_08091_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08183_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00259_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08180_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00258_ ), .CK(_08090_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08181_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00260_ ), .CK(_08090_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08179_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00262_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08177_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00261_ ), .CK(_08090_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08178_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00264_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08175_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00263_ ), .CK(_08090_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08176_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00266_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08173_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00265_ ), .CK(_08090_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08174_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00268_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08171_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00267_ ), .CK(_08089_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08172_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00269_ ), .CK(_08088_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08170_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08566_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00270_ ), .CK(_08087_ ), .Q(\ID_EX_typ [7] ), .QN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00271_ ), .CK(_08087_ ), .Q(\ID_EX_typ [6] ), .QN(_08169_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00272_ ), .CK(_08087_ ), .Q(\ID_EX_typ [5] ), .QN(_08168_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00273_ ), .CK(_08087_ ), .Q(\ID_EX_typ [4] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00274_ ), .CK(_08087_ ), .Q(\ID_EX_typ [3] ), .QN(_08167_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00275_ ), .CK(_08087_ ), .Q(\ID_EX_typ [2] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00276_ ), .CK(_08087_ ), .Q(\ID_EX_typ [1] ), .QN(_08166_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00277_ ), .CK(_08087_ ), .Q(\ID_EX_typ [0] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08086_ ), .Q(check_assert ), .QN(_08567_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08085_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08085_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08085_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08085_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08085_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08085_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08085_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08085_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08085_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08085_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08085_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08085_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08085_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08085_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08085_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08085_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08085_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08085_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08085_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08085_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08085_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08085_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08085_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08085_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08085_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08085_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08085_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08085_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08085_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08085_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08085_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08085_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08084_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08083_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08082_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08081_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08080_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08079_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08078_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08077_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08076_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08855_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08856_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08857_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08858_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08859_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08860_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08861_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08862_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08863_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08864_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08865_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08866_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08867_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08868_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08869_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08870_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08871_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08872_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08873_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08874_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08875_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08876_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08075_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08877_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08878_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08879_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08880_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08881_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08882_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08883_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08884_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08885_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08886_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08887_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08888_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08889_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08890_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08891_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08892_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08893_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08894_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08895_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08896_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08897_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08898_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08899_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08900_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08901_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08902_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08903_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08074_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08904_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08905_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08906_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08907_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08908_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08909_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08910_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08911_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08912_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08913_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08914_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08915_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08916_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08917_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08918_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08919_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08920_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08921_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08922_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08923_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08924_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08925_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08926_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08927_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08928_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08929_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08930_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08073_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08165_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00278_ ), .CK(_08072_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08164_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00279_ ), .CK(_08071_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08163_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00280_ ), .CK(_08070_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08931_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_08069_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08162_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00281_ ), .CK(_08068_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00282_ ), .CK(_08067_ ), .Q(\IF_ID_pc [30] ), .QN(_08161_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00283_ ), .CK(_08067_ ), .Q(\IF_ID_pc [21] ), .QN(_08160_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00284_ ), .CK(_08067_ ), .Q(\IF_ID_pc [20] ), .QN(_08159_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00285_ ), .CK(_08067_ ), .Q(\IF_ID_pc [19] ), .QN(_08158_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00286_ ), .CK(_08067_ ), .Q(\IF_ID_pc [18] ), .QN(_08157_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00287_ ), .CK(_08067_ ), .Q(\IF_ID_pc [17] ), .QN(_08156_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00288_ ), .CK(_08067_ ), .Q(\IF_ID_pc [16] ), .QN(_08155_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00289_ ), .CK(_08067_ ), .Q(\IF_ID_pc [15] ), .QN(_08154_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00290_ ), .CK(_08067_ ), .Q(\IF_ID_pc [14] ), .QN(_08153_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00291_ ), .CK(_08067_ ), .Q(\IF_ID_pc [13] ), .QN(_08152_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00292_ ), .CK(_08067_ ), .Q(\IF_ID_pc [12] ), .QN(_08151_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00293_ ), .CK(_08067_ ), .Q(\IF_ID_pc [29] ), .QN(_08150_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00294_ ), .CK(_08067_ ), .Q(\IF_ID_pc [11] ), .QN(_08149_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00295_ ), .CK(_08067_ ), .Q(\IF_ID_pc [10] ), .QN(_08148_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00296_ ), .CK(_08067_ ), .Q(\IF_ID_pc [9] ), .QN(_08147_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00297_ ), .CK(_08067_ ), .Q(\IF_ID_pc [8] ), .QN(_08146_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00298_ ), .CK(_08067_ ), .Q(\IF_ID_pc [7] ), .QN(_08145_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00299_ ), .CK(_08067_ ), .Q(\IF_ID_pc [6] ), .QN(_08144_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00300_ ), .CK(_08067_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00301_ ), .CK(_08067_ ), .Q(\IF_ID_pc [4] ), .QN(_08143_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00303_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08142_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00302_ ), .CK(_08067_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00305_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08140_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00304_ ), .CK(_08067_ ), .Q(\IF_ID_pc [2] ), .QN(_08141_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00306_ ), .CK(_08067_ ), .Q(\IF_ID_pc [28] ), .QN(_08139_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00307_ ), .CK(_08067_ ), .Q(\IF_ID_pc [1] ), .QN(_08138_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00308_ ), .CK(_08067_ ), .Q(\IF_ID_pc [27] ), .QN(_08137_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00309_ ), .CK(_08067_ ), .Q(\IF_ID_pc [26] ), .QN(_08136_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00310_ ), .CK(_08067_ ), .Q(\IF_ID_pc [25] ), .QN(_08135_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00311_ ), .CK(_08067_ ), .Q(\IF_ID_pc [24] ), .QN(_08134_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00312_ ), .CK(_08067_ ), .Q(\IF_ID_pc [23] ), .QN(_08133_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00313_ ), .CK(_08067_ ), .Q(\IF_ID_pc [22] ), .QN(_08132_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00314_ ), .CK(_08067_ ), .Q(\IF_ID_pc [31] ), .QN(_08131_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08933_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08130_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00315_ ), .CK(_08066_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08932_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00317_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00316_ ), .CK(_08065_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08129_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08934_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08935_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08936_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08937_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08938_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08939_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08940_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08941_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08942_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08943_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08944_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08945_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08946_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08947_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08948_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08949_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08950_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08951_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08952_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08953_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08954_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08955_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08956_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08957_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08958_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08959_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08960_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08961_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08962_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08963_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08964_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08064_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08965_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08966_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08967_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08968_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08969_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08970_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08971_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08972_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08973_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08974_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08975_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08976_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08977_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08978_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08979_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08980_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08981_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08982_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08983_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08984_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08985_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08986_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08987_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08988_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08989_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08990_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08991_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08992_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08993_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08994_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08995_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08996_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08063_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08128_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PP0P__Q ( .D(_00318_ ), .CK(_08062_ ), .Q(LS_WB_pc ), .QN(_08127_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PP0P__Q ( .D(_00319_ ), .CK(_08061_ ), .Q(\mylsu.previous_load_done ), .QN(_08997_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08998_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08999_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_09000_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(_09001_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_08064_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_08064_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_09002_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_08064_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08126_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00320_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08125_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00321_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08124_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00322_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08123_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00323_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08122_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00324_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08121_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00325_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08120_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00326_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08119_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00327_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08118_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00328_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08117_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00329_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08116_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00330_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08115_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00331_ ), .CK(_08064_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_09003_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_08064_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_09004_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_08064_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_09005_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_08064_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_09006_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_08064_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_09007_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_09008_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_09009_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_09010_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_09011_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_09012_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_09013_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_09014_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_09015_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_09016_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_09017_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_09018_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_09019_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_09020_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_09021_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_09022_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_09023_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_09024_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_09025_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_09026_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_09027_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_09028_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_09029_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_09030_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_09031_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_09032_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_09033_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_09034_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_09035_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_09036_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_09037_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_09038_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_08064_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_09039_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_09040_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_09041_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_09042_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_09043_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_09044_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_09045_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_09046_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_09047_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_09048_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_09049_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_09050_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_09051_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_09052_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_09053_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_09054_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_09055_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_09056_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_09057_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_09058_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_09059_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_09060_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_09061_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_09062_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_09063_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_09064_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_09065_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_09066_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_09067_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_09068_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_09069_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_09070_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_08060_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08114_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q ( .D(_00332_ ), .CK(_08059_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_08113_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_1 ( .D(_00333_ ), .CK(_08059_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08112_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_2 ( .D(_00334_ ), .CK(_08059_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08111_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_3 ( .D(_00335_ ), .CK(_08059_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08110_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_4 ( .D(_00336_ ), .CK(_08059_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08109_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_5 ( .D(_00337_ ), .CK(_08059_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08108_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PP0P__Q ( .D(_00338_ ), .CK(_08059_ ), .Q(LS_WB_wen_reg ), .QN(_09071_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_09072_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_09073_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08058_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08057_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08056_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08055_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08054_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08053_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08052_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08051_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08050_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08049_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08048_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08047_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08046_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08045_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08044_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_1_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_10_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_11_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_12_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_13_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_14_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_15_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_16_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_17_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_18_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_19_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_2_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_20_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_21_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_22_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_23_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_24_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_25_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_26_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_27_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_28_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_29_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_3_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_30_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_31_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_4_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_5_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_6_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_7_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_8_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[5]_$_DFFE_PP__Q_9_D ), .CK(_08043_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00339_ ), .CK(_08042_ ), .Q(loaduse_clear ), .QN(_09074_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_09075_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_09076_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08107_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(reset ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(reset ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\ID_EX_typ [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(excp_written ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_44 ) );
BUF_X8 fanout_buf_45 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_45 ) );
BUF_X8 fanout_buf_46 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_46 ) );
BUF_X8 fanout_buf_47 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_47 ) );
BUF_X8 fanout_buf_48 ( .A(\myifu.to_reset ), .Z(fanout_net_48 ) );

endmodule
