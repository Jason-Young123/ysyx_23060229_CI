//Generate the verilog at 2025-09-29T18:10:51 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire io_master_wready_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ;
wire io_master_wready_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.check_quest_$_NAND__B_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_AND__A_Y ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ;
wire \myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.check_assert_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__A_Y ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][27] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][27] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][27] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][27] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_E ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_E_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [1] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

INV_X2 _08203_ ( .A(fanout_net_1 ), .ZN(_00731_ ) );
BUF_X4 _08204_ ( .A(_00731_ ), .Z(_00732_ ) );
AND3_X4 _08205_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_00733_ ) );
AND3_X4 _08206_ ( .A1(_00733_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_00734_ ) );
AND3_X4 _08207_ ( .A1(_00734_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_00735_ ) );
AND3_X4 _08208_ ( .A1(_00735_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_00736_ ) );
AND3_X4 _08209_ ( .A1(_00736_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_00737_ ) );
AND3_X4 _08210_ ( .A1(_00737_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_00738_ ) );
AND3_X4 _08211_ ( .A1(_00738_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_00739_ ) );
AND3_X4 _08212_ ( .A1(_00739_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_00740_ ) );
AND3_X4 _08213_ ( .A1(_00740_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_00741_ ) );
AND3_X4 _08214_ ( .A1(_00741_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_00742_ ) );
AND3_X4 _08215_ ( .A1(_00742_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_00743_ ) );
AND3_X4 _08216_ ( .A1(_00743_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_00744_ ) );
AND3_X4 _08217_ ( .A1(_00744_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_00745_ ) );
AND3_X4 _08218_ ( .A1(_00745_ ), .A2(\myclint.mtime [28] ), .A3(\myclint.mtime [27] ), .ZN(_00746_ ) );
AND2_X1 _08219_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_00747_ ) );
AND4_X4 _08220_ ( .A1(\myclint.mtime [33] ), .A2(_00746_ ), .A3(\myclint.mtime [29] ), .A4(_00747_ ), .ZN(_00748_ ) );
AND3_X4 _08221_ ( .A1(_00748_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_00749_ ) );
AND2_X4 _08222_ ( .A1(_00749_ ), .A2(\myclint.mtime [35] ), .ZN(_00750_ ) );
AND2_X1 _08223_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [39] ), .ZN(_00751_ ) );
AND2_X1 _08224_ ( .A1(\myclint.mtime [36] ), .A2(\myclint.mtime [37] ), .ZN(_00752_ ) );
AND3_X4 _08225_ ( .A1(_00750_ ), .A2(_00751_ ), .A3(_00752_ ), .ZN(_00753_ ) );
NAND2_X4 _08226_ ( .A1(_00753_ ), .A2(\myclint.mtime [40] ), .ZN(_00754_ ) );
INV_X1 _08227_ ( .A(\myclint.mtime [42] ), .ZN(_00755_ ) );
INV_X1 _08228_ ( .A(\myclint.mtime [41] ), .ZN(_00756_ ) );
NOR3_X4 _08229_ ( .A1(_00754_ ), .A2(_00755_ ), .A3(_00756_ ), .ZN(_00757_ ) );
AND2_X4 _08230_ ( .A1(_00757_ ), .A2(\myclint.mtime [43] ), .ZN(_00758_ ) );
AND2_X1 _08231_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_00759_ ) );
AND3_X1 _08232_ ( .A1(_00759_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_00760_ ) );
NAND2_X4 _08233_ ( .A1(_00758_ ), .A2(_00760_ ), .ZN(_00761_ ) );
AND2_X1 _08234_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_00762_ ) );
INV_X1 _08235_ ( .A(_00762_ ), .ZN(_00763_ ) );
NOR2_X4 _08236_ ( .A1(_00761_ ), .A2(_00763_ ), .ZN(_00764_ ) );
AND2_X1 _08237_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_00765_ ) );
NAND2_X2 _08238_ ( .A1(_00764_ ), .A2(_00765_ ), .ZN(_00766_ ) );
AND2_X1 _08239_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_00767_ ) );
INV_X1 _08240_ ( .A(_00767_ ), .ZN(_00768_ ) );
NOR2_X2 _08241_ ( .A1(_00766_ ), .A2(_00768_ ), .ZN(_00769_ ) );
AND2_X1 _08242_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_00770_ ) );
NAND2_X2 _08243_ ( .A1(_00769_ ), .A2(_00770_ ), .ZN(_00771_ ) );
AND2_X1 _08244_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_00772_ ) );
INV_X1 _08245_ ( .A(_00772_ ), .ZN(_00773_ ) );
NOR2_X2 _08246_ ( .A1(_00771_ ), .A2(_00773_ ), .ZN(_00774_ ) );
AND2_X1 _08247_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_00775_ ) );
AND2_X1 _08248_ ( .A1(_00774_ ), .A2(_00775_ ), .ZN(_00776_ ) );
NAND3_X1 _08249_ ( .A1(_00776_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_00777_ ) );
NOR2_X1 _08250_ ( .A1(_00777_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00778_ ) );
OAI21_X1 _08251_ ( .A(_00732_ ), .B1(_00778_ ), .B2(\myclint.mtime [63] ), .ZN(_00779_ ) );
AND2_X4 _08252_ ( .A1(_00746_ ), .A2(\myclint.mtime [29] ), .ZN(_00780_ ) );
AND2_X1 _08253_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_00781_ ) );
AND3_X4 _08254_ ( .A1(_00780_ ), .A2(_00781_ ), .A3(_00747_ ), .ZN(_00782_ ) );
AND2_X4 _08255_ ( .A1(_00782_ ), .A2(\myclint.mtime [34] ), .ZN(_00783_ ) );
AND2_X4 _08256_ ( .A1(_00783_ ), .A2(\myclint.mtime [35] ), .ZN(_00784_ ) );
AND3_X4 _08257_ ( .A1(_00784_ ), .A2(_00751_ ), .A3(_00752_ ), .ZN(_00785_ ) );
NAND2_X4 _08258_ ( .A1(_00785_ ), .A2(\myclint.mtime [40] ), .ZN(_00786_ ) );
NOR3_X4 _08259_ ( .A1(_00786_ ), .A2(_00755_ ), .A3(_00756_ ), .ZN(_00787_ ) );
AND2_X4 _08260_ ( .A1(_00787_ ), .A2(\myclint.mtime [43] ), .ZN(_00788_ ) );
AND2_X4 _08261_ ( .A1(_00788_ ), .A2(_00760_ ), .ZN(_00789_ ) );
AND2_X4 _08262_ ( .A1(_00789_ ), .A2(_00762_ ), .ZN(_00790_ ) );
AND2_X4 _08263_ ( .A1(_00790_ ), .A2(_00765_ ), .ZN(_00791_ ) );
AND2_X4 _08264_ ( .A1(_00791_ ), .A2(_00767_ ), .ZN(_00792_ ) );
AND2_X4 _08265_ ( .A1(_00792_ ), .A2(_00770_ ), .ZN(_00793_ ) );
AND2_X4 _08266_ ( .A1(_00793_ ), .A2(_00772_ ), .ZN(_00794_ ) );
AND2_X2 _08267_ ( .A1(_00794_ ), .A2(_00775_ ), .ZN(_00795_ ) );
NAND3_X1 _08268_ ( .A1(_00795_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_00796_ ) );
NOR2_X1 _08269_ ( .A1(_00796_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00797_ ) );
AOI21_X1 _08270_ ( .A(_00779_ ), .B1(_00797_ ), .B2(\myclint.mtime [63] ), .ZN(_00000_ ) );
AND2_X2 _08271_ ( .A1(_00735_ ), .A2(\myclint.mtime [7] ), .ZN(_00798_ ) );
AND4_X1 _08272_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_00799_ ) );
AND2_X1 _08273_ ( .A1(\myclint.mtime [10] ), .A2(\myclint.mtime [11] ), .ZN(_00800_ ) );
AND4_X1 _08274_ ( .A1(\myclint.mtime [8] ), .A2(_00799_ ), .A3(\myclint.mtime [9] ), .A4(_00800_ ), .ZN(_00801_ ) );
AND2_X1 _08275_ ( .A1(_00798_ ), .A2(_00801_ ), .ZN(_00802_ ) );
AND4_X1 _08276_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [28] ), .A3(\myclint.mtime [29] ), .A4(\myclint.mtime [31] ), .ZN(_00803_ ) );
AND2_X1 _08277_ ( .A1(\myclint.mtime [26] ), .A2(\myclint.mtime [27] ), .ZN(_00804_ ) );
NAND4_X1 _08278_ ( .A1(_00803_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .A4(_00804_ ), .ZN(_00805_ ) );
NAND4_X1 _08279_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_00806_ ) );
AND2_X1 _08280_ ( .A1(\myclint.mtime [18] ), .A2(\myclint.mtime [19] ), .ZN(_00807_ ) );
NAND3_X1 _08281_ ( .A1(_00807_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_00808_ ) );
NOR3_X1 _08282_ ( .A1(_00805_ ), .A2(_00806_ ), .A3(_00808_ ), .ZN(_00809_ ) );
AND2_X1 _08283_ ( .A1(_00802_ ), .A2(_00809_ ), .ZN(_00810_ ) );
AND3_X1 _08284_ ( .A1(_00781_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_00811_ ) );
AND3_X1 _08285_ ( .A1(_00811_ ), .A2(_00751_ ), .A3(_00752_ ), .ZN(_00812_ ) );
AND2_X1 _08286_ ( .A1(\myclint.mtime [40] ), .A2(\myclint.mtime [41] ), .ZN(_00813_ ) );
AND3_X1 _08287_ ( .A1(_00813_ ), .A2(\myclint.mtime [42] ), .A3(\myclint.mtime [43] ), .ZN(_00814_ ) );
AND3_X1 _08288_ ( .A1(_00812_ ), .A2(_00760_ ), .A3(_00814_ ), .ZN(_00815_ ) );
AND2_X1 _08289_ ( .A1(_00810_ ), .A2(_00815_ ), .ZN(_00816_ ) );
AND4_X1 _08290_ ( .A1(_00770_ ), .A2(_00767_ ), .A3(_00765_ ), .A4(_00762_ ), .ZN(_00817_ ) );
AND2_X1 _08291_ ( .A1(_00816_ ), .A2(_00817_ ), .ZN(_00818_ ) );
AND4_X1 _08292_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_00819_ ) );
AND2_X1 _08293_ ( .A1(_00818_ ), .A2(_00819_ ), .ZN(_00820_ ) );
AND3_X1 _08294_ ( .A1(_00820_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_00821_ ) );
XNOR2_X1 _08295_ ( .A(_00821_ ), .B(\myclint.mtime [62] ), .ZN(_00822_ ) );
NOR2_X1 _08296_ ( .A1(_00822_ ), .A2(fanout_net_1 ), .ZN(_00001_ ) );
INV_X1 _08297_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00823_ ) );
AND3_X1 _08298_ ( .A1(_00764_ ), .A2(_00823_ ), .A3(_00765_ ), .ZN(_00824_ ) );
OAI21_X1 _08299_ ( .A(_00732_ ), .B1(_00824_ ), .B2(\myclint.mtime [53] ), .ZN(_00825_ ) );
AND3_X1 _08300_ ( .A1(_00790_ ), .A2(_00823_ ), .A3(_00765_ ), .ZN(_00826_ ) );
AOI21_X1 _08301_ ( .A(_00825_ ), .B1(_00826_ ), .B2(\myclint.mtime [53] ), .ZN(_00002_ ) );
AND2_X1 _08302_ ( .A1(_00765_ ), .A2(_00762_ ), .ZN(_00827_ ) );
AND2_X1 _08303_ ( .A1(_00816_ ), .A2(_00827_ ), .ZN(_00828_ ) );
XNOR2_X1 _08304_ ( .A(_00828_ ), .B(\myclint.mtime [52] ), .ZN(_00829_ ) );
NOR2_X1 _08305_ ( .A1(_00829_ ), .A2(fanout_net_1 ), .ZN(_00003_ ) );
BUF_X4 _08306_ ( .A(_00731_ ), .Z(_00830_ ) );
NOR3_X1 _08307_ ( .A1(_00761_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00763_ ), .ZN(_00831_ ) );
OAI21_X1 _08308_ ( .A(_00830_ ), .B1(_00831_ ), .B2(\myclint.mtime [51] ), .ZN(_00832_ ) );
INV_X1 _08309_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00833_ ) );
AND3_X1 _08310_ ( .A1(_00789_ ), .A2(_00833_ ), .A3(_00762_ ), .ZN(_00834_ ) );
AOI21_X1 _08311_ ( .A(_00832_ ), .B1(_00834_ ), .B2(\myclint.mtime [51] ), .ZN(_00004_ ) );
INV_X1 _08312_ ( .A(_00810_ ), .ZN(_00835_ ) );
INV_X1 _08313_ ( .A(_00815_ ), .ZN(_00836_ ) );
OR4_X1 _08314_ ( .A1(\myclint.mtime [50] ), .A2(_00835_ ), .A3(_00763_ ), .A4(_00836_ ), .ZN(_00837_ ) );
AND3_X1 _08315_ ( .A1(_00810_ ), .A2(_00762_ ), .A3(_00815_ ), .ZN(_00838_ ) );
INV_X1 _08316_ ( .A(_00838_ ), .ZN(_00839_ ) );
NAND2_X1 _08317_ ( .A1(_00839_ ), .A2(\myclint.mtime [50] ), .ZN(_00840_ ) );
AOI21_X1 _08318_ ( .A(fanout_net_1 ), .B1(_00837_ ), .B2(_00840_ ), .ZN(_00005_ ) );
BUF_X2 _08319_ ( .A(_00731_ ), .Z(_00841_ ) );
INV_X1 _08320_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00842_ ) );
AND3_X1 _08321_ ( .A1(_00758_ ), .A2(_00842_ ), .A3(_00760_ ), .ZN(_00843_ ) );
OAI21_X1 _08322_ ( .A(_00841_ ), .B1(_00843_ ), .B2(\myclint.mtime [49] ), .ZN(_00844_ ) );
AND4_X1 _08323_ ( .A1(\myclint.mtime [49] ), .A2(_00788_ ), .A3(_00842_ ), .A4(_00760_ ), .ZN(_00845_ ) );
NOR2_X1 _08324_ ( .A1(_00844_ ), .A2(_00845_ ), .ZN(_00006_ ) );
OR3_X1 _08325_ ( .A1(_00835_ ), .A2(\myclint.mtime [48] ), .A3(_00836_ ), .ZN(_00846_ ) );
OAI21_X1 _08326_ ( .A(\myclint.mtime [48] ), .B1(_00835_ ), .B2(_00836_ ), .ZN(_00847_ ) );
AOI21_X1 _08327_ ( .A(fanout_net_1 ), .B1(_00846_ ), .B2(_00847_ ), .ZN(_00007_ ) );
NAND3_X1 _08328_ ( .A1(_00757_ ), .A2(\myclint.mtime [43] ), .A3(_00759_ ), .ZN(_00848_ ) );
NOR2_X1 _08329_ ( .A1(_00848_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00849_ ) );
OAI21_X1 _08330_ ( .A(_00830_ ), .B1(_00849_ ), .B2(\myclint.mtime [47] ), .ZN(_00850_ ) );
NAND3_X1 _08331_ ( .A1(_00787_ ), .A2(\myclint.mtime [44] ), .A3(\myclint.mtime [43] ), .ZN(_00851_ ) );
INV_X1 _08332_ ( .A(\myclint.mtime [45] ), .ZN(_00852_ ) );
NOR3_X1 _08333_ ( .A1(_00851_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00852_ ), .ZN(_00853_ ) );
AOI21_X1 _08334_ ( .A(_00850_ ), .B1(\myclint.mtime [47] ), .B2(_00853_ ), .ZN(_00008_ ) );
AND2_X1 _08335_ ( .A1(_00810_ ), .A2(_00812_ ), .ZN(_00854_ ) );
AND3_X1 _08336_ ( .A1(_00854_ ), .A2(_00759_ ), .A3(_00814_ ), .ZN(_00855_ ) );
XNOR2_X1 _08337_ ( .A(_00855_ ), .B(\myclint.mtime [46] ), .ZN(_00856_ ) );
NOR2_X1 _08338_ ( .A1(_00856_ ), .A2(fanout_net_1 ), .ZN(_00009_ ) );
INV_X1 _08339_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00857_ ) );
NAND3_X1 _08340_ ( .A1(_00757_ ), .A2(_00857_ ), .A3(\myclint.mtime [43] ), .ZN(_00858_ ) );
AOI21_X1 _08341_ ( .A(fanout_net_1 ), .B1(_00858_ ), .B2(_00852_ ), .ZN(_00859_ ) );
NAND4_X1 _08342_ ( .A1(_00787_ ), .A2(\myclint.mtime [45] ), .A3(_00857_ ), .A4(\myclint.mtime [43] ), .ZN(_00860_ ) );
AND2_X1 _08343_ ( .A1(_00859_ ), .A2(_00860_ ), .ZN(_00010_ ) );
AND2_X1 _08344_ ( .A1(_00854_ ), .A2(_00814_ ), .ZN(_00861_ ) );
XNOR2_X1 _08345_ ( .A(_00861_ ), .B(\myclint.mtime [44] ), .ZN(_00862_ ) );
NOR2_X1 _08346_ ( .A1(_00862_ ), .A2(fanout_net_1 ), .ZN(_00011_ ) );
INV_X1 _08347_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00863_ ) );
AND3_X1 _08348_ ( .A1(_00774_ ), .A2(_00863_ ), .A3(_00775_ ), .ZN(_00864_ ) );
OAI21_X1 _08349_ ( .A(_00830_ ), .B1(_00864_ ), .B2(\myclint.mtime [61] ), .ZN(_00865_ ) );
AND3_X1 _08350_ ( .A1(_00794_ ), .A2(_00863_ ), .A3(_00775_ ), .ZN(_00866_ ) );
AOI21_X1 _08351_ ( .A(_00865_ ), .B1(_00866_ ), .B2(\myclint.mtime [61] ), .ZN(_00012_ ) );
NOR3_X1 _08352_ ( .A1(_00754_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00756_ ), .ZN(_00867_ ) );
OAI21_X1 _08353_ ( .A(_00830_ ), .B1(_00867_ ), .B2(\myclint.mtime [43] ), .ZN(_00868_ ) );
NOR3_X1 _08354_ ( .A1(_00786_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00756_ ), .ZN(_00869_ ) );
AOI21_X1 _08355_ ( .A(_00868_ ), .B1(\myclint.mtime [43] ), .B2(_00869_ ), .ZN(_00013_ ) );
AND3_X1 _08356_ ( .A1(_00753_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_00870_ ) );
OAI21_X1 _08357_ ( .A(_00841_ ), .B1(_00870_ ), .B2(\myclint.mtime [42] ), .ZN(_00871_ ) );
NOR2_X1 _08358_ ( .A1(_00871_ ), .A2(_00757_ ), .ZN(_00014_ ) );
INV_X1 _08359_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00872_ ) );
NAND2_X1 _08360_ ( .A1(_00753_ ), .A2(_00872_ ), .ZN(_00873_ ) );
AOI21_X1 _08361_ ( .A(fanout_net_1 ), .B1(_00873_ ), .B2(_00756_ ), .ZN(_00874_ ) );
AND2_X1 _08362_ ( .A1(_00784_ ), .A2(_00752_ ), .ZN(_00875_ ) );
NAND4_X1 _08363_ ( .A1(_00875_ ), .A2(\myclint.mtime [41] ), .A3(_00872_ ), .A4(_00751_ ), .ZN(_00876_ ) );
AND2_X1 _08364_ ( .A1(_00874_ ), .A2(_00876_ ), .ZN(_00015_ ) );
XNOR2_X1 _08365_ ( .A(_00854_ ), .B(\myclint.mtime [40] ), .ZN(_00877_ ) );
NOR2_X1 _08366_ ( .A1(_00877_ ), .A2(fanout_net_1 ), .ZN(_00016_ ) );
INV_X1 _08367_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00878_ ) );
AND3_X1 _08368_ ( .A1(_00750_ ), .A2(_00878_ ), .A3(_00752_ ), .ZN(_00879_ ) );
OAI21_X1 _08369_ ( .A(_00841_ ), .B1(_00879_ ), .B2(\myclint.mtime [39] ), .ZN(_00880_ ) );
AND4_X1 _08370_ ( .A1(_00878_ ), .A2(_00784_ ), .A3(\myclint.mtime [39] ), .A4(_00752_ ), .ZN(_00881_ ) );
NOR2_X1 _08371_ ( .A1(_00880_ ), .A2(_00881_ ), .ZN(_00017_ ) );
NAND3_X1 _08372_ ( .A1(_00810_ ), .A2(_00752_ ), .A3(_00811_ ), .ZN(_00882_ ) );
OR2_X1 _08373_ ( .A1(_00882_ ), .A2(\myclint.mtime [38] ), .ZN(_00883_ ) );
NAND2_X1 _08374_ ( .A1(_00882_ ), .A2(\myclint.mtime [38] ), .ZN(_00884_ ) );
AOI21_X1 _08375_ ( .A(fanout_net_1 ), .B1(_00883_ ), .B2(_00884_ ), .ZN(_00018_ ) );
BUF_X4 _08376_ ( .A(_00731_ ), .Z(_00885_ ) );
INV_X1 _08377_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00886_ ) );
AND3_X1 _08378_ ( .A1(_00749_ ), .A2(_00886_ ), .A3(\myclint.mtime [35] ), .ZN(_00887_ ) );
OAI21_X1 _08379_ ( .A(_00885_ ), .B1(_00887_ ), .B2(\myclint.mtime [37] ), .ZN(_00888_ ) );
AND4_X1 _08380_ ( .A1(\myclint.mtime [37] ), .A2(_00783_ ), .A3(_00886_ ), .A4(\myclint.mtime [35] ), .ZN(_00889_ ) );
NOR2_X1 _08381_ ( .A1(_00888_ ), .A2(_00889_ ), .ZN(_00019_ ) );
AND2_X1 _08382_ ( .A1(_00810_ ), .A2(_00811_ ), .ZN(_00890_ ) );
XNOR2_X1 _08383_ ( .A(_00890_ ), .B(\myclint.mtime [36] ), .ZN(_00891_ ) );
NOR2_X1 _08384_ ( .A1(_00891_ ), .A2(fanout_net_1 ), .ZN(_00020_ ) );
INV_X1 _08385_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00892_ ) );
AND3_X1 _08386_ ( .A1(_00782_ ), .A2(_00892_ ), .A3(\myclint.mtime [35] ), .ZN(_00893_ ) );
NAND4_X1 _08387_ ( .A1(_00746_ ), .A2(\myclint.mtime [33] ), .A3(\myclint.mtime [29] ), .A4(_00747_ ), .ZN(_00894_ ) );
INV_X1 _08388_ ( .A(\myclint.mtime [32] ), .ZN(_00895_ ) );
NOR3_X1 _08389_ ( .A1(_00894_ ), .A2(_00895_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00896_ ) );
OAI21_X1 _08390_ ( .A(_00732_ ), .B1(_00896_ ), .B2(\myclint.mtime [35] ), .ZN(_00897_ ) );
NOR2_X1 _08391_ ( .A1(_00893_ ), .A2(_00897_ ), .ZN(_00021_ ) );
NOR2_X1 _08392_ ( .A1(_00894_ ), .A2(_00895_ ), .ZN(_00898_ ) );
OAI21_X1 _08393_ ( .A(_00885_ ), .B1(_00898_ ), .B2(\myclint.mtime [34] ), .ZN(_00899_ ) );
NOR2_X1 _08394_ ( .A1(_00899_ ), .A2(_00749_ ), .ZN(_00022_ ) );
XNOR2_X1 _08395_ ( .A(_00820_ ), .B(\myclint.mtime [60] ), .ZN(_00900_ ) );
NOR2_X1 _08396_ ( .A1(_00900_ ), .A2(fanout_net_1 ), .ZN(_00023_ ) );
OR3_X1 _08397_ ( .A1(_00835_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(\myclint.mtime [33] ), .ZN(_00901_ ) );
OAI21_X1 _08398_ ( .A(\myclint.mtime [33] ), .B1(_00835_ ), .B2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_00902_ ) );
AOI21_X1 _08399_ ( .A(fanout_net_1 ), .B1(_00901_ ), .B2(_00902_ ), .ZN(_00024_ ) );
OR2_X1 _08400_ ( .A1(_00810_ ), .A2(_00895_ ), .ZN(_00903_ ) );
NAND4_X1 _08401_ ( .A1(_00798_ ), .A2(_00895_ ), .A3(_00801_ ), .A4(_00809_ ), .ZN(_00904_ ) );
AOI21_X1 _08402_ ( .A(fanout_net_1 ), .B1(_00903_ ), .B2(_00904_ ), .ZN(_00025_ ) );
NAND2_X1 _08403_ ( .A1(_00798_ ), .A2(_00801_ ), .ZN(_00905_ ) );
AND3_X1 _08404_ ( .A1(_00807_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_00906_ ) );
AND4_X1 _08405_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_00907_ ) );
NAND2_X1 _08406_ ( .A1(_00906_ ), .A2(_00907_ ), .ZN(_00908_ ) );
NOR2_X1 _08407_ ( .A1(_00905_ ), .A2(_00908_ ), .ZN(_00909_ ) );
AND3_X1 _08408_ ( .A1(_00804_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_00910_ ) );
AND2_X1 _08409_ ( .A1(_00909_ ), .A2(_00910_ ), .ZN(_00911_ ) );
NAND3_X1 _08410_ ( .A1(_00911_ ), .A2(\myclint.mtime [28] ), .A3(\myclint.mtime [29] ), .ZN(_00912_ ) );
OR3_X1 _08411_ ( .A1(_00912_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [31] ), .ZN(_00913_ ) );
OAI21_X1 _08412_ ( .A(\myclint.mtime [31] ), .B1(_00912_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00914_ ) );
AOI21_X1 _08413_ ( .A(fanout_net_1 ), .B1(_00913_ ), .B2(_00914_ ), .ZN(_00026_ ) );
OR2_X1 _08414_ ( .A1(_00912_ ), .A2(\myclint.mtime [30] ), .ZN(_00915_ ) );
NAND2_X1 _08415_ ( .A1(_00912_ ), .A2(\myclint.mtime [30] ), .ZN(_00916_ ) );
AOI21_X1 _08416_ ( .A(fanout_net_1 ), .B1(_00915_ ), .B2(_00916_ ), .ZN(_00027_ ) );
INV_X1 _08417_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00917_ ) );
AND3_X1 _08418_ ( .A1(_00745_ ), .A2(_00917_ ), .A3(\myclint.mtime [27] ), .ZN(_00918_ ) );
AND2_X1 _08419_ ( .A1(_00918_ ), .A2(\myclint.mtime [29] ), .ZN(_00919_ ) );
OAI21_X1 _08420_ ( .A(_00732_ ), .B1(_00918_ ), .B2(\myclint.mtime [29] ), .ZN(_00920_ ) );
NOR2_X1 _08421_ ( .A1(_00919_ ), .A2(_00920_ ), .ZN(_00028_ ) );
NAND2_X1 _08422_ ( .A1(_00909_ ), .A2(_00910_ ), .ZN(_00921_ ) );
OR2_X1 _08423_ ( .A1(_00921_ ), .A2(\myclint.mtime [28] ), .ZN(_00922_ ) );
NAND2_X1 _08424_ ( .A1(_00921_ ), .A2(\myclint.mtime [28] ), .ZN(_00923_ ) );
AOI21_X1 _08425_ ( .A(fanout_net_1 ), .B1(_00922_ ), .B2(_00923_ ), .ZN(_00029_ ) );
NAND3_X1 _08426_ ( .A1(_00909_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_00924_ ) );
OR3_X1 _08427_ ( .A1(_00924_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_00925_ ) );
OAI21_X1 _08428_ ( .A(\myclint.mtime [27] ), .B1(_00924_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00926_ ) );
AOI21_X1 _08429_ ( .A(fanout_net_1 ), .B1(_00925_ ), .B2(_00926_ ), .ZN(_00030_ ) );
AND2_X1 _08430_ ( .A1(_00744_ ), .A2(\myclint.mtime [25] ), .ZN(_00927_ ) );
OAI21_X1 _08431_ ( .A(_00885_ ), .B1(_00927_ ), .B2(\myclint.mtime [26] ), .ZN(_00928_ ) );
NOR2_X1 _08432_ ( .A1(_00928_ ), .A2(_00745_ ), .ZN(_00031_ ) );
OR3_X1 _08433_ ( .A1(_00905_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_00908_ ), .ZN(_00929_ ) );
NAND2_X1 _08434_ ( .A1(_00929_ ), .A2(\myclint.mtime [25] ), .ZN(_00930_ ) );
OR4_X1 _08435_ ( .A1(\myclint.mtime [25] ), .A2(_00905_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .A4(_00908_ ), .ZN(_00931_ ) );
AOI21_X1 _08436_ ( .A(fanout_net_1 ), .B1(_00930_ ), .B2(_00931_ ), .ZN(_00032_ ) );
AND2_X1 _08437_ ( .A1(_00743_ ), .A2(\myclint.mtime [23] ), .ZN(_00932_ ) );
OAI21_X1 _08438_ ( .A(_00885_ ), .B1(_00932_ ), .B2(\myclint.mtime [24] ), .ZN(_00933_ ) );
NOR2_X1 _08439_ ( .A1(_00933_ ), .A2(_00744_ ), .ZN(_00033_ ) );
NOR3_X1 _08440_ ( .A1(_00771_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00773_ ), .ZN(_00934_ ) );
OAI21_X1 _08441_ ( .A(_00830_ ), .B1(_00934_ ), .B2(\myclint.mtime [59] ), .ZN(_00935_ ) );
INV_X1 _08442_ ( .A(_00793_ ), .ZN(_00936_ ) );
NOR3_X1 _08443_ ( .A1(_00936_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00773_ ), .ZN(_00937_ ) );
AOI21_X1 _08444_ ( .A(_00935_ ), .B1(_00937_ ), .B2(\myclint.mtime [59] ), .ZN(_00034_ ) );
NOR2_X1 _08445_ ( .A1(_00905_ ), .A2(_00808_ ), .ZN(_00938_ ) );
NAND3_X1 _08446_ ( .A1(_00938_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_00939_ ) );
OR3_X1 _08447_ ( .A1(_00939_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_00940_ ) );
OAI21_X1 _08448_ ( .A(\myclint.mtime [23] ), .B1(_00939_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00941_ ) );
AOI21_X1 _08449_ ( .A(fanout_net_1 ), .B1(_00940_ ), .B2(_00941_ ), .ZN(_00035_ ) );
AND2_X1 _08450_ ( .A1(_00742_ ), .A2(\myclint.mtime [21] ), .ZN(_00942_ ) );
OAI21_X1 _08451_ ( .A(_00885_ ), .B1(_00942_ ), .B2(\myclint.mtime [22] ), .ZN(_00943_ ) );
NOR2_X1 _08452_ ( .A1(_00943_ ), .A2(_00743_ ), .ZN(_00036_ ) );
NOR3_X1 _08453_ ( .A1(_00905_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_00808_ ), .ZN(_00944_ ) );
XNOR2_X1 _08454_ ( .A(_00944_ ), .B(\myclint.mtime [21] ), .ZN(_00945_ ) );
NOR2_X1 _08455_ ( .A1(_00945_ ), .A2(fanout_net_1 ), .ZN(_00037_ ) );
AND2_X1 _08456_ ( .A1(_00741_ ), .A2(\myclint.mtime [19] ), .ZN(_00946_ ) );
OAI21_X1 _08457_ ( .A(_00885_ ), .B1(_00946_ ), .B2(\myclint.mtime [20] ), .ZN(_00947_ ) );
NOR2_X1 _08458_ ( .A1(_00947_ ), .A2(_00742_ ), .ZN(_00038_ ) );
NAND3_X1 _08459_ ( .A1(_00802_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [17] ), .ZN(_00948_ ) );
OR3_X1 _08460_ ( .A1(_00948_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_00949_ ) );
OAI21_X1 _08461_ ( .A(\myclint.mtime [19] ), .B1(_00948_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00950_ ) );
AOI21_X1 _08462_ ( .A(fanout_net_1 ), .B1(_00949_ ), .B2(_00950_ ), .ZN(_00039_ ) );
AND2_X1 _08463_ ( .A1(_00740_ ), .A2(\myclint.mtime [17] ), .ZN(_00951_ ) );
OAI21_X1 _08464_ ( .A(_00885_ ), .B1(_00951_ ), .B2(\myclint.mtime [18] ), .ZN(_00952_ ) );
NOR2_X1 _08465_ ( .A1(_00952_ ), .A2(_00741_ ), .ZN(_00040_ ) );
INV_X1 _08466_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00953_ ) );
AND3_X1 _08467_ ( .A1(_00739_ ), .A2(_00953_ ), .A3(\myclint.mtime [15] ), .ZN(_00954_ ) );
AND2_X1 _08468_ ( .A1(_00954_ ), .A2(\myclint.mtime [17] ), .ZN(_00955_ ) );
OAI21_X1 _08469_ ( .A(_00732_ ), .B1(_00954_ ), .B2(\myclint.mtime [17] ), .ZN(_00956_ ) );
NOR2_X1 _08470_ ( .A1(_00955_ ), .A2(_00956_ ), .ZN(_00041_ ) );
AND2_X1 _08471_ ( .A1(_00739_ ), .A2(\myclint.mtime [15] ), .ZN(_00957_ ) );
OAI21_X1 _08472_ ( .A(_00885_ ), .B1(_00957_ ), .B2(\myclint.mtime [16] ), .ZN(_00958_ ) );
NOR2_X1 _08473_ ( .A1(_00958_ ), .A2(_00740_ ), .ZN(_00042_ ) );
AND3_X1 _08474_ ( .A1(_00800_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_00959_ ) );
AND2_X1 _08475_ ( .A1(_00798_ ), .A2(_00959_ ), .ZN(_00960_ ) );
NAND3_X1 _08476_ ( .A1(_00960_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_00961_ ) );
OR3_X1 _08477_ ( .A1(_00961_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_00962_ ) );
OAI21_X1 _08478_ ( .A(\myclint.mtime [15] ), .B1(_00961_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00963_ ) );
AOI21_X1 _08479_ ( .A(fanout_net_1 ), .B1(_00962_ ), .B2(_00963_ ), .ZN(_00043_ ) );
AND2_X1 _08480_ ( .A1(_00738_ ), .A2(\myclint.mtime [13] ), .ZN(_00964_ ) );
OAI21_X1 _08481_ ( .A(_00885_ ), .B1(_00964_ ), .B2(\myclint.mtime [14] ), .ZN(_00965_ ) );
NOR2_X1 _08482_ ( .A1(_00965_ ), .A2(_00739_ ), .ZN(_00044_ ) );
NAND3_X1 _08483_ ( .A1(_00816_ ), .A2(_00772_ ), .A3(_00817_ ), .ZN(_00966_ ) );
OR2_X1 _08484_ ( .A1(_00966_ ), .A2(\myclint.mtime [58] ), .ZN(_00967_ ) );
NAND2_X1 _08485_ ( .A1(_00966_ ), .A2(\myclint.mtime [58] ), .ZN(_00968_ ) );
AOI21_X1 _08486_ ( .A(fanout_net_1 ), .B1(_00967_ ), .B2(_00968_ ), .ZN(_00045_ ) );
INV_X1 _08487_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00969_ ) );
AND3_X1 _08488_ ( .A1(_00737_ ), .A2(_00969_ ), .A3(\myclint.mtime [11] ), .ZN(_00970_ ) );
AND2_X1 _08489_ ( .A1(_00970_ ), .A2(\myclint.mtime [13] ), .ZN(_00971_ ) );
OAI21_X1 _08490_ ( .A(_00732_ ), .B1(_00970_ ), .B2(\myclint.mtime [13] ), .ZN(_00972_ ) );
NOR2_X1 _08491_ ( .A1(_00971_ ), .A2(_00972_ ), .ZN(_00046_ ) );
AND2_X1 _08492_ ( .A1(_00737_ ), .A2(\myclint.mtime [11] ), .ZN(_00973_ ) );
OAI21_X1 _08493_ ( .A(_00885_ ), .B1(_00973_ ), .B2(\myclint.mtime [12] ), .ZN(_00974_ ) );
NOR2_X1 _08494_ ( .A1(_00974_ ), .A2(_00738_ ), .ZN(_00047_ ) );
NAND3_X1 _08495_ ( .A1(_00798_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [9] ), .ZN(_00975_ ) );
OR3_X1 _08496_ ( .A1(_00975_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_00976_ ) );
OAI21_X1 _08497_ ( .A(\myclint.mtime [11] ), .B1(_00975_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00977_ ) );
AOI21_X1 _08498_ ( .A(fanout_net_1 ), .B1(_00976_ ), .B2(_00977_ ), .ZN(_00048_ ) );
AOI21_X1 _08499_ ( .A(\myclint.mtime [10] ), .B1(_00736_ ), .B2(\myclint.mtime [9] ), .ZN(_00978_ ) );
NOR3_X1 _08500_ ( .A1(_00737_ ), .A2(_00978_ ), .A3(fanout_net_1 ), .ZN(_00049_ ) );
INV_X1 _08501_ ( .A(_00798_ ), .ZN(_00979_ ) );
OR3_X1 _08502_ ( .A1(_00979_ ), .A2(\myclint.mtime [9] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00980_ ) );
OAI21_X1 _08503_ ( .A(\myclint.mtime [9] ), .B1(_00979_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00981_ ) );
AOI21_X1 _08504_ ( .A(fanout_net_1 ), .B1(_00980_ ), .B2(_00981_ ), .ZN(_00050_ ) );
OAI21_X1 _08505_ ( .A(_00732_ ), .B1(_00798_ ), .B2(\myclint.mtime [8] ), .ZN(_00982_ ) );
NOR2_X1 _08506_ ( .A1(_00982_ ), .A2(_00736_ ), .ZN(_00051_ ) );
AND2_X1 _08507_ ( .A1(_00734_ ), .A2(\myclint.mtime [5] ), .ZN(_00983_ ) );
INV_X1 _08508_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00984_ ) );
AND3_X1 _08509_ ( .A1(_00983_ ), .A2(_00984_ ), .A3(\myclint.mtime [7] ), .ZN(_00985_ ) );
AOI21_X1 _08510_ ( .A(\myclint.mtime [7] ), .B1(_00983_ ), .B2(_00984_ ), .ZN(_00986_ ) );
NOR3_X1 _08511_ ( .A1(_00985_ ), .A2(_00986_ ), .A3(fanout_net_1 ), .ZN(_00052_ ) );
OAI21_X1 _08512_ ( .A(_00732_ ), .B1(_00983_ ), .B2(\myclint.mtime [6] ), .ZN(_00987_ ) );
NOR2_X1 _08513_ ( .A1(_00987_ ), .A2(_00735_ ), .ZN(_00053_ ) );
AND2_X1 _08514_ ( .A1(_00733_ ), .A2(\myclint.mtime [3] ), .ZN(_00988_ ) );
INV_X1 _08515_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00989_ ) );
AND3_X1 _08516_ ( .A1(_00988_ ), .A2(\myclint.mtime [5] ), .A3(_00989_ ), .ZN(_00990_ ) );
AOI21_X1 _08517_ ( .A(\myclint.mtime [5] ), .B1(_00988_ ), .B2(_00989_ ), .ZN(_00991_ ) );
NOR3_X1 _08518_ ( .A1(_00990_ ), .A2(_00991_ ), .A3(fanout_net_1 ), .ZN(_00054_ ) );
OAI21_X1 _08519_ ( .A(_00732_ ), .B1(_00988_ ), .B2(\myclint.mtime [4] ), .ZN(_00992_ ) );
NOR2_X1 _08520_ ( .A1(_00992_ ), .A2(_00734_ ), .ZN(_00055_ ) );
INV_X1 _08521_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00993_ ) );
AND3_X1 _08522_ ( .A1(_00769_ ), .A2(_00993_ ), .A3(_00770_ ), .ZN(_00994_ ) );
OAI21_X1 _08523_ ( .A(_00830_ ), .B1(_00994_ ), .B2(\myclint.mtime [57] ), .ZN(_00995_ ) );
AND3_X1 _08524_ ( .A1(_00792_ ), .A2(_00993_ ), .A3(_00770_ ), .ZN(_00996_ ) );
AOI21_X1 _08525_ ( .A(_00995_ ), .B1(_00996_ ), .B2(\myclint.mtime [57] ), .ZN(_00056_ ) );
AND2_X1 _08526_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_00997_ ) );
INV_X1 _08527_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_00998_ ) );
AND3_X1 _08528_ ( .A1(_00997_ ), .A2(_00998_ ), .A3(\myclint.mtime [3] ), .ZN(_00999_ ) );
AOI21_X1 _08529_ ( .A(\myclint.mtime [3] ), .B1(_00997_ ), .B2(_00998_ ), .ZN(_01000_ ) );
NOR3_X1 _08530_ ( .A1(_00999_ ), .A2(_01000_ ), .A3(fanout_net_2 ), .ZN(_00057_ ) );
AOI21_X1 _08531_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01001_ ) );
NOR3_X1 _08532_ ( .A1(_00733_ ), .A2(_01001_ ), .A3(fanout_net_2 ), .ZN(_00058_ ) );
NOR2_X1 _08533_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01002_ ) );
NOR3_X1 _08534_ ( .A1(_00997_ ), .A2(_01002_ ), .A3(fanout_net_2 ), .ZN(_00059_ ) );
AND2_X1 _08535_ ( .A1(_00841_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_00060_ ) );
XNOR2_X1 _08536_ ( .A(_00818_ ), .B(\myclint.mtime [56] ), .ZN(_01003_ ) );
NOR2_X1 _08537_ ( .A1(_01003_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
NOR3_X1 _08538_ ( .A1(_00766_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00768_ ), .ZN(_01004_ ) );
OAI21_X1 _08539_ ( .A(_00830_ ), .B1(_01004_ ), .B2(\myclint.mtime [55] ), .ZN(_01005_ ) );
INV_X1 _08540_ ( .A(_00791_ ), .ZN(_01006_ ) );
NOR3_X1 _08541_ ( .A1(_01006_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00768_ ), .ZN(_01007_ ) );
AOI21_X1 _08542_ ( .A(_01005_ ), .B1(_01007_ ), .B2(\myclint.mtime [55] ), .ZN(_00062_ ) );
NAND3_X1 _08543_ ( .A1(_00816_ ), .A2(_00767_ ), .A3(_00827_ ), .ZN(_01008_ ) );
OR2_X1 _08544_ ( .A1(_01008_ ), .A2(\myclint.mtime [54] ), .ZN(_01009_ ) );
NAND2_X1 _08545_ ( .A1(_01008_ ), .A2(\myclint.mtime [54] ), .ZN(_01010_ ) );
AOI21_X1 _08546_ ( .A(fanout_net_2 ), .B1(_01009_ ), .B2(_01010_ ), .ZN(_00063_ ) );
MUX2_X1 _08547_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(fanout_net_35 ), .Z(_01011_ ) );
AND2_X1 _08548_ ( .A1(_01011_ ), .A2(fanout_net_39 ), .ZN(_01012_ ) );
INV_X8 _08549_ ( .A(fanout_net_39 ), .ZN(_01013_ ) );
BUF_X4 _08550_ ( .A(_01013_ ), .Z(_01014_ ) );
MUX2_X1 _08551_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(fanout_net_35 ), .Z(_01015_ ) );
AOI21_X1 _08552_ ( .A(_01012_ ), .B1(_01014_ ), .B2(_01015_ ), .ZN(_01016_ ) );
MUX2_X1 _08553_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_35 ), .Z(_01017_ ) );
OR2_X1 _08554_ ( .A1(_01017_ ), .A2(_01013_ ), .ZN(_01018_ ) );
MUX2_X1 _08555_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_35 ), .Z(_01019_ ) );
OAI21_X1 _08556_ ( .A(_01018_ ), .B1(fanout_net_39 ), .B2(_01019_ ), .ZN(_01020_ ) );
OAI22_X1 _08557_ ( .A1(_01016_ ), .A2(\IF_ID_pc [13] ), .B1(_01020_ ), .B2(\IF_ID_pc [15] ), .ZN(_01021_ ) );
INV_X1 _08558_ ( .A(\IF_ID_pc [5] ), .ZN(_01022_ ) );
OR2_X1 _08559_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_01023_ ) );
INV_X32 _08560_ ( .A(fanout_net_35 ), .ZN(_01024_ ) );
OAI211_X1 _08561_ ( .A(_01023_ ), .B(_01013_ ), .C1(_01024_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_01025_ ) );
OR2_X2 _08562_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[2][1] ), .ZN(_01026_ ) );
OAI211_X1 _08563_ ( .A(_01026_ ), .B(fanout_net_39 ), .C1(_01024_ ), .C2(\myifu.myicache.tag[3][1] ), .ZN(_01027_ ) );
NAND2_X1 _08564_ ( .A1(_01025_ ), .A2(_01027_ ), .ZN(_01028_ ) );
OR2_X1 _08565_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[0][12] ), .ZN(_01029_ ) );
OAI211_X1 _08566_ ( .A(_01029_ ), .B(_01013_ ), .C1(_01024_ ), .C2(\myifu.myicache.tag[1][12] ), .ZN(_01030_ ) );
OR2_X2 _08567_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[2][12] ), .ZN(_01031_ ) );
OAI211_X1 _08568_ ( .A(_01031_ ), .B(fanout_net_39 ), .C1(_01024_ ), .C2(\myifu.myicache.tag[3][12] ), .ZN(_01032_ ) );
NAND2_X1 _08569_ ( .A1(_01030_ ), .A2(_01032_ ), .ZN(_01033_ ) );
INV_X1 _08570_ ( .A(\IF_ID_pc [16] ), .ZN(_01034_ ) );
AOI22_X1 _08571_ ( .A1(_01022_ ), .A2(_01028_ ), .B1(_01033_ ), .B2(_01034_ ), .ZN(_01035_ ) );
MUX2_X1 _08572_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(fanout_net_35 ), .Z(_01036_ ) );
MUX2_X1 _08573_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_35 ), .Z(_01037_ ) );
MUX2_X1 _08574_ ( .A(_01036_ ), .B(_01037_ ), .S(fanout_net_39 ), .Z(_01038_ ) );
INV_X1 _08575_ ( .A(_01038_ ), .ZN(_01039_ ) );
OAI221_X1 _08576_ ( .A(_01035_ ), .B1(_01022_ ), .B2(_01028_ ), .C1(_01039_ ), .C2(\IF_ID_pc [24] ), .ZN(_01040_ ) );
OR2_X1 _08577_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[0][21] ), .ZN(_01041_ ) );
BUF_X4 _08578_ ( .A(_01013_ ), .Z(_01042_ ) );
BUF_X2 _08579_ ( .A(_01024_ ), .Z(_01043_ ) );
OAI211_X1 _08580_ ( .A(_01041_ ), .B(_01042_ ), .C1(_01043_ ), .C2(\myifu.myicache.tag[1][21] ), .ZN(_01044_ ) );
OR2_X1 _08581_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[2][21] ), .ZN(_01045_ ) );
OAI211_X1 _08582_ ( .A(_01045_ ), .B(fanout_net_39 ), .C1(_01043_ ), .C2(\myifu.myicache.tag[3][21] ), .ZN(_01046_ ) );
AND3_X1 _08583_ ( .A1(_01044_ ), .A2(_01046_ ), .A3(\IF_ID_pc [25] ), .ZN(_01047_ ) );
AOI21_X1 _08584_ ( .A(\IF_ID_pc [25] ), .B1(_01044_ ), .B2(_01046_ ), .ZN(_01048_ ) );
INV_X1 _08585_ ( .A(\IF_ID_pc [30] ), .ZN(_01049_ ) );
MUX2_X1 _08586_ ( .A(\myifu.myicache.tag[0][26] ), .B(\myifu.myicache.tag[1][26] ), .S(fanout_net_35 ), .Z(_01050_ ) );
MUX2_X1 _08587_ ( .A(\myifu.myicache.tag[2][26] ), .B(\myifu.myicache.tag[3][26] ), .S(fanout_net_35 ), .Z(_01051_ ) );
MUX2_X1 _08588_ ( .A(_01050_ ), .B(_01051_ ), .S(fanout_net_39 ), .Z(_01052_ ) );
MUX2_X1 _08589_ ( .A(\myifu.myicache.tag[0][3] ), .B(\myifu.myicache.tag[1][3] ), .S(fanout_net_35 ), .Z(_01053_ ) );
MUX2_X1 _08590_ ( .A(\myifu.myicache.tag[2][3] ), .B(\myifu.myicache.tag[3][3] ), .S(fanout_net_35 ), .Z(_01054_ ) );
MUX2_X1 _08591_ ( .A(_01053_ ), .B(_01054_ ), .S(fanout_net_39 ), .Z(_01055_ ) );
INV_X1 _08592_ ( .A(\IF_ID_pc [7] ), .ZN(_01056_ ) );
OAI22_X1 _08593_ ( .A1(_01049_ ), .A2(_01052_ ), .B1(_01055_ ), .B2(_01056_ ), .ZN(_01057_ ) );
OR4_X2 _08594_ ( .A1(_01040_ ), .A2(_01047_ ), .A3(_01048_ ), .A4(_01057_ ), .ZN(_01058_ ) );
OR2_X1 _08595_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[0][0] ), .ZN(_01059_ ) );
BUF_X4 _08596_ ( .A(_01043_ ), .Z(_01060_ ) );
OAI211_X1 _08597_ ( .A(_01059_ ), .B(_01014_ ), .C1(_01060_ ), .C2(\myifu.myicache.tag[1][0] ), .ZN(_01061_ ) );
OR2_X1 _08598_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[2][0] ), .ZN(_01062_ ) );
OAI211_X1 _08599_ ( .A(_01062_ ), .B(fanout_net_39 ), .C1(_01060_ ), .C2(\myifu.myicache.tag[3][0] ), .ZN(_01063_ ) );
NAND2_X1 _08600_ ( .A1(_01061_ ), .A2(_01063_ ), .ZN(_01064_ ) );
INV_X1 _08601_ ( .A(_01064_ ), .ZN(_01065_ ) );
AOI211_X2 _08602_ ( .A(_01021_ ), .B(_01058_ ), .C1(\IF_ID_pc [4] ), .C2(_01065_ ), .ZN(_01066_ ) );
OR2_X1 _08603_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[0][25] ), .ZN(_01067_ ) );
BUF_X2 _08604_ ( .A(_01024_ ), .Z(_01068_ ) );
OAI211_X1 _08605_ ( .A(_01067_ ), .B(_01042_ ), .C1(_01068_ ), .C2(\myifu.myicache.tag[1][25] ), .ZN(_01069_ ) );
OR2_X1 _08606_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[2][25] ), .ZN(_01070_ ) );
OAI211_X1 _08607_ ( .A(_01070_ ), .B(fanout_net_39 ), .C1(_01068_ ), .C2(\myifu.myicache.tag[3][25] ), .ZN(_01071_ ) );
AOI21_X1 _08608_ ( .A(\IF_ID_pc [29] ), .B1(_01069_ ), .B2(_01071_ ), .ZN(_01072_ ) );
AND2_X1 _08609_ ( .A1(_01020_ ), .A2(\IF_ID_pc [15] ), .ZN(_01073_ ) );
OR2_X1 _08610_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[0][16] ), .ZN(_01074_ ) );
OAI211_X2 _08611_ ( .A(_01074_ ), .B(_01042_ ), .C1(_01068_ ), .C2(\myifu.myicache.tag[1][16] ), .ZN(_01075_ ) );
OR2_X1 _08612_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[2][16] ), .ZN(_01076_ ) );
OAI211_X1 _08613_ ( .A(_01076_ ), .B(fanout_net_39 ), .C1(_01068_ ), .C2(\myifu.myicache.tag[3][16] ), .ZN(_01077_ ) );
AND3_X1 _08614_ ( .A1(_01075_ ), .A2(_01077_ ), .A3(\IF_ID_pc [20] ), .ZN(_01078_ ) );
OR2_X1 _08615_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[0][18] ), .ZN(_01079_ ) );
OAI211_X1 _08616_ ( .A(_01079_ ), .B(_01042_ ), .C1(_01068_ ), .C2(\myifu.myicache.tag[1][18] ), .ZN(_01080_ ) );
OR2_X1 _08617_ ( .A1(fanout_net_35 ), .A2(\myifu.myicache.tag[2][18] ), .ZN(_01081_ ) );
OAI211_X1 _08618_ ( .A(_01081_ ), .B(fanout_net_39 ), .C1(_01068_ ), .C2(\myifu.myicache.tag[3][18] ), .ZN(_01082_ ) );
AOI21_X1 _08619_ ( .A(\IF_ID_pc [22] ), .B1(_01080_ ), .B2(_01082_ ), .ZN(_01083_ ) );
OR4_X1 _08620_ ( .A1(_01072_ ), .A2(_01073_ ), .A3(_01078_ ), .A4(_01083_ ), .ZN(_01084_ ) );
MUX2_X1 _08621_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(fanout_net_35 ), .Z(_01085_ ) );
AND2_X1 _08622_ ( .A1(_01085_ ), .A2(fanout_net_39 ), .ZN(_01086_ ) );
MUX2_X1 _08623_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(fanout_net_35 ), .Z(_01087_ ) );
AOI21_X1 _08624_ ( .A(_01086_ ), .B1(_01014_ ), .B2(_01087_ ), .ZN(_01088_ ) );
MUX2_X1 _08625_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(fanout_net_35 ), .Z(_01089_ ) );
AND2_X1 _08626_ ( .A1(_01089_ ), .A2(fanout_net_39 ), .ZN(_01090_ ) );
MUX2_X1 _08627_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(fanout_net_35 ), .Z(_01091_ ) );
AOI21_X1 _08628_ ( .A(_01090_ ), .B1(_01014_ ), .B2(_01091_ ), .ZN(_01092_ ) );
OAI22_X1 _08629_ ( .A1(\IF_ID_pc [11] ), .A2(_01088_ ), .B1(_01092_ ), .B2(\IF_ID_pc [9] ), .ZN(_01093_ ) );
MUX2_X1 _08630_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(fanout_net_35 ), .Z(_01094_ ) );
AND2_X1 _08631_ ( .A1(_01094_ ), .A2(fanout_net_39 ), .ZN(_01095_ ) );
MUX2_X1 _08632_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(fanout_net_36 ), .Z(_01096_ ) );
AOI21_X1 _08633_ ( .A(_01095_ ), .B1(_01014_ ), .B2(_01096_ ), .ZN(_01097_ ) );
AND2_X1 _08634_ ( .A1(_01097_ ), .A2(\IF_ID_pc [26] ), .ZN(_01098_ ) );
MUX2_X1 _08635_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(fanout_net_36 ), .Z(_01099_ ) );
MUX2_X1 _08636_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(fanout_net_36 ), .Z(_01100_ ) );
MUX2_X1 _08637_ ( .A(_01099_ ), .B(_01100_ ), .S(fanout_net_39 ), .Z(_01101_ ) );
INV_X1 _08638_ ( .A(\IF_ID_pc [19] ), .ZN(_01102_ ) );
NOR2_X1 _08639_ ( .A1(_01101_ ), .A2(_01102_ ), .ZN(_01103_ ) );
NOR4_X1 _08640_ ( .A1(_01084_ ), .A2(_01093_ ), .A3(_01098_ ), .A4(_01103_ ), .ZN(_01104_ ) );
OR2_X1 _08641_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[0][14] ), .ZN(_01105_ ) );
OAI211_X1 _08642_ ( .A(_01105_ ), .B(_01042_ ), .C1(_01068_ ), .C2(\myifu.myicache.tag[1][14] ), .ZN(_01106_ ) );
OR2_X1 _08643_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[2][14] ), .ZN(_01107_ ) );
OAI211_X1 _08644_ ( .A(_01107_ ), .B(fanout_net_39 ), .C1(_01043_ ), .C2(\myifu.myicache.tag[3][14] ), .ZN(_01108_ ) );
NAND2_X1 _08645_ ( .A1(_01106_ ), .A2(_01108_ ), .ZN(_01109_ ) );
INV_X1 _08646_ ( .A(\IF_ID_pc [18] ), .ZN(_01110_ ) );
XNOR2_X1 _08647_ ( .A(_01109_ ), .B(_01110_ ), .ZN(_01111_ ) );
AOI221_X4 _08648_ ( .A(_01111_ ), .B1(_01049_ ), .B2(_01052_ ), .C1(\IF_ID_pc [24] ), .C2(_01039_ ), .ZN(_01112_ ) );
AND2_X1 _08649_ ( .A1(_01055_ ), .A2(_01056_ ), .ZN(_01113_ ) );
OR2_X1 _08650_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[0][27] ), .ZN(_01114_ ) );
OAI211_X1 _08651_ ( .A(_01114_ ), .B(_01014_ ), .C1(_01060_ ), .C2(\myifu.myicache.tag[1][27] ), .ZN(_01115_ ) );
OR2_X1 _08652_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[2][27] ), .ZN(_01116_ ) );
OAI211_X1 _08653_ ( .A(_01116_ ), .B(fanout_net_39 ), .C1(_01060_ ), .C2(\myifu.myicache.tag[3][27] ), .ZN(_01117_ ) );
AOI21_X1 _08654_ ( .A(\IF_ID_pc [31] ), .B1(_01115_ ), .B2(_01117_ ), .ZN(_01118_ ) );
AND3_X1 _08655_ ( .A1(_01115_ ), .A2(_01117_ ), .A3(\IF_ID_pc [31] ), .ZN(_01119_ ) );
AOI21_X1 _08656_ ( .A(\IF_ID_pc [20] ), .B1(_01075_ ), .B2(_01077_ ), .ZN(_01120_ ) );
NOR4_X1 _08657_ ( .A1(_01113_ ), .A2(_01118_ ), .A3(_01119_ ), .A4(_01120_ ), .ZN(_01121_ ) );
AND4_X2 _08658_ ( .A1(_01066_ ), .A2(_01104_ ), .A3(_01112_ ), .A4(_01121_ ), .ZN(_01122_ ) );
INV_X1 _08659_ ( .A(\IF_ID_pc [17] ), .ZN(_01123_ ) );
MUX2_X1 _08660_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(fanout_net_36 ), .Z(_01124_ ) );
MUX2_X1 _08661_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(fanout_net_36 ), .Z(_01125_ ) );
MUX2_X1 _08662_ ( .A(_01124_ ), .B(_01125_ ), .S(fanout_net_39 ), .Z(_01126_ ) );
AOI22_X1 _08663_ ( .A1(_01016_ ), .A2(\IF_ID_pc [13] ), .B1(_01123_ ), .B2(_01126_ ), .ZN(_01127_ ) );
OAI221_X1 _08664_ ( .A(_01127_ ), .B1(\IF_ID_pc [4] ), .B2(_01065_ ), .C1(_01034_ ), .C2(_01033_ ), .ZN(_01128_ ) );
MUX2_X1 _08665_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(fanout_net_36 ), .Z(_01129_ ) );
MUX2_X1 _08666_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(fanout_net_36 ), .Z(_01130_ ) );
MUX2_X1 _08667_ ( .A(_01129_ ), .B(_01130_ ), .S(fanout_net_39 ), .Z(_01131_ ) );
NAND3_X1 _08668_ ( .A1(_01080_ ), .A2(_01082_ ), .A3(\IF_ID_pc [22] ), .ZN(_01132_ ) );
AND2_X1 _08669_ ( .A1(_01131_ ), .A2(_01132_ ), .ZN(_01133_ ) );
OAI221_X1 _08670_ ( .A(_01133_ ), .B1(_01123_ ), .B2(_01126_ ), .C1(_01097_ ), .C2(\IF_ID_pc [26] ), .ZN(_01134_ ) );
NOR2_X1 _08671_ ( .A1(_01128_ ), .A2(_01134_ ), .ZN(_01135_ ) );
AND2_X1 _08672_ ( .A1(_01088_ ), .A2(\IF_ID_pc [11] ), .ZN(_01136_ ) );
OR2_X1 _08673_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[0][8] ), .ZN(_01137_ ) );
OAI211_X1 _08674_ ( .A(_01137_ ), .B(_01042_ ), .C1(_01068_ ), .C2(\myifu.myicache.tag[1][8] ), .ZN(_01138_ ) );
OR2_X1 _08675_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[2][8] ), .ZN(_01139_ ) );
OAI211_X1 _08676_ ( .A(_01139_ ), .B(fanout_net_39 ), .C1(_01068_ ), .C2(\myifu.myicache.tag[3][8] ), .ZN(_01140_ ) );
AND3_X1 _08677_ ( .A1(_01138_ ), .A2(_01140_ ), .A3(\IF_ID_pc [12] ), .ZN(_01141_ ) );
AND3_X1 _08678_ ( .A1(_01069_ ), .A2(_01071_ ), .A3(\IF_ID_pc [29] ), .ZN(_01142_ ) );
AOI21_X1 _08679_ ( .A(\IF_ID_pc [12] ), .B1(_01138_ ), .B2(_01140_ ), .ZN(_01143_ ) );
NOR4_X1 _08680_ ( .A1(_01136_ ), .A2(_01141_ ), .A3(_01142_ ), .A4(_01143_ ), .ZN(_01144_ ) );
MUX2_X1 _08681_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(fanout_net_36 ), .Z(_01145_ ) );
OR2_X1 _08682_ ( .A1(_01145_ ), .A2(_01042_ ), .ZN(_01146_ ) );
MUX2_X1 _08683_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(fanout_net_36 ), .Z(_01147_ ) );
OAI21_X1 _08684_ ( .A(_01146_ ), .B1(fanout_net_39 ), .B2(_01147_ ), .ZN(_01148_ ) );
INV_X1 _08685_ ( .A(\IF_ID_pc [28] ), .ZN(_01149_ ) );
XNOR2_X1 _08686_ ( .A(_01148_ ), .B(_01149_ ), .ZN(_01150_ ) );
AOI22_X1 _08687_ ( .A1(_01092_ ), .A2(\IF_ID_pc [9] ), .B1(_01102_ ), .B2(_01101_ ), .ZN(_01151_ ) );
AND3_X1 _08688_ ( .A1(_01144_ ), .A2(_01150_ ), .A3(_01151_ ), .ZN(_01152_ ) );
AND2_X1 _08689_ ( .A1(_01068_ ), .A2(\myifu.myicache.tag[2][17] ), .ZN(_01153_ ) );
AOI211_X1 _08690_ ( .A(_01014_ ), .B(_01153_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[3][17] ), .ZN(_01154_ ) );
AND2_X1 _08691_ ( .A1(_01043_ ), .A2(\myifu.myicache.tag[0][17] ), .ZN(_01155_ ) );
AOI211_X1 _08692_ ( .A(fanout_net_39 ), .B(_01155_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[1][17] ), .ZN(_01156_ ) );
NOR2_X1 _08693_ ( .A1(_01154_ ), .A2(_01156_ ), .ZN(_01157_ ) );
INV_X1 _08694_ ( .A(\IF_ID_pc [21] ), .ZN(_01158_ ) );
XNOR2_X1 _08695_ ( .A(_01157_ ), .B(_01158_ ), .ZN(_01159_ ) );
AND2_X1 _08696_ ( .A1(_01043_ ), .A2(\myifu.myicache.tag[2][19] ), .ZN(_01160_ ) );
AOI211_X1 _08697_ ( .A(_01042_ ), .B(_01160_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[3][19] ), .ZN(_01161_ ) );
AND2_X1 _08698_ ( .A1(_01043_ ), .A2(\myifu.myicache.tag[0][19] ), .ZN(_01162_ ) );
AOI211_X1 _08699_ ( .A(fanout_net_39 ), .B(_01162_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[1][19] ), .ZN(_01163_ ) );
NOR2_X1 _08700_ ( .A1(_01161_ ), .A2(_01163_ ), .ZN(_01164_ ) );
INV_X1 _08701_ ( .A(\IF_ID_pc [23] ), .ZN(_01165_ ) );
XNOR2_X1 _08702_ ( .A(_01164_ ), .B(_01165_ ), .ZN(_01166_ ) );
OR2_X1 _08703_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[0][10] ), .ZN(_01167_ ) );
OAI211_X1 _08704_ ( .A(_01167_ ), .B(_01014_ ), .C1(_01060_ ), .C2(\myifu.myicache.tag[1][10] ), .ZN(_01168_ ) );
OR2_X1 _08705_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[2][10] ), .ZN(_01169_ ) );
OAI211_X1 _08706_ ( .A(_01169_ ), .B(fanout_net_39 ), .C1(_01060_ ), .C2(\myifu.myicache.tag[3][10] ), .ZN(_01170_ ) );
AND3_X1 _08707_ ( .A1(_01168_ ), .A2(_01170_ ), .A3(\IF_ID_pc [14] ), .ZN(_01171_ ) );
AOI21_X1 _08708_ ( .A(\IF_ID_pc [14] ), .B1(_01168_ ), .B2(_01170_ ), .ZN(_01172_ ) );
NOR4_X1 _08709_ ( .A1(_01159_ ), .A2(_01166_ ), .A3(_01171_ ), .A4(_01172_ ), .ZN(_01173_ ) );
OR2_X1 _08710_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[0][23] ), .ZN(_01174_ ) );
OAI211_X1 _08711_ ( .A(_01174_ ), .B(_01014_ ), .C1(_01060_ ), .C2(\myifu.myicache.tag[1][23] ), .ZN(_01175_ ) );
OR2_X1 _08712_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[2][23] ), .ZN(_01176_ ) );
OAI211_X1 _08713_ ( .A(_01176_ ), .B(fanout_net_39 ), .C1(_01060_ ), .C2(\myifu.myicache.tag[3][23] ), .ZN(_01177_ ) );
NAND2_X1 _08714_ ( .A1(_01175_ ), .A2(_01177_ ), .ZN(_01178_ ) );
XNOR2_X1 _08715_ ( .A(_01178_ ), .B(\IF_ID_pc [27] ), .ZN(_01179_ ) );
AND2_X1 _08716_ ( .A1(_01043_ ), .A2(\myifu.myicache.tag[2][6] ), .ZN(_01180_ ) );
AOI211_X1 _08717_ ( .A(_01042_ ), .B(_01180_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[3][6] ), .ZN(_01181_ ) );
AND2_X1 _08718_ ( .A1(_01043_ ), .A2(\myifu.myicache.tag[0][6] ), .ZN(_01182_ ) );
AOI211_X1 _08719_ ( .A(fanout_net_39 ), .B(_01182_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[1][6] ), .ZN(_01183_ ) );
NOR2_X1 _08720_ ( .A1(_01181_ ), .A2(_01183_ ), .ZN(_01184_ ) );
XNOR2_X1 _08721_ ( .A(_01184_ ), .B(\IF_ID_pc [10] ), .ZN(_01185_ ) );
AND2_X1 _08722_ ( .A1(_01043_ ), .A2(\myifu.myicache.tag[2][2] ), .ZN(_01186_ ) );
AOI211_X1 _08723_ ( .A(_01042_ ), .B(_01186_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[3][2] ), .ZN(_01187_ ) );
AND2_X1 _08724_ ( .A1(_01024_ ), .A2(\myifu.myicache.tag[0][2] ), .ZN(_01188_ ) );
AOI211_X1 _08725_ ( .A(fanout_net_39 ), .B(_01188_ ), .C1(fanout_net_36 ), .C2(\myifu.myicache.tag[1][2] ), .ZN(_01189_ ) );
NOR2_X1 _08726_ ( .A1(_01187_ ), .A2(_01189_ ), .ZN(_01190_ ) );
XNOR2_X1 _08727_ ( .A(_01190_ ), .B(\IF_ID_pc [6] ), .ZN(_01191_ ) );
OR2_X1 _08728_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[0][4] ), .ZN(_01192_ ) );
OAI211_X1 _08729_ ( .A(_01192_ ), .B(_01014_ ), .C1(_01060_ ), .C2(\myifu.myicache.tag[1][4] ), .ZN(_01193_ ) );
OR2_X1 _08730_ ( .A1(fanout_net_36 ), .A2(\myifu.myicache.tag[2][4] ), .ZN(_01194_ ) );
OAI211_X1 _08731_ ( .A(_01194_ ), .B(fanout_net_39 ), .C1(_01060_ ), .C2(\myifu.myicache.tag[3][4] ), .ZN(_01195_ ) );
NAND2_X1 _08732_ ( .A1(_01193_ ), .A2(_01195_ ), .ZN(_01196_ ) );
XNOR2_X1 _08733_ ( .A(_01196_ ), .B(\IF_ID_pc [8] ), .ZN(_01197_ ) );
AND4_X1 _08734_ ( .A1(_01179_ ), .A2(_01185_ ), .A3(_01191_ ), .A4(_01197_ ), .ZN(_01198_ ) );
AND4_X1 _08735_ ( .A1(_01135_ ), .A2(_01152_ ), .A3(_01173_ ), .A4(_01198_ ), .ZN(_01199_ ) );
AND2_X4 _08736_ ( .A1(_01122_ ), .A2(_01199_ ), .ZN(_01200_ ) );
INV_X1 _08737_ ( .A(\myifu.state [0] ), .ZN(_01201_ ) );
NOR2_X4 _08738_ ( .A1(_01200_ ), .A2(_01201_ ), .ZN(_01202_ ) );
INV_X1 _08739_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01203_ ) );
NOR2_X4 _08740_ ( .A1(_01202_ ), .A2(_01203_ ), .ZN(_01204_ ) );
NOR2_X1 _08741_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01205_ ) );
NOR2_X4 _08742_ ( .A1(_01204_ ), .A2(_01205_ ), .ZN(_01206_ ) );
INV_X1 _08743_ ( .A(\EX_LS_flag [2] ), .ZN(_01207_ ) );
INV_X1 _08744_ ( .A(io_master_wready_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_01208_ ) );
NAND4_X1 _08745_ ( .A1(_01207_ ), .A2(_01208_ ), .A3(\EX_LS_flag [1] ), .A4(\EX_LS_flag [0] ), .ZN(_01209_ ) );
INV_X1 _08746_ ( .A(EXU_valid_LSU ), .ZN(_01210_ ) );
NOR2_X1 _08747_ ( .A1(_01209_ ), .A2(_01210_ ), .ZN(_01211_ ) );
INV_X1 _08748_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01212_ ) );
NOR2_X1 _08749_ ( .A1(_01211_ ), .A2(_01212_ ), .ZN(_01213_ ) );
NOR2_X4 _08750_ ( .A1(_01206_ ), .A2(_01213_ ), .ZN(_01214_ ) );
BUF_X4 _08751_ ( .A(_01214_ ), .Z(_01215_ ) );
CLKBUF_X2 _08752_ ( .A(_01209_ ), .Z(_01216_ ) );
CLKBUF_X2 _08753_ ( .A(_01210_ ), .Z(_01217_ ) );
OR3_X1 _08754_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(_01217_ ), .ZN(_01218_ ) );
BUF_X4 _08755_ ( .A(_01211_ ), .Z(_01219_ ) );
OAI211_X1 _08756_ ( .A(_01215_ ), .B(_01218_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01219_ ), .ZN(_01220_ ) );
INV_X4 _08757_ ( .A(_01206_ ), .ZN(_01221_ ) );
OAI21_X1 _08758_ ( .A(_01220_ ), .B1(_01102_ ), .B2(_01221_ ), .ZN(\io_master_araddr [19] ) );
CLKBUF_X2 _08759_ ( .A(_01209_ ), .Z(_01222_ ) );
CLKBUF_X2 _08760_ ( .A(_01210_ ), .Z(_01223_ ) );
OR3_X1 _08761_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(_01223_ ), .ZN(_01224_ ) );
BUF_X4 _08762_ ( .A(_01211_ ), .Z(_01225_ ) );
OAI211_X1 _08763_ ( .A(_01214_ ), .B(_01224_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01225_ ), .ZN(_01226_ ) );
OAI221_X1 _08764_ ( .A(\IF_ID_pc [20] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_01227_ ) );
AND2_X1 _08765_ ( .A1(_01226_ ), .A2(_01227_ ), .ZN(_01228_ ) );
INV_X1 _08766_ ( .A(_01228_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _08767_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(_01223_ ), .ZN(_01229_ ) );
OAI211_X1 _08768_ ( .A(_01215_ ), .B(_01229_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01225_ ), .ZN(_01230_ ) );
OAI21_X1 _08769_ ( .A(_01230_ ), .B1(_01149_ ), .B2(_01221_ ), .ZN(\io_master_araddr [28] ) );
OR3_X1 _08770_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(_01223_ ), .ZN(_01231_ ) );
OAI211_X1 _08771_ ( .A(_01215_ ), .B(_01231_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01219_ ), .ZN(_01232_ ) );
OAI21_X1 _08772_ ( .A(_01232_ ), .B1(_01110_ ), .B2(_01221_ ), .ZN(\io_master_araddr [18] ) );
OR4_X1 _08773_ ( .A1(\io_master_araddr [19] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [28] ), .A4(\io_master_araddr [18] ), .ZN(_01233_ ) );
OR3_X1 _08774_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(_01223_ ), .ZN(_01234_ ) );
OAI211_X1 _08775_ ( .A(_01214_ ), .B(_01234_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01225_ ), .ZN(_01235_ ) );
OAI221_X1 _08776_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_01236_ ) );
NAND2_X1 _08777_ ( .A1(_01235_ ), .A2(_01236_ ), .ZN(\io_master_araddr [31] ) );
OR3_X1 _08778_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(_01210_ ), .ZN(_01237_ ) );
OAI211_X1 _08779_ ( .A(_01214_ ), .B(_01237_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01211_ ), .ZN(_01238_ ) );
OAI21_X2 _08780_ ( .A(_01238_ ), .B1(_01123_ ), .B2(_01221_ ), .ZN(\io_master_araddr [17] ) );
INV_X1 _08781_ ( .A(_01213_ ), .ZN(_01239_ ) );
OR3_X1 _08782_ ( .A1(_01209_ ), .A2(\EX_LS_dest_csreg_mem [25] ), .A3(_01210_ ), .ZN(_01240_ ) );
OAI211_X1 _08783_ ( .A(_01239_ ), .B(_01240_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_01211_ ), .ZN(_01241_ ) );
INV_X1 _08784_ ( .A(\IF_ID_pc [25] ), .ZN(_01242_ ) );
MUX2_X1 _08785_ ( .A(_01241_ ), .B(_01242_ ), .S(_01206_ ), .Z(_01243_ ) );
INV_X1 _08786_ ( .A(_01243_ ), .ZN(\io_master_araddr [25] ) );
OR3_X1 _08787_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(_01210_ ), .ZN(_01244_ ) );
OAI211_X1 _08788_ ( .A(_01214_ ), .B(_01244_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01225_ ), .ZN(_01245_ ) );
OAI221_X1 _08789_ ( .A(\IF_ID_pc [22] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_01246_ ) );
NAND3_X1 _08790_ ( .A1(\io_master_araddr [25] ), .A2(_01245_ ), .A3(_01246_ ), .ZN(_01247_ ) );
NOR4_X1 _08791_ ( .A1(_01233_ ), .A2(\io_master_araddr [31] ), .A3(\io_master_araddr [17] ), .A4(_01247_ ), .ZN(_01248_ ) );
OR3_X1 _08792_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(_01223_ ), .ZN(_01249_ ) );
OAI211_X1 _08793_ ( .A(_01215_ ), .B(_01249_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01225_ ), .ZN(_01250_ ) );
OAI221_X1 _08794_ ( .A(\IF_ID_pc [23] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_01251_ ) );
AND2_X2 _08795_ ( .A1(_01250_ ), .A2(_01251_ ), .ZN(_01252_ ) );
INV_X1 _08796_ ( .A(_01252_ ), .ZN(\io_master_araddr [23] ) );
OR3_X1 _08797_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(_01210_ ), .ZN(_01253_ ) );
OAI211_X1 _08798_ ( .A(_01214_ ), .B(_01253_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01225_ ), .ZN(_01254_ ) );
OAI21_X1 _08799_ ( .A(_01254_ ), .B1(_01034_ ), .B2(_01221_ ), .ZN(\io_master_araddr [16] ) );
OR3_X1 _08800_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(_01217_ ), .ZN(_01255_ ) );
OAI211_X1 _08801_ ( .A(_01215_ ), .B(_01255_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01219_ ), .ZN(_01256_ ) );
INV_X1 _08802_ ( .A(\IF_ID_pc [29] ), .ZN(_01257_ ) );
BUF_X4 _08803_ ( .A(_01221_ ), .Z(_01258_ ) );
OAI21_X1 _08804_ ( .A(_01256_ ), .B1(_01257_ ), .B2(_01258_ ), .ZN(\io_master_araddr [29] ) );
OR3_X1 _08805_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(_01223_ ), .ZN(_01259_ ) );
OAI211_X1 _08806_ ( .A(_01215_ ), .B(_01259_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01219_ ), .ZN(_01260_ ) );
INV_X1 _08807_ ( .A(\IF_ID_pc [26] ), .ZN(_01261_ ) );
OAI21_X1 _08808_ ( .A(_01260_ ), .B1(_01261_ ), .B2(_01221_ ), .ZN(\io_master_araddr [26] ) );
NOR4_X1 _08809_ ( .A1(\io_master_araddr [23] ), .A2(\io_master_araddr [16] ), .A3(\io_master_araddr [29] ), .A4(\io_master_araddr [26] ), .ZN(_01262_ ) );
OR3_X1 _08810_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(_01223_ ), .ZN(_01263_ ) );
OAI211_X1 _08811_ ( .A(_01214_ ), .B(_01263_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01225_ ), .ZN(_01264_ ) );
OAI221_X1 _08812_ ( .A(\IF_ID_pc [21] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_01265_ ) );
AND2_X1 _08813_ ( .A1(_01264_ ), .A2(_01265_ ), .ZN(_01266_ ) );
INV_X1 _08814_ ( .A(_01266_ ), .ZN(\io_master_araddr [21] ) );
OR3_X1 _08815_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(_01223_ ), .ZN(_01267_ ) );
OAI211_X1 _08816_ ( .A(_01215_ ), .B(_01267_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01225_ ), .ZN(_01268_ ) );
OAI21_X1 _08817_ ( .A(_01268_ ), .B1(_01049_ ), .B2(_01221_ ), .ZN(\io_master_araddr [30] ) );
OR3_X1 _08818_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(_01223_ ), .ZN(_01269_ ) );
OAI211_X1 _08819_ ( .A(_01215_ ), .B(_01269_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01225_ ), .ZN(_01270_ ) );
OAI221_X1 _08820_ ( .A(\IF_ID_pc [24] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_01271_ ) );
NAND2_X1 _08821_ ( .A1(_01270_ ), .A2(_01271_ ), .ZN(\io_master_araddr [24] ) );
OR3_X1 _08822_ ( .A1(_01222_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(_01223_ ), .ZN(_01272_ ) );
OAI211_X1 _08823_ ( .A(_01214_ ), .B(_01272_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01225_ ), .ZN(_01273_ ) );
INV_X1 _08824_ ( .A(\IF_ID_pc [27] ), .ZN(_01274_ ) );
OAI21_X1 _08825_ ( .A(_01273_ ), .B1(_01274_ ), .B2(_01221_ ), .ZN(\io_master_araddr [27] ) );
NOR4_X1 _08826_ ( .A1(\io_master_araddr [21] ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [24] ), .A4(\io_master_araddr [27] ), .ZN(_01275_ ) );
AND2_X1 _08827_ ( .A1(_01262_ ), .A2(_01275_ ), .ZN(_01276_ ) );
CLKBUF_X2 _08828_ ( .A(_01206_ ), .Z(_01277_ ) );
NOR2_X1 _08829_ ( .A1(fanout_net_5 ), .A2(\EX_LS_dest_csreg_mem [1] ), .ZN(_01278_ ) );
INV_X1 _08830_ ( .A(_01278_ ), .ZN(_01279_ ) );
INV_X1 _08831_ ( .A(\EX_LS_typ [1] ), .ZN(_01280_ ) );
INV_X1 _08832_ ( .A(\EX_LS_typ [3] ), .ZN(_01281_ ) );
NAND4_X1 _08833_ ( .A1(_01279_ ), .A2(_01280_ ), .A3(_01281_ ), .A4(\EX_LS_typ [2] ), .ZN(_01282_ ) );
AND2_X1 _08834_ ( .A1(fanout_net_5 ), .A2(\EX_LS_typ [1] ), .ZN(_01283_ ) );
NOR2_X1 _08835_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_01284_ ) );
NAND2_X1 _08836_ ( .A1(_01283_ ), .A2(_01284_ ), .ZN(_01285_ ) );
AOI21_X1 _08837_ ( .A(\EX_LS_typ [0] ), .B1(_01282_ ), .B2(_01285_ ), .ZN(_01286_ ) );
AND3_X1 _08838_ ( .A1(_01283_ ), .A2(\EX_LS_typ [0] ), .A3(_01284_ ), .ZN(_01287_ ) );
OR2_X1 _08839_ ( .A1(_01286_ ), .A2(_01287_ ), .ZN(_01288_ ) );
AND2_X4 _08840_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_01289_ ) );
AND2_X1 _08841_ ( .A1(_01289_ ), .A2(_01207_ ), .ZN(_01290_ ) );
INV_X1 _08842_ ( .A(\EX_LS_typ [4] ), .ZN(_01291_ ) );
AND2_X1 _08843_ ( .A1(_01290_ ), .A2(_01291_ ), .ZN(_01292_ ) );
AND2_X1 _08844_ ( .A1(_01288_ ), .A2(_01292_ ), .ZN(_01293_ ) );
OR2_X1 _08845_ ( .A1(\EX_LS_dest_csreg_mem [24] ), .A2(\EX_LS_dest_csreg_mem [25] ), .ZN(_01294_ ) );
NOR3_X1 _08846_ ( .A1(_01294_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\EX_LS_dest_csreg_mem [26] ), .ZN(_01295_ ) );
NOR4_X1 _08847_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\EX_LS_dest_csreg_mem [29] ), .A4(\EX_LS_dest_csreg_mem [28] ), .ZN(_01296_ ) );
AND2_X1 _08848_ ( .A1(_01295_ ), .A2(_01296_ ), .ZN(_01297_ ) );
AND2_X1 _08849_ ( .A1(_01297_ ), .A2(_01290_ ), .ZN(_01298_ ) );
NOR2_X1 _08850_ ( .A1(_01293_ ), .A2(_01298_ ), .ZN(_01299_ ) );
INV_X32 _08851_ ( .A(\EX_LS_flag [1] ), .ZN(_01300_ ) );
NOR2_X4 _08852_ ( .A1(_01300_ ), .A2(\EX_LS_flag [0] ), .ZN(_01301_ ) );
BUF_X2 _08853_ ( .A(_01301_ ), .Z(_01302_ ) );
AND2_X2 _08854_ ( .A1(_01302_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_01303_ ) );
AND2_X1 _08855_ ( .A1(_01297_ ), .A2(_01303_ ), .ZN(_01304_ ) );
NAND3_X1 _08856_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_01305_ ) );
OAI21_X1 _08857_ ( .A(_01285_ ), .B1(_01278_ ), .B2(_01305_ ), .ZN(_01306_ ) );
NAND3_X1 _08858_ ( .A1(_01207_ ), .A2(_01291_ ), .A3(\EX_LS_typ [0] ), .ZN(_01307_ ) );
NOR3_X1 _08859_ ( .A1(_01307_ ), .A2(_01300_ ), .A3(\EX_LS_flag [0] ), .ZN(_01308_ ) );
AND2_X1 _08860_ ( .A1(_01306_ ), .A2(_01308_ ), .ZN(_01309_ ) );
NOR2_X1 _08861_ ( .A1(_01304_ ), .A2(_01309_ ), .ZN(_01310_ ) );
AND2_X1 _08862_ ( .A1(_01299_ ), .A2(_01310_ ), .ZN(_01311_ ) );
BUF_X4 _08863_ ( .A(_01311_ ), .Z(_01312_ ) );
AOI211_X1 _08864_ ( .A(_01212_ ), .B(_01277_ ), .C1(_01219_ ), .C2(_01312_ ), .ZN(_01313_ ) );
CLKBUF_X2 _08865_ ( .A(_01277_ ), .Z(_01314_ ) );
NOR3_X1 _08866_ ( .A1(_01200_ ), .A2(\myidu.stall_quest_fencei ), .A3(_01201_ ), .ZN(_01315_ ) );
INV_X1 _08867_ ( .A(_01315_ ), .ZN(_01316_ ) );
OAI211_X1 _08868_ ( .A(_01314_ ), .B(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .C1(fanout_net_2 ), .C2(_01316_ ), .ZN(_01317_ ) );
INV_X1 _08869_ ( .A(_01317_ ), .ZN(_01318_ ) );
NOR2_X1 _08870_ ( .A1(_01313_ ), .A2(_01318_ ), .ZN(_01319_ ) );
AND4_X1 _08871_ ( .A1(\myclint.rvalid ), .A2(_01248_ ), .A3(_01276_ ), .A4(_01319_ ), .ZN(_01320_ ) );
INV_X1 _08872_ ( .A(\myclint.rvalid ), .ZN(_01321_ ) );
NOR4_X2 _08873_ ( .A1(\io_master_araddr [29] ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [27] ), .A4(_01243_ ), .ZN(_01322_ ) );
NOR4_X1 _08874_ ( .A1(\io_master_araddr [26] ), .A2(\io_master_araddr [28] ), .A3(\io_master_araddr [24] ), .A4(\io_master_araddr [31] ), .ZN(_01323_ ) );
AND2_X4 _08875_ ( .A1(_01322_ ), .A2(_01323_ ), .ZN(_01324_ ) );
OR2_X2 _08876_ ( .A1(\io_master_araddr [16] ), .A2(\io_master_araddr [17] ), .ZN(_01325_ ) );
NOR3_X2 _08877_ ( .A1(_01325_ ), .A2(\io_master_araddr [19] ), .A3(\io_master_araddr [18] ), .ZN(_01326_ ) );
AND4_X1 _08878_ ( .A1(_01252_ ), .A2(_01324_ ), .A3(_01228_ ), .A4(_01326_ ), .ZN(_01327_ ) );
AND4_X1 _08879_ ( .A1(_01264_ ), .A2(_01245_ ), .A3(_01265_ ), .A4(_01246_ ), .ZN(_01328_ ) );
NAND2_X1 _08880_ ( .A1(_01327_ ), .A2(_01328_ ), .ZN(_01329_ ) );
AOI21_X1 _08881_ ( .A(_01314_ ), .B1(_01219_ ), .B2(_01312_ ), .ZN(_01330_ ) );
NOR2_X1 _08882_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_01331_ ) );
AOI211_X1 _08883_ ( .A(_01205_ ), .B(_01204_ ), .C1(\myifu.state [0] ), .C2(_01331_ ), .ZN(_01332_ ) );
OR3_X1 _08884_ ( .A1(_01329_ ), .A2(_01330_ ), .A3(_01332_ ), .ZN(_01333_ ) );
AOI211_X1 _08885_ ( .A(fanout_net_2 ), .B(_01320_ ), .C1(_01321_ ), .C2(_01333_ ), .ZN(_00064_ ) );
INV_X1 _08886_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_01334_ ) );
CLKBUF_X2 _08887_ ( .A(_01334_ ), .Z(_01335_ ) );
AND2_X1 _08888_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00065_ ) );
AND2_X1 _08889_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00066_ ) );
AND2_X1 _08890_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [21] ), .ZN(_00067_ ) );
AND2_X1 _08891_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [20] ), .ZN(_00068_ ) );
AND2_X1 _08892_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [19] ), .ZN(_00069_ ) );
AND2_X1 _08893_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [18] ), .ZN(_00070_ ) );
AND2_X1 _08894_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [17] ), .ZN(_00071_ ) );
AND2_X1 _08895_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00072_ ) );
INV_X1 _08896_ ( .A(\LS_WB_wdata_csreg [15] ), .ZN(_01336_ ) );
NOR2_X1 _08897_ ( .A1(_01336_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00073_ ) );
AND2_X1 _08898_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00074_ ) );
AND2_X1 _08899_ ( .A1(_01335_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00075_ ) );
CLKBUF_X2 _08900_ ( .A(_01334_ ), .Z(_01337_ ) );
AND2_X1 _08901_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00076_ ) );
AND2_X1 _08902_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00077_ ) );
AND2_X1 _08903_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00078_ ) );
AND2_X1 _08904_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00079_ ) );
AND2_X1 _08905_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [9] ), .ZN(_00080_ ) );
AND2_X1 _08906_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00081_ ) );
AND2_X1 _08907_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00082_ ) );
AND2_X1 _08908_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [6] ), .ZN(_00083_ ) );
AND2_X1 _08909_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00084_ ) );
AND2_X1 _08910_ ( .A1(_01337_ ), .A2(\LS_WB_wdata_csreg [4] ), .ZN(_00085_ ) );
AND2_X1 _08911_ ( .A1(_01334_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00086_ ) );
AND2_X1 _08912_ ( .A1(_01334_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00087_ ) );
AND2_X1 _08913_ ( .A1(_01334_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00088_ ) );
INV_X1 _08914_ ( .A(\LS_WB_wdata_csreg [25] ), .ZN(_01338_ ) );
NOR2_X1 _08915_ ( .A1(_01338_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00089_ ) );
AND2_X1 _08916_ ( .A1(_01334_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00090_ ) );
AND2_X1 _08917_ ( .A1(_01334_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00091_ ) );
AND2_X1 _08918_ ( .A1(_01334_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00092_ ) );
INV_X1 _08919_ ( .A(_01299_ ), .ZN(_01339_ ) );
INV_X1 _08920_ ( .A(exception_quest_IDU ), .ZN(_01340_ ) );
INV_X1 _08921_ ( .A(_01310_ ), .ZN(_01341_ ) );
NOR2_X1 _08922_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_01342_ ) );
NAND2_X1 _08923_ ( .A1(_01342_ ), .A2(_00830_ ), .ZN(_01343_ ) );
NOR4_X1 _08924_ ( .A1(_01339_ ), .A2(_01340_ ), .A3(_01341_ ), .A4(_01343_ ), .ZN(_00094_ ) );
BUF_X4 _08925_ ( .A(_01312_ ), .Z(_01344_ ) );
AOI21_X1 _08926_ ( .A(_01343_ ), .B1(_01344_ ), .B2(exception_quest_IDU ), .ZN(_00095_ ) );
NOR2_X1 _08927_ ( .A1(fanout_net_2 ), .A2(fanout_net_9 ), .ZN(_01345_ ) );
INV_X1 _08928_ ( .A(_01345_ ), .ZN(_01346_ ) );
INV_X1 _08929_ ( .A(IDU_valid_EXU ), .ZN(_01347_ ) );
NOR2_X1 _08930_ ( .A1(_01347_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _08931_ ( .A(\ID_EX_typ [6] ), .ZN(_01348_ ) );
INV_X1 _08932_ ( .A(fanout_net_6 ), .ZN(_01349_ ) );
BUF_X4 _08933_ ( .A(_01349_ ), .Z(_01350_ ) );
BUF_X4 _08934_ ( .A(_01350_ ), .Z(_01351_ ) );
NAND4_X1 _08935_ ( .A1(_01348_ ), .A2(_01351_ ), .A3(\ID_EX_typ [7] ), .A4(\ID_EX_typ [5] ), .ZN(_01352_ ) );
INV_X1 _08936_ ( .A(check_quest ), .ZN(_01353_ ) );
NOR2_X1 _08937_ ( .A1(_01353_ ), .A2(check_assert ), .ZN(_01354_ ) );
INV_X2 _08938_ ( .A(\ID_EX_typ [7] ), .ZN(_01355_ ) );
NOR2_X1 _08939_ ( .A1(_01355_ ), .A2(\ID_EX_typ [5] ), .ZN(_01356_ ) );
NAND2_X1 _08940_ ( .A1(_01356_ ), .A2(_01348_ ), .ZN(_01357_ ) );
MUX2_X1 _08941_ ( .A(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .B(_01354_ ), .S(_01357_ ), .Z(_01358_ ) );
INV_X1 _08942_ ( .A(\ID_EX_typ [5] ), .ZN(_01359_ ) );
NOR2_X1 _08943_ ( .A1(_01359_ ), .A2(\ID_EX_typ [6] ), .ZN(_01360_ ) );
AND2_X1 _08944_ ( .A1(_01360_ ), .A2(\ID_EX_typ [7] ), .ZN(_01361_ ) );
BUF_X4 _08945_ ( .A(_01361_ ), .Z(_01362_ ) );
OAI211_X1 _08946_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .B(_01352_ ), .C1(_01358_ ), .C2(_01362_ ), .ZN(_01363_ ) );
OAI21_X1 _08947_ ( .A(_01354_ ), .B1(EXU_valid_LSU ), .B2(_01347_ ), .ZN(_01364_ ) );
AOI21_X1 _08948_ ( .A(_01346_ ), .B1(_01363_ ), .B2(_01364_ ), .ZN(_00096_ ) );
AND2_X2 _08949_ ( .A1(_01356_ ), .A2(\ID_EX_typ [6] ), .ZN(_01365_ ) );
AND2_X1 _08950_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_01366_ ) );
AND2_X2 _08951_ ( .A1(_01366_ ), .A2(\ID_EX_typ [7] ), .ZN(_01367_ ) );
NOR2_X1 _08952_ ( .A1(_01365_ ), .A2(_01367_ ), .ZN(_01368_ ) );
INV_X1 _08953_ ( .A(_01368_ ), .ZN(_01369_ ) );
BUF_X4 _08954_ ( .A(_01369_ ), .Z(_01370_ ) );
AND2_X4 _08955_ ( .A1(_01301_ ), .A2(\EX_LS_flag [2] ), .ZN(_01371_ ) );
AND3_X1 _08956_ ( .A1(_01300_ ), .A2(\EX_LS_flag [0] ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_01372_ ) );
OR2_X4 _08957_ ( .A1(_01371_ ), .A2(_01372_ ), .ZN(_01373_ ) );
INV_X16 _08958_ ( .A(\EX_LS_flag [0] ), .ZN(_01374_ ) );
NOR2_X2 _08959_ ( .A1(_01374_ ), .A2(\EX_LS_flag [1] ), .ZN(_01375_ ) );
MUX2_X2 _08960_ ( .A(_01289_ ), .B(_01375_ ), .S(\EX_LS_flag [2] ), .Z(_01376_ ) );
NOR2_X4 _08961_ ( .A1(_01373_ ), .A2(_01376_ ), .ZN(_01377_ ) );
XOR2_X1 _08962_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .Z(_01378_ ) );
NOR4_X1 _08963_ ( .A1(\EX_LS_dest_reg [3] ), .A2(\EX_LS_dest_reg [2] ), .A3(\EX_LS_dest_reg [1] ), .A4(\EX_LS_dest_reg [0] ), .ZN(_01379_ ) );
INV_X2 _08964_ ( .A(\EX_LS_dest_reg [4] ), .ZN(_01380_ ) );
AND2_X1 _08965_ ( .A1(_01379_ ), .A2(_01380_ ), .ZN(_01381_ ) );
INV_X4 _08966_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_01382_ ) );
AND2_X1 _08967_ ( .A1(_01382_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_01383_ ) );
OR4_X4 _08968_ ( .A1(_01377_ ), .A2(_01378_ ), .A3(_01381_ ), .A4(_01383_ ), .ZN(_01384_ ) );
BUF_X8 _08969_ ( .A(_01384_ ), .Z(_01385_ ) );
BUF_X4 _08970_ ( .A(_01385_ ), .Z(_01386_ ) );
BUF_X2 _08971_ ( .A(_01386_ ), .Z(_01387_ ) );
BUF_X2 _08972_ ( .A(_01387_ ), .Z(_01388_ ) );
BUF_X2 _08973_ ( .A(_01388_ ), .Z(_01389_ ) );
XOR2_X1 _08974_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .Z(_01390_ ) );
XOR2_X1 _08975_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .Z(_01391_ ) );
INV_X1 _08976_ ( .A(\ID_EX_rs1 [3] ), .ZN(_01392_ ) );
OAI22_X1 _08977_ ( .A1(_01392_ ), .A2(\EX_LS_dest_reg [3] ), .B1(_01382_ ), .B2(\ID_EX_rs1 [1] ), .ZN(_01393_ ) );
INV_X1 _08978_ ( .A(\EX_LS_dest_reg [3] ), .ZN(_01394_ ) );
OAI21_X1 _08979_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_01394_ ), .B2(\ID_EX_rs1 [3] ), .ZN(_01395_ ) );
OR4_X4 _08980_ ( .A1(_01390_ ), .A2(_01391_ ), .A3(_01393_ ), .A4(_01395_ ), .ZN(_01396_ ) );
BUF_X4 _08981_ ( .A(_01396_ ), .Z(_01397_ ) );
BUF_X2 _08982_ ( .A(_01397_ ), .Z(_01398_ ) );
CLKBUF_X2 _08983_ ( .A(_01398_ ), .Z(_01399_ ) );
OR3_X1 _08984_ ( .A1(_01389_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_01399_ ), .ZN(_01400_ ) );
INV_X1 _08985_ ( .A(fanout_net_22 ), .ZN(_01401_ ) );
BUF_X4 _08986_ ( .A(_01401_ ), .Z(_01402_ ) );
BUF_X4 _08987_ ( .A(_01402_ ), .Z(_01403_ ) );
BUF_X4 _08988_ ( .A(_01403_ ), .Z(_01404_ ) );
INV_X1 _08989_ ( .A(fanout_net_21 ), .ZN(_01405_ ) );
BUF_X4 _08990_ ( .A(_01405_ ), .Z(_01406_ ) );
BUF_X4 _08991_ ( .A(_01406_ ), .Z(_01407_ ) );
BUF_X4 _08992_ ( .A(_01407_ ), .Z(_01408_ ) );
BUF_X4 _08993_ ( .A(_01408_ ), .Z(_01409_ ) );
BUF_X4 _08994_ ( .A(_01409_ ), .Z(_01410_ ) );
INV_X1 _08995_ ( .A(fanout_net_10 ), .ZN(_01411_ ) );
BUF_X4 _08996_ ( .A(_01411_ ), .Z(_01412_ ) );
BUF_X4 _08997_ ( .A(_01412_ ), .Z(_01413_ ) );
BUF_X4 _08998_ ( .A(_01413_ ), .Z(_01414_ ) );
BUF_X4 _08999_ ( .A(_01414_ ), .Z(_01415_ ) );
BUF_X4 _09000_ ( .A(_01415_ ), .Z(_01416_ ) );
BUF_X4 _09001_ ( .A(_01416_ ), .Z(_01417_ ) );
OAI21_X1 _09002_ ( .A(fanout_net_18 ), .B1(_01417_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01418_ ) );
NOR2_X1 _09003_ ( .A1(fanout_net_10 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01419_ ) );
NOR2_X1 _09004_ ( .A1(fanout_net_10 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01420_ ) );
INV_X1 _09005_ ( .A(fanout_net_18 ), .ZN(_01421_ ) );
BUF_X4 _09006_ ( .A(_01421_ ), .Z(_01422_ ) );
BUF_X4 _09007_ ( .A(_01422_ ), .Z(_01423_ ) );
BUF_X4 _09008_ ( .A(_01423_ ), .Z(_01424_ ) );
BUF_X4 _09009_ ( .A(_01424_ ), .Z(_01425_ ) );
BUF_X4 _09010_ ( .A(_01425_ ), .Z(_01426_ ) );
BUF_X4 _09011_ ( .A(_01426_ ), .Z(_01427_ ) );
OAI21_X1 _09012_ ( .A(_01427_ ), .B1(_01417_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01428_ ) );
OAI221_X1 _09013_ ( .A(_01410_ ), .B1(_01418_ ), .B2(_01419_ ), .C1(_01420_ ), .C2(_01428_ ), .ZN(_01429_ ) );
MUX2_X1 _09014_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01430_ ) );
MUX2_X1 _09015_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01431_ ) );
MUX2_X1 _09016_ ( .A(_01430_ ), .B(_01431_ ), .S(fanout_net_18 ), .Z(_01432_ ) );
BUF_X4 _09017_ ( .A(_01409_ ), .Z(_01433_ ) );
OAI211_X1 _09018_ ( .A(_01404_ ), .B(_01429_ ), .C1(_01432_ ), .C2(_01433_ ), .ZN(_01434_ ) );
NOR2_X1 _09019_ ( .A1(_01417_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01435_ ) );
OAI21_X1 _09020_ ( .A(fanout_net_18 ), .B1(fanout_net_10 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01436_ ) );
NOR2_X1 _09021_ ( .A1(fanout_net_10 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01437_ ) );
OAI21_X1 _09022_ ( .A(_01427_ ), .B1(_01417_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01438_ ) );
OAI221_X1 _09023_ ( .A(fanout_net_21 ), .B1(_01435_ ), .B2(_01436_ ), .C1(_01437_ ), .C2(_01438_ ), .ZN(_01439_ ) );
MUX2_X1 _09024_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01440_ ) );
MUX2_X1 _09025_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01441_ ) );
MUX2_X1 _09026_ ( .A(_01440_ ), .B(_01441_ ), .S(_01427_ ), .Z(_01442_ ) );
OAI211_X1 _09027_ ( .A(fanout_net_22 ), .B(_01439_ ), .C1(_01442_ ), .C2(fanout_net_21 ), .ZN(_01443_ ) );
BUF_X2 _09028_ ( .A(_01399_ ), .Z(_01444_ ) );
OAI211_X1 _09029_ ( .A(_01434_ ), .B(_01443_ ), .C1(_01389_ ), .C2(_01444_ ), .ZN(_01445_ ) );
AND2_X2 _09030_ ( .A1(_01400_ ), .A2(_01445_ ), .ZN(_01446_ ) );
INV_X1 _09031_ ( .A(\ID_EX_imm [30] ), .ZN(_01447_ ) );
XNOR2_X1 _09032_ ( .A(_01446_ ), .B(_01447_ ), .ZN(_01448_ ) );
OR3_X1 _09033_ ( .A1(_01389_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01444_ ), .ZN(_01449_ ) );
OR2_X1 _09034_ ( .A1(_01416_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01450_ ) );
BUF_X4 _09035_ ( .A(_01426_ ), .Z(_01451_ ) );
BUF_X4 _09036_ ( .A(_01451_ ), .Z(_01452_ ) );
OAI211_X1 _09037_ ( .A(_01450_ ), .B(_01452_ ), .C1(fanout_net_10 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01453_ ) );
OR2_X1 _09038_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01454_ ) );
BUF_X4 _09039_ ( .A(_01416_ ), .Z(_01455_ ) );
OAI211_X1 _09040_ ( .A(_01454_ ), .B(fanout_net_18 ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01456_ ) );
NAND3_X1 _09041_ ( .A1(_01453_ ), .A2(_01433_ ), .A3(_01456_ ), .ZN(_01457_ ) );
MUX2_X1 _09042_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01458_ ) );
MUX2_X1 _09043_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01459_ ) );
MUX2_X1 _09044_ ( .A(_01458_ ), .B(_01459_ ), .S(_01452_ ), .Z(_01460_ ) );
OAI211_X1 _09045_ ( .A(_01404_ ), .B(_01457_ ), .C1(_01460_ ), .C2(_01433_ ), .ZN(_01461_ ) );
OR2_X1 _09046_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01462_ ) );
OAI211_X1 _09047_ ( .A(_01462_ ), .B(_01452_ ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01463_ ) );
NOR2_X1 _09048_ ( .A1(_01455_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01464_ ) );
OAI21_X1 _09049_ ( .A(fanout_net_18 ), .B1(fanout_net_10 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01465_ ) );
OAI211_X1 _09050_ ( .A(_01463_ ), .B(fanout_net_21 ), .C1(_01464_ ), .C2(_01465_ ), .ZN(_01466_ ) );
MUX2_X1 _09051_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01467_ ) );
MUX2_X1 _09052_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01468_ ) );
MUX2_X1 _09053_ ( .A(_01467_ ), .B(_01468_ ), .S(fanout_net_18 ), .Z(_01469_ ) );
OAI211_X1 _09054_ ( .A(fanout_net_22 ), .B(_01466_ ), .C1(_01469_ ), .C2(fanout_net_21 ), .ZN(_01470_ ) );
OAI211_X1 _09055_ ( .A(_01461_ ), .B(_01470_ ), .C1(_01389_ ), .C2(_01444_ ), .ZN(_01471_ ) );
NAND2_X2 _09056_ ( .A1(_01449_ ), .A2(_01471_ ), .ZN(_01472_ ) );
INV_X1 _09057_ ( .A(\ID_EX_imm [27] ), .ZN(_01473_ ) );
XNOR2_X1 _09058_ ( .A(_01472_ ), .B(_01473_ ), .ZN(_01474_ ) );
OR3_X1 _09059_ ( .A1(_01388_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01399_ ), .ZN(_01475_ ) );
OR2_X1 _09060_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01476_ ) );
BUF_X4 _09061_ ( .A(_01416_ ), .Z(_01477_ ) );
OAI211_X1 _09062_ ( .A(_01476_ ), .B(_01451_ ), .C1(_01477_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01478_ ) );
OR2_X1 _09063_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01479_ ) );
OAI211_X1 _09064_ ( .A(_01479_ ), .B(fanout_net_18 ), .C1(_01477_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01480_ ) );
NAND3_X1 _09065_ ( .A1(_01478_ ), .A2(_01480_ ), .A3(_01410_ ), .ZN(_01481_ ) );
MUX2_X1 _09066_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01482_ ) );
MUX2_X1 _09067_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01483_ ) );
MUX2_X1 _09068_ ( .A(_01482_ ), .B(_01483_ ), .S(_01451_ ), .Z(_01484_ ) );
OAI211_X1 _09069_ ( .A(_01404_ ), .B(_01481_ ), .C1(_01484_ ), .C2(_01410_ ), .ZN(_01485_ ) );
OR2_X1 _09070_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01486_ ) );
OAI211_X1 _09071_ ( .A(_01486_ ), .B(fanout_net_18 ), .C1(_01477_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01487_ ) );
OR2_X1 _09072_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01488_ ) );
OAI211_X1 _09073_ ( .A(_01488_ ), .B(_01451_ ), .C1(_01477_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01489_ ) );
NAND3_X1 _09074_ ( .A1(_01487_ ), .A2(_01489_ ), .A3(fanout_net_21 ), .ZN(_01490_ ) );
MUX2_X1 _09075_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01491_ ) );
MUX2_X1 _09076_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01492_ ) );
MUX2_X1 _09077_ ( .A(_01491_ ), .B(_01492_ ), .S(fanout_net_18 ), .Z(_01493_ ) );
OAI211_X1 _09078_ ( .A(fanout_net_22 ), .B(_01490_ ), .C1(_01493_ ), .C2(fanout_net_21 ), .ZN(_01494_ ) );
OAI211_X1 _09079_ ( .A(_01485_ ), .B(_01494_ ), .C1(_01388_ ), .C2(_01399_ ), .ZN(_01495_ ) );
NAND2_X1 _09080_ ( .A1(_01475_ ), .A2(_01495_ ), .ZN(_01496_ ) );
INV_X1 _09081_ ( .A(\ID_EX_imm [24] ), .ZN(_01497_ ) );
XNOR2_X1 _09082_ ( .A(_01496_ ), .B(_01497_ ), .ZN(_01498_ ) );
INV_X1 _09083_ ( .A(_01498_ ), .ZN(_01499_ ) );
OR3_X1 _09084_ ( .A1(_01384_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01396_ ), .ZN(_01500_ ) );
OR2_X1 _09085_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01501_ ) );
OAI211_X1 _09086_ ( .A(_01501_ ), .B(_01423_ ), .C1(_01412_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01502_ ) );
OR2_X1 _09087_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01503_ ) );
BUF_X4 _09088_ ( .A(_01411_ ), .Z(_01504_ ) );
OAI211_X1 _09089_ ( .A(_01503_ ), .B(fanout_net_18 ), .C1(_01504_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01505_ ) );
NAND3_X1 _09090_ ( .A1(_01502_ ), .A2(_01505_ ), .A3(_01405_ ), .ZN(_01506_ ) );
MUX2_X1 _09091_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01507_ ) );
MUX2_X1 _09092_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_10 ), .Z(_01508_ ) );
MUX2_X1 _09093_ ( .A(_01507_ ), .B(_01508_ ), .S(_01422_ ), .Z(_01509_ ) );
OAI211_X1 _09094_ ( .A(fanout_net_22 ), .B(_01506_ ), .C1(_01509_ ), .C2(_01406_ ), .ZN(_01510_ ) );
OR2_X1 _09095_ ( .A1(fanout_net_10 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01511_ ) );
OAI211_X1 _09096_ ( .A(_01511_ ), .B(_01423_ ), .C1(_01412_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01512_ ) );
OR2_X1 _09097_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01513_ ) );
OAI211_X1 _09098_ ( .A(_01513_ ), .B(fanout_net_18 ), .C1(_01504_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01514_ ) );
NAND3_X1 _09099_ ( .A1(_01512_ ), .A2(_01514_ ), .A3(_01405_ ), .ZN(_01515_ ) );
MUX2_X1 _09100_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01516_ ) );
MUX2_X1 _09101_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01517_ ) );
MUX2_X1 _09102_ ( .A(_01516_ ), .B(_01517_ ), .S(_01422_ ), .Z(_01518_ ) );
OAI211_X1 _09103_ ( .A(_01401_ ), .B(_01515_ ), .C1(_01518_ ), .C2(_01406_ ), .ZN(_01519_ ) );
OAI211_X1 _09104_ ( .A(_01510_ ), .B(_01519_ ), .C1(_01385_ ), .C2(_01397_ ), .ZN(_01520_ ) );
NAND2_X2 _09105_ ( .A1(_01500_ ), .A2(_01520_ ), .ZN(_01521_ ) );
INV_X1 _09106_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_01522_ ) );
XNOR2_X2 _09107_ ( .A(_01521_ ), .B(_01522_ ), .ZN(_01523_ ) );
OR3_X2 _09108_ ( .A1(_01384_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01396_ ), .ZN(_01524_ ) );
OR2_X1 _09109_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01525_ ) );
BUF_X4 _09110_ ( .A(_01422_ ), .Z(_01526_ ) );
BUF_X4 _09111_ ( .A(_01504_ ), .Z(_01527_ ) );
OAI211_X1 _09112_ ( .A(_01525_ ), .B(_01526_ ), .C1(_01527_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01528_ ) );
OR2_X1 _09113_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01529_ ) );
OAI211_X1 _09114_ ( .A(_01529_ ), .B(fanout_net_18 ), .C1(_01412_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01530_ ) );
NAND3_X1 _09115_ ( .A1(_01528_ ), .A2(_01530_ ), .A3(_01406_ ), .ZN(_01531_ ) );
MUX2_X1 _09116_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01532_ ) );
MUX2_X1 _09117_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01533_ ) );
MUX2_X1 _09118_ ( .A(_01532_ ), .B(_01533_ ), .S(_01423_ ), .Z(_01534_ ) );
BUF_X4 _09119_ ( .A(_01405_ ), .Z(_01535_ ) );
OAI211_X1 _09120_ ( .A(_01402_ ), .B(_01531_ ), .C1(_01534_ ), .C2(_01535_ ), .ZN(_01536_ ) );
OR2_X1 _09121_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01537_ ) );
OAI211_X1 _09122_ ( .A(_01537_ ), .B(fanout_net_18 ), .C1(_01527_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01538_ ) );
OR2_X1 _09123_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01539_ ) );
OAI211_X1 _09124_ ( .A(_01539_ ), .B(_01526_ ), .C1(_01412_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01540_ ) );
NAND3_X1 _09125_ ( .A1(_01538_ ), .A2(_01540_ ), .A3(fanout_net_21 ), .ZN(_01541_ ) );
MUX2_X1 _09126_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01542_ ) );
MUX2_X1 _09127_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01543_ ) );
MUX2_X1 _09128_ ( .A(_01542_ ), .B(_01543_ ), .S(fanout_net_18 ), .Z(_01544_ ) );
OAI211_X1 _09129_ ( .A(fanout_net_22 ), .B(_01541_ ), .C1(_01544_ ), .C2(fanout_net_21 ), .ZN(_01545_ ) );
OAI211_X1 _09130_ ( .A(_01536_ ), .B(_01545_ ), .C1(_01385_ ), .C2(_01397_ ), .ZN(_01546_ ) );
NAND2_X2 _09131_ ( .A1(_01524_ ), .A2(_01546_ ), .ZN(_01547_ ) );
INV_X1 _09132_ ( .A(\ID_EX_imm [2] ), .ZN(_01548_ ) );
XNOR2_X1 _09133_ ( .A(_01547_ ), .B(_01548_ ), .ZN(_01549_ ) );
INV_X1 _09134_ ( .A(_01549_ ), .ZN(_01550_ ) );
OR3_X4 _09135_ ( .A1(_01384_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01396_ ), .ZN(_01551_ ) );
OR2_X1 _09136_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01552_ ) );
OAI211_X1 _09137_ ( .A(_01552_ ), .B(_01422_ ), .C1(_01411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01553_ ) );
OR2_X1 _09138_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01554_ ) );
OAI211_X1 _09139_ ( .A(_01554_ ), .B(fanout_net_18 ), .C1(_01411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01555_ ) );
NAND3_X1 _09140_ ( .A1(_01553_ ), .A2(_01555_ ), .A3(_01405_ ), .ZN(_01556_ ) );
MUX2_X1 _09141_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01557_ ) );
MUX2_X1 _09142_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01558_ ) );
MUX2_X1 _09143_ ( .A(_01557_ ), .B(_01558_ ), .S(_01422_ ), .Z(_01559_ ) );
OAI211_X1 _09144_ ( .A(fanout_net_22 ), .B(_01556_ ), .C1(_01559_ ), .C2(_01405_ ), .ZN(_01560_ ) );
OR2_X1 _09145_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01561_ ) );
OAI211_X1 _09146_ ( .A(_01561_ ), .B(_01422_ ), .C1(_01411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01562_ ) );
OR2_X1 _09147_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01563_ ) );
OAI211_X1 _09148_ ( .A(_01563_ ), .B(fanout_net_18 ), .C1(_01411_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01564_ ) );
NAND3_X1 _09149_ ( .A1(_01562_ ), .A2(_01564_ ), .A3(fanout_net_21 ), .ZN(_01565_ ) );
MUX2_X1 _09150_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01566_ ) );
MUX2_X1 _09151_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01567_ ) );
MUX2_X1 _09152_ ( .A(_01566_ ), .B(_01567_ ), .S(_01421_ ), .Z(_01568_ ) );
OAI211_X1 _09153_ ( .A(_01401_ ), .B(_01565_ ), .C1(_01568_ ), .C2(fanout_net_21 ), .ZN(_01569_ ) );
OAI211_X1 _09154_ ( .A(_01560_ ), .B(_01569_ ), .C1(_01384_ ), .C2(_01396_ ), .ZN(_01570_ ) );
NAND2_X4 _09155_ ( .A1(_01551_ ), .A2(_01570_ ), .ZN(_01571_ ) );
NAND2_X1 _09156_ ( .A1(_01571_ ), .A2(\ID_EX_imm [1] ), .ZN(_01572_ ) );
INV_X1 _09157_ ( .A(\ID_EX_imm [1] ), .ZN(_01573_ ) );
XNOR2_X1 _09158_ ( .A(_01571_ ), .B(_01573_ ), .ZN(_01574_ ) );
INV_X1 _09159_ ( .A(\ID_EX_imm [0] ), .ZN(_01575_ ) );
OR3_X4 _09160_ ( .A1(_01385_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_01397_ ), .ZN(_01576_ ) );
OR2_X1 _09161_ ( .A1(fanout_net_11 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01577_ ) );
OAI211_X1 _09162_ ( .A(_01577_ ), .B(_01526_ ), .C1(_01527_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01578_ ) );
OR2_X1 _09163_ ( .A1(fanout_net_11 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01579_ ) );
OAI211_X1 _09164_ ( .A(_01579_ ), .B(fanout_net_18 ), .C1(_01527_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01580_ ) );
NAND3_X1 _09165_ ( .A1(_01578_ ), .A2(_01580_ ), .A3(fanout_net_21 ), .ZN(_01581_ ) );
MUX2_X1 _09166_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01582_ ) );
MUX2_X1 _09167_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01583_ ) );
MUX2_X1 _09168_ ( .A(_01582_ ), .B(_01583_ ), .S(_01526_ ), .Z(_01584_ ) );
OAI211_X1 _09169_ ( .A(_01402_ ), .B(_01581_ ), .C1(_01584_ ), .C2(fanout_net_21 ), .ZN(_01585_ ) );
NOR2_X1 _09170_ ( .A1(_01527_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01586_ ) );
OAI21_X1 _09171_ ( .A(fanout_net_18 ), .B1(fanout_net_11 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01587_ ) );
NOR2_X1 _09172_ ( .A1(fanout_net_11 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01588_ ) );
OAI21_X1 _09173_ ( .A(_01526_ ), .B1(_01527_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01589_ ) );
OAI221_X1 _09174_ ( .A(_01406_ ), .B1(_01586_ ), .B2(_01587_ ), .C1(_01588_ ), .C2(_01589_ ), .ZN(_01590_ ) );
MUX2_X1 _09175_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01591_ ) );
MUX2_X1 _09176_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01592_ ) );
MUX2_X1 _09177_ ( .A(_01591_ ), .B(_01592_ ), .S(fanout_net_18 ), .Z(_01593_ ) );
OAI211_X1 _09178_ ( .A(fanout_net_22 ), .B(_01590_ ), .C1(_01593_ ), .C2(_01535_ ), .ZN(_01594_ ) );
OAI211_X1 _09179_ ( .A(_01585_ ), .B(_01594_ ), .C1(_01385_ ), .C2(_01397_ ), .ZN(_01595_ ) );
AOI21_X1 _09180_ ( .A(_01575_ ), .B1(_01576_ ), .B2(_01595_ ), .ZN(_01596_ ) );
NAND2_X1 _09181_ ( .A1(_01574_ ), .A2(_01596_ ), .ZN(_01597_ ) );
AOI211_X2 _09182_ ( .A(_01523_ ), .B(_01550_ ), .C1(_01572_ ), .C2(_01597_ ), .ZN(_01598_ ) );
NAND2_X1 _09183_ ( .A1(_01547_ ), .A2(\ID_EX_imm [2] ), .ZN(_01599_ ) );
OR2_X1 _09184_ ( .A1(_01523_ ), .A2(_01599_ ), .ZN(_01600_ ) );
INV_X1 _09185_ ( .A(_01521_ ), .ZN(_01601_ ) );
OAI21_X1 _09186_ ( .A(_01600_ ), .B1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ), .B2(_01601_ ), .ZN(_01602_ ) );
NOR2_X1 _09187_ ( .A1(_01598_ ), .A2(_01602_ ), .ZN(_01603_ ) );
INV_X1 _09188_ ( .A(\ID_EX_imm [4] ), .ZN(_01604_ ) );
BUF_X4 _09189_ ( .A(_01385_ ), .Z(_01605_ ) );
BUF_X4 _09190_ ( .A(_01397_ ), .Z(_01606_ ) );
OR3_X4 _09191_ ( .A1(_01605_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01606_ ), .ZN(_01607_ ) );
OR2_X1 _09192_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01608_ ) );
BUF_X4 _09193_ ( .A(_01526_ ), .Z(_01609_ ) );
BUF_X4 _09194_ ( .A(_01527_ ), .Z(_01610_ ) );
OAI211_X1 _09195_ ( .A(_01608_ ), .B(_01609_ ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01611_ ) );
OR2_X1 _09196_ ( .A1(fanout_net_11 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01612_ ) );
OAI211_X1 _09197_ ( .A(_01612_ ), .B(fanout_net_18 ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01613_ ) );
NAND3_X1 _09198_ ( .A1(_01611_ ), .A2(_01613_ ), .A3(_01407_ ), .ZN(_01614_ ) );
MUX2_X1 _09199_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_11 ), .Z(_01615_ ) );
MUX2_X1 _09200_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01616_ ) );
MUX2_X1 _09201_ ( .A(_01615_ ), .B(_01616_ ), .S(_01609_ ), .Z(_01617_ ) );
OAI211_X1 _09202_ ( .A(_01403_ ), .B(_01614_ ), .C1(_01617_ ), .C2(_01407_ ), .ZN(_01618_ ) );
OR2_X1 _09203_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01619_ ) );
OAI211_X1 _09204_ ( .A(_01619_ ), .B(fanout_net_18 ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01620_ ) );
OR2_X1 _09205_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01621_ ) );
OAI211_X1 _09206_ ( .A(_01621_ ), .B(_01609_ ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01622_ ) );
NAND3_X1 _09207_ ( .A1(_01620_ ), .A2(_01622_ ), .A3(fanout_net_21 ), .ZN(_01623_ ) );
MUX2_X1 _09208_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01624_ ) );
MUX2_X1 _09209_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01625_ ) );
MUX2_X1 _09210_ ( .A(_01624_ ), .B(_01625_ ), .S(fanout_net_18 ), .Z(_01626_ ) );
OAI211_X1 _09211_ ( .A(fanout_net_22 ), .B(_01623_ ), .C1(_01626_ ), .C2(fanout_net_21 ), .ZN(_01627_ ) );
OAI211_X1 _09212_ ( .A(_01618_ ), .B(_01627_ ), .C1(_01386_ ), .C2(_01398_ ), .ZN(_01628_ ) );
AOI21_X1 _09213_ ( .A(_01604_ ), .B1(_01607_ ), .B2(_01628_ ), .ZN(_01629_ ) );
AND3_X1 _09214_ ( .A1(_01607_ ), .A2(_01604_ ), .A3(_01628_ ), .ZN(_01630_ ) );
NOR3_X2 _09215_ ( .A1(_01603_ ), .A2(_01629_ ), .A3(_01630_ ), .ZN(_01631_ ) );
NOR2_X1 _09216_ ( .A1(_01631_ ), .A2(_01629_ ), .ZN(_01632_ ) );
NOR2_X4 _09217_ ( .A1(_01605_ ), .A2(_01606_ ), .ZN(_01633_ ) );
NAND2_X1 _09218_ ( .A1(_01633_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_01634_ ) );
OR2_X1 _09219_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01635_ ) );
OAI211_X1 _09220_ ( .A(_01635_ ), .B(_01424_ ), .C1(_01413_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01636_ ) );
OR2_X1 _09221_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01637_ ) );
BUF_X4 _09222_ ( .A(_01412_ ), .Z(_01638_ ) );
OAI211_X1 _09223_ ( .A(_01637_ ), .B(fanout_net_18 ), .C1(_01638_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01639_ ) );
NAND3_X1 _09224_ ( .A1(_01636_ ), .A2(_01639_ ), .A3(_01535_ ), .ZN(_01640_ ) );
MUX2_X1 _09225_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01641_ ) );
MUX2_X1 _09226_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01642_ ) );
MUX2_X1 _09227_ ( .A(_01641_ ), .B(_01642_ ), .S(_01526_ ), .Z(_01643_ ) );
OAI211_X1 _09228_ ( .A(_01402_ ), .B(_01640_ ), .C1(_01643_ ), .C2(_01407_ ), .ZN(_01644_ ) );
OR2_X1 _09229_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01645_ ) );
OAI211_X1 _09230_ ( .A(_01645_ ), .B(_01424_ ), .C1(_01638_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01646_ ) );
INV_X1 _09231_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01647_ ) );
NAND2_X1 _09232_ ( .A1(_01647_ ), .A2(fanout_net_12 ), .ZN(_01648_ ) );
OAI211_X1 _09233_ ( .A(_01648_ ), .B(fanout_net_18 ), .C1(fanout_net_12 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01649_ ) );
NAND3_X1 _09234_ ( .A1(_01646_ ), .A2(_01649_ ), .A3(fanout_net_21 ), .ZN(_01650_ ) );
MUX2_X1 _09235_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01651_ ) );
MUX2_X1 _09236_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01652_ ) );
MUX2_X1 _09237_ ( .A(_01651_ ), .B(_01652_ ), .S(fanout_net_18 ), .Z(_01653_ ) );
OAI211_X1 _09238_ ( .A(fanout_net_22 ), .B(_01650_ ), .C1(_01653_ ), .C2(fanout_net_21 ), .ZN(_01654_ ) );
NAND2_X1 _09239_ ( .A1(_01644_ ), .A2(_01654_ ), .ZN(_01655_ ) );
OAI21_X1 _09240_ ( .A(_01655_ ), .B1(_01605_ ), .B2(_01398_ ), .ZN(_01656_ ) );
AND2_X2 _09241_ ( .A1(_01634_ ), .A2(_01656_ ), .ZN(_01657_ ) );
XNOR2_X1 _09242_ ( .A(_01657_ ), .B(\ID_EX_imm [5] ), .ZN(_01658_ ) );
NOR2_X2 _09243_ ( .A1(_01632_ ), .A2(_01658_ ), .ZN(_01659_ ) );
INV_X1 _09244_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01660_ ) );
AND3_X1 _09245_ ( .A1(_01634_ ), .A2(_01656_ ), .A3(_01660_ ), .ZN(_01661_ ) );
NOR2_X2 _09246_ ( .A1(_01659_ ), .A2(_01661_ ), .ZN(_01662_ ) );
NAND2_X1 _09247_ ( .A1(_01633_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_01663_ ) );
OR2_X1 _09248_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01664_ ) );
OAI211_X1 _09249_ ( .A(_01664_ ), .B(_01425_ ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01665_ ) );
OR2_X1 _09250_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01666_ ) );
OAI211_X1 _09251_ ( .A(_01666_ ), .B(fanout_net_18 ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01667_ ) );
NAND3_X1 _09252_ ( .A1(_01665_ ), .A2(_01667_ ), .A3(_01407_ ), .ZN(_01668_ ) );
MUX2_X1 _09253_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01669_ ) );
MUX2_X1 _09254_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01670_ ) );
MUX2_X1 _09255_ ( .A(_01669_ ), .B(_01670_ ), .S(_01609_ ), .Z(_01671_ ) );
OAI211_X1 _09256_ ( .A(_01403_ ), .B(_01668_ ), .C1(_01671_ ), .C2(_01407_ ), .ZN(_01672_ ) );
OR2_X1 _09257_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01673_ ) );
OAI211_X1 _09258_ ( .A(_01673_ ), .B(fanout_net_18 ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01674_ ) );
OR2_X1 _09259_ ( .A1(fanout_net_12 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01675_ ) );
OAI211_X1 _09260_ ( .A(_01675_ ), .B(_01609_ ), .C1(_01610_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01676_ ) );
NAND3_X1 _09261_ ( .A1(_01674_ ), .A2(_01676_ ), .A3(fanout_net_21 ), .ZN(_01677_ ) );
MUX2_X1 _09262_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01678_ ) );
MUX2_X1 _09263_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01679_ ) );
MUX2_X1 _09264_ ( .A(_01678_ ), .B(_01679_ ), .S(fanout_net_18 ), .Z(_01680_ ) );
OAI211_X1 _09265_ ( .A(fanout_net_22 ), .B(_01677_ ), .C1(_01680_ ), .C2(fanout_net_21 ), .ZN(_01681_ ) );
NAND2_X1 _09266_ ( .A1(_01672_ ), .A2(_01681_ ), .ZN(_01682_ ) );
OAI21_X1 _09267_ ( .A(_01682_ ), .B1(_01386_ ), .B2(_01398_ ), .ZN(_01683_ ) );
AND2_X2 _09268_ ( .A1(_01663_ ), .A2(_01683_ ), .ZN(_01684_ ) );
XNOR2_X1 _09269_ ( .A(_01684_ ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_01685_ ) );
INV_X1 _09270_ ( .A(_01685_ ), .ZN(_01686_ ) );
OR3_X4 _09271_ ( .A1(_01386_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01606_ ), .ZN(_01687_ ) );
OR2_X1 _09272_ ( .A1(fanout_net_12 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01688_ ) );
OAI211_X1 _09273_ ( .A(_01688_ ), .B(_01425_ ), .C1(_01414_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01689_ ) );
OR2_X1 _09274_ ( .A1(fanout_net_12 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01690_ ) );
OAI211_X1 _09275_ ( .A(_01690_ ), .B(fanout_net_18 ), .C1(_01414_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01691_ ) );
NAND3_X1 _09276_ ( .A1(_01689_ ), .A2(_01691_ ), .A3(_01407_ ), .ZN(_01692_ ) );
MUX2_X1 _09277_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01693_ ) );
MUX2_X1 _09278_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01694_ ) );
MUX2_X1 _09279_ ( .A(_01693_ ), .B(_01694_ ), .S(_01425_ ), .Z(_01695_ ) );
OAI211_X1 _09280_ ( .A(_01403_ ), .B(_01692_ ), .C1(_01695_ ), .C2(_01408_ ), .ZN(_01696_ ) );
OR2_X1 _09281_ ( .A1(fanout_net_12 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01697_ ) );
OAI211_X1 _09282_ ( .A(_01697_ ), .B(fanout_net_19 ), .C1(_01414_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01698_ ) );
OR2_X1 _09283_ ( .A1(fanout_net_12 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01699_ ) );
OAI211_X1 _09284_ ( .A(_01699_ ), .B(_01425_ ), .C1(_01610_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01700_ ) );
NAND3_X1 _09285_ ( .A1(_01698_ ), .A2(_01700_ ), .A3(fanout_net_21 ), .ZN(_01701_ ) );
MUX2_X1 _09286_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01702_ ) );
MUX2_X1 _09287_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_12 ), .Z(_01703_ ) );
MUX2_X1 _09288_ ( .A(_01702_ ), .B(_01703_ ), .S(fanout_net_19 ), .Z(_01704_ ) );
OAI211_X1 _09289_ ( .A(fanout_net_22 ), .B(_01701_ ), .C1(_01704_ ), .C2(fanout_net_21 ), .ZN(_01705_ ) );
OAI211_X1 _09290_ ( .A(_01696_ ), .B(_01705_ ), .C1(_01386_ ), .C2(_01398_ ), .ZN(_01706_ ) );
NAND2_X4 _09291_ ( .A1(_01687_ ), .A2(_01706_ ), .ZN(_01707_ ) );
INV_X1 _09292_ ( .A(\ID_EX_imm [6] ), .ZN(_01708_ ) );
XNOR2_X1 _09293_ ( .A(_01707_ ), .B(_01708_ ), .ZN(_01709_ ) );
INV_X1 _09294_ ( .A(_01709_ ), .ZN(_01710_ ) );
NOR3_X4 _09295_ ( .A1(_01662_ ), .A2(_01686_ ), .A3(_01710_ ), .ZN(_01711_ ) );
AND2_X1 _09296_ ( .A1(_01707_ ), .A2(\ID_EX_imm [6] ), .ZN(_01712_ ) );
AND2_X1 _09297_ ( .A1(_01685_ ), .A2(_01712_ ), .ZN(_01713_ ) );
INV_X1 _09298_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_01714_ ) );
AOI21_X1 _09299_ ( .A(_01713_ ), .B1(_01714_ ), .B2(_01684_ ), .ZN(_01715_ ) );
INV_X1 _09300_ ( .A(_01715_ ), .ZN(_01716_ ) );
NOR2_X2 _09301_ ( .A1(_01711_ ), .A2(_01716_ ), .ZN(_01717_ ) );
OR3_X4 _09302_ ( .A1(_01605_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01606_ ), .ZN(_01718_ ) );
OR2_X1 _09303_ ( .A1(_01527_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01719_ ) );
OAI211_X1 _09304_ ( .A(_01719_ ), .B(fanout_net_19 ), .C1(fanout_net_13 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01720_ ) );
OR2_X1 _09305_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01721_ ) );
OAI211_X1 _09306_ ( .A(_01721_ ), .B(_01609_ ), .C1(_01413_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01722_ ) );
NAND3_X1 _09307_ ( .A1(_01720_ ), .A2(_01535_ ), .A3(_01722_ ), .ZN(_01723_ ) );
MUX2_X1 _09308_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01724_ ) );
MUX2_X1 _09309_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01725_ ) );
MUX2_X1 _09310_ ( .A(_01724_ ), .B(_01725_ ), .S(_01609_ ), .Z(_01726_ ) );
OAI211_X1 _09311_ ( .A(_01402_ ), .B(_01723_ ), .C1(_01726_ ), .C2(_01407_ ), .ZN(_01727_ ) );
OR2_X1 _09312_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01728_ ) );
OAI211_X1 _09313_ ( .A(_01728_ ), .B(fanout_net_19 ), .C1(_01610_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01729_ ) );
OR2_X1 _09314_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01730_ ) );
OAI211_X1 _09315_ ( .A(_01730_ ), .B(_01609_ ), .C1(_01413_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01731_ ) );
NAND3_X1 _09316_ ( .A1(_01729_ ), .A2(_01731_ ), .A3(fanout_net_21 ), .ZN(_01732_ ) );
MUX2_X1 _09317_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01733_ ) );
MUX2_X1 _09318_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01734_ ) );
MUX2_X1 _09319_ ( .A(_01733_ ), .B(_01734_ ), .S(fanout_net_19 ), .Z(_01735_ ) );
OAI211_X1 _09320_ ( .A(fanout_net_22 ), .B(_01732_ ), .C1(_01735_ ), .C2(fanout_net_21 ), .ZN(_01736_ ) );
OAI211_X1 _09321_ ( .A(_01727_ ), .B(_01736_ ), .C1(_01386_ ), .C2(_01398_ ), .ZN(_01737_ ) );
NAND2_X4 _09322_ ( .A1(_01718_ ), .A2(_01737_ ), .ZN(_01738_ ) );
XOR2_X1 _09323_ ( .A(_01738_ ), .B(\ID_EX_imm [14] ), .Z(_01739_ ) );
OR3_X4 _09324_ ( .A1(_01605_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01606_ ), .ZN(_01740_ ) );
OR2_X1 _09325_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01741_ ) );
OAI211_X1 _09326_ ( .A(_01741_ ), .B(_01609_ ), .C1(_01413_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01742_ ) );
OR2_X1 _09327_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01743_ ) );
OAI211_X1 _09328_ ( .A(_01743_ ), .B(fanout_net_19 ), .C1(_01413_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01744_ ) );
NAND3_X1 _09329_ ( .A1(_01742_ ), .A2(_01744_ ), .A3(fanout_net_21 ), .ZN(_01745_ ) );
MUX2_X1 _09330_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01746_ ) );
MUX2_X1 _09331_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01747_ ) );
MUX2_X1 _09332_ ( .A(_01746_ ), .B(_01747_ ), .S(_01424_ ), .Z(_01748_ ) );
OAI211_X1 _09333_ ( .A(_01402_ ), .B(_01745_ ), .C1(_01748_ ), .C2(fanout_net_21 ), .ZN(_01749_ ) );
NOR2_X1 _09334_ ( .A1(_01638_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01750_ ) );
OAI21_X1 _09335_ ( .A(fanout_net_19 ), .B1(fanout_net_13 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01751_ ) );
NOR2_X1 _09336_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01752_ ) );
OAI21_X1 _09337_ ( .A(_01424_ ), .B1(_01638_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01753_ ) );
OAI221_X1 _09338_ ( .A(_01535_ ), .B1(_01750_ ), .B2(_01751_ ), .C1(_01752_ ), .C2(_01753_ ), .ZN(_01754_ ) );
MUX2_X1 _09339_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01755_ ) );
MUX2_X1 _09340_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01756_ ) );
MUX2_X1 _09341_ ( .A(_01755_ ), .B(_01756_ ), .S(fanout_net_19 ), .Z(_01757_ ) );
OAI211_X1 _09342_ ( .A(fanout_net_22 ), .B(_01754_ ), .C1(_01757_ ), .C2(_01407_ ), .ZN(_01758_ ) );
OAI211_X1 _09343_ ( .A(_01749_ ), .B(_01758_ ), .C1(_01605_ ), .C2(_01606_ ), .ZN(_01759_ ) );
NAND2_X4 _09344_ ( .A1(_01740_ ), .A2(_01759_ ), .ZN(_01760_ ) );
INV_X1 _09345_ ( .A(\ID_EX_imm [15] ), .ZN(_01761_ ) );
XNOR2_X1 _09346_ ( .A(_01760_ ), .B(_01761_ ), .ZN(_01762_ ) );
AND2_X1 _09347_ ( .A1(_01739_ ), .A2(_01762_ ), .ZN(_01763_ ) );
OR3_X1 _09348_ ( .A1(_01385_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01397_ ), .ZN(_01764_ ) );
INV_X1 _09349_ ( .A(\ID_EX_imm [13] ), .ZN(_01765_ ) );
OR2_X1 _09350_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01766_ ) );
OAI211_X1 _09351_ ( .A(_01766_ ), .B(_01424_ ), .C1(_01638_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01767_ ) );
OR2_X1 _09352_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01768_ ) );
OAI211_X1 _09353_ ( .A(_01768_ ), .B(fanout_net_19 ), .C1(_01638_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01769_ ) );
NAND3_X1 _09354_ ( .A1(_01767_ ), .A2(_01769_ ), .A3(_01535_ ), .ZN(_01770_ ) );
MUX2_X1 _09355_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01771_ ) );
MUX2_X1 _09356_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01772_ ) );
MUX2_X1 _09357_ ( .A(_01771_ ), .B(_01772_ ), .S(_01526_ ), .Z(_01773_ ) );
OAI211_X1 _09358_ ( .A(_01402_ ), .B(_01770_ ), .C1(_01773_ ), .C2(_01535_ ), .ZN(_01774_ ) );
OR2_X1 _09359_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01775_ ) );
OAI211_X1 _09360_ ( .A(_01775_ ), .B(fanout_net_19 ), .C1(_01638_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01776_ ) );
OR2_X1 _09361_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01777_ ) );
OAI211_X1 _09362_ ( .A(_01777_ ), .B(_01424_ ), .C1(_01638_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01778_ ) );
NAND3_X1 _09363_ ( .A1(_01776_ ), .A2(_01778_ ), .A3(fanout_net_21 ), .ZN(_01779_ ) );
MUX2_X1 _09364_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01780_ ) );
MUX2_X1 _09365_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01781_ ) );
MUX2_X1 _09366_ ( .A(_01780_ ), .B(_01781_ ), .S(fanout_net_19 ), .Z(_01782_ ) );
OAI211_X1 _09367_ ( .A(fanout_net_22 ), .B(_01779_ ), .C1(_01782_ ), .C2(fanout_net_21 ), .ZN(_01783_ ) );
OAI211_X2 _09368_ ( .A(_01774_ ), .B(_01783_ ), .C1(_01605_ ), .C2(_01606_ ), .ZN(_01784_ ) );
AND3_X1 _09369_ ( .A1(_01764_ ), .A2(_01765_ ), .A3(_01784_ ), .ZN(_01785_ ) );
AOI21_X1 _09370_ ( .A(_01765_ ), .B1(_01764_ ), .B2(_01784_ ), .ZN(_01786_ ) );
NOR2_X1 _09371_ ( .A1(_01785_ ), .A2(_01786_ ), .ZN(_01787_ ) );
OR3_X1 _09372_ ( .A1(_01385_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01397_ ), .ZN(_01788_ ) );
OR2_X1 _09373_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01789_ ) );
OAI211_X1 _09374_ ( .A(_01789_ ), .B(_01424_ ), .C1(_01638_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01790_ ) );
OR2_X1 _09375_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01791_ ) );
OAI211_X1 _09376_ ( .A(_01791_ ), .B(fanout_net_19 ), .C1(_01527_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01792_ ) );
NAND3_X1 _09377_ ( .A1(_01790_ ), .A2(_01792_ ), .A3(_01535_ ), .ZN(_01793_ ) );
MUX2_X1 _09378_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01794_ ) );
MUX2_X1 _09379_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_13 ), .Z(_01795_ ) );
MUX2_X1 _09380_ ( .A(_01794_ ), .B(_01795_ ), .S(_01526_ ), .Z(_01796_ ) );
OAI211_X1 _09381_ ( .A(_01402_ ), .B(_01793_ ), .C1(_01796_ ), .C2(_01535_ ), .ZN(_01797_ ) );
OR2_X1 _09382_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01798_ ) );
OAI211_X1 _09383_ ( .A(_01798_ ), .B(fanout_net_19 ), .C1(_01638_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01799_ ) );
OR2_X1 _09384_ ( .A1(fanout_net_13 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01800_ ) );
OAI211_X1 _09385_ ( .A(_01800_ ), .B(_01526_ ), .C1(_01527_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01801_ ) );
NAND3_X1 _09386_ ( .A1(_01799_ ), .A2(_01801_ ), .A3(fanout_net_21 ), .ZN(_01802_ ) );
MUX2_X1 _09387_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01803_ ) );
MUX2_X1 _09388_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01804_ ) );
MUX2_X1 _09389_ ( .A(_01803_ ), .B(_01804_ ), .S(fanout_net_19 ), .Z(_01805_ ) );
OAI211_X1 _09390_ ( .A(fanout_net_22 ), .B(_01802_ ), .C1(_01805_ ), .C2(fanout_net_21 ), .ZN(_01806_ ) );
OAI211_X1 _09391_ ( .A(_01797_ ), .B(_01806_ ), .C1(_01605_ ), .C2(_01606_ ), .ZN(_01807_ ) );
NAND2_X4 _09392_ ( .A1(_01788_ ), .A2(_01807_ ), .ZN(_01808_ ) );
INV_X1 _09393_ ( .A(\ID_EX_imm [12] ), .ZN(_01809_ ) );
XNOR2_X1 _09394_ ( .A(_01808_ ), .B(_01809_ ), .ZN(_01810_ ) );
NAND3_X1 _09395_ ( .A1(_01763_ ), .A2(_01787_ ), .A3(_01810_ ), .ZN(_01811_ ) );
OR3_X1 _09396_ ( .A1(_01605_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01606_ ), .ZN(_01812_ ) );
OR2_X1 _09397_ ( .A1(fanout_net_14 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01813_ ) );
OAI211_X1 _09398_ ( .A(_01813_ ), .B(_01609_ ), .C1(_01413_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01814_ ) );
OR2_X1 _09399_ ( .A1(fanout_net_14 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01815_ ) );
OAI211_X1 _09400_ ( .A(_01815_ ), .B(fanout_net_19 ), .C1(_01413_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01816_ ) );
NAND3_X1 _09401_ ( .A1(_01814_ ), .A2(_01816_ ), .A3(fanout_net_21 ), .ZN(_01817_ ) );
MUX2_X1 _09402_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01818_ ) );
MUX2_X1 _09403_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01819_ ) );
MUX2_X1 _09404_ ( .A(_01818_ ), .B(_01819_ ), .S(_01424_ ), .Z(_01820_ ) );
OAI211_X1 _09405_ ( .A(_01402_ ), .B(_01817_ ), .C1(_01820_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01821_ ) );
NOR2_X1 _09406_ ( .A1(_01413_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01822_ ) );
OAI21_X1 _09407_ ( .A(fanout_net_19 ), .B1(fanout_net_14 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01823_ ) );
NOR2_X1 _09408_ ( .A1(fanout_net_14 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01824_ ) );
OAI21_X1 _09409_ ( .A(_01424_ ), .B1(_01413_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01825_ ) );
OAI221_X1 _09410_ ( .A(_01535_ ), .B1(_01822_ ), .B2(_01823_ ), .C1(_01824_ ), .C2(_01825_ ), .ZN(_01826_ ) );
MUX2_X1 _09411_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01827_ ) );
MUX2_X1 _09412_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01828_ ) );
MUX2_X1 _09413_ ( .A(_01827_ ), .B(_01828_ ), .S(fanout_net_19 ), .Z(_01829_ ) );
OAI211_X1 _09414_ ( .A(fanout_net_22 ), .B(_01826_ ), .C1(_01829_ ), .C2(_01407_ ), .ZN(_01830_ ) );
OAI211_X1 _09415_ ( .A(_01821_ ), .B(_01830_ ), .C1(_01605_ ), .C2(_01606_ ), .ZN(_01831_ ) );
NAND2_X4 _09416_ ( .A1(_01812_ ), .A2(_01831_ ), .ZN(_01832_ ) );
XOR2_X1 _09417_ ( .A(_01832_ ), .B(\ID_EX_imm [8] ), .Z(_01833_ ) );
OR3_X1 _09418_ ( .A1(_01384_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01396_ ), .ZN(_01834_ ) );
OR2_X1 _09419_ ( .A1(fanout_net_14 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01835_ ) );
OAI211_X1 _09420_ ( .A(_01835_ ), .B(_01422_ ), .C1(_01504_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01836_ ) );
OR2_X1 _09421_ ( .A1(fanout_net_14 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01837_ ) );
OAI211_X1 _09422_ ( .A(_01837_ ), .B(fanout_net_19 ), .C1(_01504_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01838_ ) );
NAND3_X1 _09423_ ( .A1(_01836_ ), .A2(_01838_ ), .A3(_01405_ ), .ZN(_01839_ ) );
MUX2_X1 _09424_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01840_ ) );
MUX2_X1 _09425_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01841_ ) );
MUX2_X1 _09426_ ( .A(_01840_ ), .B(_01841_ ), .S(_01422_ ), .Z(_01842_ ) );
OAI211_X1 _09427_ ( .A(_01401_ ), .B(_01839_ ), .C1(_01842_ ), .C2(_01406_ ), .ZN(_01843_ ) );
OR2_X1 _09428_ ( .A1(fanout_net_14 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01844_ ) );
OAI211_X1 _09429_ ( .A(_01844_ ), .B(fanout_net_19 ), .C1(_01504_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01845_ ) );
OR2_X1 _09430_ ( .A1(fanout_net_14 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01846_ ) );
OAI211_X1 _09431_ ( .A(_01846_ ), .B(_01422_ ), .C1(_01504_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01847_ ) );
NAND3_X1 _09432_ ( .A1(_01845_ ), .A2(_01847_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01848_ ) );
MUX2_X1 _09433_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01849_ ) );
MUX2_X1 _09434_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01850_ ) );
MUX2_X1 _09435_ ( .A(_01849_ ), .B(_01850_ ), .S(fanout_net_19 ), .Z(_01851_ ) );
OAI211_X1 _09436_ ( .A(fanout_net_22 ), .B(_01848_ ), .C1(_01851_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01852_ ) );
OAI211_X1 _09437_ ( .A(_01843_ ), .B(_01852_ ), .C1(_01384_ ), .C2(_01396_ ), .ZN(_01853_ ) );
NAND2_X1 _09438_ ( .A1(_01834_ ), .A2(_01853_ ), .ZN(_01854_ ) );
AND2_X1 _09439_ ( .A1(_01854_ ), .A2(\ID_EX_imm [9] ), .ZN(_01855_ ) );
INV_X1 _09440_ ( .A(_01855_ ), .ZN(_01856_ ) );
INV_X1 _09441_ ( .A(\ID_EX_imm [9] ), .ZN(_01857_ ) );
AND3_X1 _09442_ ( .A1(_01834_ ), .A2(_01857_ ), .A3(_01853_ ), .ZN(_01858_ ) );
INV_X1 _09443_ ( .A(_01858_ ), .ZN(_01859_ ) );
AND3_X1 _09444_ ( .A1(_01833_ ), .A2(_01856_ ), .A3(_01859_ ), .ZN(_01860_ ) );
OR3_X1 _09445_ ( .A1(_01384_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(_01396_ ), .ZN(_01861_ ) );
INV_X1 _09446_ ( .A(\ID_EX_imm [11] ), .ZN(_01862_ ) );
OR2_X1 _09447_ ( .A1(_01411_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01863_ ) );
OAI211_X1 _09448_ ( .A(_01863_ ), .B(_01423_ ), .C1(fanout_net_14 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01864_ ) );
OR2_X1 _09449_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01865_ ) );
OAI211_X1 _09450_ ( .A(_01865_ ), .B(fanout_net_19 ), .C1(_01412_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01866_ ) );
NAND3_X1 _09451_ ( .A1(_01864_ ), .A2(_01406_ ), .A3(_01866_ ), .ZN(_01867_ ) );
MUX2_X1 _09452_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01868_ ) );
MUX2_X1 _09453_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01869_ ) );
MUX2_X1 _09454_ ( .A(_01868_ ), .B(_01869_ ), .S(_01423_ ), .Z(_01870_ ) );
OAI211_X1 _09455_ ( .A(_01402_ ), .B(_01867_ ), .C1(_01870_ ), .C2(_01406_ ), .ZN(_01871_ ) );
OR2_X1 _09456_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01872_ ) );
OAI211_X1 _09457_ ( .A(_01872_ ), .B(fanout_net_19 ), .C1(_01412_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01873_ ) );
OR2_X1 _09458_ ( .A1(fanout_net_14 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01874_ ) );
OAI211_X1 _09459_ ( .A(_01874_ ), .B(_01423_ ), .C1(_01504_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01875_ ) );
NAND3_X1 _09460_ ( .A1(_01873_ ), .A2(_01875_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01876_ ) );
MUX2_X1 _09461_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01877_ ) );
MUX2_X1 _09462_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01878_ ) );
MUX2_X1 _09463_ ( .A(_01877_ ), .B(_01878_ ), .S(fanout_net_19 ), .Z(_01879_ ) );
OAI211_X1 _09464_ ( .A(fanout_net_22 ), .B(_01876_ ), .C1(_01879_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01880_ ) );
OAI211_X1 _09465_ ( .A(_01871_ ), .B(_01880_ ), .C1(_01385_ ), .C2(_01397_ ), .ZN(_01881_ ) );
AND3_X1 _09466_ ( .A1(_01861_ ), .A2(_01862_ ), .A3(_01881_ ), .ZN(_01882_ ) );
AOI21_X1 _09467_ ( .A(_01862_ ), .B1(_01861_ ), .B2(_01881_ ), .ZN(_01883_ ) );
NOR2_X1 _09468_ ( .A1(_01882_ ), .A2(_01883_ ), .ZN(_01884_ ) );
OR3_X1 _09469_ ( .A1(_01384_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01396_ ), .ZN(_01885_ ) );
OR2_X1 _09470_ ( .A1(fanout_net_14 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01886_ ) );
OAI211_X1 _09471_ ( .A(_01886_ ), .B(_01423_ ), .C1(_01412_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01887_ ) );
OR2_X1 _09472_ ( .A1(fanout_net_14 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01888_ ) );
OAI211_X1 _09473_ ( .A(_01888_ ), .B(fanout_net_19 ), .C1(_01504_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01889_ ) );
NAND3_X1 _09474_ ( .A1(_01887_ ), .A2(_01889_ ), .A3(_01406_ ), .ZN(_01890_ ) );
MUX2_X1 _09475_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01891_ ) );
MUX2_X1 _09476_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_14 ), .Z(_01892_ ) );
MUX2_X1 _09477_ ( .A(_01891_ ), .B(_01892_ ), .S(_01423_ ), .Z(_01893_ ) );
OAI211_X1 _09478_ ( .A(_01401_ ), .B(_01890_ ), .C1(_01893_ ), .C2(_01406_ ), .ZN(_01894_ ) );
OR2_X1 _09479_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01895_ ) );
OAI211_X1 _09480_ ( .A(_01895_ ), .B(fanout_net_19 ), .C1(_01412_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01896_ ) );
OR2_X1 _09481_ ( .A1(fanout_net_15 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01897_ ) );
OAI211_X1 _09482_ ( .A(_01897_ ), .B(_01423_ ), .C1(_01504_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01898_ ) );
NAND3_X1 _09483_ ( .A1(_01896_ ), .A2(_01898_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01899_ ) );
MUX2_X1 _09484_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01900_ ) );
MUX2_X1 _09485_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01901_ ) );
MUX2_X1 _09486_ ( .A(_01900_ ), .B(_01901_ ), .S(fanout_net_19 ), .Z(_01902_ ) );
OAI211_X1 _09487_ ( .A(fanout_net_22 ), .B(_01899_ ), .C1(_01902_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01903_ ) );
OAI211_X1 _09488_ ( .A(_01894_ ), .B(_01903_ ), .C1(_01385_ ), .C2(_01397_ ), .ZN(_01904_ ) );
NAND2_X1 _09489_ ( .A1(_01885_ ), .A2(_01904_ ), .ZN(_01905_ ) );
XOR2_X1 _09490_ ( .A(_01905_ ), .B(\ID_EX_imm [10] ), .Z(_01906_ ) );
NAND3_X1 _09491_ ( .A1(_01860_ ), .A2(_01884_ ), .A3(_01906_ ), .ZN(_01907_ ) );
NOR3_X2 _09492_ ( .A1(_01717_ ), .A2(_01811_ ), .A3(_01907_ ), .ZN(_01908_ ) );
OAI211_X1 _09493_ ( .A(\ID_EX_imm [14] ), .B(_01738_ ), .C1(_01760_ ), .C2(\ID_EX_imm [15] ), .ZN(_01909_ ) );
AND2_X1 _09494_ ( .A1(_01808_ ), .A2(\ID_EX_imm [12] ), .ZN(_01910_ ) );
AOI21_X1 _09495_ ( .A(_01786_ ), .B1(_01787_ ), .B2(_01910_ ), .ZN(_01911_ ) );
INV_X1 _09496_ ( .A(_01911_ ), .ZN(_01912_ ) );
AOI22_X1 _09497_ ( .A1(_01763_ ), .A2(_01912_ ), .B1(\ID_EX_imm [15] ), .B2(_01760_ ), .ZN(_01913_ ) );
NAND2_X1 _09498_ ( .A1(_01832_ ), .A2(\ID_EX_imm [8] ), .ZN(_01914_ ) );
NOR3_X1 _09499_ ( .A1(_01855_ ), .A2(_01858_ ), .A3(_01914_ ), .ZN(_01915_ ) );
OAI211_X1 _09500_ ( .A(_01884_ ), .B(_01906_ ), .C1(_01915_ ), .C2(_01855_ ), .ZN(_01916_ ) );
AND2_X1 _09501_ ( .A1(_01905_ ), .A2(\ID_EX_imm [10] ), .ZN(_01917_ ) );
AOI21_X1 _09502_ ( .A(_01883_ ), .B1(_01884_ ), .B2(_01917_ ), .ZN(_01918_ ) );
AND2_X1 _09503_ ( .A1(_01916_ ), .A2(_01918_ ), .ZN(_01919_ ) );
OAI211_X1 _09504_ ( .A(_01909_ ), .B(_01913_ ), .C1(_01919_ ), .C2(_01811_ ), .ZN(_01920_ ) );
NOR2_X1 _09505_ ( .A1(_01908_ ), .A2(_01920_ ), .ZN(_01921_ ) );
BUF_X2 _09506_ ( .A(_01398_ ), .Z(_01922_ ) );
OR3_X1 _09507_ ( .A1(_01387_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01922_ ), .ZN(_01923_ ) );
OR2_X1 _09508_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01924_ ) );
BUF_X4 _09509_ ( .A(_01414_ ), .Z(_01925_ ) );
OAI211_X1 _09510_ ( .A(_01924_ ), .B(_01426_ ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01926_ ) );
OR2_X1 _09511_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01927_ ) );
OAI211_X1 _09512_ ( .A(_01927_ ), .B(fanout_net_19 ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01928_ ) );
NAND3_X1 _09513_ ( .A1(_01926_ ), .A2(_01928_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01929_ ) );
MUX2_X1 _09514_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01930_ ) );
MUX2_X1 _09515_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01931_ ) );
BUF_X4 _09516_ ( .A(_01425_ ), .Z(_01932_ ) );
MUX2_X1 _09517_ ( .A(_01930_ ), .B(_01931_ ), .S(_01932_ ), .Z(_01933_ ) );
OAI211_X1 _09518_ ( .A(_01403_ ), .B(_01929_ ), .C1(_01933_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01934_ ) );
NOR2_X1 _09519_ ( .A1(_01415_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01935_ ) );
OAI21_X1 _09520_ ( .A(fanout_net_19 ), .B1(fanout_net_15 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01936_ ) );
NOR2_X1 _09521_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01937_ ) );
OAI21_X1 _09522_ ( .A(_01932_ ), .B1(_01415_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01938_ ) );
OAI221_X1 _09523_ ( .A(_01408_ ), .B1(_01935_ ), .B2(_01936_ ), .C1(_01937_ ), .C2(_01938_ ), .ZN(_01939_ ) );
MUX2_X1 _09524_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01940_ ) );
MUX2_X1 _09525_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01941_ ) );
MUX2_X1 _09526_ ( .A(_01940_ ), .B(_01941_ ), .S(fanout_net_19 ), .Z(_01942_ ) );
OAI211_X1 _09527_ ( .A(fanout_net_22 ), .B(_01939_ ), .C1(_01942_ ), .C2(_01409_ ), .ZN(_01943_ ) );
OAI211_X1 _09528_ ( .A(_01934_ ), .B(_01943_ ), .C1(_01387_ ), .C2(_01922_ ), .ZN(_01944_ ) );
NAND2_X2 _09529_ ( .A1(_01923_ ), .A2(_01944_ ), .ZN(_01945_ ) );
INV_X1 _09530_ ( .A(\ID_EX_imm [17] ), .ZN(_01946_ ) );
XNOR2_X1 _09531_ ( .A(_01945_ ), .B(_01946_ ), .ZN(_01947_ ) );
INV_X1 _09532_ ( .A(_01947_ ), .ZN(_01948_ ) );
OR3_X1 _09533_ ( .A1(_01386_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01922_ ), .ZN(_01949_ ) );
OR2_X1 _09534_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01950_ ) );
OAI211_X1 _09535_ ( .A(_01950_ ), .B(_01932_ ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01951_ ) );
OR2_X1 _09536_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01952_ ) );
OAI211_X1 _09537_ ( .A(_01952_ ), .B(fanout_net_19 ), .C1(_01415_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01953_ ) );
NAND3_X1 _09538_ ( .A1(_01951_ ), .A2(_01953_ ), .A3(_01408_ ), .ZN(_01954_ ) );
MUX2_X1 _09539_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01955_ ) );
MUX2_X1 _09540_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01956_ ) );
MUX2_X1 _09541_ ( .A(_01955_ ), .B(_01956_ ), .S(_01932_ ), .Z(_01957_ ) );
OAI211_X1 _09542_ ( .A(fanout_net_22 ), .B(_01954_ ), .C1(_01957_ ), .C2(_01409_ ), .ZN(_01958_ ) );
OR2_X1 _09543_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01959_ ) );
OAI211_X1 _09544_ ( .A(_01959_ ), .B(_01932_ ), .C1(_01415_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01960_ ) );
OR2_X1 _09545_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01961_ ) );
OAI211_X1 _09546_ ( .A(_01961_ ), .B(fanout_net_20 ), .C1(_01415_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01962_ ) );
NAND3_X1 _09547_ ( .A1(_01960_ ), .A2(_01962_ ), .A3(_01408_ ), .ZN(_01963_ ) );
MUX2_X1 _09548_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01964_ ) );
MUX2_X1 _09549_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01965_ ) );
MUX2_X1 _09550_ ( .A(_01964_ ), .B(_01965_ ), .S(_01932_ ), .Z(_01966_ ) );
OAI211_X1 _09551_ ( .A(_01403_ ), .B(_01963_ ), .C1(_01966_ ), .C2(_01409_ ), .ZN(_01967_ ) );
OAI211_X1 _09552_ ( .A(_01958_ ), .B(_01967_ ), .C1(_01387_ ), .C2(_01922_ ), .ZN(_01968_ ) );
NAND2_X2 _09553_ ( .A1(_01949_ ), .A2(_01968_ ), .ZN(_01969_ ) );
INV_X1 _09554_ ( .A(\ID_EX_imm [16] ), .ZN(_01970_ ) );
XNOR2_X1 _09555_ ( .A(_01969_ ), .B(_01970_ ), .ZN(_01971_ ) );
INV_X1 _09556_ ( .A(_01971_ ), .ZN(_01972_ ) );
NOR3_X2 _09557_ ( .A1(_01921_ ), .A2(_01948_ ), .A3(_01972_ ), .ZN(_01973_ ) );
OR3_X1 _09558_ ( .A1(_01386_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01398_ ), .ZN(_01974_ ) );
INV_X1 _09559_ ( .A(\ID_EX_imm [19] ), .ZN(_01975_ ) );
OR2_X1 _09560_ ( .A1(_01414_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01976_ ) );
OAI211_X1 _09561_ ( .A(_01976_ ), .B(fanout_net_20 ), .C1(fanout_net_15 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01977_ ) );
OR2_X1 _09562_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01978_ ) );
OAI211_X1 _09563_ ( .A(_01978_ ), .B(_01425_ ), .C1(_01414_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01979_ ) );
NAND3_X1 _09564_ ( .A1(_01977_ ), .A2(_01408_ ), .A3(_01979_ ), .ZN(_01980_ ) );
MUX2_X1 _09565_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01981_ ) );
MUX2_X1 _09566_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01982_ ) );
MUX2_X1 _09567_ ( .A(_01981_ ), .B(_01982_ ), .S(_01425_ ), .Z(_01983_ ) );
OAI211_X1 _09568_ ( .A(_01403_ ), .B(_01980_ ), .C1(_01983_ ), .C2(_01408_ ), .ZN(_01984_ ) );
OR2_X1 _09569_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01985_ ) );
OAI211_X1 _09570_ ( .A(_01985_ ), .B(fanout_net_20 ), .C1(_01414_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_01986_ ) );
OR2_X1 _09571_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01987_ ) );
OAI211_X1 _09572_ ( .A(_01987_ ), .B(_01425_ ), .C1(_01414_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01988_ ) );
NAND3_X1 _09573_ ( .A1(_01986_ ), .A2(_01988_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01989_ ) );
MUX2_X1 _09574_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01990_ ) );
MUX2_X1 _09575_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_15 ), .Z(_01991_ ) );
MUX2_X1 _09576_ ( .A(_01990_ ), .B(_01991_ ), .S(fanout_net_20 ), .Z(_01992_ ) );
OAI211_X1 _09577_ ( .A(fanout_net_22 ), .B(_01989_ ), .C1(_01992_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_01993_ ) );
OAI211_X1 _09578_ ( .A(_01984_ ), .B(_01993_ ), .C1(_01386_ ), .C2(_01398_ ), .ZN(_01994_ ) );
AND3_X1 _09579_ ( .A1(_01974_ ), .A2(_01975_ ), .A3(_01994_ ), .ZN(_01995_ ) );
AOI21_X1 _09580_ ( .A(_01975_ ), .B1(_01974_ ), .B2(_01994_ ), .ZN(_01996_ ) );
NOR2_X1 _09581_ ( .A1(_01995_ ), .A2(_01996_ ), .ZN(_01997_ ) );
OR3_X1 _09582_ ( .A1(_01386_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01398_ ), .ZN(_01998_ ) );
OR2_X1 _09583_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01999_ ) );
OAI211_X1 _09584_ ( .A(_01999_ ), .B(_01932_ ), .C1(_01415_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02000_ ) );
OR2_X1 _09585_ ( .A1(fanout_net_15 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02001_ ) );
OAI211_X1 _09586_ ( .A(_02001_ ), .B(fanout_net_20 ), .C1(_01415_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02002_ ) );
NAND3_X1 _09587_ ( .A1(_02000_ ), .A2(_02002_ ), .A3(_01408_ ), .ZN(_02003_ ) );
MUX2_X1 _09588_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02004_ ) );
MUX2_X1 _09589_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02005_ ) );
MUX2_X1 _09590_ ( .A(_02004_ ), .B(_02005_ ), .S(_01425_ ), .Z(_02006_ ) );
OAI211_X1 _09591_ ( .A(_01403_ ), .B(_02003_ ), .C1(_02006_ ), .C2(_01408_ ), .ZN(_02007_ ) );
OR2_X1 _09592_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02008_ ) );
OAI211_X1 _09593_ ( .A(_02008_ ), .B(fanout_net_20 ), .C1(_01415_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02009_ ) );
OR2_X1 _09594_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02010_ ) );
OAI211_X1 _09595_ ( .A(_02010_ ), .B(_01932_ ), .C1(_01415_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02011_ ) );
NAND3_X1 _09596_ ( .A1(_02009_ ), .A2(_02011_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02012_ ) );
MUX2_X1 _09597_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02013_ ) );
MUX2_X1 _09598_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02014_ ) );
MUX2_X1 _09599_ ( .A(_02013_ ), .B(_02014_ ), .S(fanout_net_20 ), .Z(_02015_ ) );
OAI211_X1 _09600_ ( .A(fanout_net_22 ), .B(_02012_ ), .C1(_02015_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02016_ ) );
OAI211_X1 _09601_ ( .A(_02007_ ), .B(_02016_ ), .C1(_01387_ ), .C2(_01922_ ), .ZN(_02017_ ) );
NAND2_X1 _09602_ ( .A1(_01998_ ), .A2(_02017_ ), .ZN(_02018_ ) );
INV_X1 _09603_ ( .A(\ID_EX_imm [18] ), .ZN(_02019_ ) );
XNOR2_X1 _09604_ ( .A(_02018_ ), .B(_02019_ ), .ZN(_02020_ ) );
NAND3_X1 _09605_ ( .A1(_01973_ ), .A2(_01997_ ), .A3(_02020_ ), .ZN(_02021_ ) );
OR3_X1 _09606_ ( .A1(_01387_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01922_ ), .ZN(_02022_ ) );
OR2_X1 _09607_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02023_ ) );
OAI211_X1 _09608_ ( .A(_02023_ ), .B(_01426_ ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02024_ ) );
OR2_X1 _09609_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02025_ ) );
OAI211_X1 _09610_ ( .A(_02025_ ), .B(fanout_net_20 ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02026_ ) );
NAND3_X1 _09611_ ( .A1(_02024_ ), .A2(_02026_ ), .A3(_01408_ ), .ZN(_02027_ ) );
MUX2_X1 _09612_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02028_ ) );
MUX2_X1 _09613_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02029_ ) );
MUX2_X1 _09614_ ( .A(_02028_ ), .B(_02029_ ), .S(_01932_ ), .Z(_02030_ ) );
OAI211_X1 _09615_ ( .A(_01403_ ), .B(_02027_ ), .C1(_02030_ ), .C2(_01409_ ), .ZN(_02031_ ) );
OR2_X1 _09616_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02032_ ) );
OAI211_X1 _09617_ ( .A(_02032_ ), .B(fanout_net_20 ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02033_ ) );
OR2_X1 _09618_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02034_ ) );
OAI211_X1 _09619_ ( .A(_02034_ ), .B(_01426_ ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02035_ ) );
NAND3_X1 _09620_ ( .A1(_02033_ ), .A2(_02035_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02036_ ) );
MUX2_X1 _09621_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02037_ ) );
MUX2_X1 _09622_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02038_ ) );
MUX2_X1 _09623_ ( .A(_02037_ ), .B(_02038_ ), .S(fanout_net_20 ), .Z(_02039_ ) );
OAI211_X1 _09624_ ( .A(fanout_net_22 ), .B(_02036_ ), .C1(_02039_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02040_ ) );
OAI211_X1 _09625_ ( .A(_02031_ ), .B(_02040_ ), .C1(_01387_ ), .C2(_01922_ ), .ZN(_02041_ ) );
NAND2_X1 _09626_ ( .A1(_02022_ ), .A2(_02041_ ), .ZN(_02042_ ) );
XOR2_X1 _09627_ ( .A(_02042_ ), .B(\ID_EX_imm [23] ), .Z(_02043_ ) );
OR3_X1 _09628_ ( .A1(_01387_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01922_ ), .ZN(_02044_ ) );
OR2_X1 _09629_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02045_ ) );
OAI211_X1 _09630_ ( .A(_02045_ ), .B(_01426_ ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02046_ ) );
OR2_X1 _09631_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02047_ ) );
OAI211_X1 _09632_ ( .A(_02047_ ), .B(fanout_net_20 ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02048_ ) );
NAND3_X1 _09633_ ( .A1(_02046_ ), .A2(_02048_ ), .A3(_01409_ ), .ZN(_02049_ ) );
MUX2_X1 _09634_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02050_ ) );
MUX2_X1 _09635_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02051_ ) );
MUX2_X1 _09636_ ( .A(_02050_ ), .B(_02051_ ), .S(_01932_ ), .Z(_02052_ ) );
OAI211_X1 _09637_ ( .A(_01403_ ), .B(_02049_ ), .C1(_02052_ ), .C2(_01409_ ), .ZN(_02053_ ) );
OR2_X1 _09638_ ( .A1(_01414_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02054_ ) );
OAI211_X1 _09639_ ( .A(_02054_ ), .B(fanout_net_20 ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02055_ ) );
OR2_X1 _09640_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02056_ ) );
OAI211_X1 _09641_ ( .A(_02056_ ), .B(_01426_ ), .C1(_01925_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02057_ ) );
NAND3_X1 _09642_ ( .A1(_02055_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_02057_ ), .ZN(_02058_ ) );
MUX2_X1 _09643_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02059_ ) );
MUX2_X1 _09644_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02060_ ) );
MUX2_X1 _09645_ ( .A(_02059_ ), .B(_02060_ ), .S(fanout_net_20 ), .Z(_02061_ ) );
OAI211_X1 _09646_ ( .A(fanout_net_22 ), .B(_02058_ ), .C1(_02061_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02062_ ) );
OAI211_X1 _09647_ ( .A(_02053_ ), .B(_02062_ ), .C1(_01387_ ), .C2(_01922_ ), .ZN(_02063_ ) );
NAND2_X1 _09648_ ( .A1(_02044_ ), .A2(_02063_ ), .ZN(_02064_ ) );
INV_X1 _09649_ ( .A(\ID_EX_imm [22] ), .ZN(_02065_ ) );
XNOR2_X1 _09650_ ( .A(_02064_ ), .B(_02065_ ), .ZN(_02066_ ) );
AND2_X1 _09651_ ( .A1(_02043_ ), .A2(_02066_ ), .ZN(_02067_ ) );
OR3_X1 _09652_ ( .A1(_01388_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01399_ ), .ZN(_02068_ ) );
OR2_X1 _09653_ ( .A1(_01416_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02069_ ) );
OAI211_X1 _09654_ ( .A(_02069_ ), .B(_01427_ ), .C1(fanout_net_16 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02070_ ) );
OR2_X1 _09655_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02071_ ) );
OAI211_X1 _09656_ ( .A(_02071_ ), .B(fanout_net_20 ), .C1(_01477_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02072_ ) );
NAND3_X1 _09657_ ( .A1(_02070_ ), .A2(_01410_ ), .A3(_02072_ ), .ZN(_02073_ ) );
MUX2_X1 _09658_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02074_ ) );
MUX2_X1 _09659_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02075_ ) );
MUX2_X1 _09660_ ( .A(_02074_ ), .B(_02075_ ), .S(_01451_ ), .Z(_02076_ ) );
OAI211_X1 _09661_ ( .A(_01404_ ), .B(_02073_ ), .C1(_02076_ ), .C2(_01410_ ), .ZN(_02077_ ) );
OR2_X1 _09662_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02078_ ) );
OAI211_X1 _09663_ ( .A(_02078_ ), .B(fanout_net_20 ), .C1(_01477_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02079_ ) );
OR2_X1 _09664_ ( .A1(fanout_net_16 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02080_ ) );
OAI211_X1 _09665_ ( .A(_02080_ ), .B(_01451_ ), .C1(_01477_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02081_ ) );
NAND3_X1 _09666_ ( .A1(_02079_ ), .A2(_02081_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02082_ ) );
MUX2_X1 _09667_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02083_ ) );
MUX2_X1 _09668_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_16 ), .Z(_02084_ ) );
MUX2_X1 _09669_ ( .A(_02083_ ), .B(_02084_ ), .S(fanout_net_20 ), .Z(_02085_ ) );
OAI211_X1 _09670_ ( .A(fanout_net_22 ), .B(_02082_ ), .C1(_02085_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02086_ ) );
OAI211_X1 _09671_ ( .A(_02077_ ), .B(_02086_ ), .C1(_01388_ ), .C2(_01444_ ), .ZN(_02087_ ) );
NAND2_X1 _09672_ ( .A1(_02068_ ), .A2(_02087_ ), .ZN(_02088_ ) );
INV_X1 _09673_ ( .A(\ID_EX_imm [20] ), .ZN(_02089_ ) );
XNOR2_X1 _09674_ ( .A(_02088_ ), .B(_02089_ ), .ZN(_02090_ ) );
OR3_X1 _09675_ ( .A1(_01387_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_01922_ ), .ZN(_02091_ ) );
INV_X1 _09676_ ( .A(\ID_EX_imm [21] ), .ZN(_02092_ ) );
OR2_X1 _09677_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02093_ ) );
OAI211_X1 _09678_ ( .A(_02093_ ), .B(_01426_ ), .C1(_01416_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02094_ ) );
OR2_X1 _09679_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02095_ ) );
OAI211_X1 _09680_ ( .A(_02095_ ), .B(fanout_net_20 ), .C1(_01416_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02096_ ) );
NAND3_X1 _09681_ ( .A1(_02094_ ), .A2(_02096_ ), .A3(_01409_ ), .ZN(_02097_ ) );
MUX2_X1 _09682_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02098_ ) );
MUX2_X1 _09683_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02099_ ) );
MUX2_X1 _09684_ ( .A(_02098_ ), .B(_02099_ ), .S(_01426_ ), .Z(_02100_ ) );
OAI211_X1 _09685_ ( .A(_01404_ ), .B(_02097_ ), .C1(_02100_ ), .C2(_01409_ ), .ZN(_02101_ ) );
OR2_X1 _09686_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02102_ ) );
OAI211_X1 _09687_ ( .A(_02102_ ), .B(fanout_net_20 ), .C1(_01416_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02103_ ) );
OR2_X1 _09688_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02104_ ) );
OAI211_X1 _09689_ ( .A(_02104_ ), .B(_01426_ ), .C1(_01416_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02105_ ) );
NAND3_X1 _09690_ ( .A1(_02103_ ), .A2(_02105_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02106_ ) );
MUX2_X1 _09691_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02107_ ) );
MUX2_X1 _09692_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02108_ ) );
MUX2_X1 _09693_ ( .A(_02107_ ), .B(_02108_ ), .S(fanout_net_20 ), .Z(_02109_ ) );
OAI211_X1 _09694_ ( .A(fanout_net_22 ), .B(_02106_ ), .C1(_02109_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02110_ ) );
OAI211_X1 _09695_ ( .A(_02101_ ), .B(_02110_ ), .C1(_01388_ ), .C2(_01399_ ), .ZN(_02111_ ) );
AND3_X1 _09696_ ( .A1(_02091_ ), .A2(_02092_ ), .A3(_02111_ ), .ZN(_02112_ ) );
AOI21_X1 _09697_ ( .A(_02092_ ), .B1(_02091_ ), .B2(_02111_ ), .ZN(_02113_ ) );
NOR2_X1 _09698_ ( .A1(_02112_ ), .A2(_02113_ ), .ZN(_02114_ ) );
NAND3_X1 _09699_ ( .A1(_02067_ ), .A2(_02090_ ), .A3(_02114_ ), .ZN(_02115_ ) );
NOR2_X1 _09700_ ( .A1(_02021_ ), .A2(_02115_ ), .ZN(_02116_ ) );
INV_X1 _09701_ ( .A(_02116_ ), .ZN(_02117_ ) );
AND2_X1 _09702_ ( .A1(_01969_ ), .A2(\ID_EX_imm [16] ), .ZN(_02118_ ) );
AND2_X1 _09703_ ( .A1(_01947_ ), .A2(_02118_ ), .ZN(_02119_ ) );
AOI21_X1 _09704_ ( .A(_02119_ ), .B1(\ID_EX_imm [17] ), .B2(_01945_ ), .ZN(_02120_ ) );
INV_X1 _09705_ ( .A(_02020_ ), .ZN(_02121_ ) );
NOR4_X1 _09706_ ( .A1(_02120_ ), .A2(_01996_ ), .A3(_01995_ ), .A4(_02121_ ), .ZN(_02122_ ) );
INV_X1 _09707_ ( .A(_02018_ ), .ZN(_02123_ ) );
NOR4_X1 _09708_ ( .A1(_01995_ ), .A2(_02123_ ), .A3(_01996_ ), .A4(_02019_ ), .ZN(_02124_ ) );
NOR3_X1 _09709_ ( .A1(_02122_ ), .A2(_01996_ ), .A3(_02124_ ), .ZN(_02125_ ) );
NOR2_X1 _09710_ ( .A1(_02125_ ), .A2(_02115_ ), .ZN(_02126_ ) );
AND2_X1 _09711_ ( .A1(_02042_ ), .A2(\ID_EX_imm [23] ), .ZN(_02127_ ) );
NAND2_X1 _09712_ ( .A1(_02088_ ), .A2(\ID_EX_imm [20] ), .ZN(_02128_ ) );
NOR3_X1 _09713_ ( .A1(_02128_ ), .A2(_02112_ ), .A3(_02113_ ), .ZN(_02129_ ) );
OR2_X1 _09714_ ( .A1(_02129_ ), .A2(_02113_ ), .ZN(_02130_ ) );
AND2_X1 _09715_ ( .A1(_02067_ ), .A2(_02130_ ), .ZN(_02131_ ) );
AND2_X1 _09716_ ( .A1(_02064_ ), .A2(\ID_EX_imm [22] ), .ZN(_02132_ ) );
AND2_X1 _09717_ ( .A1(_02043_ ), .A2(_02132_ ), .ZN(_02133_ ) );
NOR4_X1 _09718_ ( .A1(_02126_ ), .A2(_02127_ ), .A3(_02131_ ), .A4(_02133_ ), .ZN(_02134_ ) );
AOI21_X2 _09719_ ( .A(_01499_ ), .B1(_02117_ ), .B2(_02134_ ), .ZN(_02135_ ) );
AOI21_X1 _09720_ ( .A(_01497_ ), .B1(_01475_ ), .B2(_01495_ ), .ZN(_02136_ ) );
NOR2_X2 _09721_ ( .A1(_02135_ ), .A2(_02136_ ), .ZN(_02137_ ) );
OR3_X1 _09722_ ( .A1(_01388_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01399_ ), .ZN(_02138_ ) );
OR2_X1 _09723_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02139_ ) );
OAI211_X1 _09724_ ( .A(_02139_ ), .B(_01452_ ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02140_ ) );
OR2_X1 _09725_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02141_ ) );
OAI211_X1 _09726_ ( .A(_02141_ ), .B(fanout_net_20 ), .C1(_01417_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02142_ ) );
NAND3_X1 _09727_ ( .A1(_02140_ ), .A2(_02142_ ), .A3(_01410_ ), .ZN(_02143_ ) );
MUX2_X1 _09728_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02144_ ) );
MUX2_X1 _09729_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02145_ ) );
MUX2_X1 _09730_ ( .A(_02144_ ), .B(_02145_ ), .S(_01427_ ), .Z(_02146_ ) );
OAI211_X1 _09731_ ( .A(_01404_ ), .B(_02143_ ), .C1(_02146_ ), .C2(_01433_ ), .ZN(_02147_ ) );
OR2_X1 _09732_ ( .A1(_01416_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02148_ ) );
OAI211_X1 _09733_ ( .A(_02148_ ), .B(_01427_ ), .C1(fanout_net_17 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02149_ ) );
NOR2_X1 _09734_ ( .A1(_01455_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02150_ ) );
OAI21_X1 _09735_ ( .A(fanout_net_20 ), .B1(fanout_net_17 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02151_ ) );
OAI211_X1 _09736_ ( .A(_02149_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .C1(_02150_ ), .C2(_02151_ ), .ZN(_02152_ ) );
MUX2_X1 _09737_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02153_ ) );
MUX2_X1 _09738_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02154_ ) );
MUX2_X1 _09739_ ( .A(_02153_ ), .B(_02154_ ), .S(fanout_net_20 ), .Z(_02155_ ) );
OAI211_X1 _09740_ ( .A(_02152_ ), .B(fanout_net_22 ), .C1(_02155_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02156_ ) );
OAI211_X1 _09741_ ( .A(_02147_ ), .B(_02156_ ), .C1(_01389_ ), .C2(_01444_ ), .ZN(_02157_ ) );
NAND2_X1 _09742_ ( .A1(_02138_ ), .A2(_02157_ ), .ZN(_02158_ ) );
NAND2_X1 _09743_ ( .A1(_02158_ ), .A2(\ID_EX_imm [25] ), .ZN(_02159_ ) );
NAND2_X1 _09744_ ( .A1(_02137_ ), .A2(_02159_ ), .ZN(_02160_ ) );
OR3_X1 _09745_ ( .A1(_01388_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_01399_ ), .ZN(_02161_ ) );
OR2_X1 _09746_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02162_ ) );
OAI211_X1 _09747_ ( .A(_02162_ ), .B(_01427_ ), .C1(_01417_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02163_ ) );
INV_X1 _09748_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02164_ ) );
NAND2_X1 _09749_ ( .A1(_02164_ ), .A2(fanout_net_17 ), .ZN(_02165_ ) );
OAI211_X1 _09750_ ( .A(_02165_ ), .B(fanout_net_20 ), .C1(fanout_net_17 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02166_ ) );
NAND3_X1 _09751_ ( .A1(_02163_ ), .A2(_02166_ ), .A3(_01410_ ), .ZN(_02167_ ) );
MUX2_X1 _09752_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02168_ ) );
MUX2_X1 _09753_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02169_ ) );
MUX2_X1 _09754_ ( .A(_02168_ ), .B(_02169_ ), .S(_01451_ ), .Z(_02170_ ) );
OAI211_X1 _09755_ ( .A(fanout_net_22 ), .B(_02167_ ), .C1(_02170_ ), .C2(_01433_ ), .ZN(_02171_ ) );
OR2_X1 _09756_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02172_ ) );
OAI211_X1 _09757_ ( .A(_02172_ ), .B(_01427_ ), .C1(_01417_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02173_ ) );
OR2_X1 _09758_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02174_ ) );
OAI211_X1 _09759_ ( .A(_02174_ ), .B(fanout_net_20 ), .C1(_01417_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02175_ ) );
NAND3_X1 _09760_ ( .A1(_02173_ ), .A2(_02175_ ), .A3(_01410_ ), .ZN(_02176_ ) );
MUX2_X1 _09761_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02177_ ) );
MUX2_X1 _09762_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02178_ ) );
MUX2_X1 _09763_ ( .A(_02177_ ), .B(_02178_ ), .S(_01451_ ), .Z(_02179_ ) );
OAI211_X1 _09764_ ( .A(_01404_ ), .B(_02176_ ), .C1(_02179_ ), .C2(_01433_ ), .ZN(_02180_ ) );
OAI211_X1 _09765_ ( .A(_02171_ ), .B(_02180_ ), .C1(_01389_ ), .C2(_01444_ ), .ZN(_02181_ ) );
NAND2_X1 _09766_ ( .A1(_02161_ ), .A2(_02181_ ), .ZN(_02182_ ) );
INV_X1 _09767_ ( .A(\ID_EX_imm [26] ), .ZN(_02183_ ) );
XNOR2_X1 _09768_ ( .A(_02182_ ), .B(_02183_ ), .ZN(_02184_ ) );
INV_X1 _09769_ ( .A(\ID_EX_imm [25] ), .ZN(_02185_ ) );
NAND3_X1 _09770_ ( .A1(_02138_ ), .A2(_02185_ ), .A3(_02157_ ), .ZN(_02186_ ) );
AND4_X2 _09771_ ( .A1(_01474_ ), .A2(_02160_ ), .A3(_02184_ ), .A4(_02186_ ), .ZN(_02187_ ) );
INV_X1 _09772_ ( .A(_02187_ ), .ZN(_02188_ ) );
AND2_X1 _09773_ ( .A1(_02182_ ), .A2(\ID_EX_imm [26] ), .ZN(_02189_ ) );
AND2_X1 _09774_ ( .A1(_01474_ ), .A2(_02189_ ), .ZN(_02190_ ) );
AOI21_X1 _09775_ ( .A(_02190_ ), .B1(\ID_EX_imm [27] ), .B2(_01472_ ), .ZN(_02191_ ) );
AND2_X2 _09776_ ( .A1(_02188_ ), .A2(_02191_ ), .ZN(_02192_ ) );
OR3_X1 _09777_ ( .A1(_01389_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01444_ ), .ZN(_02193_ ) );
OR2_X1 _09778_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02194_ ) );
OAI211_X1 _09779_ ( .A(_02194_ ), .B(_01452_ ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02195_ ) );
INV_X1 _09780_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02196_ ) );
NAND2_X1 _09781_ ( .A1(_02196_ ), .A2(fanout_net_17 ), .ZN(_02197_ ) );
OAI211_X1 _09782_ ( .A(_02197_ ), .B(fanout_net_20 ), .C1(fanout_net_17 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02198_ ) );
NAND3_X1 _09783_ ( .A1(_02195_ ), .A2(_02198_ ), .A3(_01433_ ), .ZN(_02199_ ) );
MUX2_X1 _09784_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02200_ ) );
MUX2_X1 _09785_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02201_ ) );
MUX2_X1 _09786_ ( .A(_02200_ ), .B(_02201_ ), .S(_01452_ ), .Z(_02202_ ) );
OAI211_X1 _09787_ ( .A(_01404_ ), .B(_02199_ ), .C1(_02202_ ), .C2(_01433_ ), .ZN(_02203_ ) );
OR2_X1 _09788_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02204_ ) );
OAI211_X1 _09789_ ( .A(_02204_ ), .B(fanout_net_20 ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02205_ ) );
OR2_X1 _09790_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02206_ ) );
OAI211_X1 _09791_ ( .A(_02206_ ), .B(_01452_ ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02207_ ) );
NAND3_X1 _09792_ ( .A1(_02205_ ), .A2(_02207_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02208_ ) );
MUX2_X1 _09793_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02209_ ) );
MUX2_X1 _09794_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02210_ ) );
MUX2_X1 _09795_ ( .A(_02209_ ), .B(_02210_ ), .S(fanout_net_20 ), .Z(_02211_ ) );
OAI211_X1 _09796_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02208_ ), .C1(_02211_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02212_ ) );
OAI211_X1 _09797_ ( .A(_02203_ ), .B(_02212_ ), .C1(_01389_ ), .C2(_01444_ ), .ZN(_02213_ ) );
NAND2_X1 _09798_ ( .A1(_02193_ ), .A2(_02213_ ), .ZN(_02214_ ) );
XNOR2_X1 _09799_ ( .A(_02214_ ), .B(\ID_EX_imm [29] ), .ZN(_02215_ ) );
OR3_X1 _09800_ ( .A1(_01388_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_01399_ ), .ZN(_02216_ ) );
OR2_X1 _09801_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02217_ ) );
OAI211_X1 _09802_ ( .A(_02217_ ), .B(_01427_ ), .C1(_01417_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02218_ ) );
OR2_X1 _09803_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02219_ ) );
OAI211_X1 _09804_ ( .A(_02219_ ), .B(fanout_net_20 ), .C1(_01477_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02220_ ) );
NAND3_X1 _09805_ ( .A1(_02218_ ), .A2(_02220_ ), .A3(_01410_ ), .ZN(_02221_ ) );
MUX2_X1 _09806_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02222_ ) );
MUX2_X1 _09807_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02223_ ) );
MUX2_X1 _09808_ ( .A(_02222_ ), .B(_02223_ ), .S(_01451_ ), .Z(_02224_ ) );
OAI211_X1 _09809_ ( .A(_01404_ ), .B(_02221_ ), .C1(_02224_ ), .C2(_01433_ ), .ZN(_02225_ ) );
OR2_X1 _09810_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02226_ ) );
OAI211_X1 _09811_ ( .A(_02226_ ), .B(fanout_net_20 ), .C1(_01477_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02227_ ) );
OR2_X1 _09812_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02228_ ) );
OAI211_X1 _09813_ ( .A(_02228_ ), .B(_01451_ ), .C1(_01477_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02229_ ) );
NAND3_X1 _09814_ ( .A1(_02227_ ), .A2(_02229_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02230_ ) );
MUX2_X1 _09815_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02231_ ) );
MUX2_X1 _09816_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02232_ ) );
MUX2_X1 _09817_ ( .A(_02231_ ), .B(_02232_ ), .S(fanout_net_20 ), .Z(_02233_ ) );
OAI211_X1 _09818_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02230_ ), .C1(_02233_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02234_ ) );
OAI211_X1 _09819_ ( .A(_02225_ ), .B(_02234_ ), .C1(_01388_ ), .C2(_01399_ ), .ZN(_02235_ ) );
NAND2_X2 _09820_ ( .A1(_02216_ ), .A2(_02235_ ), .ZN(_02236_ ) );
XNOR2_X1 _09821_ ( .A(_02236_ ), .B(\ID_EX_imm [28] ), .ZN(_02237_ ) );
NOR3_X2 _09822_ ( .A1(_02192_ ), .A2(_02215_ ), .A3(_02237_ ), .ZN(_02238_ ) );
INV_X1 _09823_ ( .A(_02238_ ), .ZN(_02239_ ) );
INV_X1 _09824_ ( .A(_02215_ ), .ZN(_02240_ ) );
AOI21_X1 _09825_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02216_ ), .B2(_02235_ ), .ZN(_02241_ ) );
INV_X1 _09826_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02242_ ) );
AOI22_X1 _09827_ ( .A1(_02240_ ), .A2(_02241_ ), .B1(_02242_ ), .B2(_02214_ ), .ZN(_02243_ ) );
AOI21_X2 _09828_ ( .A(_01448_ ), .B1(_02239_ ), .B2(_02243_ ), .ZN(_02244_ ) );
AOI21_X1 _09829_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_01400_ ), .B2(_01445_ ), .ZN(_02245_ ) );
OR3_X1 _09830_ ( .A1(_01389_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_01444_ ), .ZN(_02246_ ) );
OR2_X1 _09831_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02247_ ) );
OAI211_X1 _09832_ ( .A(_02247_ ), .B(_01452_ ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02248_ ) );
OR2_X1 _09833_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02249_ ) );
OAI211_X1 _09834_ ( .A(_02249_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01455_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02250_ ) );
NAND3_X1 _09835_ ( .A1(_02248_ ), .A2(_02250_ ), .A3(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02251_ ) );
MUX2_X1 _09836_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02252_ ) );
MUX2_X1 _09837_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02253_ ) );
MUX2_X1 _09838_ ( .A(_02252_ ), .B(_02253_ ), .S(_01452_ ), .Z(_02254_ ) );
OAI211_X1 _09839_ ( .A(_01404_ ), .B(_02251_ ), .C1(_02254_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_02255_ ) );
NOR2_X1 _09840_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02256_ ) );
OAI21_X1 _09841_ ( .A(_01427_ ), .B1(_01417_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02257_ ) );
INV_X1 _09842_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02258_ ) );
INV_X1 _09843_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02259_ ) );
MUX2_X1 _09844_ ( .A(_02258_ ), .B(_02259_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02260_ ) );
OAI221_X1 _09845_ ( .A(_01410_ ), .B1(_02256_ ), .B2(_02257_ ), .C1(_02260_ ), .C2(_01452_ ), .ZN(_02261_ ) );
MUX2_X1 _09846_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02262_ ) );
MUX2_X1 _09847_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02263_ ) );
MUX2_X1 _09848_ ( .A(_02262_ ), .B(_02263_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02264_ ) );
OAI211_X1 _09849_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02261_ ), .C1(_02264_ ), .C2(_01433_ ), .ZN(_02265_ ) );
OAI211_X1 _09850_ ( .A(_02255_ ), .B(_02265_ ), .C1(_01389_ ), .C2(_01444_ ), .ZN(_02266_ ) );
NAND2_X1 _09851_ ( .A1(_02246_ ), .A2(_02266_ ), .ZN(_02267_ ) );
BUF_X4 _09852_ ( .A(_02267_ ), .Z(_02268_ ) );
XNOR2_X1 _09853_ ( .A(_02268_ ), .B(\ID_EX_imm [31] ), .ZN(_02269_ ) );
OR3_X1 _09854_ ( .A1(_02244_ ), .A2(_02245_ ), .A3(_02269_ ), .ZN(_02270_ ) );
OAI21_X1 _09855_ ( .A(_02269_ ), .B1(_02244_ ), .B2(_02245_ ), .ZN(_02271_ ) );
AOI21_X1 _09856_ ( .A(_01370_ ), .B1(_02270_ ), .B2(_02271_ ), .ZN(_00097_ ) );
AND3_X1 _09857_ ( .A1(_02239_ ), .A2(_02243_ ), .A3(_01448_ ), .ZN(_02272_ ) );
NOR3_X1 _09858_ ( .A1(_02272_ ), .A2(_02244_ ), .A3(_01369_ ), .ZN(_00098_ ) );
AND2_X1 _09859_ ( .A1(_02021_ ), .A2(_02125_ ), .ZN(_02273_ ) );
INV_X1 _09860_ ( .A(_02090_ ), .ZN(_02274_ ) );
NOR2_X1 _09861_ ( .A1(_02273_ ), .A2(_02274_ ), .ZN(_02275_ ) );
AND2_X1 _09862_ ( .A1(_02088_ ), .A2(\ID_EX_imm [20] ), .ZN(_02276_ ) );
OAI22_X1 _09863_ ( .A1(_02275_ ), .A2(_02276_ ), .B1(_02113_ ), .B2(_02112_ ), .ZN(_02277_ ) );
OAI211_X1 _09864_ ( .A(_02128_ ), .B(_02114_ ), .C1(_02273_ ), .C2(_02274_ ), .ZN(_02278_ ) );
AOI21_X1 _09865_ ( .A(_01370_ ), .B1(_02277_ ), .B2(_02278_ ), .ZN(_00099_ ) );
AND3_X1 _09866_ ( .A1(_02021_ ), .A2(_02274_ ), .A3(_02125_ ), .ZN(_02279_ ) );
NOR3_X1 _09867_ ( .A1(_02275_ ), .A2(_01370_ ), .A3(_02279_ ), .ZN(_00100_ ) );
INV_X1 _09868_ ( .A(_01973_ ), .ZN(_02280_ ) );
AOI21_X1 _09869_ ( .A(_02121_ ), .B1(_02280_ ), .B2(_02120_ ), .ZN(_02281_ ) );
AND2_X1 _09870_ ( .A1(_02018_ ), .A2(\ID_EX_imm [18] ), .ZN(_02282_ ) );
OR3_X1 _09871_ ( .A1(_02281_ ), .A2(_01997_ ), .A3(_02282_ ), .ZN(_02283_ ) );
BUF_X2 _09872_ ( .A(_01368_ ), .Z(_02284_ ) );
OAI21_X1 _09873_ ( .A(_01997_ ), .B1(_02281_ ), .B2(_02282_ ), .ZN(_02285_ ) );
AND3_X1 _09874_ ( .A1(_02283_ ), .A2(_02284_ ), .A3(_02285_ ), .ZN(_00101_ ) );
AND3_X1 _09875_ ( .A1(_02280_ ), .A2(_02121_ ), .A3(_02120_ ), .ZN(_02286_ ) );
NOR3_X1 _09876_ ( .A1(_02286_ ), .A2(_02281_ ), .A3(_01369_ ), .ZN(_00102_ ) );
NOR2_X1 _09877_ ( .A1(_01921_ ), .A2(_01972_ ), .ZN(_02287_ ) );
OR3_X1 _09878_ ( .A1(_02287_ ), .A2(_01948_ ), .A3(_02118_ ), .ZN(_02288_ ) );
OAI21_X1 _09879_ ( .A(_01948_ ), .B1(_02287_ ), .B2(_02118_ ), .ZN(_02289_ ) );
AOI21_X1 _09880_ ( .A(_01370_ ), .B1(_02288_ ), .B2(_02289_ ), .ZN(_00103_ ) );
NOR3_X1 _09881_ ( .A1(_01908_ ), .A2(_01920_ ), .A3(_01971_ ), .ZN(_02290_ ) );
NOR3_X1 _09882_ ( .A1(_02287_ ), .A2(_01370_ ), .A3(_02290_ ), .ZN(_00104_ ) );
NOR2_X1 _09883_ ( .A1(_01717_ ), .A2(_01907_ ), .ZN(_02291_ ) );
INV_X1 _09884_ ( .A(_01919_ ), .ZN(_02292_ ) );
NOR2_X1 _09885_ ( .A1(_02291_ ), .A2(_02292_ ), .ZN(_02293_ ) );
INV_X1 _09886_ ( .A(_01810_ ), .ZN(_02294_ ) );
NOR4_X1 _09887_ ( .A1(_02293_ ), .A2(_01785_ ), .A3(_01786_ ), .A4(_02294_ ), .ZN(_02295_ ) );
OR2_X1 _09888_ ( .A1(_02295_ ), .A2(_01912_ ), .ZN(_02296_ ) );
AND2_X1 _09889_ ( .A1(_02296_ ), .A2(_01739_ ), .ZN(_02297_ ) );
AND2_X1 _09890_ ( .A1(_01738_ ), .A2(\ID_EX_imm [14] ), .ZN(_02298_ ) );
OR3_X1 _09891_ ( .A1(_02297_ ), .A2(_01762_ ), .A3(_02298_ ), .ZN(_02299_ ) );
OAI21_X1 _09892_ ( .A(_01762_ ), .B1(_02297_ ), .B2(_02298_ ), .ZN(_02300_ ) );
AND3_X1 _09893_ ( .A1(_02299_ ), .A2(_02284_ ), .A3(_02300_ ), .ZN(_00105_ ) );
NOR3_X1 _09894_ ( .A1(_02295_ ), .A2(_01739_ ), .A3(_01912_ ), .ZN(_02301_ ) );
NOR3_X1 _09895_ ( .A1(_02297_ ), .A2(_01370_ ), .A3(_02301_ ), .ZN(_00106_ ) );
NOR2_X1 _09896_ ( .A1(_02293_ ), .A2(_02294_ ), .ZN(_02302_ ) );
OR3_X1 _09897_ ( .A1(_02302_ ), .A2(_01910_ ), .A3(_01787_ ), .ZN(_02303_ ) );
OAI21_X1 _09898_ ( .A(_01787_ ), .B1(_02302_ ), .B2(_01910_ ), .ZN(_02304_ ) );
AND3_X1 _09899_ ( .A1(_02303_ ), .A2(_02284_ ), .A3(_02304_ ), .ZN(_00107_ ) );
NOR3_X1 _09900_ ( .A1(_02291_ ), .A2(_01810_ ), .A3(_02292_ ), .ZN(_02305_ ) );
NOR3_X1 _09901_ ( .A1(_02302_ ), .A2(_01370_ ), .A3(_02305_ ), .ZN(_00108_ ) );
NOR2_X1 _09902_ ( .A1(_02192_ ), .A2(_02237_ ), .ZN(_02306_ ) );
OAI21_X1 _09903_ ( .A(_02215_ ), .B1(_02306_ ), .B2(_02241_ ), .ZN(_02307_ ) );
INV_X1 _09904_ ( .A(_02236_ ), .ZN(_02308_ ) );
OAI221_X1 _09905_ ( .A(_02240_ ), .B1(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_02308_ ), .C1(_02192_ ), .C2(_02237_ ), .ZN(_02309_ ) );
AOI21_X1 _09906_ ( .A(_01369_ ), .B1(_02307_ ), .B2(_02309_ ), .ZN(_00109_ ) );
AND3_X1 _09907_ ( .A1(_02188_ ), .A2(_02191_ ), .A3(_02237_ ), .ZN(_02310_ ) );
NOR3_X1 _09908_ ( .A1(_02306_ ), .A2(_01370_ ), .A3(_02310_ ), .ZN(_00110_ ) );
AND3_X1 _09909_ ( .A1(_02160_ ), .A2(_02184_ ), .A3(_02186_ ), .ZN(_02311_ ) );
OR3_X1 _09910_ ( .A1(_02311_ ), .A2(_02189_ ), .A3(_01474_ ), .ZN(_02312_ ) );
OAI21_X1 _09911_ ( .A(_01474_ ), .B1(_02311_ ), .B2(_02189_ ), .ZN(_02313_ ) );
AND3_X1 _09912_ ( .A1(_02312_ ), .A2(_02284_ ), .A3(_02313_ ), .ZN(_00111_ ) );
AOI21_X1 _09913_ ( .A(_02184_ ), .B1(_02160_ ), .B2(_02186_ ), .ZN(_02314_ ) );
NOR3_X1 _09914_ ( .A1(_02311_ ), .A2(_02314_ ), .A3(_01369_ ), .ZN(_00112_ ) );
NAND2_X1 _09915_ ( .A1(_02159_ ), .A2(_02186_ ), .ZN(_02315_ ) );
XNOR2_X1 _09916_ ( .A(_02137_ ), .B(_02315_ ), .ZN(_02316_ ) );
NOR2_X1 _09917_ ( .A1(_02316_ ), .A2(_01370_ ), .ZN(_00113_ ) );
AND3_X1 _09918_ ( .A1(_02117_ ), .A2(_02134_ ), .A3(_01499_ ), .ZN(_02317_ ) );
NOR3_X1 _09919_ ( .A1(_02317_ ), .A2(_02135_ ), .A3(_01369_ ), .ZN(_00114_ ) );
NOR4_X1 _09920_ ( .A1(_02273_ ), .A2(_02274_ ), .A3(_02113_ ), .A4(_02112_ ), .ZN(_02318_ ) );
OR2_X1 _09921_ ( .A1(_02318_ ), .A2(_02130_ ), .ZN(_02319_ ) );
AND2_X1 _09922_ ( .A1(_02319_ ), .A2(_02066_ ), .ZN(_02320_ ) );
OR3_X1 _09923_ ( .A1(_02320_ ), .A2(_02043_ ), .A3(_02132_ ), .ZN(_02321_ ) );
OAI21_X1 _09924_ ( .A(_02043_ ), .B1(_02320_ ), .B2(_02132_ ), .ZN(_02322_ ) );
AND3_X1 _09925_ ( .A1(_02321_ ), .A2(_02284_ ), .A3(_02322_ ), .ZN(_00115_ ) );
NOR3_X1 _09926_ ( .A1(_02318_ ), .A2(_02066_ ), .A3(_02130_ ), .ZN(_02323_ ) );
NOR3_X1 _09927_ ( .A1(_02320_ ), .A2(_01370_ ), .A3(_02323_ ), .ZN(_00116_ ) );
AND2_X1 _09928_ ( .A1(_01345_ ), .A2(\ID_EX_rd [4] ), .ZN(_00117_ ) );
AND2_X1 _09929_ ( .A1(_01345_ ), .A2(\ID_EX_rd [3] ), .ZN(_00118_ ) );
AND2_X1 _09930_ ( .A1(_01345_ ), .A2(\ID_EX_rd [2] ), .ZN(_00119_ ) );
AND2_X1 _09931_ ( .A1(_01345_ ), .A2(\ID_EX_rd [1] ), .ZN(_00120_ ) );
AND2_X1 _09932_ ( .A1(_01345_ ), .A2(\ID_EX_rd [0] ), .ZN(_00121_ ) );
INV_X1 _09933_ ( .A(\ID_EX_pc [31] ), .ZN(_02324_ ) );
NOR3_X1 _09934_ ( .A1(_02324_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00122_ ) );
INV_X1 _09935_ ( .A(\ID_EX_pc [30] ), .ZN(_02325_ ) );
NOR3_X1 _09936_ ( .A1(_02325_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00123_ ) );
INV_X1 _09937_ ( .A(\ID_EX_pc [21] ), .ZN(_02326_ ) );
NOR3_X1 _09938_ ( .A1(_02326_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00124_ ) );
INV_X1 _09939_ ( .A(\ID_EX_pc [20] ), .ZN(_02327_ ) );
NOR3_X1 _09940_ ( .A1(_02327_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00125_ ) );
INV_X1 _09941_ ( .A(\ID_EX_pc [19] ), .ZN(_02328_ ) );
NOR3_X1 _09942_ ( .A1(_02328_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00126_ ) );
INV_X1 _09943_ ( .A(\ID_EX_pc [18] ), .ZN(_02329_ ) );
NOR3_X1 _09944_ ( .A1(_02329_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00127_ ) );
INV_X1 _09945_ ( .A(\ID_EX_pc [17] ), .ZN(_02330_ ) );
NOR3_X1 _09946_ ( .A1(_02330_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00128_ ) );
INV_X1 _09947_ ( .A(\ID_EX_pc [16] ), .ZN(_02331_ ) );
NOR3_X1 _09948_ ( .A1(_02331_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00129_ ) );
INV_X1 _09949_ ( .A(\ID_EX_pc [15] ), .ZN(_02332_ ) );
NOR3_X1 _09950_ ( .A1(_02332_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00130_ ) );
INV_X1 _09951_ ( .A(\ID_EX_pc [14] ), .ZN(_02333_ ) );
NOR3_X1 _09952_ ( .A1(_02333_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00131_ ) );
INV_X1 _09953_ ( .A(\ID_EX_pc [13] ), .ZN(_02334_ ) );
NOR3_X1 _09954_ ( .A1(_02334_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00132_ ) );
INV_X1 _09955_ ( .A(\ID_EX_pc [12] ), .ZN(_02335_ ) );
NOR3_X1 _09956_ ( .A1(_02335_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00133_ ) );
INV_X1 _09957_ ( .A(\ID_EX_pc [29] ), .ZN(_02336_ ) );
NOR3_X1 _09958_ ( .A1(_02336_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00134_ ) );
INV_X1 _09959_ ( .A(\ID_EX_pc [11] ), .ZN(_02337_ ) );
NOR3_X1 _09960_ ( .A1(_02337_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00135_ ) );
INV_X1 _09961_ ( .A(\ID_EX_pc [10] ), .ZN(_02338_ ) );
NOR3_X1 _09962_ ( .A1(_02338_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00136_ ) );
INV_X1 _09963_ ( .A(\ID_EX_pc [9] ), .ZN(_02339_ ) );
NOR3_X1 _09964_ ( .A1(_02339_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00137_ ) );
INV_X1 _09965_ ( .A(\ID_EX_pc [8] ), .ZN(_02340_ ) );
NOR3_X1 _09966_ ( .A1(_02340_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00138_ ) );
INV_X1 _09967_ ( .A(\ID_EX_pc [7] ), .ZN(_02341_ ) );
NOR3_X1 _09968_ ( .A1(_02341_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00139_ ) );
AND2_X1 _09969_ ( .A1(_01345_ ), .A2(\ID_EX_pc [6] ), .ZN(_00140_ ) );
INV_X1 _09970_ ( .A(\ID_EX_pc [5] ), .ZN(_02342_ ) );
NOR3_X1 _09971_ ( .A1(_02342_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00141_ ) );
INV_X1 _09972_ ( .A(\ID_EX_pc [4] ), .ZN(_02343_ ) );
NOR3_X1 _09973_ ( .A1(_02343_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00142_ ) );
INV_X1 _09974_ ( .A(\ID_EX_pc [3] ), .ZN(_02344_ ) );
NOR3_X1 _09975_ ( .A1(_02344_ ), .A2(fanout_net_2 ), .A3(fanout_net_9 ), .ZN(_00143_ ) );
INV_X1 _09976_ ( .A(\ID_EX_pc [2] ), .ZN(_02345_ ) );
NOR3_X1 _09977_ ( .A1(_02345_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00144_ ) );
INV_X1 _09978_ ( .A(\ID_EX_pc [28] ), .ZN(_02346_ ) );
NOR3_X1 _09979_ ( .A1(_02346_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00145_ ) );
INV_X1 _09980_ ( .A(\ID_EX_pc [1] ), .ZN(_02347_ ) );
NOR3_X1 _09981_ ( .A1(_02347_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00146_ ) );
INV_X1 _09982_ ( .A(\ID_EX_pc [0] ), .ZN(_02348_ ) );
NOR3_X1 _09983_ ( .A1(_02348_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00147_ ) );
INV_X1 _09984_ ( .A(\ID_EX_pc [27] ), .ZN(_02349_ ) );
NOR3_X1 _09985_ ( .A1(_02349_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00148_ ) );
INV_X1 _09986_ ( .A(\ID_EX_pc [26] ), .ZN(_02350_ ) );
NOR3_X1 _09987_ ( .A1(_02350_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00149_ ) );
INV_X1 _09988_ ( .A(\ID_EX_pc [25] ), .ZN(_02351_ ) );
NOR3_X1 _09989_ ( .A1(_02351_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00150_ ) );
INV_X1 _09990_ ( .A(\ID_EX_pc [24] ), .ZN(_02352_ ) );
NOR3_X1 _09991_ ( .A1(_02352_ ), .A2(fanout_net_3 ), .A3(fanout_net_9 ), .ZN(_00151_ ) );
INV_X1 _09992_ ( .A(\ID_EX_pc [23] ), .ZN(_02353_ ) );
NOR3_X1 _09993_ ( .A1(_02353_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00152_ ) );
INV_X1 _09994_ ( .A(\ID_EX_pc [22] ), .ZN(_02354_ ) );
NOR3_X1 _09995_ ( .A1(_02354_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00153_ ) );
NOR3_X1 _09996_ ( .A1(_01355_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00154_ ) );
INV_X4 _09997_ ( .A(_01324_ ), .ZN(_02355_ ) );
AND2_X1 _09998_ ( .A1(_01245_ ), .A2(_01246_ ), .ZN(_02356_ ) );
AND4_X2 _09999_ ( .A1(_01252_ ), .A2(_01266_ ), .A3(_01228_ ), .A4(_02356_ ), .ZN(_02357_ ) );
NAND2_X4 _10000_ ( .A1(_01326_ ), .A2(_02357_ ), .ZN(_02358_ ) );
NOR2_X4 _10001_ ( .A1(_02355_ ), .A2(_02358_ ), .ZN(_02359_ ) );
BUF_X8 _10002_ ( .A(_02359_ ), .Z(_02360_ ) );
BUF_X16 _10003_ ( .A(_02360_ ), .Z(_02361_ ) );
MUX2_X1 _10004_ ( .A(io_master_arready ), .B(_01321_ ), .S(_02361_ ), .Z(_02362_ ) );
BUF_X2 _10005_ ( .A(_01215_ ), .Z(_02363_ ) );
BUF_X2 _10006_ ( .A(_02363_ ), .Z(_02364_ ) );
BUF_X2 _10007_ ( .A(_02364_ ), .Z(\io_master_arid [1] ) );
AND2_X1 _10008_ ( .A1(_02362_ ), .A2(\io_master_arid [1] ), .ZN(_02365_ ) );
INV_X1 _10009_ ( .A(_01290_ ), .ZN(_02366_ ) );
NOR3_X1 _10010_ ( .A1(_02365_ ), .A2(_01217_ ), .A3(_02366_ ), .ZN(_02367_ ) );
INV_X1 _10011_ ( .A(_02367_ ), .ZN(_02368_ ) );
INV_X1 _10012_ ( .A(io_master_awready ), .ZN(_02369_ ) );
NAND4_X1 _10013_ ( .A1(_01374_ ), .A2(_02369_ ), .A3(\EX_LS_flag [1] ), .A4(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02370_ ) );
OAI21_X1 _10014_ ( .A(_02370_ ), .B1(\mylsu.state [4] ), .B2(\mylsu.state [0] ), .ZN(_02371_ ) );
AOI21_X1 _10015_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .B1(_02371_ ), .B2(EXU_valid_LSU ), .ZN(_02372_ ) );
AOI21_X1 _10016_ ( .A(_01346_ ), .B1(_02368_ ), .B2(_02372_ ), .ZN(_00155_ ) );
NOR3_X1 _10017_ ( .A1(_01348_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00156_ ) );
NOR3_X1 _10018_ ( .A1(_01359_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00157_ ) );
INV_X1 _10019_ ( .A(fanout_net_8 ), .ZN(_02373_ ) );
BUF_X4 _10020_ ( .A(_02373_ ), .Z(_02374_ ) );
BUF_X4 _10021_ ( .A(_02374_ ), .Z(_02375_ ) );
BUF_X2 _10022_ ( .A(_02375_ ), .Z(_02376_ ) );
NOR3_X1 _10023_ ( .A1(_02376_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00158_ ) );
INV_X1 _10024_ ( .A(\ID_EX_typ [3] ), .ZN(_02377_ ) );
NOR3_X1 _10025_ ( .A1(_02377_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00159_ ) );
INV_X1 _10026_ ( .A(fanout_net_7 ), .ZN(_02378_ ) );
BUF_X4 _10027_ ( .A(_02378_ ), .Z(_02379_ ) );
NOR3_X1 _10028_ ( .A1(_02379_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00160_ ) );
INV_X1 _10029_ ( .A(\ID_EX_typ [1] ), .ZN(_02380_ ) );
NOR3_X1 _10030_ ( .A1(_02380_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00161_ ) );
BUF_X4 _10031_ ( .A(_01350_ ), .Z(_02381_ ) );
NOR3_X1 _10032_ ( .A1(_02381_ ), .A2(fanout_net_3 ), .A3(excp_written ), .ZN(_00162_ ) );
AND2_X1 _10033_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_02382_ ) );
NOR2_X1 _10034_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_02383_ ) );
AND2_X2 _10035_ ( .A1(_02382_ ), .A2(_02383_ ), .ZN(_02384_ ) );
AND2_X1 _10036_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_02385_ ) );
INV_X1 _10037_ ( .A(\IF_ID_inst [6] ), .ZN(_02386_ ) );
NOR2_X1 _10038_ ( .A1(_02386_ ), .A2(\IF_ID_inst [12] ), .ZN(_02387_ ) );
AND3_X1 _10039_ ( .A1(_02384_ ), .A2(_02385_ ), .A3(_02387_ ), .ZN(_02388_ ) );
AND2_X2 _10040_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_02389_ ) );
NAND2_X1 _10041_ ( .A1(_02388_ ), .A2(_02389_ ), .ZN(_02390_ ) );
CLKBUF_X2 _10042_ ( .A(_02384_ ), .Z(_02391_ ) );
INV_X1 _10043_ ( .A(\IF_ID_inst [13] ), .ZN(_02392_ ) );
NOR2_X1 _10044_ ( .A1(_02392_ ), .A2(\IF_ID_inst [14] ), .ZN(_02393_ ) );
NAND4_X1 _10045_ ( .A1(_02391_ ), .A2(_02385_ ), .A3(_02387_ ), .A4(_02393_ ), .ZN(_02394_ ) );
NAND2_X1 _10046_ ( .A1(_02390_ ), .A2(_02394_ ), .ZN(_02395_ ) );
AND2_X1 _10047_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_02396_ ) );
AND3_X1 _10048_ ( .A1(_02382_ ), .A2(_02396_ ), .A3(_02383_ ), .ZN(_02397_ ) );
AND2_X1 _10049_ ( .A1(_02397_ ), .A2(_02385_ ), .ZN(_02398_ ) );
NOR2_X1 _10050_ ( .A1(_02395_ ), .A2(_02398_ ), .ZN(_02399_ ) );
BUF_X4 _10051_ ( .A(_02399_ ), .Z(_02400_ ) );
INV_X1 _10052_ ( .A(\IF_ID_inst [31] ), .ZN(_02401_ ) );
AND2_X2 _10053_ ( .A1(_01342_ ), .A2(_01345_ ), .ZN(_02402_ ) );
INV_X2 _10054_ ( .A(_02402_ ), .ZN(_02403_ ) );
BUF_X4 _10055_ ( .A(_02403_ ), .Z(_02404_ ) );
NOR3_X1 _10056_ ( .A1(_02400_ ), .A2(_02401_ ), .A3(_02404_ ), .ZN(_00163_ ) );
INV_X1 _10057_ ( .A(\IF_ID_inst [30] ), .ZN(_02405_ ) );
NOR3_X1 _10058_ ( .A1(_02400_ ), .A2(_02405_ ), .A3(_02404_ ), .ZN(_00164_ ) );
INV_X1 _10059_ ( .A(\IF_ID_inst [21] ), .ZN(_02406_ ) );
NOR3_X1 _10060_ ( .A1(_02400_ ), .A2(_02406_ ), .A3(_02404_ ), .ZN(_00165_ ) );
BUF_X4 _10061_ ( .A(_02403_ ), .Z(_02407_ ) );
INV_X2 _10062_ ( .A(_02399_ ), .ZN(_02408_ ) );
INV_X1 _10063_ ( .A(\IF_ID_inst [20] ), .ZN(_02409_ ) );
AOI21_X1 _10064_ ( .A(_02407_ ), .B1(_02408_ ), .B2(_02409_ ), .ZN(_00166_ ) );
INV_X1 _10065_ ( .A(\IF_ID_inst [29] ), .ZN(_02410_ ) );
AOI21_X1 _10066_ ( .A(_02407_ ), .B1(_02408_ ), .B2(_02410_ ), .ZN(_00167_ ) );
INV_X1 _10067_ ( .A(\IF_ID_inst [28] ), .ZN(_02411_ ) );
AOI21_X1 _10068_ ( .A(_02407_ ), .B1(_02408_ ), .B2(_02411_ ), .ZN(_00168_ ) );
INV_X1 _10069_ ( .A(\IF_ID_inst [27] ), .ZN(_02412_ ) );
NOR3_X1 _10070_ ( .A1(_02400_ ), .A2(_02412_ ), .A3(_02404_ ), .ZN(_00169_ ) );
INV_X1 _10071_ ( .A(\IF_ID_inst [26] ), .ZN(_02413_ ) );
AOI21_X1 _10072_ ( .A(_02407_ ), .B1(_02408_ ), .B2(_02413_ ), .ZN(_00170_ ) );
INV_X1 _10073_ ( .A(\IF_ID_inst [25] ), .ZN(_02414_ ) );
NOR3_X1 _10074_ ( .A1(_02400_ ), .A2(_02414_ ), .A3(_02404_ ), .ZN(_00171_ ) );
INV_X1 _10075_ ( .A(\IF_ID_inst [24] ), .ZN(_02415_ ) );
NOR3_X1 _10076_ ( .A1(_02400_ ), .A2(_02415_ ), .A3(_02404_ ), .ZN(_00172_ ) );
INV_X1 _10077_ ( .A(\IF_ID_inst [23] ), .ZN(_02416_ ) );
NOR3_X1 _10078_ ( .A1(_02400_ ), .A2(_02416_ ), .A3(_02403_ ), .ZN(_00173_ ) );
INV_X1 _10079_ ( .A(\IF_ID_inst [22] ), .ZN(_02417_ ) );
NOR3_X1 _10080_ ( .A1(_02400_ ), .A2(_02417_ ), .A3(_02403_ ), .ZN(_00174_ ) );
AND3_X1 _10081_ ( .A1(_01342_ ), .A2(_01345_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00175_ ) );
AND3_X1 _10082_ ( .A1(_01342_ ), .A2(_01345_ ), .A3(\myidu.state [2] ), .ZN(_00176_ ) );
INV_X1 _10083_ ( .A(\IF_ID_inst [5] ), .ZN(_02418_ ) );
NOR2_X4 _10084_ ( .A1(_02418_ ), .A2(\IF_ID_inst [4] ), .ZN(_02419_ ) );
NOR2_X1 _10085_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_02420_ ) );
AND3_X1 _10086_ ( .A1(_02387_ ), .A2(_02419_ ), .A3(_02420_ ), .ZN(_02421_ ) );
AND2_X1 _10087_ ( .A1(_02421_ ), .A2(_02391_ ), .ZN(_02422_ ) );
INV_X1 _10088_ ( .A(_02422_ ), .ZN(_02423_ ) );
NOR2_X1 _10089_ ( .A1(\IF_ID_inst [7] ), .A2(\IF_ID_inst [15] ), .ZN(_02424_ ) );
AND4_X1 _10090_ ( .A1(_02385_ ), .A2(_02387_ ), .A3(_02420_ ), .A4(_02424_ ), .ZN(_02425_ ) );
OR3_X1 _10091_ ( .A1(\IF_ID_inst [11] ), .A2(\IF_ID_inst [10] ), .A3(\IF_ID_inst [9] ), .ZN(_02426_ ) );
NOR2_X1 _10092_ ( .A1(_02426_ ), .A2(\IF_ID_inst [8] ), .ZN(_02427_ ) );
AND3_X1 _10093_ ( .A1(_02425_ ), .A2(_02384_ ), .A3(_02427_ ), .ZN(_02428_ ) );
INV_X1 _10094_ ( .A(_02428_ ), .ZN(_02429_ ) );
NOR2_X1 _10095_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [18] ), .ZN(_02430_ ) );
NOR2_X1 _10096_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_02431_ ) );
AND2_X1 _10097_ ( .A1(_02430_ ), .A2(_02431_ ), .ZN(_02432_ ) );
NOR2_X1 _10098_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [31] ), .ZN(_02433_ ) );
AND3_X1 _10099_ ( .A1(_02433_ ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_02434_ ) );
NOR2_X1 _10100_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_02435_ ) );
AND3_X1 _10101_ ( .A1(_02435_ ), .A2(\IF_ID_inst [21] ), .A3(_02409_ ), .ZN(_02436_ ) );
NOR2_X1 _10102_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_02437_ ) );
NOR2_X1 _10103_ ( .A1(\IF_ID_inst [27] ), .A2(\IF_ID_inst [24] ), .ZN(_02438_ ) );
AND2_X1 _10104_ ( .A1(_02437_ ), .A2(_02438_ ), .ZN(_02439_ ) );
AND4_X1 _10105_ ( .A1(_02432_ ), .A2(_02434_ ), .A3(_02436_ ), .A4(_02439_ ), .ZN(_02440_ ) );
INV_X1 _10106_ ( .A(_02440_ ), .ZN(_02441_ ) );
OAI21_X1 _10107_ ( .A(_02423_ ), .B1(_02429_ ), .B2(_02441_ ), .ZN(_02442_ ) );
AND2_X1 _10108_ ( .A1(_02387_ ), .A2(_02419_ ), .ZN(_02443_ ) );
AND2_X1 _10109_ ( .A1(_02443_ ), .A2(_02391_ ), .ZN(_02444_ ) );
AND2_X1 _10110_ ( .A1(_02444_ ), .A2(\IF_ID_inst [14] ), .ZN(_02445_ ) );
AND3_X1 _10111_ ( .A1(_02397_ ), .A2(_02392_ ), .A3(_02419_ ), .ZN(_02446_ ) );
OR2_X1 _10112_ ( .A1(_02445_ ), .A2(_02446_ ), .ZN(_02447_ ) );
AND2_X1 _10113_ ( .A1(_02397_ ), .A2(_02419_ ), .ZN(_02448_ ) );
AOI211_X1 _10114_ ( .A(_02442_ ), .B(_02447_ ), .C1(_02389_ ), .C2(_02448_ ), .ZN(_02449_ ) );
BUF_X2 _10115_ ( .A(_02402_ ), .Z(_02450_ ) );
NOR2_X1 _10116_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_02451_ ) );
AND3_X1 _10117_ ( .A1(_02384_ ), .A2(_02419_ ), .A3(_02451_ ), .ZN(_02452_ ) );
BUF_X2 _10118_ ( .A(_02420_ ), .Z(_02453_ ) );
AND2_X1 _10119_ ( .A1(_02452_ ), .A2(_02453_ ), .ZN(_02454_ ) );
INV_X1 _10120_ ( .A(\IF_ID_inst [12] ), .ZN(_02455_ ) );
NOR2_X1 _10121_ ( .A1(_02455_ ), .A2(\IF_ID_inst [6] ), .ZN(_02456_ ) );
AND3_X1 _10122_ ( .A1(_02384_ ), .A2(_02419_ ), .A3(_02456_ ), .ZN(_02457_ ) );
AND2_X1 _10123_ ( .A1(_02457_ ), .A2(_02420_ ), .ZN(_02458_ ) );
OR2_X1 _10124_ ( .A1(_02454_ ), .A2(_02458_ ), .ZN(_02459_ ) );
AND3_X1 _10125_ ( .A1(_02430_ ), .A2(_02431_ ), .A3(_02435_ ), .ZN(_02460_ ) );
AND3_X1 _10126_ ( .A1(_02460_ ), .A2(_02406_ ), .A3(\IF_ID_inst [20] ), .ZN(_02461_ ) );
NOR4_X1 _10127_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .A4(\IF_ID_inst [31] ), .ZN(_02462_ ) );
AND2_X1 _10128_ ( .A1(_02462_ ), .A2(_02439_ ), .ZN(_02463_ ) );
AND3_X1 _10129_ ( .A1(_02428_ ), .A2(_02461_ ), .A3(_02463_ ), .ZN(_02464_ ) );
AND2_X2 _10130_ ( .A1(_02452_ ), .A2(_02393_ ), .ZN(_02465_ ) );
AND3_X1 _10131_ ( .A1(_02382_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_02466_ ) );
INV_X1 _10132_ ( .A(_02466_ ), .ZN(_02467_ ) );
NOR2_X1 _10133_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_02468_ ) );
NAND4_X1 _10134_ ( .A1(_02453_ ), .A2(_02468_ ), .A3(\IF_ID_inst [12] ), .A4(_02386_ ), .ZN(_02469_ ) );
NOR2_X1 _10135_ ( .A1(_02467_ ), .A2(_02469_ ), .ZN(_02470_ ) );
NOR4_X1 _10136_ ( .A1(_02459_ ), .A2(_02464_ ), .A3(_02465_ ), .A4(_02470_ ), .ZN(_02471_ ) );
AND4_X1 _10137_ ( .A1(\IF_ID_inst [11] ), .A2(_02449_ ), .A3(_02450_ ), .A4(_02471_ ), .ZN(_00177_ ) );
CLKBUF_X2 _10138_ ( .A(_02402_ ), .Z(_02472_ ) );
AND4_X1 _10139_ ( .A1(\IF_ID_inst [10] ), .A2(_02449_ ), .A3(_02472_ ), .A4(_02471_ ), .ZN(_00178_ ) );
AND4_X1 _10140_ ( .A1(\IF_ID_inst [9] ), .A2(_02449_ ), .A3(_02472_ ), .A4(_02471_ ), .ZN(_00179_ ) );
AND4_X1 _10141_ ( .A1(\IF_ID_inst [8] ), .A2(_02449_ ), .A3(_02472_ ), .A4(_02471_ ), .ZN(_00180_ ) );
AND4_X1 _10142_ ( .A1(\IF_ID_inst [7] ), .A2(_02449_ ), .A3(_02472_ ), .A4(_02471_ ), .ZN(_00181_ ) );
INV_X1 _10143_ ( .A(\IF_ID_inst [7] ), .ZN(_02473_ ) );
AND4_X1 _10144_ ( .A1(\IF_ID_inst [6] ), .A2(_02384_ ), .A3(_02473_ ), .A4(_02385_ ), .ZN(_02474_ ) );
NOR4_X1 _10145_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_02475_ ) );
AND3_X1 _10146_ ( .A1(_02474_ ), .A2(_02427_ ), .A3(_02475_ ), .ZN(_02476_ ) );
AND2_X1 _10147_ ( .A1(_02461_ ), .A2(_02463_ ), .ZN(_02477_ ) );
AND2_X1 _10148_ ( .A1(_02476_ ), .A2(_02477_ ), .ZN(_02478_ ) );
AND3_X1 _10149_ ( .A1(_02468_ ), .A2(\IF_ID_inst [12] ), .A3(_02386_ ), .ZN(_02479_ ) );
AND2_X1 _10150_ ( .A1(_02466_ ), .A2(_02479_ ), .ZN(_02480_ ) );
AOI21_X1 _10151_ ( .A(_02478_ ), .B1(_02453_ ), .B2(_02480_ ), .ZN(_02481_ ) );
AND2_X1 _10152_ ( .A1(_02428_ ), .A2(_02440_ ), .ZN(_02482_ ) );
INV_X1 _10153_ ( .A(_02419_ ), .ZN(_02483_ ) );
NOR2_X2 _10154_ ( .A1(_02483_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02484_ ) );
AND2_X2 _10155_ ( .A1(_02484_ ), .A2(_02466_ ), .ZN(_02485_ ) );
CLKBUF_X2 _10156_ ( .A(_02485_ ), .Z(_02486_ ) );
BUF_X2 _10157_ ( .A(_02486_ ), .Z(_02487_ ) );
INV_X1 _10158_ ( .A(\IF_ID_inst [2] ), .ZN(_02488_ ) );
NOR2_X1 _10159_ ( .A1(_02488_ ), .A2(\IF_ID_inst [3] ), .ZN(_02489_ ) );
AND2_X1 _10160_ ( .A1(_02489_ ), .A2(_02382_ ), .ZN(_02490_ ) );
INV_X1 _10161_ ( .A(\IF_ID_inst [4] ), .ZN(_02491_ ) );
NOR2_X1 _10162_ ( .A1(_02491_ ), .A2(\IF_ID_inst [6] ), .ZN(_02492_ ) );
AND2_X2 _10163_ ( .A1(_02490_ ), .A2(_02492_ ), .ZN(_02493_ ) );
NOR3_X1 _10164_ ( .A1(_02482_ ), .A2(_02487_ ), .A3(_02493_ ), .ZN(_02494_ ) );
AND4_X1 _10165_ ( .A1(\IF_ID_inst [19] ), .A2(_02481_ ), .A3(_02472_ ), .A4(_02494_ ), .ZN(_00182_ ) );
AND4_X1 _10166_ ( .A1(\IF_ID_inst [18] ), .A2(_02481_ ), .A3(_02472_ ), .A4(_02494_ ), .ZN(_00183_ ) );
AND4_X1 _10167_ ( .A1(\IF_ID_inst [17] ), .A2(_02481_ ), .A3(_02472_ ), .A4(_02494_ ), .ZN(_00184_ ) );
AND2_X1 _10168_ ( .A1(_02481_ ), .A2(_02494_ ), .ZN(_02495_ ) );
NAND2_X1 _10169_ ( .A1(_02495_ ), .A2(\IF_ID_inst [18] ), .ZN(_02496_ ) );
NOR4_X1 _10170_ ( .A1(\IF_ID_pc [15] ), .A2(\IF_ID_pc [14] ), .A3(\IF_ID_pc [5] ), .A4(\IF_ID_pc [4] ), .ZN(_02497_ ) );
NOR2_X1 _10171_ ( .A1(\IF_ID_pc [0] ), .A2(\IF_ID_pc [1] ), .ZN(_02498_ ) );
NOR2_X1 _10172_ ( .A1(\IF_ID_pc [24] ), .A2(\IF_ID_pc [23] ), .ZN(_02499_ ) );
AND3_X1 _10173_ ( .A1(_02497_ ), .A2(_02498_ ), .A3(_02499_ ), .ZN(_02500_ ) );
NOR4_X1 _10174_ ( .A1(\IF_ID_pc [29] ), .A2(\IF_ID_pc [28] ), .A3(\IF_ID_pc [27] ), .A4(\IF_ID_pc [26] ), .ZN(_02501_ ) );
INV_X1 _10175_ ( .A(\IF_ID_pc [3] ), .ZN(_02502_ ) );
INV_X1 _10176_ ( .A(\IF_ID_pc [2] ), .ZN(_02503_ ) );
AND4_X1 _10177_ ( .A1(_02502_ ), .A2(_02503_ ), .A3(_01049_ ), .A4(\IF_ID_pc [31] ), .ZN(_02504_ ) );
NAND3_X1 _10178_ ( .A1(_02500_ ), .A2(_02501_ ), .A3(_02504_ ), .ZN(_02505_ ) );
INV_X1 _10179_ ( .A(\IF_ID_pc [13] ), .ZN(_02506_ ) );
INV_X1 _10180_ ( .A(\IF_ID_pc [22] ), .ZN(_02507_ ) );
INV_X1 _10181_ ( .A(\IF_ID_pc [20] ), .ZN(_02508_ ) );
NAND4_X1 _10182_ ( .A1(_02506_ ), .A2(_02507_ ), .A3(_01158_ ), .A4(_02508_ ), .ZN(_02509_ ) );
NAND2_X1 _10183_ ( .A1(_01123_ ), .A2(_01034_ ), .ZN(_02510_ ) );
NOR4_X1 _10184_ ( .A1(_02509_ ), .A2(_02510_ ), .A3(\IF_ID_pc [19] ), .A4(\IF_ID_pc [18] ), .ZN(_02511_ ) );
INV_X1 _10185_ ( .A(\IF_ID_pc [12] ), .ZN(_02512_ ) );
INV_X1 _10186_ ( .A(\IF_ID_pc [11] ), .ZN(_02513_ ) );
INV_X1 _10187_ ( .A(\IF_ID_pc [10] ), .ZN(_02514_ ) );
NAND4_X1 _10188_ ( .A1(_01242_ ), .A2(_02512_ ), .A3(_02513_ ), .A4(_02514_ ), .ZN(_02515_ ) );
INV_X1 _10189_ ( .A(\IF_ID_pc [9] ), .ZN(_02516_ ) );
INV_X1 _10190_ ( .A(\IF_ID_pc [6] ), .ZN(_02517_ ) );
NAND2_X1 _10191_ ( .A1(_02516_ ), .A2(_02517_ ), .ZN(_02518_ ) );
NOR4_X1 _10192_ ( .A1(_02515_ ), .A2(_02518_ ), .A3(\IF_ID_pc [8] ), .A4(\IF_ID_pc [7] ), .ZN(_02519_ ) );
NAND2_X1 _10193_ ( .A1(_02511_ ), .A2(_02519_ ), .ZN(_02520_ ) );
NOR2_X1 _10194_ ( .A1(_02505_ ), .A2(_02520_ ), .ZN(_02521_ ) );
NOR2_X2 _10195_ ( .A1(_02521_ ), .A2(_01353_ ), .ZN(_02522_ ) );
INV_X1 _10196_ ( .A(fanout_net_42 ), .ZN(_02523_ ) );
NAND2_X1 _10197_ ( .A1(_02523_ ), .A2(\myifu.state [1] ), .ZN(_02524_ ) );
NOR2_X1 _10198_ ( .A1(_02522_ ), .A2(_02524_ ), .ZN(_02525_ ) );
AND2_X2 _10199_ ( .A1(_02525_ ), .A2(IDU_ready_IFU ), .ZN(_02526_ ) );
AND2_X1 _10200_ ( .A1(_02384_ ), .A2(_02451_ ), .ZN(_02527_ ) );
NOR2_X1 _10201_ ( .A1(_02491_ ), .A2(\IF_ID_inst [5] ), .ZN(_02528_ ) );
AND2_X1 _10202_ ( .A1(_02527_ ), .A2(_02528_ ), .ZN(_02529_ ) );
INV_X1 _10203_ ( .A(_02529_ ), .ZN(_02530_ ) );
INV_X1 _10204_ ( .A(\IF_ID_inst [14] ), .ZN(_02531_ ) );
AOI21_X1 _10205_ ( .A(_02530_ ), .B1(\IF_ID_inst [13] ), .B2(_02531_ ), .ZN(_02532_ ) );
AND3_X1 _10206_ ( .A1(_02528_ ), .A2(_02382_ ), .A3(_02383_ ), .ZN(_02533_ ) );
AND2_X2 _10207_ ( .A1(_02533_ ), .A2(_02456_ ), .ZN(_02534_ ) );
AOI21_X1 _10208_ ( .A(_02532_ ), .B1(_02389_ ), .B2(_02534_ ), .ZN(_02535_ ) );
AND2_X1 _10209_ ( .A1(_02527_ ), .A2(_02385_ ), .ZN(_02536_ ) );
INV_X1 _10210_ ( .A(_02536_ ), .ZN(_02537_ ) );
NAND3_X1 _10211_ ( .A1(_02411_ ), .A2(_02412_ ), .A3(\IF_ID_inst [30] ), .ZN(_02538_ ) );
INV_X1 _10212_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02539_ ) );
NOR3_X1 _10213_ ( .A1(_02538_ ), .A2(\IF_ID_inst [29] ), .A3(_02539_ ), .ZN(_02540_ ) );
AND2_X2 _10214_ ( .A1(_02453_ ), .A2(_02437_ ), .ZN(_02541_ ) );
NOR3_X1 _10215_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_02542_ ) );
AND2_X2 _10216_ ( .A1(_02542_ ), .A2(_02412_ ), .ZN(_02543_ ) );
AND4_X1 _10217_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02437_ ), .A3(\IF_ID_inst [13] ), .A4(_02531_ ), .ZN(_02544_ ) );
AOI22_X1 _10218_ ( .A1(_02540_ ), .A2(_02541_ ), .B1(_02543_ ), .B2(_02544_ ), .ZN(_02545_ ) );
OR2_X1 _10219_ ( .A1(_02537_ ), .A2(_02545_ ), .ZN(_02546_ ) );
NOR2_X1 _10220_ ( .A1(_02531_ ), .A2(\IF_ID_inst [13] ), .ZN(_02547_ ) );
AND2_X1 _10221_ ( .A1(_02547_ ), .A2(_02437_ ), .ZN(_02548_ ) );
AND2_X2 _10222_ ( .A1(_02540_ ), .A2(_02548_ ), .ZN(_02549_ ) );
AND4_X1 _10223_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A2(_02437_ ), .A3(_02392_ ), .A4(\IF_ID_inst [14] ), .ZN(_02550_ ) );
AND2_X1 _10224_ ( .A1(_02543_ ), .A2(_02550_ ), .ZN(_02551_ ) );
OAI21_X1 _10225_ ( .A(_02534_ ), .B1(_02549_ ), .B2(_02551_ ), .ZN(_02552_ ) );
AND3_X1 _10226_ ( .A1(_02535_ ), .A2(_02546_ ), .A3(_02552_ ), .ZN(_02553_ ) );
AND4_X1 _10227_ ( .A1(\IF_ID_inst [4] ), .A2(_02386_ ), .A3(\IF_ID_inst [5] ), .A4(\IF_ID_inst [12] ), .ZN(_02554_ ) );
AND2_X2 _10228_ ( .A1(_02391_ ), .A2(_02554_ ), .ZN(_02555_ ) );
AND2_X1 _10229_ ( .A1(_02543_ ), .A2(_02544_ ), .ZN(_02556_ ) );
OR2_X1 _10230_ ( .A1(_02556_ ), .A2(_02551_ ), .ZN(_02557_ ) );
AND3_X1 _10231_ ( .A1(_02420_ ), .A2(_02437_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02558_ ) );
AND2_X1 _10232_ ( .A1(_02543_ ), .A2(_02558_ ), .ZN(_02559_ ) );
OAI21_X1 _10233_ ( .A(_02555_ ), .B1(_02557_ ), .B2(_02559_ ), .ZN(_02560_ ) );
BUF_X2 _10234_ ( .A(_02385_ ), .Z(_02561_ ) );
BUF_X2 _10235_ ( .A(_02527_ ), .Z(_02562_ ) );
OAI211_X1 _10236_ ( .A(_02561_ ), .B(_02562_ ), .C1(_02559_ ), .C2(_02551_ ), .ZN(_02563_ ) );
NAND2_X1 _10237_ ( .A1(_02560_ ), .A2(_02563_ ), .ZN(_02564_ ) );
AND2_X1 _10238_ ( .A1(_02549_ ), .A2(_02555_ ), .ZN(_02565_ ) );
AND3_X1 _10239_ ( .A1(_02543_ ), .A2(_02389_ ), .A3(_02437_ ), .ZN(_02566_ ) );
NAND3_X1 _10240_ ( .A1(_02536_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02566_ ), .ZN(_02567_ ) );
NAND3_X1 _10241_ ( .A1(_02566_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02555_ ), .ZN(_02568_ ) );
NAND2_X1 _10242_ ( .A1(_02567_ ), .A2(_02568_ ), .ZN(_02569_ ) );
NOR3_X1 _10243_ ( .A1(_02564_ ), .A2(_02565_ ), .A3(_02569_ ), .ZN(_02570_ ) );
OAI21_X1 _10244_ ( .A(_02393_ ), .B1(_02529_ ), .B2(_02534_ ), .ZN(_02571_ ) );
AND3_X1 _10245_ ( .A1(_02391_ ), .A2(_02451_ ), .A3(_02468_ ), .ZN(_02572_ ) );
NAND2_X1 _10246_ ( .A1(_02572_ ), .A2(_02393_ ), .ZN(_02573_ ) );
AND3_X1 _10247_ ( .A1(_02571_ ), .A2(_02423_ ), .A3(_02573_ ), .ZN(_02574_ ) );
NAND4_X1 _10248_ ( .A1(_02553_ ), .A2(_02495_ ), .A3(_02570_ ), .A4(_02574_ ), .ZN(_02575_ ) );
NOR2_X1 _10249_ ( .A1(_02459_ ), .A2(_02465_ ), .ZN(_02576_ ) );
INV_X1 _10250_ ( .A(_02576_ ), .ZN(_02577_ ) );
OAI21_X1 _10251_ ( .A(_02572_ ), .B1(_02453_ ), .B2(_02547_ ), .ZN(_02578_ ) );
AND2_X1 _10252_ ( .A1(_02479_ ), .A2(_02391_ ), .ZN(_02579_ ) );
NAND2_X1 _10253_ ( .A1(_02579_ ), .A2(_02392_ ), .ZN(_02580_ ) );
NAND2_X1 _10254_ ( .A1(_02578_ ), .A2(_02580_ ), .ZN(_02581_ ) );
INV_X1 _10255_ ( .A(_02581_ ), .ZN(_02582_ ) );
NAND3_X1 _10256_ ( .A1(_02397_ ), .A2(_02389_ ), .A3(_02419_ ), .ZN(_02583_ ) );
AND2_X1 _10257_ ( .A1(_02421_ ), .A2(_02490_ ), .ZN(_02584_ ) );
INV_X1 _10258_ ( .A(_02584_ ), .ZN(_02585_ ) );
NAND2_X1 _10259_ ( .A1(_02534_ ), .A2(_02559_ ), .ZN(_02586_ ) );
NAND4_X1 _10260_ ( .A1(_02582_ ), .A2(_02583_ ), .A3(_02585_ ), .A4(_02586_ ), .ZN(_02587_ ) );
OR4_X2 _10261_ ( .A1(_02408_ ), .A2(_02577_ ), .A3(_02447_ ), .A4(_02587_ ), .ZN(_02588_ ) );
OAI211_X1 _10262_ ( .A(_02496_ ), .B(_02526_ ), .C1(_02575_ ), .C2(_02588_ ), .ZN(_02589_ ) );
INV_X1 _10263_ ( .A(_02589_ ), .ZN(_02590_ ) );
NOR2_X2 _10264_ ( .A1(_02575_ ), .A2(_02588_ ), .ZN(_02591_ ) );
INV_X1 _10265_ ( .A(_02526_ ), .ZN(_02592_ ) );
NOR2_X1 _10266_ ( .A1(_02591_ ), .A2(_02592_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _10267_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_02593_ ) );
AOI211_X1 _10268_ ( .A(_02403_ ), .B(_02590_ ), .C1(_02593_ ), .C2(_01392_ ), .ZN(_00185_ ) );
AND4_X1 _10269_ ( .A1(\IF_ID_inst [16] ), .A2(_02481_ ), .A3(_02472_ ), .A4(_02494_ ), .ZN(_00186_ ) );
OAI21_X1 _10270_ ( .A(_02450_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [2] ), .ZN(_02594_ ) );
INV_X1 _10271_ ( .A(\IF_ID_inst [17] ), .ZN(_02595_ ) );
INV_X1 _10272_ ( .A(_02495_ ), .ZN(_02596_ ) );
OAI221_X1 _10273_ ( .A(_02526_ ), .B1(_02595_ ), .B2(_02596_ ), .C1(_02575_ ), .C2(_02588_ ), .ZN(_02597_ ) );
INV_X1 _10274_ ( .A(_02597_ ), .ZN(_02598_ ) );
NOR2_X1 _10275_ ( .A1(_02594_ ), .A2(_02598_ ), .ZN(_00187_ ) );
AND4_X1 _10276_ ( .A1(\IF_ID_inst [15] ), .A2(_02481_ ), .A3(_02472_ ), .A4(_02494_ ), .ZN(_00188_ ) );
INV_X1 _10277_ ( .A(_02591_ ), .ZN(_02599_ ) );
AOI21_X1 _10278_ ( .A(\ID_EX_rs1 [1] ), .B1(_02599_ ), .B2(_02526_ ), .ZN(_02600_ ) );
NAND2_X1 _10279_ ( .A1(_02495_ ), .A2(\IF_ID_inst [16] ), .ZN(_02601_ ) );
AOI211_X1 _10280_ ( .A(_02403_ ), .B(_02600_ ), .C1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .C2(_02601_ ), .ZN(_00189_ ) );
AND3_X1 _10281_ ( .A1(_02533_ ), .A2(\IF_ID_inst [13] ), .A3(_02456_ ), .ZN(_02602_ ) );
OR2_X1 _10282_ ( .A1(_02532_ ), .A2(_02602_ ), .ZN(_02603_ ) );
AND2_X1 _10283_ ( .A1(_02562_ ), .A2(_02468_ ), .ZN(_02604_ ) );
AND2_X1 _10284_ ( .A1(_02604_ ), .A2(_02393_ ), .ZN(_02605_ ) );
OR3_X1 _10285_ ( .A1(_02605_ ), .A2(_02581_ ), .A3(_02584_ ), .ZN(_02606_ ) );
NOR2_X1 _10286_ ( .A1(_02464_ ), .A2(_02487_ ), .ZN(_02607_ ) );
INV_X1 _10287_ ( .A(_02607_ ), .ZN(_02608_ ) );
INV_X1 _10288_ ( .A(_02482_ ), .ZN(_02609_ ) );
INV_X1 _10289_ ( .A(_02470_ ), .ZN(_02610_ ) );
NAND3_X1 _10290_ ( .A1(_02609_ ), .A2(_02399_ ), .A3(_02610_ ), .ZN(_02611_ ) );
NOR4_X1 _10291_ ( .A1(_02603_ ), .A2(_02606_ ), .A3(_02608_ ), .A4(_02611_ ), .ZN(_02612_ ) );
AND2_X1 _10292_ ( .A1(_02529_ ), .A2(_02393_ ), .ZN(_02613_ ) );
NOR2_X1 _10293_ ( .A1(_02613_ ), .A2(_02493_ ), .ZN(_02614_ ) );
AND4_X1 _10294_ ( .A1(\IF_ID_inst [4] ), .A2(_02418_ ), .A3(_02386_ ), .A4(\IF_ID_inst [12] ), .ZN(_02615_ ) );
AND2_X1 _10295_ ( .A1(_02391_ ), .A2(_02615_ ), .ZN(_02616_ ) );
AND3_X1 _10296_ ( .A1(_02542_ ), .A2(_02412_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02617_ ) );
AND2_X1 _10297_ ( .A1(_02617_ ), .A2(_02548_ ), .ZN(_02618_ ) );
OAI21_X1 _10298_ ( .A(_02616_ ), .B1(_02618_ ), .B2(_02549_ ), .ZN(_02619_ ) );
NAND3_X1 _10299_ ( .A1(_02616_ ), .A2(_02617_ ), .A3(_02541_ ), .ZN(_02620_ ) );
AND2_X1 _10300_ ( .A1(_02619_ ), .A2(_02620_ ), .ZN(_02621_ ) );
AND2_X2 _10301_ ( .A1(_02614_ ), .A2(_02621_ ), .ZN(_02622_ ) );
AND4_X1 _10302_ ( .A1(\IF_ID_inst [24] ), .A2(_02612_ ), .A3(_02472_ ), .A4(_02622_ ), .ZN(_00190_ ) );
OAI21_X1 _10303_ ( .A(_02450_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [0] ), .ZN(_02623_ ) );
INV_X1 _10304_ ( .A(\IF_ID_inst [15] ), .ZN(_02624_ ) );
OAI221_X1 _10305_ ( .A(_02526_ ), .B1(_02624_ ), .B2(_02596_ ), .C1(_02575_ ), .C2(_02588_ ), .ZN(_02625_ ) );
INV_X1 _10306_ ( .A(_02625_ ), .ZN(_02626_ ) );
NOR2_X1 _10307_ ( .A1(_02623_ ), .A2(_02626_ ), .ZN(_00191_ ) );
AND4_X1 _10308_ ( .A1(\IF_ID_inst [23] ), .A2(_02612_ ), .A3(_02402_ ), .A4(_02622_ ), .ZN(_00192_ ) );
AND4_X1 _10309_ ( .A1(\IF_ID_inst [22] ), .A2(_02612_ ), .A3(_02402_ ), .A4(_02622_ ), .ZN(_00193_ ) );
AND2_X1 _10310_ ( .A1(_02612_ ), .A2(_02622_ ), .ZN(_02627_ ) );
AOI211_X1 _10311_ ( .A(_02592_ ), .B(_02591_ ), .C1(\IF_ID_inst [23] ), .C2(_02627_ ), .ZN(_02628_ ) );
INV_X16 _10312_ ( .A(\ID_EX_rs2 [3] ), .ZN(_02629_ ) );
AOI211_X1 _10313_ ( .A(_02403_ ), .B(_02628_ ), .C1(_02629_ ), .C2(_02593_ ), .ZN(_00194_ ) );
AND4_X1 _10314_ ( .A1(\IF_ID_inst [21] ), .A2(_02612_ ), .A3(_02402_ ), .A4(_02622_ ), .ZN(_00195_ ) );
NAND4_X1 _10315_ ( .A1(_02599_ ), .A2(\IF_ID_inst [22] ), .A3(_02526_ ), .A4(_02627_ ), .ZN(_02630_ ) );
OAI21_X1 _10316_ ( .A(\ID_EX_rs2 [2] ), .B1(_02591_ ), .B2(_02592_ ), .ZN(_02631_ ) );
AOI21_X1 _10317_ ( .A(_02407_ ), .B1(_02630_ ), .B2(_02631_ ), .ZN(_00196_ ) );
AND4_X1 _10318_ ( .A1(\IF_ID_inst [20] ), .A2(_02612_ ), .A3(_02402_ ), .A4(_02622_ ), .ZN(_00197_ ) );
NAND4_X1 _10319_ ( .A1(_02599_ ), .A2(\IF_ID_inst [21] ), .A3(_02526_ ), .A4(_02627_ ), .ZN(_02632_ ) );
OAI21_X1 _10320_ ( .A(\ID_EX_rs2 [1] ), .B1(_02591_ ), .B2(_02592_ ), .ZN(_02633_ ) );
AOI21_X1 _10321_ ( .A(_02407_ ), .B1(_02632_ ), .B2(_02633_ ), .ZN(_00198_ ) );
NOR4_X1 _10322_ ( .A1(_02467_ ), .A2(_02403_ ), .A3(IDU_valid_EXU ), .A4(_02469_ ), .ZN(_00199_ ) );
AOI211_X1 _10323_ ( .A(_02592_ ), .B(_02591_ ), .C1(\IF_ID_inst [20] ), .C2(_02627_ ), .ZN(_02634_ ) );
OAI21_X1 _10324_ ( .A(_02450_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs2 [0] ), .ZN(_02635_ ) );
NOR2_X1 _10325_ ( .A1(_02634_ ), .A2(_02635_ ), .ZN(_00200_ ) );
NAND3_X1 _10326_ ( .A1(_02535_ ), .A2(_02578_ ), .A3(_02571_ ), .ZN(_02636_ ) );
AND4_X1 _10327_ ( .A1(_02382_ ), .A2(_02387_ ), .A3(_02419_ ), .A4(_02489_ ), .ZN(_02637_ ) );
NAND2_X1 _10328_ ( .A1(_02637_ ), .A2(_02453_ ), .ZN(_02638_ ) );
NAND3_X1 _10329_ ( .A1(_02573_ ), .A2(_02580_ ), .A3(_02638_ ), .ZN(_02639_ ) );
NOR2_X1 _10330_ ( .A1(_02636_ ), .A2(_02639_ ), .ZN(_02640_ ) );
BUF_X4 _10331_ ( .A(_02640_ ), .Z(_02641_ ) );
XNOR2_X1 _10332_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_02642_ ) );
XNOR2_X1 _10333_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_02643_ ) );
XNOR2_X1 _10334_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_02644_ ) );
XNOR2_X1 _10335_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_02645_ ) );
NAND4_X1 _10336_ ( .A1(_02642_ ), .A2(_02643_ ), .A3(_02644_ ), .A4(_02645_ ), .ZN(_02646_ ) );
XOR2_X1 _10337_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .Z(_02647_ ) );
NOR2_X1 _10338_ ( .A1(_02646_ ), .A2(_02647_ ), .ZN(_02648_ ) );
AND2_X1 _10339_ ( .A1(_01366_ ), .A2(_01355_ ), .ZN(_02649_ ) );
AND2_X1 _10340_ ( .A1(_02648_ ), .A2(_02649_ ), .ZN(_02650_ ) );
INV_X1 _10341_ ( .A(_02650_ ), .ZN(_02651_ ) );
XNOR2_X1 _10342_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_02652_ ) );
XNOR2_X1 _10343_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_02653_ ) );
XNOR2_X1 _10344_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_02654_ ) );
AND4_X1 _10345_ ( .A1(_02649_ ), .A2(_02652_ ), .A3(_02653_ ), .A4(_02654_ ), .ZN(_02655_ ) );
XNOR2_X1 _10346_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_02656_ ) );
XNOR2_X1 _10347_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_02657_ ) );
NAND3_X1 _10348_ ( .A1(_02655_ ), .A2(_02656_ ), .A3(_02657_ ), .ZN(_02658_ ) );
AND2_X1 _10349_ ( .A1(_02651_ ), .A2(_02658_ ), .ZN(_02659_ ) );
OAI211_X1 _10350_ ( .A(_02399_ ), .B(_02641_ ), .C1(_02596_ ), .C2(_02659_ ), .ZN(_02660_ ) );
NAND3_X1 _10351_ ( .A1(_02660_ ), .A2(IDU_ready_IFU ), .A3(_02450_ ), .ZN(_02661_ ) );
AOI21_X1 _10352_ ( .A(_02650_ ), .B1(_02641_ ), .B2(_02399_ ), .ZN(_02662_ ) );
NOR2_X1 _10353_ ( .A1(_02661_ ), .A2(_02662_ ), .ZN(_00201_ ) );
AND4_X1 _10354_ ( .A1(_02561_ ), .A2(_02387_ ), .A3(_02453_ ), .A4(_02424_ ), .ZN(_02663_ ) );
AND3_X1 _10355_ ( .A1(_02663_ ), .A2(_02391_ ), .A3(_02427_ ), .ZN(_02664_ ) );
AND4_X1 _10356_ ( .A1(_02432_ ), .A2(_02434_ ), .A3(_02436_ ), .A4(_02439_ ), .ZN(_02665_ ) );
AND2_X1 _10357_ ( .A1(_02664_ ), .A2(_02665_ ), .ZN(_02666_ ) );
NOR2_X1 _10358_ ( .A1(_02666_ ), .A2(_02470_ ), .ZN(_02667_ ) );
AND3_X1 _10359_ ( .A1(_02460_ ), .A2(_02406_ ), .A3(_02409_ ), .ZN(_02668_ ) );
NAND3_X1 _10360_ ( .A1(_02664_ ), .A2(_02463_ ), .A3(_02668_ ), .ZN(_02669_ ) );
AND2_X1 _10361_ ( .A1(_02399_ ), .A2(_02669_ ), .ZN(_02670_ ) );
INV_X1 _10362_ ( .A(_02487_ ), .ZN(_02671_ ) );
AND4_X1 _10363_ ( .A1(_02667_ ), .A2(_02670_ ), .A3(_02671_ ), .A4(_02585_ ), .ZN(_02672_ ) );
OAI21_X1 _10364_ ( .A(\IF_ID_inst [14] ), .B1(_02444_ ), .B2(_02448_ ), .ZN(_02673_ ) );
AND3_X1 _10365_ ( .A1(_02397_ ), .A2(_02453_ ), .A3(_02419_ ), .ZN(_02674_ ) );
NOR2_X1 _10366_ ( .A1(_02422_ ), .A2(_02674_ ), .ZN(_02675_ ) );
AND2_X1 _10367_ ( .A1(_02673_ ), .A2(_02675_ ), .ZN(_02676_ ) );
AOI21_X1 _10368_ ( .A(_02407_ ), .B1(_02672_ ), .B2(_02676_ ), .ZN(_00202_ ) );
AND3_X1 _10369_ ( .A1(_02479_ ), .A2(_02391_ ), .A3(_02453_ ), .ZN(_02677_ ) );
AND2_X1 _10370_ ( .A1(_02572_ ), .A2(_02547_ ), .ZN(_02678_ ) );
AOI211_X1 _10371_ ( .A(_02677_ ), .B(_02678_ ), .C1(_02453_ ), .C2(_02572_ ), .ZN(_02679_ ) );
NAND2_X1 _10372_ ( .A1(_02579_ ), .A2(_02547_ ), .ZN(_02680_ ) );
AND4_X1 _10373_ ( .A1(_02576_ ), .A2(_02679_ ), .A3(_02680_ ), .A4(_02573_ ), .ZN(_02681_ ) );
AOI21_X1 _10374_ ( .A(_02407_ ), .B1(_02681_ ), .B2(_02670_ ), .ZN(_00203_ ) );
AND3_X1 _10375_ ( .A1(_02389_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02437_ ), .ZN(_02682_ ) );
NAND3_X1 _10376_ ( .A1(_02536_ ), .A2(_02543_ ), .A3(_02682_ ), .ZN(_02683_ ) );
AND3_X1 _10377_ ( .A1(_02555_ ), .A2(_02543_ ), .A3(_02682_ ), .ZN(_02684_ ) );
INV_X1 _10378_ ( .A(_02684_ ), .ZN(_02685_ ) );
NAND4_X1 _10379_ ( .A1(_02562_ ), .A2(_02561_ ), .A3(_02617_ ), .A4(_02541_ ), .ZN(_02686_ ) );
NAND3_X1 _10380_ ( .A1(_02618_ ), .A2(_02561_ ), .A3(_02562_ ), .ZN(_02687_ ) );
NAND4_X1 _10381_ ( .A1(_02683_ ), .A2(_02685_ ), .A3(_02686_ ), .A4(_02687_ ), .ZN(_02688_ ) );
INV_X1 _10382_ ( .A(_02555_ ), .ZN(_02689_ ) );
INV_X1 _10383_ ( .A(_02618_ ), .ZN(_02690_ ) );
AOI22_X1 _10384_ ( .A1(_02617_ ), .A2(_02541_ ), .B1(_02543_ ), .B2(_02544_ ), .ZN(_02691_ ) );
AOI21_X1 _10385_ ( .A(_02689_ ), .B1(_02690_ ), .B2(_02691_ ), .ZN(_02692_ ) );
NOR2_X1 _10386_ ( .A1(_02688_ ), .A2(_02692_ ), .ZN(_02693_ ) );
AOI21_X1 _10387_ ( .A(_02565_ ), .B1(_02393_ ), .B2(_02604_ ), .ZN(_02694_ ) );
NAND2_X1 _10388_ ( .A1(_02694_ ), .A2(_02669_ ), .ZN(_02695_ ) );
NOR4_X1 _10389_ ( .A1(_02603_ ), .A2(_02487_ ), .A3(_02695_ ), .A4(_02584_ ), .ZN(_02696_ ) );
NAND3_X1 _10390_ ( .A1(_02556_ ), .A2(_02561_ ), .A3(_02562_ ), .ZN(_02697_ ) );
NAND4_X1 _10391_ ( .A1(_02562_ ), .A2(_02561_ ), .A3(_02540_ ), .A4(_02541_ ), .ZN(_02698_ ) );
AND2_X1 _10392_ ( .A1(_02697_ ), .A2(_02698_ ), .ZN(_02699_ ) );
AND4_X1 _10393_ ( .A1(_02693_ ), .A2(_02696_ ), .A3(_02582_ ), .A4(_02699_ ), .ZN(_02700_ ) );
AOI21_X1 _10394_ ( .A(_02407_ ), .B1(_02700_ ), .B2(_02622_ ), .ZN(_00204_ ) );
NOR3_X1 _10395_ ( .A1(_02532_ ), .A2(_02470_ ), .A3(_02602_ ), .ZN(_02701_ ) );
AOI21_X1 _10396_ ( .A(_02407_ ), .B1(_02622_ ), .B2(_02701_ ), .ZN(_00205_ ) );
AND3_X1 _10397_ ( .A1(_02556_ ), .A2(_02561_ ), .A3(_02562_ ), .ZN(_02702_ ) );
AND4_X1 _10398_ ( .A1(_02561_ ), .A2(_02562_ ), .A3(_02540_ ), .A4(_02541_ ), .ZN(_02703_ ) );
NOR4_X1 _10399_ ( .A1(_02666_ ), .A2(_02702_ ), .A3(_02703_ ), .A4(_02465_ ), .ZN(_02704_ ) );
AOI21_X1 _10400_ ( .A(_02404_ ), .B1(_02704_ ), .B2(_02614_ ), .ZN(_00206_ ) );
INV_X1 _10401_ ( .A(_02493_ ), .ZN(_02705_ ) );
NAND2_X1 _10402_ ( .A1(_02549_ ), .A2(_02534_ ), .ZN(_02706_ ) );
NAND4_X1 _10403_ ( .A1(_02533_ ), .A2(_02543_ ), .A3(_02550_ ), .A4(_02456_ ), .ZN(_02707_ ) );
NAND3_X1 _10404_ ( .A1(_02706_ ), .A2(_02586_ ), .A3(_02707_ ), .ZN(_02708_ ) );
AOI221_X4 _10405_ ( .A(_02708_ ), .B1(\IF_ID_inst [13] ), .B2(_02398_ ), .C1(\IF_ID_inst [14] ), .C2(_02448_ ), .ZN(_02709_ ) );
OAI21_X1 _10406_ ( .A(_02393_ ), .B1(_02604_ ), .B2(_02534_ ), .ZN(_02710_ ) );
INV_X1 _10407_ ( .A(_02565_ ), .ZN(_02711_ ) );
AND2_X1 _10408_ ( .A1(_02560_ ), .A2(_02711_ ), .ZN(_02712_ ) );
AND4_X1 _10409_ ( .A1(_02705_ ), .A2(_02709_ ), .A3(_02710_ ), .A4(_02712_ ), .ZN(_02713_ ) );
INV_X1 _10410_ ( .A(_02465_ ), .ZN(_02714_ ) );
AOI21_X1 _10411_ ( .A(_02404_ ), .B1(_02713_ ), .B2(_02714_ ), .ZN(_00207_ ) );
NOR2_X1 _10412_ ( .A1(_02445_ ), .A2(_02395_ ), .ZN(_02715_ ) );
NAND2_X1 _10413_ ( .A1(_02529_ ), .A2(\IF_ID_inst [14] ), .ZN(_02716_ ) );
AND4_X1 _10414_ ( .A1(_02714_ ), .A2(_02715_ ), .A3(_02683_ ), .A4(_02716_ ), .ZN(_02717_ ) );
AND3_X1 _10415_ ( .A1(_02386_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_02718_ ) );
AOI21_X1 _10416_ ( .A(_02458_ ), .B1(_02490_ ), .B2(_02718_ ), .ZN(_02719_ ) );
AND4_X1 _10417_ ( .A1(_02687_ ), .A2(_02717_ ), .A3(_02580_ ), .A4(_02719_ ), .ZN(_02720_ ) );
OAI22_X1 _10418_ ( .A1(_02618_ ), .A2(_02549_ ), .B1(_02555_ ), .B2(_02616_ ), .ZN(_02721_ ) );
AOI21_X1 _10419_ ( .A(_02404_ ), .B1(_02720_ ), .B2(_02721_ ), .ZN(_00208_ ) );
AOI22_X1 _10420_ ( .A1(_02536_ ), .A2(_02556_ ), .B1(_02534_ ), .B2(_02559_ ), .ZN(_02722_ ) );
NAND3_X1 _10421_ ( .A1(_02533_ ), .A2(_02389_ ), .A3(_02456_ ), .ZN(_02723_ ) );
OAI21_X1 _10422_ ( .A(_02389_ ), .B1(_02444_ ), .B2(_02398_ ), .ZN(_02724_ ) );
OAI21_X1 _10423_ ( .A(_02555_ ), .B1(_02549_ ), .B2(_02559_ ), .ZN(_02725_ ) );
NAND4_X1 _10424_ ( .A1(_02722_ ), .A2(_02723_ ), .A3(_02724_ ), .A4(_02725_ ), .ZN(_02726_ ) );
NAND2_X1 _10425_ ( .A1(_02529_ ), .A2(_02547_ ), .ZN(_02727_ ) );
NAND3_X1 _10426_ ( .A1(_02551_ ), .A2(_02561_ ), .A3(_02562_ ), .ZN(_02728_ ) );
NAND3_X1 _10427_ ( .A1(_02727_ ), .A2(_02568_ ), .A3(_02728_ ), .ZN(_02729_ ) );
OR2_X1 _10428_ ( .A1(_02465_ ), .A2(_02674_ ), .ZN(_02730_ ) );
NAND3_X1 _10429_ ( .A1(_02562_ ), .A2(_02547_ ), .A3(_02468_ ), .ZN(_02731_ ) );
NAND3_X1 _10430_ ( .A1(_02397_ ), .A2(_02561_ ), .A3(_02547_ ), .ZN(_02732_ ) );
NAND4_X1 _10431_ ( .A1(_02731_ ), .A2(_02390_ ), .A3(_02732_ ), .A4(_02680_ ), .ZN(_02733_ ) );
NOR4_X1 _10432_ ( .A1(_02726_ ), .A2(_02729_ ), .A3(_02730_ ), .A4(_02733_ ), .ZN(_02734_ ) );
INV_X1 _10433_ ( .A(_02459_ ), .ZN(_02735_ ) );
AND2_X1 _10434_ ( .A1(_02549_ ), .A2(_02534_ ), .ZN(_02736_ ) );
AND4_X1 _10435_ ( .A1(_02391_ ), .A2(_02461_ ), .A3(_02427_ ), .A4(_02425_ ), .ZN(_02737_ ) );
AOI21_X1 _10436_ ( .A(_02736_ ), .B1(_02737_ ), .B2(_02463_ ), .ZN(_02738_ ) );
AND4_X1 _10437_ ( .A1(_02735_ ), .A2(_02583_ ), .A3(_02585_ ), .A4(_02738_ ), .ZN(_02739_ ) );
AOI21_X1 _10438_ ( .A(_02404_ ), .B1(_02734_ ), .B2(_02739_ ), .ZN(_00209_ ) );
NOR2_X1 _10439_ ( .A1(_02522_ ), .A2(fanout_net_42 ), .ZN(_02740_ ) );
BUF_X4 _10440_ ( .A(_02740_ ), .Z(_02741_ ) );
NOR4_X1 _10441_ ( .A1(_02401_ ), .A2(_02418_ ), .A3(\IF_ID_inst [4] ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02742_ ) );
AND2_X2 _10442_ ( .A1(_02742_ ), .A2(_02384_ ), .ZN(_02743_ ) );
AOI21_X1 _10443_ ( .A(_02743_ ), .B1(_02486_ ), .B2(\IF_ID_inst [31] ), .ZN(_02744_ ) );
AND2_X2 _10444_ ( .A1(_02743_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02745_ ) );
OR3_X1 _10445_ ( .A1(_02744_ ), .A2(_01257_ ), .A3(_02745_ ), .ZN(_02746_ ) );
NOR2_X2 _10446_ ( .A1(_02744_ ), .A2(_02745_ ), .ZN(_02747_ ) );
XNOR2_X1 _10447_ ( .A(_02747_ ), .B(\IF_ID_pc [24] ), .ZN(_02748_ ) );
INV_X1 _10448_ ( .A(_02748_ ), .ZN(_02749_ ) );
AND2_X1 _10449_ ( .A1(_02485_ ), .A2(\IF_ID_inst [26] ), .ZN(_02750_ ) );
INV_X1 _10450_ ( .A(_02750_ ), .ZN(_02751_ ) );
AND2_X1 _10451_ ( .A1(_02484_ ), .A2(_02384_ ), .ZN(_02752_ ) );
NAND2_X2 _10452_ ( .A1(_02752_ ), .A2(\IF_ID_inst [31] ), .ZN(_02753_ ) );
MUX2_X1 _10453_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B(_02751_ ), .S(_02753_ ), .Z(_02754_ ) );
NOR2_X1 _10454_ ( .A1(_02754_ ), .A2(_02517_ ), .ZN(_02755_ ) );
INV_X1 _10455_ ( .A(_02755_ ), .ZN(_02756_ ) );
AND2_X4 _10456_ ( .A1(_02485_ ), .A2(\IF_ID_inst [21] ), .ZN(_02757_ ) );
INV_X1 _10457_ ( .A(_02757_ ), .ZN(_02758_ ) );
MUX2_X1 _10458_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B(_02758_ ), .S(_02753_ ), .Z(_02759_ ) );
INV_X2 _10459_ ( .A(_02759_ ), .ZN(_02760_ ) );
AND3_X1 _10460_ ( .A1(_02484_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .A3(_02466_ ), .ZN(_02761_ ) );
AND3_X1 _10461_ ( .A1(_02742_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02384_ ), .ZN(_02762_ ) );
OR3_X1 _10462_ ( .A1(_02761_ ), .A2(_02503_ ), .A3(_02762_ ), .ZN(_02763_ ) );
OAI21_X1 _10463_ ( .A(_02503_ ), .B1(_02761_ ), .B2(_02762_ ), .ZN(_02764_ ) );
AND2_X1 _10464_ ( .A1(_02763_ ), .A2(_02764_ ), .ZN(_02765_ ) );
NAND3_X1 _10465_ ( .A1(_02760_ ), .A2(\IF_ID_pc [1] ), .A3(_02765_ ), .ZN(_02766_ ) );
NAND2_X1 _10466_ ( .A1(_02766_ ), .A2(_02763_ ), .ZN(_02767_ ) );
AND2_X1 _10467_ ( .A1(_02485_ ), .A2(\IF_ID_inst [23] ), .ZN(_02768_ ) );
INV_X1 _10468_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_02769_ ) );
AOI21_X1 _10469_ ( .A(_02768_ ), .B1(_02769_ ), .B2(_02743_ ), .ZN(_02770_ ) );
XNOR2_X1 _10470_ ( .A(_02770_ ), .B(\IF_ID_pc [3] ), .ZN(_02771_ ) );
NAND2_X1 _10471_ ( .A1(_02767_ ), .A2(_02771_ ), .ZN(_02772_ ) );
OR2_X1 _10472_ ( .A1(_02770_ ), .A2(_02502_ ), .ZN(_02773_ ) );
INV_X1 _10473_ ( .A(\IF_ID_pc [4] ), .ZN(_02774_ ) );
AND2_X1 _10474_ ( .A1(_02485_ ), .A2(\IF_ID_inst [24] ), .ZN(_02775_ ) );
INV_X1 _10475_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_02776_ ) );
AOI21_X1 _10476_ ( .A(_02775_ ), .B1(_02776_ ), .B2(_02743_ ), .ZN(_02777_ ) );
AOI22_X1 _10477_ ( .A1(_02772_ ), .A2(_02773_ ), .B1(_02774_ ), .B2(_02777_ ), .ZN(_02778_ ) );
NOR2_X1 _10478_ ( .A1(_02777_ ), .A2(_02774_ ), .ZN(_02779_ ) );
OR2_X2 _10479_ ( .A1(_02778_ ), .A2(_02779_ ), .ZN(_02780_ ) );
NAND2_X1 _10480_ ( .A1(_02485_ ), .A2(\IF_ID_inst [25] ), .ZN(_02781_ ) );
MUX2_X1 _10481_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(_02781_ ), .S(_02753_ ), .Z(_02782_ ) );
XNOR2_X1 _10482_ ( .A(_02782_ ), .B(\IF_ID_pc [5] ), .ZN(_02783_ ) );
AND2_X1 _10483_ ( .A1(_02780_ ), .A2(_02783_ ), .ZN(_02784_ ) );
NOR2_X1 _10484_ ( .A1(_02782_ ), .A2(_01022_ ), .ZN(_02785_ ) );
NOR2_X2 _10485_ ( .A1(_02784_ ), .A2(_02785_ ), .ZN(_02786_ ) );
AND2_X1 _10486_ ( .A1(_02754_ ), .A2(_02517_ ), .ZN(_02787_ ) );
OAI21_X1 _10487_ ( .A(_02756_ ), .B1(_02786_ ), .B2(_02787_ ), .ZN(_02788_ ) );
AND2_X1 _10488_ ( .A1(_02485_ ), .A2(\IF_ID_inst [27] ), .ZN(_02789_ ) );
INV_X1 _10489_ ( .A(_02789_ ), .ZN(_02790_ ) );
MUX2_X1 _10490_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(_02790_ ), .S(_02753_ ), .Z(_02791_ ) );
XNOR2_X1 _10491_ ( .A(_02791_ ), .B(\IF_ID_pc [7] ), .ZN(_02792_ ) );
AND2_X2 _10492_ ( .A1(_02788_ ), .A2(_02792_ ), .ZN(_02793_ ) );
NOR2_X1 _10493_ ( .A1(_02791_ ), .A2(_01056_ ), .ZN(_02794_ ) );
AND2_X1 _10494_ ( .A1(_02486_ ), .A2(\IF_ID_inst [28] ), .ZN(_02795_ ) );
INV_X1 _10495_ ( .A(_02795_ ), .ZN(_02796_ ) );
MUX2_X1 _10496_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B(_02796_ ), .S(_02753_ ), .Z(_02797_ ) );
INV_X1 _10497_ ( .A(_02797_ ), .ZN(_02798_ ) );
OAI22_X1 _10498_ ( .A1(_02793_ ), .A2(_02794_ ), .B1(\IF_ID_pc [8] ), .B2(_02798_ ), .ZN(_02799_ ) );
INV_X1 _10499_ ( .A(\IF_ID_pc [8] ), .ZN(_02800_ ) );
NOR2_X1 _10500_ ( .A1(_02797_ ), .A2(_02800_ ), .ZN(_02801_ ) );
INV_X1 _10501_ ( .A(_02801_ ), .ZN(_02802_ ) );
NAND2_X2 _10502_ ( .A1(_02799_ ), .A2(_02802_ ), .ZN(_02803_ ) );
AND2_X1 _10503_ ( .A1(_02486_ ), .A2(\IF_ID_inst [14] ), .ZN(_02804_ ) );
INV_X2 _10504_ ( .A(_02743_ ), .ZN(_02805_ ) );
MUX2_X1 _10505_ ( .A(_02539_ ), .B(_02804_ ), .S(_02805_ ), .Z(_02806_ ) );
INV_X1 _10506_ ( .A(\IF_ID_pc [14] ), .ZN(_02807_ ) );
XNOR2_X1 _10507_ ( .A(_02806_ ), .B(_02807_ ), .ZN(_02808_ ) );
AND2_X1 _10508_ ( .A1(_02486_ ), .A2(\IF_ID_inst [13] ), .ZN(_02809_ ) );
MUX2_X1 _10509_ ( .A(_02539_ ), .B(_02809_ ), .S(_02805_ ), .Z(_02810_ ) );
XNOR2_X1 _10510_ ( .A(_02810_ ), .B(_02506_ ), .ZN(_02811_ ) );
AND2_X1 _10511_ ( .A1(_02808_ ), .A2(_02811_ ), .ZN(_02812_ ) );
AND2_X1 _10512_ ( .A1(_02486_ ), .A2(\IF_ID_inst [16] ), .ZN(_02813_ ) );
MUX2_X1 _10513_ ( .A(_02539_ ), .B(_02813_ ), .S(_02805_ ), .Z(_02814_ ) );
XNOR2_X1 _10514_ ( .A(_02814_ ), .B(_01034_ ), .ZN(_02815_ ) );
AND2_X1 _10515_ ( .A1(_02486_ ), .A2(\IF_ID_inst [15] ), .ZN(_02816_ ) );
MUX2_X1 _10516_ ( .A(_02539_ ), .B(_02816_ ), .S(_02805_ ), .Z(_02817_ ) );
INV_X1 _10517_ ( .A(\IF_ID_pc [15] ), .ZN(_02818_ ) );
XNOR2_X1 _10518_ ( .A(_02817_ ), .B(_02818_ ), .ZN(_02819_ ) );
AND3_X1 _10519_ ( .A1(_02812_ ), .A2(_02815_ ), .A3(_02819_ ), .ZN(_02820_ ) );
AND2_X1 _10520_ ( .A1(_02485_ ), .A2(\IF_ID_inst [20] ), .ZN(_02821_ ) );
INV_X1 _10521_ ( .A(_02821_ ), .ZN(_02822_ ) );
MUX2_X1 _10522_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(_02822_ ), .S(_02753_ ), .Z(_02823_ ) );
XNOR2_X1 _10523_ ( .A(_02823_ ), .B(\IF_ID_pc [11] ), .ZN(_02824_ ) );
AND2_X1 _10524_ ( .A1(_02485_ ), .A2(\IF_ID_inst [12] ), .ZN(_02825_ ) );
MUX2_X1 _10525_ ( .A(_02539_ ), .B(_02825_ ), .S(_02805_ ), .Z(_02826_ ) );
XNOR2_X1 _10526_ ( .A(_02826_ ), .B(_02512_ ), .ZN(_02827_ ) );
NAND2_X1 _10527_ ( .A1(_02824_ ), .A2(_02827_ ), .ZN(_02828_ ) );
AND2_X1 _10528_ ( .A1(_02485_ ), .A2(\IF_ID_inst [30] ), .ZN(_02829_ ) );
INV_X1 _10529_ ( .A(_02829_ ), .ZN(_02830_ ) );
MUX2_X1 _10530_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B(_02830_ ), .S(_02753_ ), .Z(_02831_ ) );
XNOR2_X1 _10531_ ( .A(_02831_ ), .B(\IF_ID_pc [10] ), .ZN(_02832_ ) );
AND2_X1 _10532_ ( .A1(_02486_ ), .A2(\IF_ID_inst [29] ), .ZN(_02833_ ) );
INV_X1 _10533_ ( .A(_02833_ ), .ZN(_02834_ ) );
OAI21_X1 _10534_ ( .A(_02834_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B2(_02805_ ), .ZN(_02835_ ) );
XNOR2_X1 _10535_ ( .A(_02835_ ), .B(_02516_ ), .ZN(_02836_ ) );
NAND2_X1 _10536_ ( .A1(_02832_ ), .A2(_02836_ ), .ZN(_02837_ ) );
NOR2_X1 _10537_ ( .A1(_02828_ ), .A2(_02837_ ), .ZN(_02838_ ) );
NAND3_X1 _10538_ ( .A1(_02803_ ), .A2(_02820_ ), .A3(_02838_ ), .ZN(_02839_ ) );
NOR2_X1 _10539_ ( .A1(_02831_ ), .A2(_02514_ ), .ZN(_02840_ ) );
AND2_X1 _10540_ ( .A1(_02831_ ), .A2(_02514_ ), .ZN(_02841_ ) );
INV_X1 _10541_ ( .A(_02841_ ), .ZN(_02842_ ) );
MUX2_X1 _10542_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(_02834_ ), .S(_02753_ ), .Z(_02843_ ) );
NOR2_X1 _10543_ ( .A1(_02843_ ), .A2(_02516_ ), .ZN(_02844_ ) );
AOI21_X1 _10544_ ( .A(_02840_ ), .B1(_02842_ ), .B2(_02844_ ), .ZN(_02845_ ) );
OR2_X1 _10545_ ( .A1(_02845_ ), .A2(_02828_ ), .ZN(_02846_ ) );
AND2_X1 _10546_ ( .A1(_02826_ ), .A2(\IF_ID_pc [12] ), .ZN(_02847_ ) );
INV_X1 _10547_ ( .A(_02847_ ), .ZN(_02848_ ) );
NOR2_X1 _10548_ ( .A1(_02823_ ), .A2(_02513_ ), .ZN(_02849_ ) );
NAND2_X1 _10549_ ( .A1(_02827_ ), .A2(_02849_ ), .ZN(_02850_ ) );
NAND3_X1 _10550_ ( .A1(_02846_ ), .A2(_02848_ ), .A3(_02850_ ), .ZN(_02851_ ) );
NAND2_X1 _10551_ ( .A1(_02851_ ), .A2(_02820_ ), .ZN(_02852_ ) );
AND2_X1 _10552_ ( .A1(_02814_ ), .A2(\IF_ID_pc [16] ), .ZN(_02853_ ) );
AND2_X1 _10553_ ( .A1(_02817_ ), .A2(\IF_ID_pc [15] ), .ZN(_02854_ ) );
AOI21_X1 _10554_ ( .A(_02853_ ), .B1(_02815_ ), .B2(_02854_ ), .ZN(_02855_ ) );
AND2_X1 _10555_ ( .A1(_02810_ ), .A2(\IF_ID_pc [13] ), .ZN(_02856_ ) );
AND2_X1 _10556_ ( .A1(_02808_ ), .A2(_02856_ ), .ZN(_02857_ ) );
AND2_X1 _10557_ ( .A1(_02806_ ), .A2(\IF_ID_pc [14] ), .ZN(_02858_ ) );
OAI211_X1 _10558_ ( .A(_02815_ ), .B(_02819_ ), .C1(_02857_ ), .C2(_02858_ ), .ZN(_02859_ ) );
AND3_X1 _10559_ ( .A1(_02852_ ), .A2(_02855_ ), .A3(_02859_ ), .ZN(_02860_ ) );
NAND2_X2 _10560_ ( .A1(_02839_ ), .A2(_02860_ ), .ZN(_02861_ ) );
AND2_X1 _10561_ ( .A1(_02486_ ), .A2(\IF_ID_inst [18] ), .ZN(_02862_ ) );
MUX2_X1 _10562_ ( .A(_02539_ ), .B(_02862_ ), .S(_02805_ ), .Z(_02863_ ) );
XNOR2_X1 _10563_ ( .A(_02863_ ), .B(_01110_ ), .ZN(_02864_ ) );
AND2_X1 _10564_ ( .A1(_02486_ ), .A2(\IF_ID_inst [17] ), .ZN(_02865_ ) );
MUX2_X1 _10565_ ( .A(_02539_ ), .B(_02865_ ), .S(_02805_ ), .Z(_02866_ ) );
XNOR2_X1 _10566_ ( .A(_02866_ ), .B(_01123_ ), .ZN(_02867_ ) );
AND2_X1 _10567_ ( .A1(_02864_ ), .A2(_02867_ ), .ZN(_02868_ ) );
XNOR2_X1 _10568_ ( .A(_02747_ ), .B(_02508_ ), .ZN(_02869_ ) );
AND2_X1 _10569_ ( .A1(_02487_ ), .A2(\IF_ID_inst [19] ), .ZN(_02870_ ) );
MUX2_X1 _10570_ ( .A(_02539_ ), .B(_02870_ ), .S(_02805_ ), .Z(_02871_ ) );
XNOR2_X1 _10571_ ( .A(_02871_ ), .B(_01102_ ), .ZN(_02872_ ) );
NAND4_X1 _10572_ ( .A1(_02861_ ), .A2(_02868_ ), .A3(_02869_ ), .A4(_02872_ ), .ZN(_02873_ ) );
AND2_X1 _10573_ ( .A1(_02866_ ), .A2(\IF_ID_pc [17] ), .ZN(_02874_ ) );
AND2_X1 _10574_ ( .A1(_02864_ ), .A2(_02874_ ), .ZN(_02875_ ) );
AND2_X1 _10575_ ( .A1(_02863_ ), .A2(\IF_ID_pc [18] ), .ZN(_02876_ ) );
OAI211_X1 _10576_ ( .A(_02869_ ), .B(_02872_ ), .C1(_02875_ ), .C2(_02876_ ), .ZN(_02877_ ) );
AND3_X1 _10577_ ( .A1(_02869_ ), .A2(\IF_ID_pc [19] ), .A3(_02871_ ), .ZN(_02878_ ) );
AOI21_X1 _10578_ ( .A(_02878_ ), .B1(\IF_ID_pc [20] ), .B2(_02747_ ), .ZN(_02879_ ) );
AND2_X1 _10579_ ( .A1(_02877_ ), .A2(_02879_ ), .ZN(_02880_ ) );
NAND2_X2 _10580_ ( .A1(_02873_ ), .A2(_02880_ ), .ZN(_02881_ ) );
XNOR2_X1 _10581_ ( .A(_02747_ ), .B(_01165_ ), .ZN(_02882_ ) );
XNOR2_X1 _10582_ ( .A(_02747_ ), .B(_02507_ ), .ZN(_02883_ ) );
XNOR2_X1 _10583_ ( .A(_02747_ ), .B(_01158_ ), .ZN(_02884_ ) );
AND2_X1 _10584_ ( .A1(_02883_ ), .A2(_02884_ ), .ZN(_02885_ ) );
AND4_X1 _10585_ ( .A1(_02749_ ), .A2(_02881_ ), .A3(_02882_ ), .A4(_02885_ ), .ZN(_02886_ ) );
NOR4_X1 _10586_ ( .A1(_02744_ ), .A2(_02745_ ), .A3(\IF_ID_pc [22] ), .A4(_01158_ ), .ZN(_02887_ ) );
NOR3_X1 _10587_ ( .A1(_02744_ ), .A2(_02745_ ), .A3(_02507_ ), .ZN(_02888_ ) );
NOR2_X1 _10588_ ( .A1(_02887_ ), .A2(_02888_ ), .ZN(_02889_ ) );
BUF_X4 _10589_ ( .A(_02747_ ), .Z(_02890_ ) );
INV_X1 _10590_ ( .A(_02890_ ), .ZN(_02891_ ) );
OAI21_X1 _10591_ ( .A(_02889_ ), .B1(_02891_ ), .B2(_02499_ ), .ZN(_02892_ ) );
NOR2_X1 _10592_ ( .A1(_02886_ ), .A2(_02892_ ), .ZN(_02893_ ) );
INV_X1 _10593_ ( .A(_02893_ ), .ZN(_02894_ ) );
XNOR2_X1 _10594_ ( .A(_02747_ ), .B(_01149_ ), .ZN(_02895_ ) );
XNOR2_X1 _10595_ ( .A(_02747_ ), .B(_01274_ ), .ZN(_02896_ ) );
AND2_X1 _10596_ ( .A1(_02895_ ), .A2(_02896_ ), .ZN(_02897_ ) );
XNOR2_X1 _10597_ ( .A(_02890_ ), .B(_01261_ ), .ZN(_02898_ ) );
XNOR2_X1 _10598_ ( .A(_02890_ ), .B(_01242_ ), .ZN(_02899_ ) );
NAND4_X1 _10599_ ( .A1(_02894_ ), .A2(_02897_ ), .A3(_02898_ ), .A4(_02899_ ), .ZN(_02900_ ) );
AND2_X1 _10600_ ( .A1(_02747_ ), .A2(\IF_ID_pc [27] ), .ZN(_02901_ ) );
OAI21_X1 _10601_ ( .A(_02890_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_02902_ ) );
INV_X1 _10602_ ( .A(_02902_ ), .ZN(_02903_ ) );
AOI221_X4 _10603_ ( .A(_02901_ ), .B1(\IF_ID_pc [28] ), .B2(_02890_ ), .C1(_02897_ ), .C2(_02903_ ), .ZN(_02904_ ) );
AND2_X1 _10604_ ( .A1(_02900_ ), .A2(_02904_ ), .ZN(_02905_ ) );
INV_X2 _10605_ ( .A(_02905_ ), .ZN(_02906_ ) );
XNOR2_X1 _10606_ ( .A(_02890_ ), .B(_01257_ ), .ZN(_02907_ ) );
NAND2_X1 _10607_ ( .A1(_02906_ ), .A2(_02907_ ), .ZN(_02908_ ) );
AND2_X1 _10608_ ( .A1(_02890_ ), .A2(\IF_ID_pc [30] ), .ZN(_02909_ ) );
INV_X1 _10609_ ( .A(_02909_ ), .ZN(_02910_ ) );
OAI21_X1 _10610_ ( .A(_01049_ ), .B1(_02744_ ), .B2(_02745_ ), .ZN(_02911_ ) );
AND4_X1 _10611_ ( .A1(_02746_ ), .A2(_02908_ ), .A3(_02910_ ), .A4(_02911_ ), .ZN(_02912_ ) );
AOI22_X1 _10612_ ( .A1(_02908_ ), .A2(_02746_ ), .B1(_02910_ ), .B2(_02911_ ), .ZN(_02913_ ) );
OAI21_X1 _10613_ ( .A(_02741_ ), .B1(_02912_ ), .B2(_02913_ ), .ZN(_02914_ ) );
NAND2_X1 _10614_ ( .A1(\mtvec [30] ), .A2(fanout_net_42 ), .ZN(_02915_ ) );
AOI21_X1 _10615_ ( .A(fanout_net_3 ), .B1(_02914_ ), .B2(_02915_ ), .ZN(_00213_ ) );
BUF_X4 _10616_ ( .A(_02522_ ), .Z(_02916_ ) );
AOI211_X1 _10617_ ( .A(fanout_net_42 ), .B(_02916_ ), .C1(_02906_ ), .C2(_02907_ ), .ZN(_02917_ ) );
OAI21_X1 _10618_ ( .A(_02917_ ), .B1(_02907_ ), .B2(_02906_ ), .ZN(_02918_ ) );
NAND2_X1 _10619_ ( .A1(\mtvec [29] ), .A2(fanout_net_42 ), .ZN(_02919_ ) );
AOI21_X1 _10620_ ( .A(fanout_net_3 ), .B1(_02918_ ), .B2(_02919_ ), .ZN(_00214_ ) );
INV_X1 _10621_ ( .A(_02872_ ), .ZN(_02920_ ) );
NAND2_X1 _10622_ ( .A1(_02861_ ), .A2(_02868_ ), .ZN(_02921_ ) );
AOI21_X1 _10623_ ( .A(_02876_ ), .B1(_02864_ ), .B2(_02874_ ), .ZN(_02922_ ) );
AOI21_X1 _10624_ ( .A(_02920_ ), .B1(_02921_ ), .B2(_02922_ ), .ZN(_02923_ ) );
AND2_X1 _10625_ ( .A1(_02871_ ), .A2(\IF_ID_pc [19] ), .ZN(_02924_ ) );
OR3_X1 _10626_ ( .A1(_02923_ ), .A2(_02924_ ), .A3(_02869_ ), .ZN(_02925_ ) );
OAI21_X1 _10627_ ( .A(_02869_ ), .B1(_02923_ ), .B2(_02924_ ), .ZN(_02926_ ) );
NAND3_X1 _10628_ ( .A1(_02925_ ), .A2(_02741_ ), .A3(_02926_ ), .ZN(_02927_ ) );
NAND2_X1 _10629_ ( .A1(\mtvec [20] ), .A2(fanout_net_42 ), .ZN(_02928_ ) );
AOI21_X1 _10630_ ( .A(fanout_net_3 ), .B1(_02927_ ), .B2(_02928_ ), .ZN(_00215_ ) );
NOR3_X1 _10631_ ( .A1(_02923_ ), .A2(fanout_net_42 ), .A3(_02916_ ), .ZN(_02929_ ) );
AND2_X1 _10632_ ( .A1(_02921_ ), .A2(_02922_ ), .ZN(_02930_ ) );
INV_X1 _10633_ ( .A(_02930_ ), .ZN(_02931_ ) );
OAI21_X1 _10634_ ( .A(_02929_ ), .B1(_02872_ ), .B2(_02931_ ), .ZN(_02932_ ) );
NAND2_X1 _10635_ ( .A1(\mtvec [19] ), .A2(fanout_net_42 ), .ZN(_02933_ ) );
AOI21_X1 _10636_ ( .A(fanout_net_3 ), .B1(_02932_ ), .B2(_02933_ ), .ZN(_00216_ ) );
AND2_X1 _10637_ ( .A1(_02861_ ), .A2(_02867_ ), .ZN(_02934_ ) );
OR3_X1 _10638_ ( .A1(_02934_ ), .A2(_02864_ ), .A3(_02874_ ), .ZN(_02935_ ) );
OAI21_X1 _10639_ ( .A(_02864_ ), .B1(_02934_ ), .B2(_02874_ ), .ZN(_02936_ ) );
NAND3_X1 _10640_ ( .A1(_02935_ ), .A2(_02741_ ), .A3(_02936_ ), .ZN(_02937_ ) );
NAND2_X1 _10641_ ( .A1(\mtvec [18] ), .A2(fanout_net_42 ), .ZN(_02938_ ) );
AOI21_X1 _10642_ ( .A(fanout_net_3 ), .B1(_02937_ ), .B2(_02938_ ), .ZN(_00217_ ) );
AOI211_X1 _10643_ ( .A(fanout_net_42 ), .B(_02916_ ), .C1(_02861_ ), .C2(_02867_ ), .ZN(_02939_ ) );
OAI21_X1 _10644_ ( .A(_02939_ ), .B1(_02861_ ), .B2(_02867_ ), .ZN(_02940_ ) );
NAND2_X1 _10645_ ( .A1(\mtvec [17] ), .A2(fanout_net_42 ), .ZN(_02941_ ) );
AOI21_X1 _10646_ ( .A(fanout_net_3 ), .B1(_02940_ ), .B2(_02941_ ), .ZN(_00218_ ) );
NAND2_X1 _10647_ ( .A1(_02808_ ), .A2(_02856_ ), .ZN(_02942_ ) );
INV_X1 _10648_ ( .A(_02858_ ), .ZN(_02943_ ) );
AND2_X1 _10649_ ( .A1(_02942_ ), .A2(_02943_ ), .ZN(_02944_ ) );
INV_X1 _10650_ ( .A(_02944_ ), .ZN(_02945_ ) );
AOI211_X1 _10651_ ( .A(_02837_ ), .B(_02828_ ), .C1(_02799_ ), .C2(_02802_ ), .ZN(_02946_ ) );
OR2_X1 _10652_ ( .A1(_02946_ ), .A2(_02851_ ), .ZN(_02947_ ) );
AOI21_X1 _10653_ ( .A(_02945_ ), .B1(_02947_ ), .B2(_02812_ ), .ZN(_02948_ ) );
INV_X1 _10654_ ( .A(_02948_ ), .ZN(_02949_ ) );
AND2_X1 _10655_ ( .A1(_02949_ ), .A2(_02819_ ), .ZN(_02950_ ) );
OR3_X1 _10656_ ( .A1(_02950_ ), .A2(_02854_ ), .A3(_02815_ ), .ZN(_02951_ ) );
OAI21_X1 _10657_ ( .A(_02815_ ), .B1(_02950_ ), .B2(_02854_ ), .ZN(_02952_ ) );
NAND3_X1 _10658_ ( .A1(_02951_ ), .A2(_02741_ ), .A3(_02952_ ), .ZN(_02953_ ) );
NAND2_X1 _10659_ ( .A1(\mtvec [16] ), .A2(fanout_net_42 ), .ZN(_02954_ ) );
AOI21_X1 _10660_ ( .A(fanout_net_3 ), .B1(_02953_ ), .B2(_02954_ ), .ZN(_00219_ ) );
AOI211_X1 _10661_ ( .A(fanout_net_42 ), .B(_02916_ ), .C1(_02949_ ), .C2(_02819_ ), .ZN(_02955_ ) );
OAI21_X1 _10662_ ( .A(_02955_ ), .B1(_02819_ ), .B2(_02949_ ), .ZN(_02956_ ) );
NAND2_X1 _10663_ ( .A1(\mtvec [15] ), .A2(fanout_net_42 ), .ZN(_02957_ ) );
AOI21_X1 _10664_ ( .A(fanout_net_3 ), .B1(_02956_ ), .B2(_02957_ ), .ZN(_00220_ ) );
NAND3_X1 _10665_ ( .A1(_02803_ ), .A2(_02836_ ), .A3(_02832_ ), .ZN(_02958_ ) );
NAND2_X1 _10666_ ( .A1(_02958_ ), .A2(_02845_ ), .ZN(_02959_ ) );
AND2_X1 _10667_ ( .A1(_02959_ ), .A2(_02824_ ), .ZN(_02960_ ) );
NOR2_X1 _10668_ ( .A1(_02960_ ), .A2(_02849_ ), .ZN(_02961_ ) );
NOR2_X1 _10669_ ( .A1(_02826_ ), .A2(\IF_ID_pc [12] ), .ZN(_02962_ ) );
OAI21_X1 _10670_ ( .A(_02848_ ), .B1(_02961_ ), .B2(_02962_ ), .ZN(_02963_ ) );
AND2_X1 _10671_ ( .A1(_02963_ ), .A2(_02811_ ), .ZN(_02964_ ) );
OR3_X1 _10672_ ( .A1(_02964_ ), .A2(_02856_ ), .A3(_02808_ ), .ZN(_02965_ ) );
OAI21_X1 _10673_ ( .A(_02808_ ), .B1(_02964_ ), .B2(_02856_ ), .ZN(_02966_ ) );
NAND3_X1 _10674_ ( .A1(_02965_ ), .A2(_02741_ ), .A3(_02966_ ), .ZN(_02967_ ) );
NAND2_X1 _10675_ ( .A1(\mtvec [14] ), .A2(fanout_net_42 ), .ZN(_02968_ ) );
AOI21_X1 _10676_ ( .A(fanout_net_3 ), .B1(_02967_ ), .B2(_02968_ ), .ZN(_00221_ ) );
AOI21_X1 _10677_ ( .A(_02962_ ), .B1(_02961_ ), .B2(_02848_ ), .ZN(_02969_ ) );
NAND2_X1 _10678_ ( .A1(_02969_ ), .A2(_02811_ ), .ZN(_02970_ ) );
OAI211_X1 _10679_ ( .A(_02970_ ), .B(_02740_ ), .C1(_02811_ ), .C2(_02947_ ), .ZN(_02971_ ) );
NAND2_X1 _10680_ ( .A1(\mtvec [13] ), .A2(fanout_net_42 ), .ZN(_02972_ ) );
AOI21_X1 _10681_ ( .A(fanout_net_3 ), .B1(_02971_ ), .B2(_02972_ ), .ZN(_00222_ ) );
XNOR2_X1 _10682_ ( .A(_02961_ ), .B(_02827_ ), .ZN(_02973_ ) );
AOI22_X1 _10683_ ( .A1(_02973_ ), .A2(_02741_ ), .B1(\mtvec [12] ), .B2(fanout_net_42 ), .ZN(_02974_ ) );
NOR2_X1 _10684_ ( .A1(_02974_ ), .A2(fanout_net_3 ), .ZN(_00223_ ) );
AOI211_X1 _10685_ ( .A(fanout_net_42 ), .B(_02916_ ), .C1(_02959_ ), .C2(_02824_ ), .ZN(_02975_ ) );
OAI21_X1 _10686_ ( .A(_02975_ ), .B1(_02824_ ), .B2(_02959_ ), .ZN(_02976_ ) );
NAND2_X1 _10687_ ( .A1(\mtvec [11] ), .A2(fanout_net_42 ), .ZN(_02977_ ) );
AOI21_X1 _10688_ ( .A(fanout_net_3 ), .B1(_02976_ ), .B2(_02977_ ), .ZN(_00224_ ) );
INV_X1 _10689_ ( .A(_02899_ ), .ZN(_02978_ ) );
NOR2_X1 _10690_ ( .A1(_02893_ ), .A2(_02978_ ), .ZN(_02979_ ) );
AOI21_X1 _10691_ ( .A(_02903_ ), .B1(_02979_ ), .B2(_02898_ ), .ZN(_02980_ ) );
INV_X1 _10692_ ( .A(_02980_ ), .ZN(_02981_ ) );
AOI21_X1 _10693_ ( .A(_02901_ ), .B1(_02981_ ), .B2(_02896_ ), .ZN(_02982_ ) );
INV_X1 _10694_ ( .A(_02982_ ), .ZN(_02983_ ) );
AND2_X1 _10695_ ( .A1(_02983_ ), .A2(_02895_ ), .ZN(_02984_ ) );
OAI21_X1 _10696_ ( .A(_02740_ ), .B1(_02983_ ), .B2(_02895_ ), .ZN(_02985_ ) );
OR2_X1 _10697_ ( .A1(_02984_ ), .A2(_02985_ ), .ZN(_02986_ ) );
NAND2_X1 _10698_ ( .A1(\mtvec [28] ), .A2(fanout_net_42 ), .ZN(_02987_ ) );
AOI21_X1 _10699_ ( .A(fanout_net_4 ), .B1(_02986_ ), .B2(_02987_ ), .ZN(_00225_ ) );
NAND2_X1 _10700_ ( .A1(_02803_ ), .A2(_02836_ ), .ZN(_02988_ ) );
INV_X1 _10701_ ( .A(_02844_ ), .ZN(_02989_ ) );
NAND2_X1 _10702_ ( .A1(_02988_ ), .A2(_02989_ ), .ZN(_02990_ ) );
AND2_X1 _10703_ ( .A1(_02990_ ), .A2(_02832_ ), .ZN(_02991_ ) );
OAI21_X1 _10704_ ( .A(_02740_ ), .B1(_02990_ ), .B2(_02832_ ), .ZN(_02992_ ) );
OR2_X1 _10705_ ( .A1(_02991_ ), .A2(_02992_ ), .ZN(_02993_ ) );
NAND2_X1 _10706_ ( .A1(\mtvec [10] ), .A2(fanout_net_42 ), .ZN(_02994_ ) );
AOI21_X1 _10707_ ( .A(fanout_net_4 ), .B1(_02993_ ), .B2(_02994_ ), .ZN(_00226_ ) );
AOI211_X1 _10708_ ( .A(fanout_net_42 ), .B(_02916_ ), .C1(_02803_ ), .C2(_02836_ ), .ZN(_02995_ ) );
OAI21_X1 _10709_ ( .A(_02995_ ), .B1(_02803_ ), .B2(_02836_ ), .ZN(_02996_ ) );
NAND2_X1 _10710_ ( .A1(\mtvec [9] ), .A2(fanout_net_42 ), .ZN(_02997_ ) );
AOI21_X1 _10711_ ( .A(fanout_net_4 ), .B1(_02996_ ), .B2(_02997_ ), .ZN(_00227_ ) );
XNOR2_X1 _10712_ ( .A(_02797_ ), .B(\IF_ID_pc [8] ), .ZN(_02998_ ) );
OR3_X1 _10713_ ( .A1(_02793_ ), .A2(_02794_ ), .A3(_02998_ ), .ZN(_02999_ ) );
OAI21_X1 _10714_ ( .A(_02998_ ), .B1(_02793_ ), .B2(_02794_ ), .ZN(_03000_ ) );
NAND3_X1 _10715_ ( .A1(_02999_ ), .A2(_02741_ ), .A3(_03000_ ), .ZN(_03001_ ) );
NAND2_X1 _10716_ ( .A1(\mtvec [8] ), .A2(fanout_net_42 ), .ZN(_03002_ ) );
AOI21_X1 _10717_ ( .A(fanout_net_4 ), .B1(_03001_ ), .B2(_03002_ ), .ZN(_00228_ ) );
AOI211_X1 _10718_ ( .A(fanout_net_42 ), .B(_02916_ ), .C1(_02788_ ), .C2(_02792_ ), .ZN(_03003_ ) );
OAI21_X1 _10719_ ( .A(_03003_ ), .B1(_02792_ ), .B2(_02788_ ), .ZN(_03004_ ) );
NAND2_X1 _10720_ ( .A1(\mtvec [7] ), .A2(fanout_net_42 ), .ZN(_03005_ ) );
AOI21_X1 _10721_ ( .A(fanout_net_4 ), .B1(_03004_ ), .B2(_03005_ ), .ZN(_00229_ ) );
INV_X1 _10722_ ( .A(_02786_ ), .ZN(_03006_ ) );
XNOR2_X1 _10723_ ( .A(_02754_ ), .B(\IF_ID_pc [6] ), .ZN(_03007_ ) );
OAI21_X1 _10724_ ( .A(_02740_ ), .B1(_03006_ ), .B2(_03007_ ), .ZN(_03008_ ) );
NOR3_X1 _10725_ ( .A1(_02786_ ), .A2(_02755_ ), .A3(_02787_ ), .ZN(_03009_ ) );
OR2_X1 _10726_ ( .A1(_03008_ ), .A2(_03009_ ), .ZN(_03010_ ) );
NAND2_X1 _10727_ ( .A1(\mtvec [6] ), .A2(fanout_net_42 ), .ZN(_03011_ ) );
AOI21_X1 _10728_ ( .A(fanout_net_4 ), .B1(_03010_ ), .B2(_03011_ ), .ZN(_00230_ ) );
AOI211_X1 _10729_ ( .A(fanout_net_42 ), .B(_02522_ ), .C1(_02780_ ), .C2(_02783_ ), .ZN(_03012_ ) );
OAI21_X1 _10730_ ( .A(_03012_ ), .B1(_02780_ ), .B2(_02783_ ), .ZN(_03013_ ) );
NAND2_X1 _10731_ ( .A1(\mtvec [5] ), .A2(fanout_net_42 ), .ZN(_03014_ ) );
AOI21_X1 _10732_ ( .A(fanout_net_4 ), .B1(_03013_ ), .B2(_03014_ ), .ZN(_00231_ ) );
AND2_X1 _10733_ ( .A1(_02772_ ), .A2(_02773_ ), .ZN(_03015_ ) );
XNOR2_X1 _10734_ ( .A(_02777_ ), .B(\IF_ID_pc [4] ), .ZN(_03016_ ) );
XNOR2_X1 _10735_ ( .A(_03015_ ), .B(_03016_ ), .ZN(_03017_ ) );
OAI211_X1 _10736_ ( .A(_03017_ ), .B(_02523_ ), .C1(_01353_ ), .C2(_02521_ ), .ZN(_03018_ ) );
NAND2_X1 _10737_ ( .A1(\mtvec [4] ), .A2(fanout_net_42 ), .ZN(_03019_ ) );
AOI21_X1 _10738_ ( .A(fanout_net_4 ), .B1(_03018_ ), .B2(_03019_ ), .ZN(_00232_ ) );
OR2_X1 _10739_ ( .A1(_02767_ ), .A2(_02771_ ), .ZN(_03020_ ) );
AND3_X1 _10740_ ( .A1(_03020_ ), .A2(_02740_ ), .A3(_02772_ ), .ZN(_03021_ ) );
AOI21_X1 _10741_ ( .A(_03021_ ), .B1(\mtvec [3] ), .B2(\myifu.to_reset ), .ZN(_03022_ ) );
NOR2_X1 _10742_ ( .A1(_03022_ ), .A2(fanout_net_4 ), .ZN(_00233_ ) );
AND2_X1 _10743_ ( .A1(_02760_ ), .A2(\IF_ID_pc [1] ), .ZN(_03023_ ) );
XNOR2_X1 _10744_ ( .A(_03023_ ), .B(_02765_ ), .ZN(_03024_ ) );
INV_X1 _10745_ ( .A(_02521_ ), .ZN(_03025_ ) );
AOI211_X1 _10746_ ( .A(\myifu.to_reset ), .B(_03024_ ), .C1(check_quest ), .C2(_03025_ ), .ZN(_03026_ ) );
AOI21_X1 _10747_ ( .A(_03026_ ), .B1(\mtvec [2] ), .B2(\myifu.to_reset ), .ZN(_03027_ ) );
NOR2_X1 _10748_ ( .A1(_03027_ ), .A2(fanout_net_4 ), .ZN(_00234_ ) );
AND2_X1 _10749_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _10750_ ( .A(_00830_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_E ), .B2(\IF_ID_pc [3] ), .ZN(_03028_ ) );
AOI21_X1 _10751_ ( .A(_03028_ ), .B1(_03022_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_E ), .ZN(_00235_ ) );
AOI211_X1 _10752_ ( .A(\myifu.to_reset ), .B(_02522_ ), .C1(_02760_ ), .C2(\IF_ID_pc [1] ), .ZN(_03029_ ) );
OAI21_X1 _10753_ ( .A(_03029_ ), .B1(\IF_ID_pc [1] ), .B2(_02760_ ), .ZN(_03030_ ) );
NAND2_X1 _10754_ ( .A1(\mtvec [1] ), .A2(\myifu.to_reset ), .ZN(_03031_ ) );
AOI21_X1 _10755_ ( .A(fanout_net_4 ), .B1(_03030_ ), .B2(_03031_ ), .ZN(_00236_ ) );
OAI21_X1 _10756_ ( .A(_00830_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_E ), .B2(\IF_ID_pc [2] ), .ZN(_03032_ ) );
AOI21_X1 _10757_ ( .A(_03032_ ), .B1(_03027_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_E ), .ZN(_00237_ ) );
AOI211_X1 _10758_ ( .A(\myifu.to_reset ), .B(_02522_ ), .C1(_02981_ ), .C2(_02896_ ), .ZN(_03033_ ) );
OAI21_X1 _10759_ ( .A(_03033_ ), .B1(_02896_ ), .B2(_02981_ ), .ZN(_03034_ ) );
NAND2_X1 _10760_ ( .A1(\mtvec [27] ), .A2(\myifu.to_reset ), .ZN(_03035_ ) );
AOI21_X1 _10761_ ( .A(fanout_net_4 ), .B1(_03034_ ), .B2(_03035_ ), .ZN(_00238_ ) );
AND3_X1 _10762_ ( .A1(_00841_ ), .A2(\mtvec [0] ), .A3(\myifu.to_reset ), .ZN(_00239_ ) );
INV_X1 _10763_ ( .A(_02979_ ), .ZN(_03036_ ) );
OAI21_X1 _10764_ ( .A(_03036_ ), .B1(_01242_ ), .B2(_02891_ ), .ZN(_03037_ ) );
AND2_X1 _10765_ ( .A1(_03037_ ), .A2(_02898_ ), .ZN(_03038_ ) );
OAI21_X1 _10766_ ( .A(_02740_ ), .B1(_03037_ ), .B2(_02898_ ), .ZN(_03039_ ) );
OR2_X1 _10767_ ( .A1(_03038_ ), .A2(_03039_ ), .ZN(_03040_ ) );
NAND2_X1 _10768_ ( .A1(\mtvec [26] ), .A2(\myifu.to_reset ), .ZN(_03041_ ) );
AOI21_X1 _10769_ ( .A(fanout_net_4 ), .B1(_03040_ ), .B2(_03041_ ), .ZN(_00240_ ) );
NOR3_X1 _10770_ ( .A1(_02979_ ), .A2(\myifu.to_reset ), .A3(_02916_ ), .ZN(_03042_ ) );
OAI21_X1 _10771_ ( .A(_03042_ ), .B1(_02894_ ), .B2(_02899_ ), .ZN(_03043_ ) );
NAND2_X1 _10772_ ( .A1(\mtvec [25] ), .A2(\myifu.to_reset ), .ZN(_03044_ ) );
AOI21_X1 _10773_ ( .A(fanout_net_4 ), .B1(_03043_ ), .B2(_03044_ ), .ZN(_00241_ ) );
NOR3_X1 _10774_ ( .A1(_02744_ ), .A2(_02745_ ), .A3(_01165_ ), .ZN(_03045_ ) );
NAND2_X1 _10775_ ( .A1(_02881_ ), .A2(_02885_ ), .ZN(_03046_ ) );
NAND2_X1 _10776_ ( .A1(_03046_ ), .A2(_02889_ ), .ZN(_03047_ ) );
AOI21_X1 _10777_ ( .A(_03045_ ), .B1(_03047_ ), .B2(_02882_ ), .ZN(_03048_ ) );
AOI211_X1 _10778_ ( .A(\myifu.to_reset ), .B(_02522_ ), .C1(_03048_ ), .C2(_02748_ ), .ZN(_03049_ ) );
OAI21_X1 _10779_ ( .A(_03049_ ), .B1(_02748_ ), .B2(_03048_ ), .ZN(_03050_ ) );
NAND2_X1 _10780_ ( .A1(\mtvec [24] ), .A2(\myifu.to_reset ), .ZN(_03051_ ) );
AOI21_X1 _10781_ ( .A(fanout_net_4 ), .B1(_03050_ ), .B2(_03051_ ), .ZN(_00242_ ) );
AOI211_X1 _10782_ ( .A(\myifu.to_reset ), .B(_02522_ ), .C1(_03047_ ), .C2(_02882_ ), .ZN(_03052_ ) );
OAI21_X1 _10783_ ( .A(_03052_ ), .B1(_02882_ ), .B2(_03047_ ), .ZN(_03053_ ) );
NAND2_X1 _10784_ ( .A1(\mtvec [23] ), .A2(\myifu.to_reset ), .ZN(_03054_ ) );
AOI21_X1 _10785_ ( .A(fanout_net_4 ), .B1(_03053_ ), .B2(_03054_ ), .ZN(_00243_ ) );
AND2_X1 _10786_ ( .A1(_02881_ ), .A2(_02884_ ), .ZN(_03055_ ) );
AND2_X1 _10787_ ( .A1(_02890_ ), .A2(\IF_ID_pc [21] ), .ZN(_03056_ ) );
OR3_X1 _10788_ ( .A1(_03055_ ), .A2(_03056_ ), .A3(_02883_ ), .ZN(_03057_ ) );
OAI21_X1 _10789_ ( .A(_02883_ ), .B1(_03055_ ), .B2(_03056_ ), .ZN(_03058_ ) );
NAND3_X1 _10790_ ( .A1(_03057_ ), .A2(_02741_ ), .A3(_03058_ ), .ZN(_03059_ ) );
NAND2_X1 _10791_ ( .A1(\mtvec [22] ), .A2(\myifu.to_reset ), .ZN(_03060_ ) );
AOI21_X1 _10792_ ( .A(fanout_net_4 ), .B1(_03059_ ), .B2(_03060_ ), .ZN(_00244_ ) );
AOI211_X1 _10793_ ( .A(\myifu.to_reset ), .B(_02522_ ), .C1(_02881_ ), .C2(_02884_ ), .ZN(_03061_ ) );
OAI21_X1 _10794_ ( .A(_03061_ ), .B1(_02884_ ), .B2(_02881_ ), .ZN(_03062_ ) );
NAND2_X1 _10795_ ( .A1(\mtvec [21] ), .A2(\myifu.to_reset ), .ZN(_03063_ ) );
AOI21_X1 _10796_ ( .A(fanout_net_4 ), .B1(_03062_ ), .B2(_03063_ ), .ZN(_00245_ ) );
NAND4_X1 _10797_ ( .A1(_02906_ ), .A2(_02907_ ), .A3(_02910_ ), .A4(_02911_ ), .ZN(_03064_ ) );
NAND3_X1 _10798_ ( .A1(_02890_ ), .A2(_01049_ ), .A3(\IF_ID_pc [29] ), .ZN(_03065_ ) );
AND3_X1 _10799_ ( .A1(_03064_ ), .A2(_02910_ ), .A3(_03065_ ), .ZN(_03066_ ) );
INV_X1 _10800_ ( .A(_03066_ ), .ZN(_03067_ ) );
XNOR2_X1 _10801_ ( .A(_02890_ ), .B(\IF_ID_pc [31] ), .ZN(_03068_ ) );
AOI211_X1 _10802_ ( .A(\myifu.to_reset ), .B(_02522_ ), .C1(_03067_ ), .C2(_03068_ ), .ZN(_03069_ ) );
OAI21_X1 _10803_ ( .A(_03069_ ), .B1(_03067_ ), .B2(_03068_ ), .ZN(_03070_ ) );
OAI211_X1 _10804_ ( .A(_03070_ ), .B(_00732_ ), .C1(\mtvec [31] ), .C2(_02523_ ), .ZN(_03071_ ) );
NAND2_X1 _10805_ ( .A1(_03071_ ), .A2(_00841_ ), .ZN(_00246_ ) );
NOR3_X1 _10806_ ( .A1(fanout_net_4 ), .A2(\myifu.state [1] ), .A3(fanout_net_41 ), .ZN(_00247_ ) );
INV_X1 _10807_ ( .A(\myifu.state [1] ), .ZN(_03072_ ) );
AND3_X1 _10808_ ( .A1(_01342_ ), .A2(_03072_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_03073_ ) );
INV_X1 _10809_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_03074_ ) );
MUX2_X1 _10810_ ( .A(_01342_ ), .B(_03074_ ), .S(\myifu.to_reset ), .Z(_03075_ ) );
AOI211_X1 _10811_ ( .A(fanout_net_4 ), .B(_03073_ ), .C1(_03075_ ), .C2(\myifu.state [1] ), .ZN(_00248_ ) );
INV_X1 _10812_ ( .A(\myec.state [0] ), .ZN(_03076_ ) );
NOR2_X1 _10813_ ( .A1(_03076_ ), .A2(\myec.state [1] ), .ZN(_03077_ ) );
INV_X1 _10814_ ( .A(\EX_LS_pc [2] ), .ZN(_03078_ ) );
NOR3_X1 _10815_ ( .A1(_01346_ ), .A2(_03077_ ), .A3(_03078_ ), .ZN(_00249_ ) );
NOR2_X1 _10816_ ( .A1(_01346_ ), .A2(_03077_ ), .ZN(_03079_ ) );
AND2_X1 _10817_ ( .A1(_03079_ ), .A2(fanout_net_43 ), .ZN(_00250_ ) );
AOI21_X1 _10818_ ( .A(\LS_WB_waddr_csreg [11] ), .B1(_01302_ ), .B2(\EX_LS_flag [2] ), .ZN(_03080_ ) );
INV_X1 _10819_ ( .A(_01303_ ), .ZN(_03081_ ) );
NOR2_X1 _10820_ ( .A1(_01310_ ), .A2(_03081_ ), .ZN(_03082_ ) );
BUF_X4 _10821_ ( .A(_01207_ ), .Z(_03083_ ) );
NOR2_X1 _10822_ ( .A1(_03083_ ), .A2(\EX_LS_flag [1] ), .ZN(_03084_ ) );
NOR2_X1 _10823_ ( .A1(_03084_ ), .A2(_01289_ ), .ZN(_03085_ ) );
INV_X1 _10824_ ( .A(_03085_ ), .ZN(_03086_ ) );
NOR2_X1 _10825_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_03087_ ) );
AND2_X1 _10826_ ( .A1(_03087_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_03088_ ) );
NOR2_X2 _10827_ ( .A1(_03086_ ), .A2(_03088_ ), .ZN(_03089_ ) );
INV_X1 _10828_ ( .A(_03089_ ), .ZN(_03090_ ) );
OR2_X1 _10829_ ( .A1(_03082_ ), .A2(_03090_ ), .ZN(_03091_ ) );
BUF_X4 _10830_ ( .A(_03091_ ), .Z(_03092_ ) );
BUF_X4 _10831_ ( .A(_03092_ ), .Z(_03093_ ) );
INV_X1 _10832_ ( .A(\EX_LS_dest_csreg_mem [11] ), .ZN(_03094_ ) );
BUF_X4 _10833_ ( .A(_01371_ ), .Z(_03095_ ) );
BUF_X4 _10834_ ( .A(_03095_ ), .Z(_03096_ ) );
BUF_X4 _10835_ ( .A(_03096_ ), .Z(_03097_ ) );
AOI211_X1 _10836_ ( .A(_03080_ ), .B(_03093_ ), .C1(_03094_ ), .C2(_03097_ ), .ZN(_00251_ ) );
INV_X1 _10837_ ( .A(_03082_ ), .ZN(_03098_ ) );
NOR2_X1 _10838_ ( .A1(_01290_ ), .A2(_03088_ ), .ZN(_03099_ ) );
AND2_X1 _10839_ ( .A1(_03098_ ), .A2(_03099_ ), .ZN(_03100_ ) );
INV_X1 _10840_ ( .A(_03100_ ), .ZN(_03101_ ) );
NAND3_X1 _10841_ ( .A1(_01302_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_03102_ ) );
NAND2_X1 _10842_ ( .A1(_03083_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03103_ ) );
AOI21_X1 _10843_ ( .A(_03101_ ), .B1(_03102_ ), .B2(_03103_ ), .ZN(_00252_ ) );
NAND3_X1 _10844_ ( .A1(_01302_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_03104_ ) );
NAND2_X1 _10845_ ( .A1(_03083_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_03105_ ) );
AOI21_X1 _10846_ ( .A(_03101_ ), .B1(_03104_ ), .B2(_03105_ ), .ZN(_00253_ ) );
NAND3_X1 _10847_ ( .A1(_01302_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_03106_ ) );
NAND2_X1 _10848_ ( .A1(_03083_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_03107_ ) );
AOI21_X1 _10849_ ( .A(_03101_ ), .B1(_03106_ ), .B2(_03107_ ), .ZN(_00254_ ) );
NAND3_X1 _10850_ ( .A1(_01302_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_03108_ ) );
NAND2_X1 _10851_ ( .A1(_03083_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03109_ ) );
AOI21_X1 _10852_ ( .A(_03101_ ), .B1(_03108_ ), .B2(_03109_ ), .ZN(_00255_ ) );
NAND3_X1 _10853_ ( .A1(_01302_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_03110_ ) );
NAND2_X1 _10854_ ( .A1(_03083_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_03111_ ) );
AOI21_X1 _10855_ ( .A(_03101_ ), .B1(_03110_ ), .B2(_03111_ ), .ZN(_00256_ ) );
NAND3_X1 _10856_ ( .A1(_01302_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_03112_ ) );
NAND2_X1 _10857_ ( .A1(_03083_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_03113_ ) );
AOI21_X1 _10858_ ( .A(_03101_ ), .B1(_03112_ ), .B2(_03113_ ), .ZN(_00257_ ) );
NAND3_X1 _10859_ ( .A1(_01302_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_flag [2] ), .ZN(_03114_ ) );
NAND2_X1 _10860_ ( .A1(_03083_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_03115_ ) );
AOI21_X1 _10861_ ( .A(_03101_ ), .B1(_03114_ ), .B2(_03115_ ), .ZN(_00258_ ) );
INV_X1 _10862_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_03116_ ) );
AND4_X1 _10863_ ( .A1(_03116_ ), .A2(_01374_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03117_ ) );
NOR2_X1 _10864_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_03118_ ) );
BUF_X2 _10865_ ( .A(_01310_ ), .Z(_03119_ ) );
OAI221_X1 _10866_ ( .A(_03099_ ), .B1(_03117_ ), .B2(_03118_ ), .C1(_03119_ ), .C2(_03081_ ), .ZN(_00259_ ) );
INV_X1 _10867_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_03120_ ) );
AND4_X1 _10868_ ( .A1(_03120_ ), .A2(_01374_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03121_ ) );
NOR2_X1 _10869_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_03122_ ) );
OAI221_X1 _10870_ ( .A(_03099_ ), .B1(_03121_ ), .B2(_03122_ ), .C1(_03119_ ), .C2(_03081_ ), .ZN(_00260_ ) );
NOR4_X1 _10871_ ( .A1(_03083_ ), .A2(_01300_ ), .A3(\EX_LS_dest_csreg_mem [6] ), .A4(\EX_LS_flag [0] ), .ZN(_03123_ ) );
NOR2_X1 _10872_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_03124_ ) );
OAI221_X1 _10873_ ( .A(_03099_ ), .B1(_03123_ ), .B2(_03124_ ), .C1(_03119_ ), .C2(_03081_ ), .ZN(_00261_ ) );
INV_X1 _10874_ ( .A(fanout_net_5 ), .ZN(_03125_ ) );
AND4_X1 _10875_ ( .A1(_03125_ ), .A2(_01374_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03126_ ) );
NOR2_X1 _10876_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_03127_ ) );
OAI221_X1 _10877_ ( .A(_03099_ ), .B1(_03126_ ), .B2(_03127_ ), .C1(_03119_ ), .C2(_03081_ ), .ZN(_00262_ ) );
INV_X1 _10878_ ( .A(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_03128_ ) );
AND2_X1 _10879_ ( .A1(_03079_ ), .A2(_03128_ ), .ZN(_03129_ ) );
NOR2_X1 _10880_ ( .A1(fanout_net_43 ), .A2(\mylsu.state [1] ), .ZN(_03130_ ) );
NAND2_X1 _10881_ ( .A1(_03129_ ), .A2(_03130_ ), .ZN(_03131_ ) );
NOR2_X1 _10882_ ( .A1(_03082_ ), .A2(_03088_ ), .ZN(_03132_ ) );
NAND2_X1 _10883_ ( .A1(\EX_LS_flag [2] ), .A2(\EX_LS_flag [1] ), .ZN(_03133_ ) );
AOI21_X1 _10884_ ( .A(_03131_ ), .B1(_03132_ ), .B2(_03133_ ), .ZN(_03134_ ) );
NOR2_X1 _10885_ ( .A1(_01299_ ), .A2(_03131_ ), .ZN(_03135_ ) );
OR2_X1 _10886_ ( .A1(_03134_ ), .A2(_03135_ ), .ZN(_00263_ ) );
OR2_X1 _10887_ ( .A1(_01299_ ), .A2(_03131_ ), .ZN(_03136_ ) );
INV_X1 _10888_ ( .A(_03132_ ), .ZN(_03137_ ) );
AND2_X1 _10889_ ( .A1(_01289_ ), .A2(\EX_LS_flag [2] ), .ZN(_03138_ ) );
OAI211_X1 _10890_ ( .A(_03128_ ), .B(_03130_ ), .C1(_03137_ ), .C2(_03138_ ), .ZN(_03139_ ) );
BUF_X2 _10891_ ( .A(_03079_ ), .Z(_03140_ ) );
INV_X1 _10892_ ( .A(_03140_ ), .ZN(_03141_ ) );
OAI21_X1 _10893_ ( .A(_03136_ ), .B1(_03139_ ), .B2(_03141_ ), .ZN(_00264_ ) );
AND4_X1 _10894_ ( .A1(_03128_ ), .A2(_03140_ ), .A3(_03138_ ), .A4(_03130_ ), .ZN(_00265_ ) );
BUF_X4 _10895_ ( .A(_03098_ ), .Z(_03142_ ) );
AOI21_X1 _10896_ ( .A(_03131_ ), .B1(_03142_ ), .B2(_01299_ ), .ZN(_00266_ ) );
NOR2_X1 _10897_ ( .A1(_03139_ ), .A2(_03141_ ), .ZN(_00267_ ) );
INV_X1 _10898_ ( .A(_01309_ ), .ZN(_03143_ ) );
INV_X1 _10899_ ( .A(_01298_ ), .ZN(_03144_ ) );
AOI21_X1 _10900_ ( .A(_03144_ ), .B1(_01288_ ), .B2(_01292_ ), .ZN(_03145_ ) );
OR3_X1 _10901_ ( .A1(_03145_ ), .A2(_01304_ ), .A3(_03138_ ), .ZN(_03146_ ) );
AND4_X1 _10902_ ( .A1(_03143_ ), .A2(_03146_ ), .A3(_03130_ ), .A4(_03129_ ), .ZN(_00268_ ) );
INV_X1 _10903_ ( .A(_00250_ ), .ZN(_03147_ ) );
AND3_X1 _10904_ ( .A1(_03140_ ), .A2(EXU_valid_LSU ), .A3(_03130_ ), .ZN(_03148_ ) );
OAI21_X1 _10905_ ( .A(_03148_ ), .B1(_03097_ ), .B2(_01375_ ), .ZN(_03149_ ) );
OAI21_X1 _10906_ ( .A(_03147_ ), .B1(_01304_ ), .B2(_03149_ ), .ZN(_00269_ ) );
INV_X1 _10907_ ( .A(\mysc.state [2] ), .ZN(_03150_ ) );
NOR2_X1 _10908_ ( .A1(_03150_ ), .A2(fanout_net_4 ), .ZN(_00270_ ) );
AND3_X1 _10909_ ( .A1(_00731_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00093_ ) );
CLKBUF_X2 _10910_ ( .A(_01331_ ), .Z(_03151_ ) );
AND2_X1 _10911_ ( .A1(_03151_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y ) );
AND4_X1 _10912_ ( .A1(_02502_ ), .A2(_03151_ ), .A3(_02503_ ), .A4(\myifu.myicache.valid_data_in ), .ZN(_00210_ ) );
AND4_X1 _10913_ ( .A1(_02502_ ), .A2(_03151_ ), .A3(\IF_ID_pc [2] ), .A4(\myifu.myicache.valid_data_in ), .ZN(_00211_ ) );
AND4_X1 _10914_ ( .A1(\IF_ID_pc [3] ), .A2(_03151_ ), .A3(_02503_ ), .A4(\myifu.myicache.valid_data_in ), .ZN(_00212_ ) );
CLKBUF_X2 _10915_ ( .A(_01314_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _10916_ ( .A(_01216_ ), .Z(_03152_ ) );
CLKBUF_X2 _10917_ ( .A(_01217_ ), .Z(_03153_ ) );
NOR3_X1 _10918_ ( .A1(_03152_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(_03153_ ), .ZN(_03154_ ) );
INV_X1 _10919_ ( .A(_02363_ ), .ZN(_03155_ ) );
BUF_X2 _10920_ ( .A(_03155_ ), .Z(_03156_ ) );
BUF_X4 _10921_ ( .A(_03156_ ), .Z(_03157_ ) );
BUF_X4 _10922_ ( .A(_03157_ ), .Z(_03158_ ) );
INV_X1 _10923_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_03159_ ) );
BUF_X4 _10924_ ( .A(_01219_ ), .Z(_03160_ ) );
INV_X1 _10925_ ( .A(_03160_ ), .ZN(_03161_ ) );
AOI211_X1 _10926_ ( .A(_03154_ ), .B(_03158_ ), .C1(_03159_ ), .C2(_03161_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _10927_ ( .A1(_03152_ ), .A2(fanout_net_5 ), .A3(_03153_ ), .ZN(_03162_ ) );
INV_X1 _10928_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_03163_ ) );
AOI211_X1 _10929_ ( .A(_03162_ ), .B(_03158_ ), .C1(_03163_ ), .C2(_03161_ ), .ZN(\io_master_araddr [0] ) );
BUF_X4 _10930_ ( .A(_03158_ ), .Z(_03164_ ) );
OR3_X1 _10931_ ( .A1(_03152_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(_03153_ ), .ZN(_03165_ ) );
OAI21_X1 _10932_ ( .A(_03165_ ), .B1(\mylsu.araddr_tmp [15] ), .B2(_03160_ ), .ZN(_03166_ ) );
BUF_X4 _10933_ ( .A(_01258_ ), .Z(_03167_ ) );
BUF_X4 _10934_ ( .A(_03167_ ), .Z(_03168_ ) );
OAI22_X1 _10935_ ( .A1(_03164_ ), .A2(_03166_ ), .B1(_02818_ ), .B2(_03168_ ), .ZN(\io_master_araddr [15] ) );
AND2_X1 _10936_ ( .A1(_01219_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .ZN(_03169_ ) );
AOI21_X1 _10937_ ( .A(_03169_ ), .B1(\mylsu.araddr_tmp [14] ), .B2(_03161_ ), .ZN(_03170_ ) );
OAI22_X1 _10938_ ( .A1(_03164_ ), .A2(_03170_ ), .B1(_02807_ ), .B2(_03168_ ), .ZN(\io_master_araddr [14] ) );
OR3_X1 _10939_ ( .A1(_03152_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(_03153_ ), .ZN(_03171_ ) );
OAI21_X1 _10940_ ( .A(_03171_ ), .B1(\mylsu.araddr_tmp [5] ), .B2(_03160_ ), .ZN(_03172_ ) );
OAI22_X1 _10941_ ( .A1(_03164_ ), .A2(_03172_ ), .B1(_01022_ ), .B2(_03168_ ), .ZN(\io_master_araddr [5] ) );
OR3_X1 _10942_ ( .A1(_03152_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(_03153_ ), .ZN(_03173_ ) );
OAI21_X1 _10943_ ( .A(_03173_ ), .B1(\mylsu.araddr_tmp [4] ), .B2(_03160_ ), .ZN(_03174_ ) );
OAI22_X1 _10944_ ( .A1(_03164_ ), .A2(_03174_ ), .B1(_02774_ ), .B2(_03168_ ), .ZN(\io_master_araddr [4] ) );
AND2_X1 _10945_ ( .A1(_01219_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .ZN(_03175_ ) );
AOI21_X1 _10946_ ( .A(_03175_ ), .B1(\mylsu.araddr_tmp [3] ), .B2(_03161_ ), .ZN(_03176_ ) );
OAI22_X1 _10947_ ( .A1(_03164_ ), .A2(_03176_ ), .B1(_02502_ ), .B2(_03168_ ), .ZN(\io_master_araddr [3] ) );
OR3_X1 _10948_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(_01217_ ), .ZN(_03177_ ) );
OAI211_X1 _10949_ ( .A(_01215_ ), .B(_03177_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01219_ ), .ZN(_03178_ ) );
OAI221_X1 _10950_ ( .A(\IF_ID_pc [2] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01202_ ), .C2(_01203_ ), .ZN(_03179_ ) );
NAND2_X2 _10951_ ( .A1(_03178_ ), .A2(_03179_ ), .ZN(_03180_ ) );
BUF_X4 _10952_ ( .A(_03180_ ), .Z(_03181_ ) );
BUF_X4 _10953_ ( .A(_03181_ ), .Z(_03182_ ) );
BUF_X4 _10954_ ( .A(_03182_ ), .Z(\io_master_araddr [2] ) );
OR3_X1 _10955_ ( .A1(_03152_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(_03153_ ), .ZN(_03183_ ) );
OAI21_X1 _10956_ ( .A(_03183_ ), .B1(\mylsu.araddr_tmp [13] ), .B2(_03160_ ), .ZN(_03184_ ) );
OAI22_X1 _10957_ ( .A1(_03164_ ), .A2(_03184_ ), .B1(_02506_ ), .B2(_03168_ ), .ZN(\io_master_araddr [13] ) );
INV_X1 _10958_ ( .A(_02356_ ), .ZN(\io_master_araddr [22] ) );
OR3_X1 _10959_ ( .A1(_03152_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(_03153_ ), .ZN(_03185_ ) );
OAI21_X1 _10960_ ( .A(_03185_ ), .B1(\mylsu.araddr_tmp [12] ), .B2(_03160_ ), .ZN(_03186_ ) );
OAI22_X1 _10961_ ( .A1(_03164_ ), .A2(_03186_ ), .B1(_02512_ ), .B2(_03168_ ), .ZN(\io_master_araddr [12] ) );
NOR3_X1 _10962_ ( .A1(_03152_ ), .A2(_03094_ ), .A3(_03153_ ), .ZN(_03187_ ) );
AOI21_X1 _10963_ ( .A(_03187_ ), .B1(_03161_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_03188_ ) );
OAI22_X1 _10964_ ( .A1(_03164_ ), .A2(_03188_ ), .B1(_02513_ ), .B2(_03168_ ), .ZN(\io_master_araddr [11] ) );
OR3_X1 _10965_ ( .A1(_03152_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(_01217_ ), .ZN(_03189_ ) );
OAI21_X1 _10966_ ( .A(_03189_ ), .B1(\mylsu.araddr_tmp [10] ), .B2(_03160_ ), .ZN(_03190_ ) );
OAI22_X1 _10967_ ( .A1(_03164_ ), .A2(_03190_ ), .B1(_02514_ ), .B2(_03168_ ), .ZN(\io_master_araddr [10] ) );
NOR3_X1 _10968_ ( .A1(_03152_ ), .A2(_03116_ ), .A3(_03153_ ), .ZN(_03191_ ) );
AOI21_X1 _10969_ ( .A(_03191_ ), .B1(_03161_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_03192_ ) );
OAI22_X1 _10970_ ( .A1(_03164_ ), .A2(_03192_ ), .B1(_02516_ ), .B2(_03168_ ), .ZN(\io_master_araddr [9] ) );
OR3_X1 _10971_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [8] ), .A3(_01217_ ), .ZN(_03193_ ) );
OAI21_X1 _10972_ ( .A(_03193_ ), .B1(\mylsu.araddr_tmp [8] ), .B2(_03160_ ), .ZN(_03194_ ) );
OAI22_X1 _10973_ ( .A1(_03158_ ), .A2(_03194_ ), .B1(_02800_ ), .B2(_03167_ ), .ZN(\io_master_araddr [8] ) );
OR3_X1 _10974_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(_01217_ ), .ZN(_03195_ ) );
OAI21_X1 _10975_ ( .A(_03195_ ), .B1(\mylsu.araddr_tmp [7] ), .B2(_03160_ ), .ZN(_03196_ ) );
OAI22_X1 _10976_ ( .A1(_03158_ ), .A2(_03196_ ), .B1(_01056_ ), .B2(_03167_ ), .ZN(\io_master_araddr [7] ) );
OR3_X1 _10977_ ( .A1(_01216_ ), .A2(\EX_LS_dest_csreg_mem [6] ), .A3(_01217_ ), .ZN(_03197_ ) );
OAI21_X1 _10978_ ( .A(_03197_ ), .B1(\mylsu.araddr_tmp [6] ), .B2(_03160_ ), .ZN(_03198_ ) );
OAI22_X1 _10979_ ( .A1(_03158_ ), .A2(_03198_ ), .B1(_02517_ ), .B2(_03167_ ), .ZN(\io_master_araddr [6] ) );
NOR3_X1 _10980_ ( .A1(\io_master_arburst [0] ), .A2(_01281_ ), .A3(_01213_ ), .ZN(\io_master_arsize [2] ) );
NOR3_X1 _10981_ ( .A1(\io_master_arburst [0] ), .A2(_01280_ ), .A3(_01213_ ), .ZN(\io_master_arsize [0] ) );
INV_X1 _10982_ ( .A(\EX_LS_typ [2] ), .ZN(_03199_ ) );
OAI22_X1 _10983_ ( .A1(_01204_ ), .A2(_01205_ ), .B1(_03199_ ), .B2(_01213_ ), .ZN(\io_master_arsize [1] ) );
BUF_X4 _10984_ ( .A(_02359_ ), .Z(_03200_ ) );
CLKBUF_X2 _10985_ ( .A(_03200_ ), .Z(_03201_ ) );
BUF_X2 _10986_ ( .A(_03201_ ), .Z(_03202_ ) );
NOR3_X1 _10987_ ( .A1(_03202_ ), .A2(_01330_ ), .A3(_01332_ ), .ZN(io_master_arvalid ) );
AND2_X1 _10988_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ) );
AND2_X1 _10989_ ( .A1(_01303_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_03203_ ) );
BUF_X4 _10990_ ( .A(_03203_ ), .Z(_03204_ ) );
BUF_X4 _10991_ ( .A(_03204_ ), .Z(_03205_ ) );
MUX2_X1 _10992_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_03205_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _10993_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_03205_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _10994_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_03205_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _10995_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_03205_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _10996_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_03205_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _10997_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_03205_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _10998_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_03205_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _10999_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_03205_ ), .Z(\io_master_awaddr [16] ) );
BUF_X4 _11000_ ( .A(_03204_ ), .Z(_03206_ ) );
MUX2_X1 _11001_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_03206_ ), .Z(\io_master_awaddr [15] ) );
MUX2_X1 _11002_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_03206_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _11003_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_03206_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _11004_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_03206_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _11005_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_03206_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _11006_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_03206_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _11007_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_03206_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _11008_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_03206_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _11009_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_03206_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _11010_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_03206_ ), .Z(\io_master_awaddr [7] ) );
BUF_X4 _11011_ ( .A(_03204_ ), .Z(_03207_ ) );
MUX2_X1 _11012_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_03207_ ), .Z(\io_master_awaddr [6] ) );
MUX2_X1 _11013_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_03207_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _11014_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_03207_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _11015_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_03207_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _11016_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_03207_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _11017_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_03207_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _11018_ ( .A(\mylsu.awaddr_tmp [1] ), .B(\EX_LS_dest_csreg_mem [1] ), .S(_03207_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _11019_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_5 ), .S(_03207_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _11020_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_03207_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _11021_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_03207_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _11022_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_03204_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _11023_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_03204_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _11024_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_03204_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _11025_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_03204_ ), .Z(\io_master_awaddr [22] ) );
NAND3_X1 _11026_ ( .A1(_01291_ ), .A2(_01374_ ), .A3(\EX_LS_flag [1] ), .ZN(_03208_ ) );
NOR2_X1 _11027_ ( .A1(_03208_ ), .A2(\EX_LS_flag [2] ), .ZN(_03209_ ) );
AND4_X1 _11028_ ( .A1(\EX_LS_typ [1] ), .A2(_03209_ ), .A3(\EX_LS_typ [0] ), .A4(_01284_ ), .ZN(\io_master_awsize [0] ) );
NAND3_X1 _11029_ ( .A1(_03209_ ), .A2(\EX_LS_typ [0] ), .A3(_01284_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _11030_ ( .A1(_01299_ ), .A2(_03119_ ), .A3(_03205_ ), .ZN(_03210_ ) );
INV_X1 _11031_ ( .A(\mylsu.state [4] ), .ZN(_03211_ ) );
NAND2_X1 _11032_ ( .A1(_03210_ ), .A2(_03211_ ), .ZN(io_master_awvalid ) );
INV_X1 _11033_ ( .A(\mylsu.state [2] ), .ZN(_03212_ ) );
INV_X1 _11034_ ( .A(\mylsu.state [1] ), .ZN(_03213_ ) );
NAND4_X1 _11035_ ( .A1(_03210_ ), .A2(_03212_ ), .A3(_03211_ ), .A4(_03213_ ), .ZN(io_master_bready ) );
NOR3_X1 _11036_ ( .A1(_01212_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_03214_ ) );
NAND2_X1 _11037_ ( .A1(\io_master_bid [1] ), .A2(\io_master_bid [0] ), .ZN(_03215_ ) );
OR3_X1 _11038_ ( .A1(_03215_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bid [2] ), .ZN(_03216_ ) );
NOR2_X1 _11039_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_03217_ ) );
NAND2_X1 _11040_ ( .A1(_03217_ ), .A2(io_master_bvalid ), .ZN(_03218_ ) );
OR2_X1 _11041_ ( .A1(_03216_ ), .A2(_03218_ ), .ZN(_03219_ ) );
OR2_X2 _11042_ ( .A1(_01329_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .ZN(_03220_ ) );
NAND2_X1 _11043_ ( .A1(_01329_ ), .A2(io_master_rvalid ), .ZN(_03221_ ) );
AND2_X1 _11044_ ( .A1(_03220_ ), .A2(_03221_ ), .ZN(_03222_ ) );
INV_X1 _11045_ ( .A(_03222_ ), .ZN(_03223_ ) );
AND2_X1 _11046_ ( .A1(_01248_ ), .A2(_01276_ ), .ZN(_03224_ ) );
NOR2_X1 _11047_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_03225_ ) );
NOR2_X1 _11048_ ( .A1(_03224_ ), .A2(_03225_ ), .ZN(_03226_ ) );
INV_X1 _11049_ ( .A(_03224_ ), .ZN(_03227_ ) );
NOR2_X1 _11050_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_03228_ ) );
INV_X1 _11051_ ( .A(\io_master_rid [0] ), .ZN(_03229_ ) );
NAND4_X1 _11052_ ( .A1(_03228_ ), .A2(\io_master_rid [1] ), .A3(_03229_ ), .A4(io_master_rlast ), .ZN(_03230_ ) );
AOI21_X1 _11053_ ( .A(_03226_ ), .B1(_03227_ ), .B2(_03230_ ), .ZN(_03231_ ) );
AND3_X1 _11054_ ( .A1(_03223_ ), .A2(\io_master_arid [1] ), .A3(_03231_ ), .ZN(_03232_ ) );
INV_X1 _11055_ ( .A(_03232_ ), .ZN(_03233_ ) );
AOI221_X4 _11056_ ( .A(_03214_ ), .B1(\mylsu.state [1] ), .B2(_03219_ ), .C1(_03233_ ), .C2(fanout_net_43 ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
NOR3_X1 _11057_ ( .A1(_03202_ ), .A2(_01313_ ), .A3(_01318_ ), .ZN(io_master_rready ) );
MUX2_X1 _11058_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_5 ), .Z(_03234_ ) );
INV_X1 _11059_ ( .A(\EX_LS_dest_csreg_mem [1] ), .ZN(_03235_ ) );
CLKBUF_X2 _11060_ ( .A(_03235_ ), .Z(_03236_ ) );
AND2_X1 _11061_ ( .A1(_03234_ ), .A2(_03236_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _11062_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_5 ), .Z(_03237_ ) );
AND2_X1 _11063_ ( .A1(_03237_ ), .A2(_03236_ ), .ZN(\io_master_wdata [14] ) );
INV_X1 _11064_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_03238_ ) );
NOR3_X1 _11065_ ( .A1(_03238_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [5] ) );
INV_X1 _11066_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_03239_ ) );
NOR3_X1 _11067_ ( .A1(_03239_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [4] ) );
INV_X1 _11068_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_03240_ ) );
NOR3_X1 _11069_ ( .A1(_03240_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [3] ) );
INV_X1 _11070_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_03241_ ) );
NOR3_X1 _11071_ ( .A1(_03241_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _11072_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_03242_ ) );
NOR3_X1 _11073_ ( .A1(_03242_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _11074_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_03243_ ) );
NOR3_X1 _11075_ ( .A1(_03243_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _11076_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_5 ), .Z(_03244_ ) );
AND2_X1 _11077_ ( .A1(_03244_ ), .A2(_03236_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _11078_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_5 ), .Z(_03245_ ) );
AND2_X1 _11079_ ( .A1(_03245_ ), .A2(_03236_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _11080_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_5 ), .Z(_03246_ ) );
AND2_X1 _11081_ ( .A1(_03246_ ), .A2(_03236_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _11082_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_5 ), .Z(_03247_ ) );
AND2_X1 _11083_ ( .A1(_03247_ ), .A2(_03236_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _11084_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_5 ), .Z(_03248_ ) );
AND2_X1 _11085_ ( .A1(_03248_ ), .A2(_03236_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _11086_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_5 ), .Z(_03249_ ) );
AND2_X1 _11087_ ( .A1(_03249_ ), .A2(_03236_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _11088_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_03250_ ) );
NOR3_X1 _11089_ ( .A1(_03250_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [7] ) );
INV_X1 _11090_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_03251_ ) );
NOR3_X1 _11091_ ( .A1(_03251_ ), .A2(fanout_net_5 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _11092_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_5 ), .Z(_03252_ ) );
MUX2_X1 _11093_ ( .A(_03252_ ), .B(_03234_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _11094_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_5 ), .Z(_03253_ ) );
MUX2_X1 _11095_ ( .A(_03253_ ), .B(_03237_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [30] ) );
BUF_X4 _11096_ ( .A(_03235_ ), .Z(_03254_ ) );
NOR2_X1 _11097_ ( .A1(_03254_ ), .A2(fanout_net_5 ), .ZN(_03255_ ) );
INV_X1 _11098_ ( .A(_03255_ ), .ZN(_03256_ ) );
BUF_X2 _11099_ ( .A(_03125_ ), .Z(_03257_ ) );
OAI21_X1 _11100_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [13] ), .ZN(_03258_ ) );
NOR2_X1 _11101_ ( .A1(fanout_net_5 ), .A2(\EX_LS_result_csreg_mem [21] ), .ZN(_03259_ ) );
OAI22_X1 _11102_ ( .A1(_03256_ ), .A2(_03238_ ), .B1(_03258_ ), .B2(_03259_ ), .ZN(\io_master_wdata [21] ) );
OAI21_X1 _11103_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [12] ), .ZN(_03260_ ) );
NOR2_X1 _11104_ ( .A1(fanout_net_5 ), .A2(\EX_LS_result_csreg_mem [20] ), .ZN(_03261_ ) );
OAI22_X1 _11105_ ( .A1(_03256_ ), .A2(_03239_ ), .B1(_03260_ ), .B2(_03261_ ), .ZN(\io_master_wdata [20] ) );
OAI21_X1 _11106_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_03262_ ) );
NOR2_X1 _11107_ ( .A1(fanout_net_5 ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_03263_ ) );
OAI22_X1 _11108_ ( .A1(_03256_ ), .A2(_03240_ ), .B1(_03262_ ), .B2(_03263_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _11109_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_03264_ ) );
NOR2_X1 _11110_ ( .A1(fanout_net_5 ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_03265_ ) );
OAI22_X1 _11111_ ( .A1(_03256_ ), .A2(_03241_ ), .B1(_03264_ ), .B2(_03265_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _11112_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_03266_ ) );
NOR2_X1 _11113_ ( .A1(fanout_net_5 ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_03267_ ) );
OAI22_X1 _11114_ ( .A1(_03256_ ), .A2(_03242_ ), .B1(_03266_ ), .B2(_03267_ ), .ZN(\io_master_wdata [17] ) );
OAI21_X1 _11115_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [8] ), .ZN(_03268_ ) );
NOR2_X1 _11116_ ( .A1(fanout_net_5 ), .A2(\EX_LS_result_csreg_mem [16] ), .ZN(_03269_ ) );
OAI22_X1 _11117_ ( .A1(_03256_ ), .A2(_03243_ ), .B1(_03268_ ), .B2(_03269_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _11118_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03270_ ) );
MUX2_X1 _11119_ ( .A(_03270_ ), .B(_03244_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _11120_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03271_ ) );
MUX2_X1 _11121_ ( .A(_03271_ ), .B(_03245_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _11122_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03272_ ) );
MUX2_X1 _11123_ ( .A(_03272_ ), .B(_03246_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _11124_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03273_ ) );
MUX2_X1 _11125_ ( .A(_03273_ ), .B(_03247_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _11126_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03274_ ) );
MUX2_X1 _11127_ ( .A(_03274_ ), .B(_03248_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _11128_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03275_ ) );
MUX2_X1 _11129_ ( .A(_03275_ ), .B(_03249_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [24] ) );
OAI21_X1 _11130_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [15] ), .ZN(_03276_ ) );
NOR2_X1 _11131_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [23] ), .ZN(_03277_ ) );
OAI22_X1 _11132_ ( .A1(_03256_ ), .A2(_03250_ ), .B1(_03276_ ), .B2(_03277_ ), .ZN(\io_master_wdata [23] ) );
OAI21_X1 _11133_ ( .A(_03254_ ), .B1(_03257_ ), .B2(\EX_LS_result_csreg_mem [14] ), .ZN(_03278_ ) );
NOR2_X1 _11134_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [22] ), .ZN(_03279_ ) );
OAI22_X1 _11135_ ( .A1(_03256_ ), .A2(_03251_ ), .B1(_03278_ ), .B2(_03279_ ), .ZN(\io_master_wdata [22] ) );
NAND2_X1 _11136_ ( .A1(_01303_ ), .A2(EXU_valid_LSU ), .ZN(_03280_ ) );
INV_X1 _11137_ ( .A(io_master_wready ), .ZN(_03281_ ) );
AOI211_X1 _11138_ ( .A(io_master_wready_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ), .B(_03280_ ), .C1(_03281_ ), .C2(_02369_ ), .ZN(_03282_ ) );
AND3_X1 _11139_ ( .A1(_03119_ ), .A2(_03140_ ), .A3(_03282_ ), .ZN(io_master_wready_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _11140_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03283_ ) );
AND2_X1 _11141_ ( .A1(_03283_ ), .A2(_03236_ ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _11142_ ( .A1(_03257_ ), .A2(_03236_ ), .A3(\EX_LS_typ [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _11143_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_03284_ ) );
MUX2_X1 _11144_ ( .A(_03284_ ), .B(_03283_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _11145_ ( .A1(_03254_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_03285_ ) );
NAND3_X1 _11146_ ( .A1(_03257_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_typ [0] ), .ZN(_03286_ ) );
OAI211_X1 _11147_ ( .A(_03285_ ), .B(_03286_ ), .C1(_01279_ ), .C2(_03199_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _11148_ ( .A1(_03210_ ), .A2(_03212_ ), .ZN(io_master_wvalid ) );
MUX2_X1 _11149_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _11150_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _11151_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _11152_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
NOR2_X1 _11153_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03287_ ) );
INV_X1 _11154_ ( .A(\LS_WB_waddr_csreg [7] ), .ZN(_03288_ ) );
INV_X1 _11155_ ( .A(\LS_WB_waddr_csreg [6] ), .ZN(_03289_ ) );
NAND3_X1 _11156_ ( .A1(_03287_ ), .A2(_03288_ ), .A3(_03289_ ), .ZN(_03290_ ) );
OR2_X1 _11157_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03291_ ) );
NAND2_X1 _11158_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_03292_ ) );
NOR3_X1 _11159_ ( .A1(_03290_ ), .A2(_03291_ ), .A3(_03292_ ), .ZN(_03293_ ) );
AND2_X1 _11160_ ( .A1(_00731_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(_03294_ ) );
INV_X1 _11161_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_03295_ ) );
NOR3_X1 _11162_ ( .A1(_03295_ ), .A2(\LS_WB_waddr_csreg [3] ), .A3(\LS_WB_waddr_csreg [1] ), .ZN(_03296_ ) );
AND4_X1 _11163_ ( .A1(\LS_WB_waddr_csreg [2] ), .A2(_03293_ ), .A3(_03294_ ), .A4(_03296_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ) );
AND3_X1 _11164_ ( .A1(_03287_ ), .A2(_03288_ ), .A3(\LS_WB_waddr_csreg [6] ), .ZN(_03297_ ) );
NOR2_X1 _11165_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_03298_ ) );
AND2_X1 _11166_ ( .A1(_03297_ ), .A2(_03298_ ), .ZN(_03299_ ) );
INV_X1 _11167_ ( .A(_03299_ ), .ZN(_03300_ ) );
NOR2_X1 _11168_ ( .A1(_03291_ ), .A2(_03292_ ), .ZN(_03301_ ) );
NAND2_X1 _11169_ ( .A1(_03301_ ), .A2(_03294_ ), .ZN(_03302_ ) );
NOR4_X1 _11170_ ( .A1(_03300_ ), .A2(\LS_WB_waddr_csreg [1] ), .A3(_03295_ ), .A4(_03302_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ) );
AND3_X1 _11171_ ( .A1(_03297_ ), .A2(_03301_ ), .A3(_03298_ ), .ZN(_03303_ ) );
AND4_X1 _11172_ ( .A1(\LS_WB_waddr_csreg [1] ), .A2(_03303_ ), .A3(_03295_ ), .A4(_03294_ ), .ZN(_03304_ ) );
OR2_X1 _11173_ ( .A1(_03304_ ), .A2(_00093_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OR3_X1 _11174_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .A3(\LS_WB_waddr_csreg [1] ), .ZN(_03305_ ) );
NOR4_X1 _11175_ ( .A1(_03302_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(_03290_ ), .A4(_03305_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
MUX2_X1 _11176_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _11177_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _11178_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _11179_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _11180_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _11181_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _11182_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _11183_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_01344_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
BUF_X4 _11184_ ( .A(_01312_ ), .Z(_03306_ ) );
MUX2_X1 _11185_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _11186_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
MUX2_X1 _11187_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _11188_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _11189_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _11190_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _11191_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _11192_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _11193_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _11194_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_03306_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
BUF_X4 _11195_ ( .A(_01312_ ), .Z(_03307_ ) );
MUX2_X1 _11196_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _11197_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
MUX2_X1 _11198_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _11199_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _11200_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _11201_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _11202_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _11203_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _11204_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _11205_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_03307_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _11206_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_01312_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _11207_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_01312_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _11208_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_01312_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _11209_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_01312_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
NAND4_X1 _11210_ ( .A1(_01299_ ), .A2(_01340_ ), .A3(_03119_ ), .A4(_01342_ ), .ZN(_03308_ ) );
XNOR2_X1 _11211_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_03309_ ) );
XNOR2_X1 _11212_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_03310_ ) );
XNOR2_X1 _11213_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_03311_ ) );
XNOR2_X1 _11214_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_03312_ ) );
AND4_X1 _11215_ ( .A1(_03309_ ), .A2(_03310_ ), .A3(_03311_ ), .A4(_03312_ ), .ZN(_03313_ ) );
XNOR2_X1 _11216_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_03314_ ) );
XNOR2_X1 _11217_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_03315_ ) );
XNOR2_X1 _11218_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_03316_ ) );
XNOR2_X1 _11219_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_03317_ ) );
AND4_X1 _11220_ ( .A1(_03314_ ), .A2(_03315_ ), .A3(_03316_ ), .A4(_03317_ ), .ZN(_03318_ ) );
XNOR2_X1 _11221_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_03319_ ) );
XNOR2_X1 _11222_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_03320_ ) );
XNOR2_X1 _11223_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_03321_ ) );
XNOR2_X1 _11224_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_03322_ ) );
AND4_X1 _11225_ ( .A1(_03319_ ), .A2(_03320_ ), .A3(_03321_ ), .A4(_03322_ ), .ZN(_03323_ ) );
XNOR2_X1 _11226_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_03324_ ) );
XNOR2_X1 _11227_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_03325_ ) );
XNOR2_X1 _11228_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_03326_ ) );
XNOR2_X1 _11229_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_03327_ ) );
AND4_X1 _11230_ ( .A1(_03324_ ), .A2(_03325_ ), .A3(_03326_ ), .A4(_03327_ ), .ZN(_03328_ ) );
AND4_X1 _11231_ ( .A1(_03313_ ), .A2(_03318_ ), .A3(_03323_ ), .A4(_03328_ ), .ZN(_03329_ ) );
XNOR2_X1 _11232_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_03330_ ) );
XNOR2_X1 _11233_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_03331_ ) );
XNOR2_X1 _11234_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_03332_ ) );
XNOR2_X1 _11235_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_03333_ ) );
AND4_X1 _11236_ ( .A1(_03330_ ), .A2(_03331_ ), .A3(_03332_ ), .A4(_03333_ ), .ZN(_03334_ ) );
XNOR2_X1 _11237_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_03335_ ) );
XNOR2_X1 _11238_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_03336_ ) );
XNOR2_X1 _11239_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_03337_ ) );
XNOR2_X1 _11240_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_03338_ ) );
AND4_X1 _11241_ ( .A1(_03335_ ), .A2(_03336_ ), .A3(_03337_ ), .A4(_03338_ ), .ZN(_03339_ ) );
XNOR2_X1 _11242_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_03340_ ) );
XNOR2_X1 _11243_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_03341_ ) );
XNOR2_X1 _11244_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_03342_ ) );
XNOR2_X1 _11245_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_03343_ ) );
AND4_X1 _11246_ ( .A1(_03340_ ), .A2(_03341_ ), .A3(_03342_ ), .A4(_03343_ ), .ZN(_03344_ ) );
XNOR2_X1 _11247_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_03345_ ) );
XNOR2_X1 _11248_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_03346_ ) );
XNOR2_X1 _11249_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_03347_ ) );
XNOR2_X1 _11250_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_03348_ ) );
AND4_X1 _11251_ ( .A1(_03345_ ), .A2(_03346_ ), .A3(_03347_ ), .A4(_03348_ ), .ZN(_03349_ ) );
AND4_X1 _11252_ ( .A1(_03334_ ), .A2(_03339_ ), .A3(_03344_ ), .A4(_03349_ ), .ZN(_03350_ ) );
NAND3_X1 _11253_ ( .A1(_03329_ ), .A2(_03350_ ), .A3(excp_written ), .ZN(_03351_ ) );
OAI21_X1 _11254_ ( .A(_03351_ ), .B1(\myec.state [0] ), .B2(\myec.state [1] ), .ZN(_03352_ ) );
AND2_X1 _11255_ ( .A1(_03308_ ), .A2(_03352_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _11256_ ( .A1(_02502_ ), .A2(_03151_ ), .A3(_02503_ ), .A4(\myifu.myicache.valid_data_in ), .ZN(\myexu.check_quest_$_NAND__B_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_AND__A_Y ) );
NAND2_X1 _11257_ ( .A1(_01597_ ), .A2(_02284_ ), .ZN(_03353_ ) );
NOR2_X1 _11258_ ( .A1(_01574_ ), .A2(_01596_ ), .ZN(_03354_ ) );
INV_X1 _11259_ ( .A(\ID_EX_csr [1] ), .ZN(_03355_ ) );
INV_X2 _11260_ ( .A(_01365_ ), .ZN(_03356_ ) );
BUF_X4 _11261_ ( .A(_03356_ ), .Z(_03357_ ) );
BUF_X4 _11262_ ( .A(_03357_ ), .Z(_03358_ ) );
OAI22_X1 _11263_ ( .A1(_03353_ ), .A2(_03354_ ), .B1(_03355_ ), .B2(_03358_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
NAND2_X4 _11264_ ( .A1(_01576_ ), .A2(_01595_ ), .ZN(_03359_ ) );
XNOR2_X1 _11265_ ( .A(_03359_ ), .B(\ID_EX_imm [0] ), .ZN(_03360_ ) );
INV_X1 _11266_ ( .A(_01367_ ), .ZN(_03361_ ) );
BUF_X4 _11267_ ( .A(_03361_ ), .Z(_03362_ ) );
NAND2_X1 _11268_ ( .A1(_03360_ ), .A2(_03362_ ), .ZN(_03363_ ) );
BUF_X4 _11269_ ( .A(_03356_ ), .Z(_03364_ ) );
MUX2_X1 _11270_ ( .A(\ID_EX_csr [0] ), .B(_03363_ ), .S(_03364_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
OAI21_X1 _11271_ ( .A(_01860_ ), .B1(_01711_ ), .B2(_01716_ ), .ZN(_03365_ ) );
OR3_X1 _11272_ ( .A1(_01855_ ), .A2(_01858_ ), .A3(_01914_ ), .ZN(_03366_ ) );
AND3_X1 _11273_ ( .A1(_03365_ ), .A2(_01856_ ), .A3(_03366_ ), .ZN(_03367_ ) );
INV_X1 _11274_ ( .A(_03367_ ), .ZN(_03368_ ) );
OR2_X1 _11275_ ( .A1(_03368_ ), .A2(_01906_ ), .ZN(_03369_ ) );
BUF_X4 _11276_ ( .A(_03361_ ), .Z(_03370_ ) );
NAND2_X1 _11277_ ( .A1(_03368_ ), .A2(_01906_ ), .ZN(_03371_ ) );
AND3_X1 _11278_ ( .A1(_03369_ ), .A2(_03370_ ), .A3(_03371_ ), .ZN(_03372_ ) );
MUX2_X1 _11279_ ( .A(\ID_EX_csr [10] ), .B(_03372_ ), .S(_03364_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
OAI21_X1 _11280_ ( .A(_01833_ ), .B1(_01711_ ), .B2(_01716_ ), .ZN(_03373_ ) );
AND2_X1 _11281_ ( .A1(_03373_ ), .A2(_01914_ ), .ZN(_03374_ ) );
XNOR2_X1 _11282_ ( .A(_01854_ ), .B(\ID_EX_imm [9] ), .ZN(_03375_ ) );
XNOR2_X1 _11283_ ( .A(_03374_ ), .B(_03375_ ), .ZN(_03376_ ) );
INV_X1 _11284_ ( .A(\ID_EX_csr [9] ), .ZN(_03377_ ) );
BUF_X4 _11285_ ( .A(_01365_ ), .Z(_03378_ ) );
BUF_X4 _11286_ ( .A(_03378_ ), .Z(_03379_ ) );
AOI22_X1 _11287_ ( .A1(_03376_ ), .A2(_02284_ ), .B1(_03377_ ), .B2(_03379_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
XOR2_X1 _11288_ ( .A(_01717_ ), .B(_01833_ ), .Z(_03380_ ) );
INV_X1 _11289_ ( .A(\ID_EX_csr [8] ), .ZN(_03381_ ) );
AOI22_X1 _11290_ ( .A1(_03380_ ), .A2(_02284_ ), .B1(_03381_ ), .B2(_03379_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
OAI21_X1 _11291_ ( .A(_01709_ ), .B1(_01659_ ), .B2(_01661_ ), .ZN(_03382_ ) );
INV_X1 _11292_ ( .A(_01712_ ), .ZN(_03383_ ) );
AND3_X1 _11293_ ( .A1(_03382_ ), .A2(_03383_ ), .A3(_01686_ ), .ZN(_03384_ ) );
AOI21_X1 _11294_ ( .A(_01686_ ), .B1(_03382_ ), .B2(_03383_ ), .ZN(_03385_ ) );
OR3_X1 _11295_ ( .A1(_03384_ ), .A2(_03385_ ), .A3(_01369_ ), .ZN(_03386_ ) );
INV_X1 _11296_ ( .A(\ID_EX_csr [7] ), .ZN(_03387_ ) );
OAI21_X1 _11297_ ( .A(_03386_ ), .B1(_03387_ ), .B2(_03358_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
XNOR2_X1 _11298_ ( .A(_01662_ ), .B(_01710_ ), .ZN(_03388_ ) );
NAND2_X1 _11299_ ( .A1(_03388_ ), .A2(_03362_ ), .ZN(_03389_ ) );
BUF_X4 _11300_ ( .A(_03356_ ), .Z(_03390_ ) );
MUX2_X1 _11301_ ( .A(\ID_EX_csr [6] ), .B(_03389_ ), .S(_03390_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
AND2_X1 _11302_ ( .A1(_01632_ ), .A2(_01658_ ), .ZN(_03391_ ) );
OR3_X1 _11303_ ( .A1(_03391_ ), .A2(_01659_ ), .A3(_01369_ ), .ZN(_03392_ ) );
INV_X1 _11304_ ( .A(\ID_EX_csr [5] ), .ZN(_03393_ ) );
OAI21_X1 _11305_ ( .A(_03392_ ), .B1(_03393_ ), .B2(_03358_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND2_X4 _11306_ ( .A1(_01607_ ), .A2(_01628_ ), .ZN(_03394_ ) );
XNOR2_X1 _11307_ ( .A(_03394_ ), .B(_01604_ ), .ZN(_03395_ ) );
NOR3_X1 _11308_ ( .A1(_01598_ ), .A2(_01602_ ), .A3(_03395_ ), .ZN(_03396_ ) );
NOR3_X1 _11309_ ( .A1(_01631_ ), .A2(_01367_ ), .A3(_03396_ ), .ZN(_03397_ ) );
MUX2_X1 _11310_ ( .A(\ID_EX_csr [4] ), .B(_03397_ ), .S(_03390_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
AND2_X1 _11311_ ( .A1(_01597_ ), .A2(_01572_ ), .ZN(_03398_ ) );
OR2_X1 _11312_ ( .A1(_03398_ ), .A2(_01550_ ), .ZN(_03399_ ) );
AND3_X1 _11313_ ( .A1(_03399_ ), .A2(_01599_ ), .A3(_01523_ ), .ZN(_03400_ ) );
AOI21_X1 _11314_ ( .A(_01523_ ), .B1(_03399_ ), .B2(_01599_ ), .ZN(_03401_ ) );
OR3_X1 _11315_ ( .A1(_03400_ ), .A2(_03401_ ), .A3(_01369_ ), .ZN(_03402_ ) );
INV_X1 _11316_ ( .A(\ID_EX_csr [3] ), .ZN(_03403_ ) );
OAI21_X1 _11317_ ( .A(_03402_ ), .B1(_03403_ ), .B2(_03358_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
OAI21_X1 _11318_ ( .A(_02284_ ), .B1(_03398_ ), .B2(_01550_ ), .ZN(_03404_ ) );
AND3_X1 _11319_ ( .A1(_01597_ ), .A2(_01572_ ), .A3(_01550_ ), .ZN(_03405_ ) );
INV_X1 _11320_ ( .A(\ID_EX_csr [2] ), .ZN(_03406_ ) );
BUF_X4 _11321_ ( .A(_03357_ ), .Z(_03407_ ) );
OAI22_X1 _11322_ ( .A1(_03404_ ), .A2(_03405_ ), .B1(_03406_ ), .B2(_03407_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
INV_X1 _11323_ ( .A(_01917_ ), .ZN(_03408_ ) );
INV_X1 _11324_ ( .A(_01884_ ), .ZN(_03409_ ) );
NAND3_X1 _11325_ ( .A1(_03371_ ), .A2(_03408_ ), .A3(_03409_ ), .ZN(_03410_ ) );
NAND2_X1 _11326_ ( .A1(_03410_ ), .A2(_02284_ ), .ZN(_03411_ ) );
AOI21_X1 _11327_ ( .A(_03409_ ), .B1(_03371_ ), .B2(_03408_ ), .ZN(_03412_ ) );
INV_X1 _11328_ ( .A(\ID_EX_csr [11] ), .ZN(_03413_ ) );
OAI22_X1 _11329_ ( .A1(_03411_ ), .A2(_03412_ ), .B1(_03413_ ), .B2(_03407_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
AOI22_X1 _11330_ ( .A1(\EX_LS_dest_csreg_mem [9] ), .A2(_03377_ ), .B1(_03381_ ), .B2(\EX_LS_dest_csreg_mem [8] ), .ZN(_03414_ ) );
AOI22_X1 _11331_ ( .A1(_03116_ ), .A2(\ID_EX_csr [9] ), .B1(_03120_ ), .B2(\ID_EX_csr [8] ), .ZN(_03415_ ) );
XNOR2_X1 _11332_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .ZN(_03416_ ) );
AND4_X1 _11333_ ( .A1(_03095_ ), .A2(_03414_ ), .A3(_03415_ ), .A4(_03416_ ), .ZN(_03417_ ) );
XNOR2_X1 _11334_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_03418_ ) );
XNOR2_X1 _11335_ ( .A(\EX_LS_dest_csreg_mem [1] ), .B(\ID_EX_csr [1] ), .ZN(_03419_ ) );
XNOR2_X1 _11336_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_03420_ ) );
XNOR2_X1 _11337_ ( .A(\EX_LS_dest_csreg_mem [0] ), .B(\ID_EX_csr [0] ), .ZN(_03421_ ) );
AND4_X1 _11338_ ( .A1(_03418_ ), .A2(_03419_ ), .A3(_03420_ ), .A4(_03421_ ), .ZN(_03422_ ) );
NAND2_X1 _11339_ ( .A1(_03417_ ), .A2(_03422_ ), .ZN(_03423_ ) );
CLKBUF_X2 _11340_ ( .A(_03423_ ), .Z(_03424_ ) );
XNOR2_X1 _11341_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_03425_ ) );
XNOR2_X1 _11342_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_03426_ ) );
AND2_X1 _11343_ ( .A1(_03425_ ), .A2(_03426_ ), .ZN(_03427_ ) );
XNOR2_X1 _11344_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_03428_ ) );
XNOR2_X1 _11345_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_03429_ ) );
XNOR2_X1 _11346_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_03430_ ) );
NAND4_X1 _11347_ ( .A1(_03427_ ), .A2(_03428_ ), .A3(_03429_ ), .A4(_03430_ ), .ZN(_03431_ ) );
CLKBUF_X2 _11348_ ( .A(_03431_ ), .Z(_03432_ ) );
NOR3_X1 _11349_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [21] ), .A3(_03432_ ), .ZN(_03433_ ) );
INV_X1 _11350_ ( .A(_03433_ ), .ZN(_03434_ ) );
AND4_X1 _11351_ ( .A1(\ID_EX_csr [10] ), .A2(_03393_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_03435_ ) );
AND2_X1 _11352_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_03436_ ) );
NOR2_X1 _11353_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_03437_ ) );
AND3_X1 _11354_ ( .A1(_03435_ ), .A2(_03436_ ), .A3(_03437_ ), .ZN(_03438_ ) );
NAND3_X1 _11355_ ( .A1(_03355_ ), .A2(_03403_ ), .A3(\ID_EX_csr [0] ), .ZN(_03439_ ) );
NOR2_X1 _11356_ ( .A1(_03439_ ), .A2(\ID_EX_csr [2] ), .ZN(_03440_ ) );
AND2_X1 _11357_ ( .A1(_03438_ ), .A2(_03440_ ), .ZN(_03441_ ) );
INV_X1 _11358_ ( .A(_03441_ ), .ZN(_03442_ ) );
BUF_X2 _11359_ ( .A(_03442_ ), .Z(_03443_ ) );
NOR2_X1 _11360_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_03444_ ) );
NAND3_X1 _11361_ ( .A1(_03444_ ), .A2(_03387_ ), .A3(\ID_EX_csr [6] ), .ZN(_03445_ ) );
NAND3_X1 _11362_ ( .A1(_03413_ ), .A2(\ID_EX_csr [9] ), .A3(\ID_EX_csr [8] ), .ZN(_03446_ ) );
NOR3_X1 _11363_ ( .A1(_03445_ ), .A2(\ID_EX_csr [10] ), .A3(_03446_ ), .ZN(_03447_ ) );
BUF_X4 _11364_ ( .A(_03447_ ), .Z(_03448_ ) );
BUF_X4 _11365_ ( .A(_03448_ ), .Z(_03449_ ) );
NAND3_X1 _11366_ ( .A1(_03403_ ), .A2(_03406_ ), .A3(\ID_EX_csr [1] ), .ZN(_03450_ ) );
NOR2_X1 _11367_ ( .A1(_03450_ ), .A2(\ID_EX_csr [0] ), .ZN(_03451_ ) );
BUF_X4 _11368_ ( .A(_03451_ ), .Z(_03452_ ) );
NAND3_X1 _11369_ ( .A1(_03449_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_03452_ ), .ZN(_03453_ ) );
OAI211_X1 _11370_ ( .A(_03443_ ), .B(_03453_ ), .C1(_03424_ ), .C2(_03432_ ), .ZN(_03454_ ) );
AND2_X1 _11371_ ( .A1(_03437_ ), .A2(_03444_ ), .ZN(_03455_ ) );
BUF_X4 _11372_ ( .A(_03455_ ), .Z(_03456_ ) );
AND4_X2 _11373_ ( .A1(_03355_ ), .A2(_03456_ ), .A3(\ID_EX_csr [0] ), .A4(_03403_ ), .ZN(_03457_ ) );
NOR2_X2 _11374_ ( .A1(_03446_ ), .A2(\ID_EX_csr [10] ), .ZN(_03458_ ) );
BUF_X4 _11375_ ( .A(_03458_ ), .Z(_03459_ ) );
BUF_X4 _11376_ ( .A(_03459_ ), .Z(_03460_ ) );
NAND4_X1 _11377_ ( .A1(_03457_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [21] ), .A4(_03460_ ), .ZN(_03461_ ) );
BUF_X4 _11378_ ( .A(_03440_ ), .Z(_03462_ ) );
BUF_X2 _11379_ ( .A(_03462_ ), .Z(_03463_ ) );
NAND3_X1 _11380_ ( .A1(_03449_ ), .A2(\mepc [21] ), .A3(_03463_ ), .ZN(_03464_ ) );
NOR2_X1 _11381_ ( .A1(\ID_EX_csr [1] ), .A2(\ID_EX_csr [0] ), .ZN(_03465_ ) );
AND3_X1 _11382_ ( .A1(_03465_ ), .A2(_03403_ ), .A3(_03406_ ), .ZN(_03466_ ) );
AND2_X2 _11383_ ( .A1(_03466_ ), .A2(_03456_ ), .ZN(_03467_ ) );
NAND3_X1 _11384_ ( .A1(_03467_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_03460_ ), .ZN(_03468_ ) );
NAND3_X1 _11385_ ( .A1(_03461_ ), .A2(_03464_ ), .A3(_03468_ ), .ZN(_03469_ ) );
OAI21_X1 _11386_ ( .A(_03434_ ), .B1(_03454_ ), .B2(_03469_ ), .ZN(_03470_ ) );
AOI22_X1 _11387_ ( .A1(_03470_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_02092_ ), .ZN(_03471_ ) );
NAND2_X1 _11388_ ( .A1(_02091_ ), .A2(_02111_ ), .ZN(_03472_ ) );
OAI21_X1 _11389_ ( .A(_03471_ ), .B1(_03472_ ), .B2(fanout_net_6 ), .ZN(_03473_ ) );
NOR2_X2 _11390_ ( .A1(_02380_ ), .A2(fanout_net_7 ), .ZN(_03474_ ) );
OAI211_X1 _11391_ ( .A(_03434_ ), .B(_03474_ ), .C1(_03454_ ), .C2(_03469_ ), .ZN(_03475_ ) );
NAND2_X1 _11392_ ( .A1(_03473_ ), .A2(_03475_ ), .ZN(_03476_ ) );
MUX2_X1 _11393_ ( .A(\myreg.Reg[14][21] ), .B(\myreg.Reg[15][21] ), .S(fanout_net_23 ), .Z(_03477_ ) );
MUX2_X1 _11394_ ( .A(\myreg.Reg[12][21] ), .B(\myreg.Reg[13][21] ), .S(fanout_net_23 ), .Z(_03478_ ) );
INV_X1 _11395_ ( .A(fanout_net_31 ), .ZN(_03479_ ) );
BUF_X4 _11396_ ( .A(_03479_ ), .Z(_03480_ ) );
BUF_X4 _11397_ ( .A(_03480_ ), .Z(_03481_ ) );
BUF_X4 _11398_ ( .A(_03481_ ), .Z(_03482_ ) );
MUX2_X1 _11399_ ( .A(_03477_ ), .B(_03478_ ), .S(_03482_ ), .Z(_03483_ ) );
MUX2_X1 _11400_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_23 ), .Z(_03484_ ) );
MUX2_X1 _11401_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_23 ), .Z(_03485_ ) );
MUX2_X1 _11402_ ( .A(_03484_ ), .B(_03485_ ), .S(_03482_ ), .Z(_03486_ ) );
INV_X1 _11403_ ( .A(fanout_net_33 ), .ZN(_03487_ ) );
BUF_X4 _11404_ ( .A(_03487_ ), .Z(_03488_ ) );
BUF_X4 _11405_ ( .A(_03488_ ), .Z(_03489_ ) );
BUF_X4 _11406_ ( .A(_03489_ ), .Z(_03490_ ) );
MUX2_X1 _11407_ ( .A(_03483_ ), .B(_03486_ ), .S(_03490_ ), .Z(_03491_ ) );
INV_X1 _11408_ ( .A(fanout_net_34 ), .ZN(_03492_ ) );
BUF_X4 _11409_ ( .A(_03492_ ), .Z(_03493_ ) );
BUF_X4 _11410_ ( .A(_03493_ ), .Z(_03494_ ) );
OR2_X1 _11411_ ( .A1(_03491_ ), .A2(_03494_ ), .ZN(_03495_ ) );
CLKBUF_X2 _11412_ ( .A(_01377_ ), .Z(_03496_ ) );
BUF_X2 _11413_ ( .A(_03496_ ), .Z(_03497_ ) );
BUF_X2 _11414_ ( .A(_03497_ ), .Z(_03498_ ) );
AOI22_X4 _11415_ ( .A1(_01380_ ), .A2(\ID_EX_rs2 [4] ), .B1(_02629_ ), .B2(\EX_LS_dest_reg [3] ), .ZN(_03499_ ) );
INV_X1 _11416_ ( .A(\EX_LS_dest_reg [2] ), .ZN(_03500_ ) );
NAND2_X1 _11417_ ( .A1(_03500_ ), .A2(\ID_EX_rs2 [2] ), .ZN(_03501_ ) );
OAI211_X2 _11418_ ( .A(_03499_ ), .B(_03501_ ), .C1(_01380_ ), .C2(\ID_EX_rs2 [4] ), .ZN(_03502_ ) );
XOR2_X1 _11419_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .Z(_03503_ ) );
OAI21_X1 _11420_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_03500_ ), .B2(\ID_EX_rs2 [2] ), .ZN(_03504_ ) );
OR3_X4 _11421_ ( .A1(_03502_ ), .A2(_03503_ ), .A3(_03504_ ), .ZN(_03505_ ) );
AND2_X1 _11422_ ( .A1(_01382_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_03506_ ) );
NAND2_X1 _11423_ ( .A1(_01394_ ), .A2(\ID_EX_rs2 [3] ), .ZN(_03507_ ) );
OAI21_X1 _11424_ ( .A(_03507_ ), .B1(_01382_ ), .B2(\ID_EX_rs2 [1] ), .ZN(_03508_ ) );
OR4_X4 _11425_ ( .A1(_01381_ ), .A2(_03505_ ), .A3(_03506_ ), .A4(_03508_ ), .ZN(_03509_ ) );
BUF_X8 _11426_ ( .A(_03509_ ), .Z(_03510_ ) );
BUF_X8 _11427_ ( .A(_03510_ ), .Z(_03511_ ) );
BUF_X8 _11428_ ( .A(_03511_ ), .Z(_03512_ ) );
MUX2_X1 _11429_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_23 ), .Z(_03513_ ) );
MUX2_X1 _11430_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_23 ), .Z(_03514_ ) );
MUX2_X1 _11431_ ( .A(_03513_ ), .B(_03514_ ), .S(_03482_ ), .Z(_03515_ ) );
MUX2_X1 _11432_ ( .A(\myreg.Reg[2][21] ), .B(\myreg.Reg[3][21] ), .S(fanout_net_23 ), .Z(_03516_ ) );
MUX2_X1 _11433_ ( .A(\myreg.Reg[0][21] ), .B(\myreg.Reg[1][21] ), .S(fanout_net_23 ), .Z(_03517_ ) );
MUX2_X1 _11434_ ( .A(_03516_ ), .B(_03517_ ), .S(_03482_ ), .Z(_03518_ ) );
BUF_X4 _11435_ ( .A(_03490_ ), .Z(_03519_ ) );
MUX2_X1 _11436_ ( .A(_03515_ ), .B(_03518_ ), .S(_03519_ ), .Z(_03520_ ) );
OAI221_X1 _11437_ ( .A(_03495_ ), .B1(_03498_ ), .B2(_03512_ ), .C1(_03520_ ), .C2(fanout_net_34 ), .ZN(_03521_ ) );
INV_X1 _11438_ ( .A(\EX_LS_result_reg [21] ), .ZN(_03522_ ) );
OR3_X1 _11439_ ( .A1(_03512_ ), .A2(_03498_ ), .A3(_03522_ ), .ZN(_03523_ ) );
NAND2_X1 _11440_ ( .A1(_03521_ ), .A2(_03523_ ), .ZN(_03524_ ) );
MUX2_X1 _11441_ ( .A(\ID_EX_pc [21] ), .B(_03524_ ), .S(_03370_ ), .Z(_03525_ ) );
MUX2_X1 _11442_ ( .A(_03476_ ), .B(_03525_ ), .S(_03390_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
AND3_X1 _11443_ ( .A1(_02068_ ), .A2(_01350_ ), .A3(_02087_ ), .ZN(_03526_ ) );
AND2_X1 _11444_ ( .A1(_03438_ ), .A2(_03451_ ), .ZN(_03527_ ) );
NOR2_X1 _11445_ ( .A1(_03441_ ), .A2(_03527_ ), .ZN(_03528_ ) );
NOR3_X1 _11446_ ( .A1(_03445_ ), .A2(\ID_EX_csr [0] ), .A3(_03450_ ), .ZN(_03529_ ) );
BUF_X4 _11447_ ( .A(_03458_ ), .Z(_03530_ ) );
NAND3_X1 _11448_ ( .A1(_03529_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_03530_ ), .ZN(_03531_ ) );
NAND3_X1 _11449_ ( .A1(_03447_ ), .A2(\mepc [20] ), .A3(_03440_ ), .ZN(_03532_ ) );
NOR2_X1 _11450_ ( .A1(_03439_ ), .A2(_03406_ ), .ZN(_03533_ ) );
NAND4_X1 _11451_ ( .A1(_03533_ ), .A2(_03458_ ), .A3(\mtvec [20] ), .A4(_03456_ ), .ZN(_03534_ ) );
NAND4_X1 _11452_ ( .A1(_03466_ ), .A2(_03458_ ), .A3(\mycsreg.CSReg[0][20] ), .A4(_03456_ ), .ZN(_03535_ ) );
AND3_X1 _11453_ ( .A1(_03532_ ), .A2(_03534_ ), .A3(_03535_ ), .ZN(_03536_ ) );
NAND3_X1 _11454_ ( .A1(_03528_ ), .A2(_03531_ ), .A3(_03536_ ), .ZN(_03537_ ) );
INV_X2 _11455_ ( .A(_03095_ ), .ZN(_03538_ ) );
AND4_X1 _11456_ ( .A1(_03429_ ), .A2(_03419_ ), .A3(_03430_ ), .A4(_03421_ ), .ZN(_03539_ ) );
AND4_X2 _11457_ ( .A1(_03418_ ), .A2(_03539_ ), .A3(_03420_ ), .A4(_03427_ ), .ZN(_03540_ ) );
AND4_X2 _11458_ ( .A1(_03428_ ), .A2(_03414_ ), .A3(_03416_ ), .A4(_03415_ ), .ZN(_03541_ ) );
NAND2_X1 _11459_ ( .A1(_03540_ ), .A2(_03541_ ), .ZN(_03542_ ) );
OAI21_X1 _11460_ ( .A(_03537_ ), .B1(_03538_ ), .B2(_03542_ ), .ZN(_03543_ ) );
NAND4_X1 _11461_ ( .A1(_03540_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_03095_ ), .A4(_03541_ ), .ZN(_03544_ ) );
AND2_X1 _11462_ ( .A1(_03543_ ), .A2(_03544_ ), .ZN(_03545_ ) );
AOI221_X4 _11463_ ( .A(_03526_ ), .B1(fanout_net_6 ), .B2(_02089_ ), .C1(fanout_net_7 ), .C2(_03545_ ), .ZN(_03546_ ) );
INV_X1 _11464_ ( .A(_03474_ ), .ZN(_03547_ ) );
BUF_X2 _11465_ ( .A(_03547_ ), .Z(_03548_ ) );
AOI21_X1 _11466_ ( .A(_03548_ ), .B1(_03543_ ), .B2(_03544_ ), .ZN(_03549_ ) );
OAI21_X1 _11467_ ( .A(_03379_ ), .B1(_03546_ ), .B2(_03549_ ), .ZN(_03550_ ) );
BUF_X4 _11468_ ( .A(_01365_ ), .Z(_03551_ ) );
BUF_X4 _11469_ ( .A(_03551_ ), .Z(_03552_ ) );
BUF_X4 _11470_ ( .A(_03512_ ), .Z(_03553_ ) );
CLKBUF_X2 _11471_ ( .A(_03498_ ), .Z(_03554_ ) );
OR3_X1 _11472_ ( .A1(_03553_ ), .A2(_03554_ ), .A3(\EX_LS_result_reg [20] ), .ZN(_03555_ ) );
BUF_X4 _11473_ ( .A(_03494_ ), .Z(_03556_ ) );
INV_X1 _11474_ ( .A(fanout_net_23 ), .ZN(_03557_ ) );
BUF_X2 _11475_ ( .A(_03557_ ), .Z(_03558_ ) );
BUF_X4 _11476_ ( .A(_03558_ ), .Z(_03559_ ) );
BUF_X4 _11477_ ( .A(_03559_ ), .Z(_03560_ ) );
BUF_X4 _11478_ ( .A(_03560_ ), .Z(_03561_ ) );
CLKBUF_X2 _11479_ ( .A(_03561_ ), .Z(_03562_ ) );
OR2_X1 _11480_ ( .A1(_03562_ ), .A2(\myreg.Reg[3][20] ), .ZN(_03563_ ) );
OAI211_X1 _11481_ ( .A(_03563_ ), .B(fanout_net_31 ), .C1(fanout_net_23 ), .C2(\myreg.Reg[2][20] ), .ZN(_03564_ ) );
BUF_X4 _11482_ ( .A(_03490_ ), .Z(_03565_ ) );
OR2_X1 _11483_ ( .A1(fanout_net_23 ), .A2(\myreg.Reg[0][20] ), .ZN(_03566_ ) );
BUF_X4 _11484_ ( .A(_03482_ ), .Z(_03567_ ) );
BUF_X4 _11485_ ( .A(_03562_ ), .Z(_03568_ ) );
OAI211_X1 _11486_ ( .A(_03566_ ), .B(_03567_ ), .C1(_03568_ ), .C2(\myreg.Reg[1][20] ), .ZN(_03569_ ) );
NAND3_X1 _11487_ ( .A1(_03564_ ), .A2(_03565_ ), .A3(_03569_ ), .ZN(_03570_ ) );
MUX2_X1 _11488_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_23 ), .Z(_03571_ ) );
MUX2_X1 _11489_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_23 ), .Z(_03572_ ) );
BUF_X4 _11490_ ( .A(_03482_ ), .Z(_03573_ ) );
MUX2_X1 _11491_ ( .A(_03571_ ), .B(_03572_ ), .S(_03573_ ), .Z(_03574_ ) );
BUF_X4 _11492_ ( .A(_03519_ ), .Z(_03575_ ) );
OAI211_X1 _11493_ ( .A(_03556_ ), .B(_03570_ ), .C1(_03574_ ), .C2(_03575_ ), .ZN(_03576_ ) );
OR2_X1 _11494_ ( .A1(_03562_ ), .A2(\myreg.Reg[15][20] ), .ZN(_03577_ ) );
OAI211_X1 _11495_ ( .A(_03577_ ), .B(fanout_net_31 ), .C1(fanout_net_23 ), .C2(\myreg.Reg[14][20] ), .ZN(_03578_ ) );
OR2_X1 _11496_ ( .A1(_03562_ ), .A2(\myreg.Reg[13][20] ), .ZN(_03579_ ) );
OAI211_X1 _11497_ ( .A(_03579_ ), .B(_03567_ ), .C1(fanout_net_23 ), .C2(\myreg.Reg[12][20] ), .ZN(_03580_ ) );
NAND3_X1 _11498_ ( .A1(_03578_ ), .A2(_03580_ ), .A3(fanout_net_33 ), .ZN(_03581_ ) );
MUX2_X1 _11499_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_23 ), .Z(_03582_ ) );
MUX2_X1 _11500_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_23 ), .Z(_03583_ ) );
MUX2_X1 _11501_ ( .A(_03582_ ), .B(_03583_ ), .S(fanout_net_31 ), .Z(_03584_ ) );
OAI211_X1 _11502_ ( .A(fanout_net_34 ), .B(_03581_ ), .C1(_03584_ ), .C2(fanout_net_33 ), .ZN(_03585_ ) );
BUF_X4 _11503_ ( .A(_03512_ ), .Z(_03586_ ) );
BUF_X4 _11504_ ( .A(_03498_ ), .Z(_03587_ ) );
OAI211_X1 _11505_ ( .A(_03576_ ), .B(_03585_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_03588_ ) );
NAND2_X1 _11506_ ( .A1(_03555_ ), .A2(_03588_ ), .ZN(_03589_ ) );
BUF_X4 _11507_ ( .A(_03361_ ), .Z(_03590_ ) );
MUX2_X1 _11508_ ( .A(_02327_ ), .B(_03589_ ), .S(_03590_ ), .Z(_03591_ ) );
OAI21_X1 _11509_ ( .A(_03550_ ), .B1(_03552_ ), .B2(_03591_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
BUF_X4 _11510_ ( .A(_03448_ ), .Z(_03592_ ) );
NAND3_X1 _11511_ ( .A1(_03592_ ), .A2(\mepc [19] ), .A3(_03462_ ), .ZN(_03593_ ) );
BUF_X4 _11512_ ( .A(_03466_ ), .Z(_03594_ ) );
BUF_X4 _11513_ ( .A(_03456_ ), .Z(_03595_ ) );
NAND4_X1 _11514_ ( .A1(_03594_ ), .A2(_03530_ ), .A3(\mycsreg.CSReg[0][19] ), .A4(_03595_ ), .ZN(_03596_ ) );
AND2_X1 _11515_ ( .A1(_03593_ ), .A2(_03596_ ), .ZN(_03597_ ) );
AND4_X1 _11516_ ( .A1(\mtvec [19] ), .A2(_03533_ ), .A3(_03459_ ), .A4(_03456_ ), .ZN(_03598_ ) );
BUF_X4 _11517_ ( .A(_03451_ ), .Z(_03599_ ) );
AOI21_X1 _11518_ ( .A(_03598_ ), .B1(_03438_ ), .B2(_03599_ ), .ZN(_03600_ ) );
AND3_X1 _11519_ ( .A1(_03448_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_03451_ ), .ZN(_03601_ ) );
INV_X1 _11520_ ( .A(_03601_ ), .ZN(_03602_ ) );
NAND3_X1 _11521_ ( .A1(_03597_ ), .A2(_03600_ ), .A3(_03602_ ), .ZN(_03603_ ) );
OAI21_X1 _11522_ ( .A(_03603_ ), .B1(_03542_ ), .B2(_03538_ ), .ZN(_03604_ ) );
BUF_X4 _11523_ ( .A(_03540_ ), .Z(_03605_ ) );
BUF_X4 _11524_ ( .A(_03541_ ), .Z(_03606_ ) );
NAND4_X1 _11525_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_03096_ ), .A4(_03606_ ), .ZN(_03607_ ) );
AOI21_X1 _11526_ ( .A(_03547_ ), .B1(_03604_ ), .B2(_03607_ ), .ZN(_03608_ ) );
NAND2_X1 _11527_ ( .A1(_03604_ ), .A2(_03607_ ), .ZN(_03609_ ) );
INV_X1 _11528_ ( .A(_03609_ ), .ZN(_03610_ ) );
AOI22_X1 _11529_ ( .A1(_03610_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01975_ ), .ZN(_03611_ ) );
NAND3_X1 _11530_ ( .A1(_01974_ ), .A2(_01994_ ), .A3(_01351_ ), .ZN(_03612_ ) );
AOI211_X1 _11531_ ( .A(_03357_ ), .B(_03608_ ), .C1(_03611_ ), .C2(_03612_ ), .ZN(_03613_ ) );
OR3_X1 _11532_ ( .A1(_03512_ ), .A2(_03498_ ), .A3(\EX_LS_result_reg [19] ), .ZN(_03614_ ) );
OR2_X1 _11533_ ( .A1(fanout_net_23 ), .A2(\myreg.Reg[8][19] ), .ZN(_03615_ ) );
BUF_X4 _11534_ ( .A(_03482_ ), .Z(_03616_ ) );
BUF_X4 _11535_ ( .A(_03561_ ), .Z(_03617_ ) );
OAI211_X1 _11536_ ( .A(_03615_ ), .B(_03616_ ), .C1(_03617_ ), .C2(\myreg.Reg[9][19] ), .ZN(_03618_ ) );
OR2_X1 _11537_ ( .A1(fanout_net_23 ), .A2(\myreg.Reg[10][19] ), .ZN(_03619_ ) );
OAI211_X1 _11538_ ( .A(_03619_ ), .B(fanout_net_31 ), .C1(_03617_ ), .C2(\myreg.Reg[11][19] ), .ZN(_03620_ ) );
NAND3_X1 _11539_ ( .A1(_03618_ ), .A2(_03620_ ), .A3(_03519_ ), .ZN(_03621_ ) );
MUX2_X1 _11540_ ( .A(\myreg.Reg[14][19] ), .B(\myreg.Reg[15][19] ), .S(fanout_net_23 ), .Z(_03622_ ) );
MUX2_X1 _11541_ ( .A(\myreg.Reg[12][19] ), .B(\myreg.Reg[13][19] ), .S(fanout_net_23 ), .Z(_03623_ ) );
BUF_X4 _11542_ ( .A(_03482_ ), .Z(_03624_ ) );
MUX2_X1 _11543_ ( .A(_03622_ ), .B(_03623_ ), .S(_03624_ ), .Z(_03625_ ) );
OAI211_X1 _11544_ ( .A(fanout_net_34 ), .B(_03621_ ), .C1(_03625_ ), .C2(_03565_ ), .ZN(_03626_ ) );
BUF_X2 _11545_ ( .A(_03561_ ), .Z(_03627_ ) );
NOR2_X1 _11546_ ( .A1(_03627_ ), .A2(\myreg.Reg[3][19] ), .ZN(_03628_ ) );
OAI21_X1 _11547_ ( .A(fanout_net_31 ), .B1(fanout_net_23 ), .B2(\myreg.Reg[2][19] ), .ZN(_03629_ ) );
NOR2_X1 _11548_ ( .A1(fanout_net_23 ), .A2(\myreg.Reg[0][19] ), .ZN(_03630_ ) );
OAI21_X1 _11549_ ( .A(_03624_ ), .B1(_03627_ ), .B2(\myreg.Reg[1][19] ), .ZN(_03631_ ) );
OAI221_X1 _11550_ ( .A(_03519_ ), .B1(_03628_ ), .B2(_03629_ ), .C1(_03630_ ), .C2(_03631_ ), .ZN(_03632_ ) );
MUX2_X1 _11551_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_23 ), .Z(_03633_ ) );
MUX2_X1 _11552_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_23 ), .Z(_03634_ ) );
MUX2_X1 _11553_ ( .A(_03633_ ), .B(_03634_ ), .S(_03624_ ), .Z(_03635_ ) );
OAI211_X1 _11554_ ( .A(_03494_ ), .B(_03632_ ), .C1(_03635_ ), .C2(_03565_ ), .ZN(_03636_ ) );
OAI211_X1 _11555_ ( .A(_03626_ ), .B(_03636_ ), .C1(_03553_ ), .C2(_03554_ ), .ZN(_03637_ ) );
NAND2_X1 _11556_ ( .A1(_03614_ ), .A2(_03637_ ), .ZN(_03638_ ) );
MUX2_X1 _11557_ ( .A(_02328_ ), .B(_03638_ ), .S(_03590_ ), .Z(_03639_ ) );
AOI21_X1 _11558_ ( .A(_03613_ ), .B1(_03358_ ), .B2(_03639_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
NOR2_X1 _11559_ ( .A1(_01350_ ), .A2(\ID_EX_imm [18] ), .ZN(_03640_ ) );
AND4_X1 _11560_ ( .A1(_03420_ ), .A2(_03421_ ), .A3(_03416_ ), .A4(_03426_ ), .ZN(_03641_ ) );
AND4_X1 _11561_ ( .A1(_03095_ ), .A2(_03641_ ), .A3(_03419_ ), .A4(_03430_ ), .ZN(_03642_ ) );
AND4_X1 _11562_ ( .A1(_03414_ ), .A2(_03418_ ), .A3(_03429_ ), .A4(_03415_ ), .ZN(_03643_ ) );
AND3_X1 _11563_ ( .A1(_03643_ ), .A2(_03428_ ), .A3(_03425_ ), .ZN(_03644_ ) );
AND2_X1 _11564_ ( .A1(_03642_ ), .A2(_03644_ ), .ZN(_03645_ ) );
INV_X1 _11565_ ( .A(_03645_ ), .ZN(_03646_ ) );
AND3_X1 _11566_ ( .A1(_03447_ ), .A2(\mepc [18] ), .A3(_03462_ ), .ZN(_03647_ ) );
OR2_X1 _11567_ ( .A1(_03527_ ), .A2(_03647_ ), .ZN(_03648_ ) );
NAND3_X1 _11568_ ( .A1(_03448_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_03451_ ), .ZN(_03649_ ) );
BUF_X4 _11569_ ( .A(_03456_ ), .Z(_03650_ ) );
NAND4_X1 _11570_ ( .A1(_03594_ ), .A2(_03459_ ), .A3(\mycsreg.CSReg[0][18] ), .A4(_03650_ ), .ZN(_03651_ ) );
BUF_X4 _11571_ ( .A(_03533_ ), .Z(_03652_ ) );
NAND4_X1 _11572_ ( .A1(_03652_ ), .A2(_03459_ ), .A3(\mtvec [18] ), .A4(_03650_ ), .ZN(_03653_ ) );
NAND3_X1 _11573_ ( .A1(_03649_ ), .A2(_03651_ ), .A3(_03653_ ), .ZN(_03654_ ) );
OAI21_X1 _11574_ ( .A(_03646_ ), .B1(_03648_ ), .B2(_03654_ ), .ZN(_03655_ ) );
NAND4_X1 _11575_ ( .A1(_03540_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_03095_ ), .A4(_03541_ ), .ZN(_03656_ ) );
AND2_X1 _11576_ ( .A1(_03655_ ), .A2(_03656_ ), .ZN(_03657_ ) );
AOI221_X4 _11577_ ( .A(_03640_ ), .B1(_02123_ ), .B2(_01350_ ), .C1(_03657_ ), .C2(fanout_net_7 ), .ZN(_03658_ ) );
AOI21_X1 _11578_ ( .A(_03548_ ), .B1(_03655_ ), .B2(_03656_ ), .ZN(_03659_ ) );
OAI21_X1 _11579_ ( .A(_03379_ ), .B1(_03658_ ), .B2(_03659_ ), .ZN(_03660_ ) );
OR3_X1 _11580_ ( .A1(_03553_ ), .A2(_03554_ ), .A3(\EX_LS_result_reg [18] ), .ZN(_03661_ ) );
OR2_X1 _11581_ ( .A1(_03627_ ), .A2(\myreg.Reg[1][18] ), .ZN(_03662_ ) );
BUF_X4 _11582_ ( .A(_03482_ ), .Z(_03663_ ) );
OAI211_X1 _11583_ ( .A(_03662_ ), .B(_03663_ ), .C1(fanout_net_23 ), .C2(\myreg.Reg[0][18] ), .ZN(_03664_ ) );
BUF_X4 _11584_ ( .A(_03490_ ), .Z(_03665_ ) );
OR2_X1 _11585_ ( .A1(fanout_net_23 ), .A2(\myreg.Reg[2][18] ), .ZN(_03666_ ) );
OAI211_X1 _11586_ ( .A(_03666_ ), .B(fanout_net_31 ), .C1(_03568_ ), .C2(\myreg.Reg[3][18] ), .ZN(_03667_ ) );
NAND3_X1 _11587_ ( .A1(_03664_ ), .A2(_03665_ ), .A3(_03667_ ), .ZN(_03668_ ) );
MUX2_X1 _11588_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_23 ), .Z(_03669_ ) );
MUX2_X1 _11589_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_23 ), .Z(_03670_ ) );
MUX2_X1 _11590_ ( .A(_03669_ ), .B(_03670_ ), .S(_03567_ ), .Z(_03671_ ) );
OAI211_X1 _11591_ ( .A(_03556_ ), .B(_03668_ ), .C1(_03671_ ), .C2(_03575_ ), .ZN(_03672_ ) );
OR2_X1 _11592_ ( .A1(_03562_ ), .A2(\myreg.Reg[15][18] ), .ZN(_03673_ ) );
OAI211_X1 _11593_ ( .A(_03673_ ), .B(fanout_net_31 ), .C1(fanout_net_23 ), .C2(\myreg.Reg[14][18] ), .ZN(_03674_ ) );
OR2_X1 _11594_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[12][18] ), .ZN(_03675_ ) );
OAI211_X1 _11595_ ( .A(_03675_ ), .B(_03663_ ), .C1(_03568_ ), .C2(\myreg.Reg[13][18] ), .ZN(_03676_ ) );
NAND3_X1 _11596_ ( .A1(_03674_ ), .A2(fanout_net_33 ), .A3(_03676_ ), .ZN(_03677_ ) );
MUX2_X1 _11597_ ( .A(\myreg.Reg[8][18] ), .B(\myreg.Reg[9][18] ), .S(fanout_net_24 ), .Z(_03678_ ) );
MUX2_X1 _11598_ ( .A(\myreg.Reg[10][18] ), .B(\myreg.Reg[11][18] ), .S(fanout_net_24 ), .Z(_03679_ ) );
MUX2_X1 _11599_ ( .A(_03678_ ), .B(_03679_ ), .S(fanout_net_31 ), .Z(_03680_ ) );
OAI211_X1 _11600_ ( .A(fanout_net_34 ), .B(_03677_ ), .C1(_03680_ ), .C2(fanout_net_33 ), .ZN(_03681_ ) );
OAI211_X1 _11601_ ( .A(_03672_ ), .B(_03681_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_03682_ ) );
NAND2_X1 _11602_ ( .A1(_03661_ ), .A2(_03682_ ), .ZN(_03683_ ) );
MUX2_X1 _11603_ ( .A(_02329_ ), .B(_03683_ ), .S(_03590_ ), .Z(_03684_ ) );
OAI21_X1 _11604_ ( .A(_03660_ ), .B1(_03552_ ), .B2(_03684_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
BUF_X2 _11605_ ( .A(_03530_ ), .Z(_03685_ ) );
AND3_X1 _11606_ ( .A1(_03467_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_03685_ ), .ZN(_03686_ ) );
NAND3_X1 _11607_ ( .A1(_03449_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_03452_ ), .ZN(_03687_ ) );
NOR3_X1 _11608_ ( .A1(_03445_ ), .A2(\ID_EX_csr [2] ), .A3(_03439_ ), .ZN(_03688_ ) );
NAND3_X1 _11609_ ( .A1(_03688_ ), .A2(\mepc [17] ), .A3(_03460_ ), .ZN(_03689_ ) );
BUF_X4 _11610_ ( .A(_03652_ ), .Z(_03690_ ) );
BUF_X4 _11611_ ( .A(_03650_ ), .Z(_03691_ ) );
NAND4_X1 _11612_ ( .A1(_03690_ ), .A2(_03460_ ), .A3(\mtvec [17] ), .A4(_03691_ ), .ZN(_03692_ ) );
NAND4_X1 _11613_ ( .A1(_03528_ ), .A2(_03687_ ), .A3(_03689_ ), .A4(_03692_ ), .ZN(_03693_ ) );
OAI21_X1 _11614_ ( .A(_03646_ ), .B1(_03686_ ), .B2(_03693_ ), .ZN(_03694_ ) );
NAND4_X1 _11615_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_03096_ ), .A4(_03606_ ), .ZN(_03695_ ) );
AND2_X1 _11616_ ( .A1(_03694_ ), .A2(_03695_ ), .ZN(_03696_ ) );
AOI22_X1 _11617_ ( .A1(_03696_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01946_ ), .ZN(_03697_ ) );
BUF_X4 _11618_ ( .A(_01365_ ), .Z(_03698_ ) );
OAI211_X1 _11619_ ( .A(_03697_ ), .B(_03698_ ), .C1(fanout_net_6 ), .C2(_01945_ ), .ZN(_03699_ ) );
BUF_X2 _11620_ ( .A(_03356_ ), .Z(_03700_ ) );
AOI21_X1 _11621_ ( .A(_03700_ ), .B1(_03694_ ), .B2(_03695_ ), .ZN(_03701_ ) );
BUF_X4 _11622_ ( .A(_03474_ ), .Z(_03702_ ) );
NAND2_X1 _11623_ ( .A1(_03701_ ), .A2(_03702_ ), .ZN(_03703_ ) );
OR3_X4 _11624_ ( .A1(_03553_ ), .A2(_03554_ ), .A3(\EX_LS_result_reg [17] ), .ZN(_03704_ ) );
OR2_X1 _11625_ ( .A1(_03562_ ), .A2(\myreg.Reg[1][17] ), .ZN(_03705_ ) );
OAI211_X1 _11626_ ( .A(_03705_ ), .B(_03663_ ), .C1(fanout_net_24 ), .C2(\myreg.Reg[0][17] ), .ZN(_03706_ ) );
OR2_X1 _11627_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[2][17] ), .ZN(_03707_ ) );
OAI211_X1 _11628_ ( .A(_03707_ ), .B(fanout_net_31 ), .C1(_03568_ ), .C2(\myreg.Reg[3][17] ), .ZN(_03708_ ) );
NAND3_X1 _11629_ ( .A1(_03706_ ), .A2(_03565_ ), .A3(_03708_ ), .ZN(_03709_ ) );
MUX2_X1 _11630_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_24 ), .Z(_03710_ ) );
MUX2_X1 _11631_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_24 ), .Z(_03711_ ) );
MUX2_X1 _11632_ ( .A(_03710_ ), .B(_03711_ ), .S(_03573_ ), .Z(_03712_ ) );
OAI211_X1 _11633_ ( .A(_03556_ ), .B(_03709_ ), .C1(_03712_ ), .C2(_03575_ ), .ZN(_03713_ ) );
OR2_X1 _11634_ ( .A1(_03562_ ), .A2(\myreg.Reg[13][17] ), .ZN(_03714_ ) );
OAI211_X1 _11635_ ( .A(_03714_ ), .B(_03663_ ), .C1(fanout_net_24 ), .C2(\myreg.Reg[12][17] ), .ZN(_03715_ ) );
OR2_X1 _11636_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[14][17] ), .ZN(_03716_ ) );
OAI211_X1 _11637_ ( .A(_03716_ ), .B(fanout_net_31 ), .C1(_03568_ ), .C2(\myreg.Reg[15][17] ), .ZN(_03717_ ) );
NAND3_X1 _11638_ ( .A1(_03715_ ), .A2(fanout_net_33 ), .A3(_03717_ ), .ZN(_03718_ ) );
MUX2_X1 _11639_ ( .A(\myreg.Reg[8][17] ), .B(\myreg.Reg[9][17] ), .S(fanout_net_24 ), .Z(_03719_ ) );
MUX2_X1 _11640_ ( .A(\myreg.Reg[10][17] ), .B(\myreg.Reg[11][17] ), .S(fanout_net_24 ), .Z(_03720_ ) );
MUX2_X1 _11641_ ( .A(_03719_ ), .B(_03720_ ), .S(fanout_net_31 ), .Z(_03721_ ) );
OAI211_X1 _11642_ ( .A(fanout_net_34 ), .B(_03718_ ), .C1(_03721_ ), .C2(fanout_net_33 ), .ZN(_03722_ ) );
OAI211_X1 _11643_ ( .A(_03713_ ), .B(_03722_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_03723_ ) );
NAND2_X1 _11644_ ( .A1(_03704_ ), .A2(_03723_ ), .ZN(_03724_ ) );
MUX2_X1 _11645_ ( .A(_02330_ ), .B(_03724_ ), .S(_03370_ ), .Z(_03725_ ) );
OAI211_X1 _11646_ ( .A(_03699_ ), .B(_03703_ ), .C1(_03552_ ), .C2(_03725_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _11647_ ( .A1(_03529_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_03685_ ), .ZN(_03726_ ) );
NAND3_X1 _11648_ ( .A1(_03448_ ), .A2(\mepc [16] ), .A3(_03462_ ), .ZN(_03727_ ) );
NAND4_X1 _11649_ ( .A1(_03652_ ), .A2(_03530_ ), .A3(\mtvec [16] ), .A4(_03650_ ), .ZN(_03728_ ) );
NAND4_X1 _11650_ ( .A1(_03594_ ), .A2(_03459_ ), .A3(\mycsreg.CSReg[0][16] ), .A4(_03650_ ), .ZN(_03729_ ) );
AND3_X1 _11651_ ( .A1(_03727_ ), .A2(_03728_ ), .A3(_03729_ ), .ZN(_03730_ ) );
NAND3_X1 _11652_ ( .A1(_03528_ ), .A2(_03726_ ), .A3(_03730_ ), .ZN(_03731_ ) );
OAI21_X1 _11653_ ( .A(_03731_ ), .B1(_03538_ ), .B2(_03542_ ), .ZN(_03732_ ) );
NAND4_X1 _11654_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [16] ), .A3(_03096_ ), .A4(_03606_ ), .ZN(_03733_ ) );
AOI21_X1 _11655_ ( .A(_03357_ ), .B1(_03732_ ), .B2(_03733_ ), .ZN(_03734_ ) );
NAND2_X1 _11656_ ( .A1(_03734_ ), .A2(_03702_ ), .ZN(_03735_ ) );
AND2_X1 _11657_ ( .A1(_03732_ ), .A2(_03733_ ), .ZN(_03736_ ) );
AOI22_X1 _11658_ ( .A1(_03736_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01970_ ), .ZN(_03737_ ) );
OAI211_X1 _11659_ ( .A(_03737_ ), .B(_03551_ ), .C1(fanout_net_6 ), .C2(_01969_ ), .ZN(_03738_ ) );
OR3_X1 _11660_ ( .A1(_03512_ ), .A2(_03498_ ), .A3(\EX_LS_result_reg [16] ), .ZN(_03739_ ) );
OR2_X1 _11661_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[0][16] ), .ZN(_03740_ ) );
BUF_X4 _11662_ ( .A(_03561_ ), .Z(_03741_ ) );
OAI211_X1 _11663_ ( .A(_03740_ ), .B(_03567_ ), .C1(_03741_ ), .C2(\myreg.Reg[1][16] ), .ZN(_03742_ ) );
OR2_X1 _11664_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[2][16] ), .ZN(_03743_ ) );
OAI211_X1 _11665_ ( .A(_03743_ ), .B(fanout_net_31 ), .C1(_03741_ ), .C2(\myreg.Reg[3][16] ), .ZN(_03744_ ) );
NAND3_X1 _11666_ ( .A1(_03742_ ), .A2(_03744_ ), .A3(_03565_ ), .ZN(_03745_ ) );
MUX2_X1 _11667_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_24 ), .Z(_03746_ ) );
MUX2_X1 _11668_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_24 ), .Z(_03747_ ) );
MUX2_X1 _11669_ ( .A(_03746_ ), .B(_03747_ ), .S(_03616_ ), .Z(_03748_ ) );
OAI211_X1 _11670_ ( .A(_03556_ ), .B(_03745_ ), .C1(_03748_ ), .C2(_03665_ ), .ZN(_03749_ ) );
OR2_X1 _11671_ ( .A1(_03561_ ), .A2(\myreg.Reg[15][16] ), .ZN(_03750_ ) );
OAI211_X1 _11672_ ( .A(_03750_ ), .B(fanout_net_31 ), .C1(fanout_net_24 ), .C2(\myreg.Reg[14][16] ), .ZN(_03751_ ) );
OR2_X1 _11673_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[12][16] ), .ZN(_03752_ ) );
OAI211_X1 _11674_ ( .A(_03752_ ), .B(_03616_ ), .C1(_03741_ ), .C2(\myreg.Reg[13][16] ), .ZN(_03753_ ) );
NAND3_X1 _11675_ ( .A1(_03751_ ), .A2(fanout_net_33 ), .A3(_03753_ ), .ZN(_03754_ ) );
MUX2_X1 _11676_ ( .A(\myreg.Reg[8][16] ), .B(\myreg.Reg[9][16] ), .S(fanout_net_24 ), .Z(_03755_ ) );
MUX2_X1 _11677_ ( .A(\myreg.Reg[10][16] ), .B(\myreg.Reg[11][16] ), .S(fanout_net_24 ), .Z(_03756_ ) );
MUX2_X1 _11678_ ( .A(_03755_ ), .B(_03756_ ), .S(fanout_net_31 ), .Z(_03757_ ) );
OAI211_X1 _11679_ ( .A(fanout_net_34 ), .B(_03754_ ), .C1(_03757_ ), .C2(fanout_net_33 ), .ZN(_03758_ ) );
OAI211_X1 _11680_ ( .A(_03749_ ), .B(_03758_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_03759_ ) );
NAND2_X1 _11681_ ( .A1(_03739_ ), .A2(_03759_ ), .ZN(_03760_ ) );
MUX2_X1 _11682_ ( .A(_02331_ ), .B(_03760_ ), .S(_03590_ ), .Z(_03761_ ) );
BUF_X4 _11683_ ( .A(_03378_ ), .Z(_03762_ ) );
OAI211_X1 _11684_ ( .A(_03735_ ), .B(_03738_ ), .C1(_03761_ ), .C2(_03762_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
AND4_X1 _11685_ ( .A1(\mtvec [15] ), .A2(_03652_ ), .A3(_03459_ ), .A4(_03650_ ), .ZN(_03763_ ) );
OR2_X1 _11686_ ( .A1(_03527_ ), .A2(_03763_ ), .ZN(_03764_ ) );
BUF_X4 _11687_ ( .A(_03448_ ), .Z(_03765_ ) );
NAND3_X1 _11688_ ( .A1(_03765_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_03599_ ), .ZN(_03766_ ) );
NAND3_X1 _11689_ ( .A1(_03449_ ), .A2(\mepc [15] ), .A3(_03463_ ), .ZN(_03767_ ) );
BUF_X4 _11690_ ( .A(_03594_ ), .Z(_03768_ ) );
NAND4_X1 _11691_ ( .A1(_03768_ ), .A2(_03460_ ), .A3(\mycsreg.CSReg[0][15] ), .A4(_03691_ ), .ZN(_03769_ ) );
NAND3_X1 _11692_ ( .A1(_03766_ ), .A2(_03767_ ), .A3(_03769_ ), .ZN(_03770_ ) );
OAI21_X1 _11693_ ( .A(_03646_ ), .B1(_03764_ ), .B2(_03770_ ), .ZN(_03771_ ) );
NAND4_X1 _11694_ ( .A1(_03540_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_03096_ ), .A4(_03541_ ), .ZN(_03772_ ) );
AOI21_X1 _11695_ ( .A(_03547_ ), .B1(_03771_ ), .B2(_03772_ ), .ZN(_03773_ ) );
AND2_X1 _11696_ ( .A1(_03771_ ), .A2(_03772_ ), .ZN(_03774_ ) );
AOI22_X1 _11697_ ( .A1(_03774_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01761_ ), .ZN(_03775_ ) );
NAND3_X1 _11698_ ( .A1(_01740_ ), .A2(_01759_ ), .A3(_01350_ ), .ZN(_03776_ ) );
AOI211_X1 _11699_ ( .A(_03357_ ), .B(_03773_ ), .C1(_03775_ ), .C2(_03776_ ), .ZN(_03777_ ) );
OR3_X4 _11700_ ( .A1(_03511_ ), .A2(_03497_ ), .A3(\EX_LS_result_reg [15] ), .ZN(_03778_ ) );
BUF_X2 _11701_ ( .A(_03558_ ), .Z(_03779_ ) );
OR2_X1 _11702_ ( .A1(_03779_ ), .A2(\myreg.Reg[3][15] ), .ZN(_03780_ ) );
OAI211_X1 _11703_ ( .A(_03780_ ), .B(fanout_net_31 ), .C1(fanout_net_24 ), .C2(\myreg.Reg[2][15] ), .ZN(_03781_ ) );
BUF_X4 _11704_ ( .A(_03488_ ), .Z(_03782_ ) );
OR2_X1 _11705_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[0][15] ), .ZN(_03783_ ) );
BUF_X4 _11706_ ( .A(_03480_ ), .Z(_03784_ ) );
BUF_X4 _11707_ ( .A(_03784_ ), .Z(_03785_ ) );
OAI211_X1 _11708_ ( .A(_03783_ ), .B(_03785_ ), .C1(_03560_ ), .C2(\myreg.Reg[1][15] ), .ZN(_03786_ ) );
NAND3_X1 _11709_ ( .A1(_03781_ ), .A2(_03782_ ), .A3(_03786_ ), .ZN(_03787_ ) );
MUX2_X1 _11710_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_24 ), .Z(_03788_ ) );
MUX2_X1 _11711_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_24 ), .Z(_03789_ ) );
MUX2_X1 _11712_ ( .A(_03788_ ), .B(_03789_ ), .S(_03785_ ), .Z(_03790_ ) );
OAI211_X1 _11713_ ( .A(_03494_ ), .B(_03787_ ), .C1(_03790_ ), .C2(_03490_ ), .ZN(_03791_ ) );
OR2_X1 _11714_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[14][15] ), .ZN(_03792_ ) );
OAI211_X1 _11715_ ( .A(_03792_ ), .B(fanout_net_31 ), .C1(_03560_ ), .C2(\myreg.Reg[15][15] ), .ZN(_03793_ ) );
OR2_X1 _11716_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[12][15] ), .ZN(_03794_ ) );
OAI211_X1 _11717_ ( .A(_03794_ ), .B(_03785_ ), .C1(_03560_ ), .C2(\myreg.Reg[13][15] ), .ZN(_03795_ ) );
NAND3_X1 _11718_ ( .A1(_03793_ ), .A2(_03795_ ), .A3(fanout_net_33 ), .ZN(_03796_ ) );
MUX2_X1 _11719_ ( .A(\myreg.Reg[8][15] ), .B(\myreg.Reg[9][15] ), .S(fanout_net_24 ), .Z(_03797_ ) );
MUX2_X1 _11720_ ( .A(\myreg.Reg[10][15] ), .B(\myreg.Reg[11][15] ), .S(fanout_net_24 ), .Z(_03798_ ) );
MUX2_X1 _11721_ ( .A(_03797_ ), .B(_03798_ ), .S(fanout_net_31 ), .Z(_03799_ ) );
OAI211_X1 _11722_ ( .A(fanout_net_34 ), .B(_03796_ ), .C1(_03799_ ), .C2(fanout_net_33 ), .ZN(_03800_ ) );
OAI211_X1 _11723_ ( .A(_03791_ ), .B(_03800_ ), .C1(_03511_ ), .C2(_03497_ ), .ZN(_03801_ ) );
NAND2_X2 _11724_ ( .A1(_03778_ ), .A2(_03801_ ), .ZN(_03802_ ) );
MUX2_X1 _11725_ ( .A(_02332_ ), .B(_03802_ ), .S(_03590_ ), .Z(_03803_ ) );
AOI21_X1 _11726_ ( .A(_03777_ ), .B1(_03358_ ), .B2(_03803_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
NOR2_X1 _11727_ ( .A1(_01350_ ), .A2(\ID_EX_imm [14] ), .ZN(_03804_ ) );
NAND4_X1 _11728_ ( .A1(_03533_ ), .A2(_03459_ ), .A3(\mtvec [14] ), .A4(_03456_ ), .ZN(_03805_ ) );
NAND3_X1 _11729_ ( .A1(_03447_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_03451_ ), .ZN(_03806_ ) );
NAND3_X1 _11730_ ( .A1(_03447_ ), .A2(\mepc [14] ), .A3(_03440_ ), .ZN(_03807_ ) );
NAND4_X1 _11731_ ( .A1(_03466_ ), .A2(_03458_ ), .A3(\mycsreg.CSReg[0][14] ), .A4(_03456_ ), .ZN(_03808_ ) );
AND3_X1 _11732_ ( .A1(_03806_ ), .A2(_03807_ ), .A3(_03808_ ), .ZN(_03809_ ) );
NAND3_X1 _11733_ ( .A1(_03528_ ), .A2(_03805_ ), .A3(_03809_ ), .ZN(_03810_ ) );
OAI21_X1 _11734_ ( .A(_03810_ ), .B1(_03538_ ), .B2(_03542_ ), .ZN(_03811_ ) );
NAND4_X1 _11735_ ( .A1(_03540_ ), .A2(\EX_LS_result_csreg_mem [14] ), .A3(_03095_ ), .A4(_03541_ ), .ZN(_03812_ ) );
AND2_X1 _11736_ ( .A1(_03811_ ), .A2(_03812_ ), .ZN(_03813_ ) );
INV_X1 _11737_ ( .A(_01738_ ), .ZN(_03814_ ) );
AOI221_X4 _11738_ ( .A(_03804_ ), .B1(_03813_ ), .B2(fanout_net_7 ), .C1(_01350_ ), .C2(_03814_ ), .ZN(_03815_ ) );
AOI21_X1 _11739_ ( .A(_03548_ ), .B1(_03811_ ), .B2(_03812_ ), .ZN(_03816_ ) );
OAI21_X1 _11740_ ( .A(_03379_ ), .B1(_03815_ ), .B2(_03816_ ), .ZN(_03817_ ) );
OR3_X2 _11741_ ( .A1(_03511_ ), .A2(_03497_ ), .A3(\EX_LS_result_reg [14] ), .ZN(_03818_ ) );
OR2_X1 _11742_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[0][14] ), .ZN(_03819_ ) );
OAI211_X1 _11743_ ( .A(_03819_ ), .B(_03785_ ), .C1(_03560_ ), .C2(\myreg.Reg[1][14] ), .ZN(_03820_ ) );
OR2_X1 _11744_ ( .A1(fanout_net_24 ), .A2(\myreg.Reg[2][14] ), .ZN(_03821_ ) );
OAI211_X1 _11745_ ( .A(_03821_ ), .B(fanout_net_31 ), .C1(_03560_ ), .C2(\myreg.Reg[3][14] ), .ZN(_03822_ ) );
NAND3_X1 _11746_ ( .A1(_03820_ ), .A2(_03822_ ), .A3(_03782_ ), .ZN(_03823_ ) );
MUX2_X1 _11747_ ( .A(\myreg.Reg[6][14] ), .B(\myreg.Reg[7][14] ), .S(fanout_net_24 ), .Z(_03824_ ) );
MUX2_X1 _11748_ ( .A(\myreg.Reg[4][14] ), .B(\myreg.Reg[5][14] ), .S(fanout_net_25 ), .Z(_03825_ ) );
MUX2_X1 _11749_ ( .A(_03824_ ), .B(_03825_ ), .S(_03785_ ), .Z(_03826_ ) );
OAI211_X1 _11750_ ( .A(_03494_ ), .B(_03823_ ), .C1(_03826_ ), .C2(_03490_ ), .ZN(_03827_ ) );
OR2_X1 _11751_ ( .A1(_03779_ ), .A2(\myreg.Reg[15][14] ), .ZN(_03828_ ) );
OAI211_X1 _11752_ ( .A(_03828_ ), .B(fanout_net_31 ), .C1(fanout_net_25 ), .C2(\myreg.Reg[14][14] ), .ZN(_03829_ ) );
OR2_X1 _11753_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[12][14] ), .ZN(_03830_ ) );
OAI211_X1 _11754_ ( .A(_03830_ ), .B(_03785_ ), .C1(_03560_ ), .C2(\myreg.Reg[13][14] ), .ZN(_03831_ ) );
NAND3_X1 _11755_ ( .A1(_03829_ ), .A2(fanout_net_33 ), .A3(_03831_ ), .ZN(_03832_ ) );
MUX2_X1 _11756_ ( .A(\myreg.Reg[8][14] ), .B(\myreg.Reg[9][14] ), .S(fanout_net_25 ), .Z(_03833_ ) );
MUX2_X1 _11757_ ( .A(\myreg.Reg[10][14] ), .B(\myreg.Reg[11][14] ), .S(fanout_net_25 ), .Z(_03834_ ) );
MUX2_X1 _11758_ ( .A(_03833_ ), .B(_03834_ ), .S(fanout_net_31 ), .Z(_03835_ ) );
OAI211_X1 _11759_ ( .A(fanout_net_34 ), .B(_03832_ ), .C1(_03835_ ), .C2(fanout_net_33 ), .ZN(_03836_ ) );
OAI211_X1 _11760_ ( .A(_03827_ ), .B(_03836_ ), .C1(_03511_ ), .C2(_03497_ ), .ZN(_03837_ ) );
NAND2_X2 _11761_ ( .A1(_03818_ ), .A2(_03837_ ), .ZN(_03838_ ) );
MUX2_X1 _11762_ ( .A(_02333_ ), .B(_03838_ ), .S(_03370_ ), .Z(_03839_ ) );
OAI21_X1 _11763_ ( .A(_03817_ ), .B1(_03552_ ), .B2(_03839_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OR3_X1 _11764_ ( .A1(_03423_ ), .A2(\EX_LS_result_csreg_mem [13] ), .A3(_03431_ ), .ZN(_03840_ ) );
NAND3_X1 _11765_ ( .A1(_03449_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_03452_ ), .ZN(_03841_ ) );
BUF_X4 _11766_ ( .A(_03458_ ), .Z(_03842_ ) );
NAND4_X1 _11767_ ( .A1(_03457_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [13] ), .A4(_03842_ ), .ZN(_03843_ ) );
NAND3_X1 _11768_ ( .A1(_03443_ ), .A2(_03841_ ), .A3(_03843_ ), .ZN(_03844_ ) );
NAND3_X1 _11769_ ( .A1(_03592_ ), .A2(\mepc [13] ), .A3(_03463_ ), .ZN(_03845_ ) );
NAND3_X1 _11770_ ( .A1(_03467_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_03842_ ), .ZN(_03846_ ) );
OAI211_X1 _11771_ ( .A(_03845_ ), .B(_03846_ ), .C1(_03424_ ), .C2(_03432_ ), .ZN(_03847_ ) );
OAI21_X1 _11772_ ( .A(_03840_ ), .B1(_03844_ ), .B2(_03847_ ), .ZN(_03848_ ) );
AOI221_X4 _11773_ ( .A(_03356_ ), .B1(fanout_net_6 ), .B2(_01765_ ), .C1(_03848_ ), .C2(fanout_net_7 ), .ZN(_03849_ ) );
NAND2_X2 _11774_ ( .A1(_01764_ ), .A2(_01784_ ), .ZN(_03850_ ) );
OAI21_X1 _11775_ ( .A(_03849_ ), .B1(_03850_ ), .B2(fanout_net_6 ), .ZN(_03851_ ) );
OR3_X1 _11776_ ( .A1(_03848_ ), .A2(_03700_ ), .A3(_03548_ ), .ZN(_03852_ ) );
OR3_X4 _11777_ ( .A1(_03510_ ), .A2(_03496_ ), .A3(\EX_LS_result_reg [13] ), .ZN(_03853_ ) );
OR2_X1 _11778_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[0][13] ), .ZN(_03854_ ) );
BUF_X4 _11779_ ( .A(_03480_ ), .Z(_03855_ ) );
OAI211_X1 _11780_ ( .A(_03854_ ), .B(_03855_ ), .C1(_03779_ ), .C2(\myreg.Reg[1][13] ), .ZN(_03856_ ) );
OR2_X1 _11781_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[2][13] ), .ZN(_03857_ ) );
OAI211_X1 _11782_ ( .A(_03857_ ), .B(fanout_net_31 ), .C1(_03779_ ), .C2(\myreg.Reg[3][13] ), .ZN(_03858_ ) );
NAND3_X1 _11783_ ( .A1(_03856_ ), .A2(_03858_ ), .A3(_03489_ ), .ZN(_03859_ ) );
MUX2_X1 _11784_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_25 ), .Z(_03860_ ) );
MUX2_X1 _11785_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_25 ), .Z(_03861_ ) );
MUX2_X1 _11786_ ( .A(_03860_ ), .B(_03861_ ), .S(_03784_ ), .Z(_03862_ ) );
OAI211_X1 _11787_ ( .A(_03493_ ), .B(_03859_ ), .C1(_03862_ ), .C2(_03489_ ), .ZN(_03863_ ) );
OR2_X1 _11788_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[14][13] ), .ZN(_03864_ ) );
OAI211_X1 _11789_ ( .A(_03864_ ), .B(fanout_net_31 ), .C1(_03779_ ), .C2(\myreg.Reg[15][13] ), .ZN(_03865_ ) );
OR2_X1 _11790_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[12][13] ), .ZN(_03866_ ) );
OAI211_X1 _11791_ ( .A(_03866_ ), .B(_03784_ ), .C1(_03779_ ), .C2(\myreg.Reg[13][13] ), .ZN(_03867_ ) );
NAND3_X1 _11792_ ( .A1(_03865_ ), .A2(_03867_ ), .A3(fanout_net_33 ), .ZN(_03868_ ) );
MUX2_X1 _11793_ ( .A(\myreg.Reg[8][13] ), .B(\myreg.Reg[9][13] ), .S(fanout_net_25 ), .Z(_03869_ ) );
MUX2_X1 _11794_ ( .A(\myreg.Reg[10][13] ), .B(\myreg.Reg[11][13] ), .S(fanout_net_25 ), .Z(_03870_ ) );
MUX2_X1 _11795_ ( .A(_03869_ ), .B(_03870_ ), .S(fanout_net_31 ), .Z(_03871_ ) );
OAI211_X1 _11796_ ( .A(fanout_net_34 ), .B(_03868_ ), .C1(_03871_ ), .C2(fanout_net_33 ), .ZN(_03872_ ) );
BUF_X4 _11797_ ( .A(_03509_ ), .Z(_03873_ ) );
BUF_X2 _11798_ ( .A(_01377_ ), .Z(_03874_ ) );
OAI211_X2 _11799_ ( .A(_03863_ ), .B(_03872_ ), .C1(_03873_ ), .C2(_03874_ ), .ZN(_03875_ ) );
NAND2_X1 _11800_ ( .A1(_03853_ ), .A2(_03875_ ), .ZN(_03876_ ) );
MUX2_X1 _11801_ ( .A(_02334_ ), .B(_03876_ ), .S(_03590_ ), .Z(_03877_ ) );
OAI211_X1 _11802_ ( .A(_03851_ ), .B(_03852_ ), .C1(_03877_ ), .C2(_03762_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
INV_X1 _11803_ ( .A(_03527_ ), .ZN(_03878_ ) );
NAND4_X1 _11804_ ( .A1(_03690_ ), .A2(_03460_ ), .A3(\mtvec [12] ), .A4(_03691_ ), .ZN(_03879_ ) );
NAND3_X1 _11805_ ( .A1(_03443_ ), .A2(_03878_ ), .A3(_03879_ ), .ZN(_03880_ ) );
NAND3_X1 _11806_ ( .A1(_03765_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_03599_ ), .ZN(_03881_ ) );
NAND3_X1 _11807_ ( .A1(_03765_ ), .A2(\mepc [12] ), .A3(_03463_ ), .ZN(_03882_ ) );
NAND4_X1 _11808_ ( .A1(_03768_ ), .A2(_03460_ ), .A3(\mycsreg.CSReg[0][12] ), .A4(_03691_ ), .ZN(_03883_ ) );
NAND3_X1 _11809_ ( .A1(_03881_ ), .A2(_03882_ ), .A3(_03883_ ), .ZN(_03884_ ) );
OAI21_X1 _11810_ ( .A(_03646_ ), .B1(_03880_ ), .B2(_03884_ ), .ZN(_03885_ ) );
NAND4_X1 _11811_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [12] ), .A3(_03096_ ), .A4(_03606_ ), .ZN(_03886_ ) );
AND2_X1 _11812_ ( .A1(_03885_ ), .A2(_03886_ ), .ZN(_03887_ ) );
AOI22_X1 _11813_ ( .A1(_03887_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01809_ ), .ZN(_03888_ ) );
OAI211_X1 _11814_ ( .A(_03888_ ), .B(_03551_ ), .C1(fanout_net_6 ), .C2(_01808_ ), .ZN(_03889_ ) );
AOI21_X1 _11815_ ( .A(_03700_ ), .B1(_03885_ ), .B2(_03886_ ), .ZN(_03890_ ) );
NAND2_X1 _11816_ ( .A1(_03890_ ), .A2(_03702_ ), .ZN(_03891_ ) );
OR3_X2 _11817_ ( .A1(_03873_ ), .A2(_03496_ ), .A3(\EX_LS_result_reg [12] ), .ZN(_03892_ ) );
OR2_X1 _11818_ ( .A1(_03559_ ), .A2(\myreg.Reg[3][12] ), .ZN(_03893_ ) );
OAI211_X1 _11819_ ( .A(_03893_ ), .B(fanout_net_31 ), .C1(fanout_net_25 ), .C2(\myreg.Reg[2][12] ), .ZN(_03894_ ) );
OR2_X1 _11820_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[0][12] ), .ZN(_03895_ ) );
BUF_X4 _11821_ ( .A(_03559_ ), .Z(_03896_ ) );
OAI211_X1 _11822_ ( .A(_03895_ ), .B(_03855_ ), .C1(_03896_ ), .C2(\myreg.Reg[1][12] ), .ZN(_03897_ ) );
NAND3_X1 _11823_ ( .A1(_03894_ ), .A2(_03489_ ), .A3(_03897_ ), .ZN(_03898_ ) );
MUX2_X1 _11824_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_25 ), .Z(_03899_ ) );
MUX2_X1 _11825_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_25 ), .Z(_03900_ ) );
MUX2_X1 _11826_ ( .A(_03899_ ), .B(_03900_ ), .S(_03855_ ), .Z(_03901_ ) );
OAI211_X1 _11827_ ( .A(_03493_ ), .B(_03898_ ), .C1(_03901_ ), .C2(_03782_ ), .ZN(_03902_ ) );
OR2_X1 _11828_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[14][12] ), .ZN(_03903_ ) );
OAI211_X1 _11829_ ( .A(_03903_ ), .B(fanout_net_31 ), .C1(_03896_ ), .C2(\myreg.Reg[15][12] ), .ZN(_03904_ ) );
OR2_X1 _11830_ ( .A1(fanout_net_25 ), .A2(\myreg.Reg[12][12] ), .ZN(_03905_ ) );
OAI211_X1 _11831_ ( .A(_03905_ ), .B(_03855_ ), .C1(_03896_ ), .C2(\myreg.Reg[13][12] ), .ZN(_03906_ ) );
NAND3_X1 _11832_ ( .A1(_03904_ ), .A2(_03906_ ), .A3(fanout_net_33 ), .ZN(_03907_ ) );
MUX2_X1 _11833_ ( .A(\myreg.Reg[8][12] ), .B(\myreg.Reg[9][12] ), .S(fanout_net_25 ), .Z(_03908_ ) );
MUX2_X1 _11834_ ( .A(\myreg.Reg[10][12] ), .B(\myreg.Reg[11][12] ), .S(fanout_net_25 ), .Z(_03909_ ) );
MUX2_X1 _11835_ ( .A(_03908_ ), .B(_03909_ ), .S(fanout_net_31 ), .Z(_03910_ ) );
OAI211_X1 _11836_ ( .A(fanout_net_34 ), .B(_03907_ ), .C1(_03910_ ), .C2(fanout_net_33 ), .ZN(_03911_ ) );
OAI211_X4 _11837_ ( .A(_03902_ ), .B(_03911_ ), .C1(_03873_ ), .C2(_03497_ ), .ZN(_03912_ ) );
NAND2_X2 _11838_ ( .A1(_03892_ ), .A2(_03912_ ), .ZN(_03913_ ) );
MUX2_X1 _11839_ ( .A(_02335_ ), .B(_03913_ ), .S(_03370_ ), .Z(_03914_ ) );
OAI211_X1 _11840_ ( .A(_03889_ ), .B(_03891_ ), .C1(_03552_ ), .C2(_03914_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
OR3_X1 _11841_ ( .A1(_03553_ ), .A2(_03554_ ), .A3(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_03915_ ) );
OR2_X1 _11842_ ( .A1(_03562_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03916_ ) );
OAI211_X1 _11843_ ( .A(_03916_ ), .B(_03663_ ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03917_ ) );
OR2_X1 _11844_ ( .A1(_03562_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03918_ ) );
OAI211_X1 _11845_ ( .A(_03918_ ), .B(fanout_net_31 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03919_ ) );
NAND3_X1 _11846_ ( .A1(_03917_ ), .A2(_03919_ ), .A3(fanout_net_33 ), .ZN(_03920_ ) );
MUX2_X1 _11847_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03921_ ) );
MUX2_X1 _11848_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03922_ ) );
MUX2_X1 _11849_ ( .A(_03921_ ), .B(_03922_ ), .S(_03573_ ), .Z(_03923_ ) );
OAI211_X1 _11850_ ( .A(_03556_ ), .B(_03920_ ), .C1(_03923_ ), .C2(fanout_net_33 ), .ZN(_03924_ ) );
NOR2_X1 _11851_ ( .A1(_03617_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03925_ ) );
OAI21_X1 _11852_ ( .A(fanout_net_31 ), .B1(fanout_net_25 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03926_ ) );
NOR2_X1 _11853_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03927_ ) );
OAI21_X1 _11854_ ( .A(_03573_ ), .B1(_03741_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03928_ ) );
OAI221_X1 _11855_ ( .A(_03565_ ), .B1(_03925_ ), .B2(_03926_ ), .C1(_03927_ ), .C2(_03928_ ), .ZN(_03929_ ) );
MUX2_X1 _11856_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03930_ ) );
MUX2_X1 _11857_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_03931_ ) );
MUX2_X1 _11858_ ( .A(_03930_ ), .B(_03931_ ), .S(fanout_net_31 ), .Z(_03932_ ) );
OAI211_X1 _11859_ ( .A(fanout_net_34 ), .B(_03929_ ), .C1(_03932_ ), .C2(_03575_ ), .ZN(_03933_ ) );
OAI211_X1 _11860_ ( .A(_03924_ ), .B(_03933_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_03934_ ) );
NAND2_X1 _11861_ ( .A1(_03915_ ), .A2(_03934_ ), .ZN(_03935_ ) );
MUX2_X1 _11862_ ( .A(\ID_EX_pc [30] ), .B(_03935_ ), .S(_03370_ ), .Z(_03936_ ) );
NOR3_X1 _11863_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_03432_ ), .ZN(_03937_ ) );
INV_X1 _11864_ ( .A(_03937_ ), .ZN(_03938_ ) );
NOR2_X1 _11865_ ( .A1(_03423_ ), .A2(_03431_ ), .ZN(_03939_ ) );
AND4_X1 _11866_ ( .A1(\ID_EX_csr [2] ), .A2(_03457_ ), .A3(\mtvec [30] ), .A4(_03459_ ), .ZN(_03940_ ) );
NOR2_X1 _11867_ ( .A1(_03939_ ), .A2(_03940_ ), .ZN(_03941_ ) );
INV_X1 _11868_ ( .A(_03941_ ), .ZN(_03942_ ) );
NAND3_X1 _11869_ ( .A1(_03449_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_03452_ ), .ZN(_03943_ ) );
NAND3_X1 _11870_ ( .A1(_03467_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_03842_ ), .ZN(_03944_ ) );
NAND3_X1 _11871_ ( .A1(_03592_ ), .A2(\mepc [30] ), .A3(_03463_ ), .ZN(_03945_ ) );
NAND4_X1 _11872_ ( .A1(_03442_ ), .A2(_03943_ ), .A3(_03944_ ), .A4(_03945_ ), .ZN(_03946_ ) );
OAI21_X1 _11873_ ( .A(_03938_ ), .B1(_03942_ ), .B2(_03946_ ), .ZN(_03947_ ) );
AOI22_X1 _11874_ ( .A1(_03947_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01447_ ), .ZN(_03948_ ) );
INV_X1 _11875_ ( .A(_01446_ ), .ZN(_03949_ ) );
OAI21_X1 _11876_ ( .A(_03948_ ), .B1(_03949_ ), .B2(fanout_net_6 ), .ZN(_03950_ ) );
OAI211_X1 _11877_ ( .A(_03474_ ), .B(_03938_ ), .C1(_03942_ ), .C2(_03946_ ), .ZN(_03951_ ) );
NAND2_X1 _11878_ ( .A1(_03950_ ), .A2(_03951_ ), .ZN(_03952_ ) );
MUX2_X1 _11879_ ( .A(_03936_ ), .B(_03952_ ), .S(_03551_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _11880_ ( .A1(_03529_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_03685_ ), .ZN(_03953_ ) );
NAND3_X1 _11881_ ( .A1(_03448_ ), .A2(\mepc [11] ), .A3(_03462_ ), .ZN(_03954_ ) );
NAND4_X1 _11882_ ( .A1(_03652_ ), .A2(_03459_ ), .A3(\mtvec [11] ), .A4(_03650_ ), .ZN(_03955_ ) );
NAND4_X1 _11883_ ( .A1(_03594_ ), .A2(_03459_ ), .A3(\mycsreg.CSReg[0][11] ), .A4(_03650_ ), .ZN(_03956_ ) );
AND3_X1 _11884_ ( .A1(_03954_ ), .A2(_03955_ ), .A3(_03956_ ), .ZN(_03957_ ) );
NAND3_X1 _11885_ ( .A1(_03528_ ), .A2(_03953_ ), .A3(_03957_ ), .ZN(_03958_ ) );
OAI21_X1 _11886_ ( .A(_03958_ ), .B1(_03538_ ), .B2(_03542_ ), .ZN(_03959_ ) );
NAND4_X1 _11887_ ( .A1(_03540_ ), .A2(\EX_LS_result_csreg_mem [11] ), .A3(_03095_ ), .A4(_03541_ ), .ZN(_03960_ ) );
AOI21_X1 _11888_ ( .A(_03547_ ), .B1(_03959_ ), .B2(_03960_ ), .ZN(_03961_ ) );
AND2_X1 _11889_ ( .A1(_03959_ ), .A2(_03960_ ), .ZN(_03962_ ) );
AOI22_X1 _11890_ ( .A1(_03962_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01862_ ), .ZN(_03963_ ) );
NAND3_X1 _11891_ ( .A1(_01861_ ), .A2(_01881_ ), .A3(_01350_ ), .ZN(_03964_ ) );
AOI211_X1 _11892_ ( .A(_03357_ ), .B(_03961_ ), .C1(_03963_ ), .C2(_03964_ ), .ZN(_03965_ ) );
OR3_X4 _11893_ ( .A1(_03510_ ), .A2(_03496_ ), .A3(\EX_LS_result_reg [11] ), .ZN(_03966_ ) );
OR2_X1 _11894_ ( .A1(_03558_ ), .A2(\myreg.Reg[3][11] ), .ZN(_03967_ ) );
OAI211_X1 _11895_ ( .A(_03967_ ), .B(fanout_net_32 ), .C1(fanout_net_25 ), .C2(\myreg.Reg[2][11] ), .ZN(_03968_ ) );
OR2_X1 _11896_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[0][11] ), .ZN(_03969_ ) );
OAI211_X1 _11897_ ( .A(_03969_ ), .B(_03784_ ), .C1(_03559_ ), .C2(\myreg.Reg[1][11] ), .ZN(_03970_ ) );
NAND3_X1 _11898_ ( .A1(_03968_ ), .A2(_03488_ ), .A3(_03970_ ), .ZN(_03971_ ) );
MUX2_X1 _11899_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_26 ), .Z(_03972_ ) );
MUX2_X1 _11900_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_26 ), .Z(_03973_ ) );
MUX2_X1 _11901_ ( .A(_03972_ ), .B(_03973_ ), .S(_03784_ ), .Z(_03974_ ) );
OAI211_X1 _11902_ ( .A(_03493_ ), .B(_03971_ ), .C1(_03974_ ), .C2(_03489_ ), .ZN(_03975_ ) );
OR2_X1 _11903_ ( .A1(_03558_ ), .A2(\myreg.Reg[13][11] ), .ZN(_03976_ ) );
OAI211_X1 _11904_ ( .A(_03976_ ), .B(_03784_ ), .C1(fanout_net_26 ), .C2(\myreg.Reg[12][11] ), .ZN(_03977_ ) );
OR2_X1 _11905_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[14][11] ), .ZN(_03978_ ) );
OAI211_X1 _11906_ ( .A(_03978_ ), .B(fanout_net_32 ), .C1(_03559_ ), .C2(\myreg.Reg[15][11] ), .ZN(_03979_ ) );
NAND3_X1 _11907_ ( .A1(_03977_ ), .A2(fanout_net_33 ), .A3(_03979_ ), .ZN(_03980_ ) );
MUX2_X1 _11908_ ( .A(\myreg.Reg[8][11] ), .B(\myreg.Reg[9][11] ), .S(fanout_net_26 ), .Z(_03981_ ) );
MUX2_X1 _11909_ ( .A(\myreg.Reg[10][11] ), .B(\myreg.Reg[11][11] ), .S(fanout_net_26 ), .Z(_03982_ ) );
MUX2_X1 _11910_ ( .A(_03981_ ), .B(_03982_ ), .S(fanout_net_32 ), .Z(_03983_ ) );
OAI211_X1 _11911_ ( .A(fanout_net_34 ), .B(_03980_ ), .C1(_03983_ ), .C2(fanout_net_33 ), .ZN(_03984_ ) );
OAI211_X1 _11912_ ( .A(_03975_ ), .B(_03984_ ), .C1(_03510_ ), .C2(_03874_ ), .ZN(_03985_ ) );
NAND2_X2 _11913_ ( .A1(_03966_ ), .A2(_03985_ ), .ZN(_03986_ ) );
MUX2_X1 _11914_ ( .A(_02337_ ), .B(_03986_ ), .S(_03590_ ), .Z(_03987_ ) );
AOI21_X1 _11915_ ( .A(_03965_ ), .B1(_03358_ ), .B2(_03987_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
AOI21_X1 _11916_ ( .A(fanout_net_6 ), .B1(_01885_ ), .B2(_01904_ ), .ZN(_03988_ ) );
AND2_X1 _11917_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [10] ), .ZN(_03989_ ) );
AND2_X1 _11918_ ( .A1(_03592_ ), .A2(_03463_ ), .ZN(_03990_ ) );
AOI22_X1 _11919_ ( .A1(_03990_ ), .A2(\mepc [10] ), .B1(_03438_ ), .B2(_03599_ ), .ZN(_03991_ ) );
NAND3_X1 _11920_ ( .A1(_03592_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_03452_ ), .ZN(_03992_ ) );
NAND4_X1 _11921_ ( .A1(_03594_ ), .A2(_03842_ ), .A3(\mycsreg.CSReg[0][10] ), .A4(_03595_ ), .ZN(_03993_ ) );
NAND4_X1 _11922_ ( .A1(_03652_ ), .A2(_03530_ ), .A3(\mtvec [10] ), .A4(_03595_ ), .ZN(_03994_ ) );
AND3_X1 _11923_ ( .A1(_03992_ ), .A2(_03993_ ), .A3(_03994_ ), .ZN(_03995_ ) );
NAND2_X1 _11924_ ( .A1(_03991_ ), .A2(_03995_ ), .ZN(_03996_ ) );
OAI21_X1 _11925_ ( .A(_03996_ ), .B1(_03542_ ), .B2(_03538_ ), .ZN(_03997_ ) );
NAND4_X1 _11926_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_03096_ ), .A4(_03606_ ), .ZN(_03998_ ) );
AND2_X1 _11927_ ( .A1(_03997_ ), .A2(_03998_ ), .ZN(_03999_ ) );
INV_X1 _11928_ ( .A(_03999_ ), .ZN(_04000_ ) );
OAI221_X1 _11929_ ( .A(_03378_ ), .B1(_03988_ ), .B2(_03989_ ), .C1(_04000_ ), .C2(_02379_ ), .ZN(_04001_ ) );
AOI21_X1 _11930_ ( .A(_03357_ ), .B1(_03997_ ), .B2(_03998_ ), .ZN(_04002_ ) );
NAND2_X1 _11931_ ( .A1(_04002_ ), .A2(_03702_ ), .ZN(_04003_ ) );
OR3_X2 _11932_ ( .A1(_03510_ ), .A2(_03496_ ), .A3(\EX_LS_result_reg [10] ), .ZN(_04004_ ) );
CLKBUF_X2 _11933_ ( .A(_03557_ ), .Z(_04005_ ) );
OR2_X1 _11934_ ( .A1(_04005_ ), .A2(\myreg.Reg[3][10] ), .ZN(_04006_ ) );
OAI211_X1 _11935_ ( .A(_04006_ ), .B(fanout_net_32 ), .C1(fanout_net_26 ), .C2(\myreg.Reg[2][10] ), .ZN(_04007_ ) );
OR2_X1 _11936_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[0][10] ), .ZN(_04008_ ) );
OAI211_X1 _11937_ ( .A(_04008_ ), .B(_03784_ ), .C1(_03779_ ), .C2(\myreg.Reg[1][10] ), .ZN(_04009_ ) );
NAND3_X1 _11938_ ( .A1(_04007_ ), .A2(_03488_ ), .A3(_04009_ ), .ZN(_04010_ ) );
MUX2_X1 _11939_ ( .A(\myreg.Reg[6][10] ), .B(\myreg.Reg[7][10] ), .S(fanout_net_26 ), .Z(_04011_ ) );
MUX2_X1 _11940_ ( .A(\myreg.Reg[4][10] ), .B(\myreg.Reg[5][10] ), .S(fanout_net_26 ), .Z(_04012_ ) );
MUX2_X1 _11941_ ( .A(_04011_ ), .B(_04012_ ), .S(_03784_ ), .Z(_04013_ ) );
OAI211_X1 _11942_ ( .A(_03493_ ), .B(_04010_ ), .C1(_04013_ ), .C2(_03489_ ), .ZN(_04014_ ) );
OR2_X1 _11943_ ( .A1(_03558_ ), .A2(\myreg.Reg[15][10] ), .ZN(_04015_ ) );
OAI211_X1 _11944_ ( .A(_04015_ ), .B(fanout_net_32 ), .C1(fanout_net_26 ), .C2(\myreg.Reg[14][10] ), .ZN(_04016_ ) );
OR2_X1 _11945_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[12][10] ), .ZN(_04017_ ) );
OAI211_X1 _11946_ ( .A(_04017_ ), .B(_03784_ ), .C1(_03779_ ), .C2(\myreg.Reg[13][10] ), .ZN(_04018_ ) );
NAND3_X1 _11947_ ( .A1(_04016_ ), .A2(fanout_net_33 ), .A3(_04018_ ), .ZN(_04019_ ) );
MUX2_X1 _11948_ ( .A(\myreg.Reg[8][10] ), .B(\myreg.Reg[9][10] ), .S(fanout_net_26 ), .Z(_04020_ ) );
MUX2_X1 _11949_ ( .A(\myreg.Reg[10][10] ), .B(\myreg.Reg[11][10] ), .S(fanout_net_26 ), .Z(_04021_ ) );
MUX2_X1 _11950_ ( .A(_04020_ ), .B(_04021_ ), .S(fanout_net_32 ), .Z(_04022_ ) );
OAI211_X1 _11951_ ( .A(fanout_net_34 ), .B(_04019_ ), .C1(_04022_ ), .C2(fanout_net_33 ), .ZN(_04023_ ) );
OAI211_X1 _11952_ ( .A(_04014_ ), .B(_04023_ ), .C1(_03873_ ), .C2(_03874_ ), .ZN(_04024_ ) );
NAND2_X2 _11953_ ( .A1(_04004_ ), .A2(_04024_ ), .ZN(_04025_ ) );
MUX2_X1 _11954_ ( .A(_02338_ ), .B(_04025_ ), .S(_03370_ ), .Z(_04026_ ) );
OAI211_X1 _11955_ ( .A(_04001_ ), .B(_04003_ ), .C1(_03552_ ), .C2(_04026_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
NAND3_X1 _11956_ ( .A1(_03448_ ), .A2(\mepc [9] ), .A3(_03462_ ), .ZN(_04027_ ) );
NAND4_X1 _11957_ ( .A1(_03594_ ), .A2(_03530_ ), .A3(\mycsreg.CSReg[0][9] ), .A4(_03595_ ), .ZN(_04028_ ) );
AND2_X1 _11958_ ( .A1(_04027_ ), .A2(_04028_ ), .ZN(_04029_ ) );
AND4_X1 _11959_ ( .A1(\mtvec [9] ), .A2(_03533_ ), .A3(_03458_ ), .A4(_03456_ ), .ZN(_04030_ ) );
AOI21_X1 _11960_ ( .A(_04030_ ), .B1(_03438_ ), .B2(_03599_ ), .ZN(_04031_ ) );
NAND3_X1 _11961_ ( .A1(_03765_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_03599_ ), .ZN(_04032_ ) );
NAND3_X1 _11962_ ( .A1(_04029_ ), .A2(_04031_ ), .A3(_04032_ ), .ZN(_04033_ ) );
OAI21_X1 _11963_ ( .A(_04033_ ), .B1(_03538_ ), .B2(_03542_ ), .ZN(_04034_ ) );
NAND4_X1 _11964_ ( .A1(_03540_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_03095_ ), .A4(_03541_ ), .ZN(_04035_ ) );
AOI21_X1 _11965_ ( .A(_03547_ ), .B1(_04034_ ), .B2(_04035_ ), .ZN(_04036_ ) );
AND2_X1 _11966_ ( .A1(_04034_ ), .A2(_04035_ ), .ZN(_04037_ ) );
AOI22_X1 _11967_ ( .A1(_04037_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01857_ ), .ZN(_04038_ ) );
NAND3_X1 _11968_ ( .A1(_01834_ ), .A2(_01853_ ), .A3(_01350_ ), .ZN(_04039_ ) );
AOI211_X1 _11969_ ( .A(_03357_ ), .B(_04036_ ), .C1(_04038_ ), .C2(_04039_ ), .ZN(_04040_ ) );
OR3_X4 _11970_ ( .A1(_03510_ ), .A2(_03496_ ), .A3(\EX_LS_result_reg [9] ), .ZN(_04041_ ) );
OR2_X1 _11971_ ( .A1(_03558_ ), .A2(\myreg.Reg[3][9] ), .ZN(_04042_ ) );
OAI211_X1 _11972_ ( .A(_04042_ ), .B(fanout_net_32 ), .C1(fanout_net_26 ), .C2(\myreg.Reg[2][9] ), .ZN(_04043_ ) );
OR2_X1 _11973_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[0][9] ), .ZN(_04044_ ) );
OAI211_X1 _11974_ ( .A(_04044_ ), .B(_03784_ ), .C1(_03559_ ), .C2(\myreg.Reg[1][9] ), .ZN(_04045_ ) );
NAND3_X1 _11975_ ( .A1(_04043_ ), .A2(_03488_ ), .A3(_04045_ ), .ZN(_04046_ ) );
MUX2_X1 _11976_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_26 ), .Z(_04047_ ) );
MUX2_X1 _11977_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_26 ), .Z(_04048_ ) );
MUX2_X1 _11978_ ( .A(_04047_ ), .B(_04048_ ), .S(_03480_ ), .Z(_04049_ ) );
OAI211_X1 _11979_ ( .A(_03492_ ), .B(_04046_ ), .C1(_04049_ ), .C2(_03488_ ), .ZN(_04050_ ) );
OR2_X1 _11980_ ( .A1(_03558_ ), .A2(\myreg.Reg[15][9] ), .ZN(_04051_ ) );
OAI211_X1 _11981_ ( .A(_04051_ ), .B(fanout_net_32 ), .C1(fanout_net_26 ), .C2(\myreg.Reg[14][9] ), .ZN(_04052_ ) );
OR2_X1 _11982_ ( .A1(_03558_ ), .A2(\myreg.Reg[13][9] ), .ZN(_04053_ ) );
OAI211_X1 _11983_ ( .A(_04053_ ), .B(_03480_ ), .C1(fanout_net_26 ), .C2(\myreg.Reg[12][9] ), .ZN(_04054_ ) );
NAND3_X1 _11984_ ( .A1(_04052_ ), .A2(_04054_ ), .A3(fanout_net_33 ), .ZN(_04055_ ) );
MUX2_X1 _11985_ ( .A(\myreg.Reg[8][9] ), .B(\myreg.Reg[9][9] ), .S(fanout_net_26 ), .Z(_04056_ ) );
MUX2_X1 _11986_ ( .A(\myreg.Reg[10][9] ), .B(\myreg.Reg[11][9] ), .S(fanout_net_26 ), .Z(_04057_ ) );
MUX2_X1 _11987_ ( .A(_04056_ ), .B(_04057_ ), .S(fanout_net_32 ), .Z(_04058_ ) );
OAI211_X1 _11988_ ( .A(fanout_net_34 ), .B(_04055_ ), .C1(_04058_ ), .C2(fanout_net_33 ), .ZN(_04059_ ) );
OAI211_X2 _11989_ ( .A(_04050_ ), .B(_04059_ ), .C1(_03510_ ), .C2(_03496_ ), .ZN(_04060_ ) );
NAND2_X2 _11990_ ( .A1(_04041_ ), .A2(_04060_ ), .ZN(_04061_ ) );
MUX2_X1 _11991_ ( .A(_02339_ ), .B(_04061_ ), .S(_03590_ ), .Z(_04062_ ) );
AOI21_X1 _11992_ ( .A(_04040_ ), .B1(_03358_ ), .B2(_04062_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _11993_ ( .A(fanout_net_6 ), .B1(_01812_ ), .B2(_01831_ ), .ZN(_04063_ ) );
AND2_X1 _11994_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [8] ), .ZN(_04064_ ) );
BUF_X4 _11995_ ( .A(_03592_ ), .Z(_04065_ ) );
BUF_X4 _11996_ ( .A(_03462_ ), .Z(_04066_ ) );
NAND3_X1 _11997_ ( .A1(_04065_ ), .A2(\mepc [8] ), .A3(_04066_ ), .ZN(_04067_ ) );
NAND3_X1 _11998_ ( .A1(_03443_ ), .A2(_03878_ ), .A3(_04067_ ), .ZN(_04068_ ) );
BUF_X4 _11999_ ( .A(_03452_ ), .Z(_04069_ ) );
NAND3_X1 _12000_ ( .A1(_04065_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_04069_ ), .ZN(_04070_ ) );
BUF_X4 _12001_ ( .A(_03842_ ), .Z(_04071_ ) );
BUF_X4 _12002_ ( .A(_03595_ ), .Z(_04072_ ) );
NAND4_X1 _12003_ ( .A1(_03768_ ), .A2(_04071_ ), .A3(\mycsreg.CSReg[0][8] ), .A4(_04072_ ), .ZN(_04073_ ) );
NAND4_X1 _12004_ ( .A1(_03690_ ), .A2(_03685_ ), .A3(\mtvec [8] ), .A4(_04072_ ), .ZN(_04074_ ) );
NAND3_X1 _12005_ ( .A1(_04070_ ), .A2(_04073_ ), .A3(_04074_ ), .ZN(_04075_ ) );
OAI21_X1 _12006_ ( .A(_03646_ ), .B1(_04068_ ), .B2(_04075_ ), .ZN(_04076_ ) );
BUF_X4 _12007_ ( .A(_03095_ ), .Z(_04077_ ) );
NAND4_X1 _12008_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [8] ), .A3(_04077_ ), .A4(_03606_ ), .ZN(_04078_ ) );
AND2_X1 _12009_ ( .A1(_04076_ ), .A2(_04078_ ), .ZN(_04079_ ) );
INV_X1 _12010_ ( .A(_04079_ ), .ZN(_04080_ ) );
OAI221_X1 _12011_ ( .A(_03378_ ), .B1(_04063_ ), .B2(_04064_ ), .C1(_04080_ ), .C2(_02379_ ), .ZN(_04081_ ) );
AOI21_X1 _12012_ ( .A(_03700_ ), .B1(_04076_ ), .B2(_04078_ ), .ZN(_04082_ ) );
NAND2_X1 _12013_ ( .A1(_04082_ ), .A2(_03702_ ), .ZN(_04083_ ) );
OR3_X2 _12014_ ( .A1(_03873_ ), .A2(_03874_ ), .A3(\EX_LS_result_reg [8] ), .ZN(_04084_ ) );
OR2_X1 _12015_ ( .A1(_03559_ ), .A2(\myreg.Reg[3][8] ), .ZN(_04085_ ) );
OAI211_X1 _12016_ ( .A(_04085_ ), .B(fanout_net_32 ), .C1(fanout_net_26 ), .C2(\myreg.Reg[2][8] ), .ZN(_04086_ ) );
OR2_X1 _12017_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[0][8] ), .ZN(_04087_ ) );
OAI211_X1 _12018_ ( .A(_04087_ ), .B(_03481_ ), .C1(_03560_ ), .C2(\myreg.Reg[1][8] ), .ZN(_04088_ ) );
NAND3_X1 _12019_ ( .A1(_04086_ ), .A2(_03782_ ), .A3(_04088_ ), .ZN(_04089_ ) );
MUX2_X1 _12020_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_26 ), .Z(_04090_ ) );
MUX2_X1 _12021_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_26 ), .Z(_04091_ ) );
MUX2_X1 _12022_ ( .A(_04090_ ), .B(_04091_ ), .S(_03481_ ), .Z(_04092_ ) );
OAI211_X1 _12023_ ( .A(_03493_ ), .B(_04089_ ), .C1(_04092_ ), .C2(_03782_ ), .ZN(_04093_ ) );
OR2_X1 _12024_ ( .A1(_03559_ ), .A2(\myreg.Reg[13][8] ), .ZN(_04094_ ) );
OAI211_X1 _12025_ ( .A(_04094_ ), .B(_03785_ ), .C1(fanout_net_26 ), .C2(\myreg.Reg[12][8] ), .ZN(_04095_ ) );
OR2_X1 _12026_ ( .A1(fanout_net_26 ), .A2(\myreg.Reg[14][8] ), .ZN(_04096_ ) );
OAI211_X1 _12027_ ( .A(_04096_ ), .B(fanout_net_32 ), .C1(_03896_ ), .C2(\myreg.Reg[15][8] ), .ZN(_04097_ ) );
NAND3_X1 _12028_ ( .A1(_04095_ ), .A2(fanout_net_33 ), .A3(_04097_ ), .ZN(_04098_ ) );
MUX2_X1 _12029_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_26 ), .Z(_04099_ ) );
MUX2_X1 _12030_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_27 ), .Z(_04100_ ) );
MUX2_X1 _12031_ ( .A(_04099_ ), .B(_04100_ ), .S(fanout_net_32 ), .Z(_04101_ ) );
OAI211_X1 _12032_ ( .A(fanout_net_34 ), .B(_04098_ ), .C1(_04101_ ), .C2(fanout_net_33 ), .ZN(_04102_ ) );
OAI211_X1 _12033_ ( .A(_04093_ ), .B(_04102_ ), .C1(_03511_ ), .C2(_03497_ ), .ZN(_04103_ ) );
NAND2_X2 _12034_ ( .A1(_04084_ ), .A2(_04103_ ), .ZN(_04104_ ) );
MUX2_X1 _12035_ ( .A(_02340_ ), .B(_04104_ ), .S(_03370_ ), .Z(_04105_ ) );
OAI211_X1 _12036_ ( .A(_04081_ ), .B(_04083_ ), .C1(_03552_ ), .C2(_04105_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
BUF_X2 _12037_ ( .A(_03642_ ), .Z(_04106_ ) );
BUF_X2 _12038_ ( .A(_03644_ ), .Z(_04107_ ) );
NAND3_X1 _12039_ ( .A1(_04106_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_04107_ ), .ZN(_04108_ ) );
NAND3_X1 _12040_ ( .A1(_03448_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_03452_ ), .ZN(_04109_ ) );
NAND3_X1 _12041_ ( .A1(_03448_ ), .A2(\mepc [7] ), .A3(_03462_ ), .ZN(_04110_ ) );
NAND4_X1 _12042_ ( .A1(_03652_ ), .A2(_03530_ ), .A3(\mtvec [7] ), .A4(_03595_ ), .ZN(_04111_ ) );
NAND4_X1 _12043_ ( .A1(_03594_ ), .A2(_03530_ ), .A3(\mycsreg.CSReg[0][7] ), .A4(_03650_ ), .ZN(_04112_ ) );
AND4_X1 _12044_ ( .A1(_04109_ ), .A2(_04110_ ), .A3(_04111_ ), .A4(_04112_ ), .ZN(_04113_ ) );
OAI21_X1 _12045_ ( .A(_04108_ ), .B1(_03645_ ), .B2(_04113_ ), .ZN(_04114_ ) );
AOI22_X1 _12046_ ( .A1(_04114_ ), .A2(_03474_ ), .B1(fanout_net_6 ), .B2(\ID_EX_imm [7] ), .ZN(_04115_ ) );
INV_X1 _12047_ ( .A(_01684_ ), .ZN(_04116_ ) );
OAI21_X1 _12048_ ( .A(_04115_ ), .B1(_04116_ ), .B2(fanout_net_6 ), .ZN(_04117_ ) );
OR3_X1 _12049_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_03432_ ), .ZN(_04118_ ) );
BUF_X4 _12050_ ( .A(_03457_ ), .Z(_04119_ ) );
BUF_X4 _12051_ ( .A(_03842_ ), .Z(_04120_ ) );
NAND4_X1 _12052_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [7] ), .A4(_04120_ ), .ZN(_04121_ ) );
BUF_X2 _12053_ ( .A(_03467_ ), .Z(_04122_ ) );
NAND3_X1 _12054_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_04120_ ), .ZN(_04123_ ) );
NAND4_X1 _12055_ ( .A1(_04121_ ), .A2(_04109_ ), .A3(_04110_ ), .A4(_04123_ ), .ZN(_04124_ ) );
OAI21_X1 _12056_ ( .A(_04118_ ), .B1(_04124_ ), .B2(_03939_ ), .ZN(_04125_ ) );
AOI21_X1 _12057_ ( .A(_03356_ ), .B1(_04125_ ), .B2(fanout_net_7 ), .ZN(_04126_ ) );
AND2_X1 _12058_ ( .A1(_04117_ ), .A2(_04126_ ), .ZN(_04127_ ) );
AND4_X1 _12059_ ( .A1(_02341_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_04128_ ) );
OR3_X4 _12060_ ( .A1(_03873_ ), .A2(_03874_ ), .A3(\EX_LS_result_reg [7] ), .ZN(_04129_ ) );
OR2_X1 _12061_ ( .A1(_03559_ ), .A2(\myreg.Reg[11][7] ), .ZN(_04130_ ) );
OAI211_X1 _12062_ ( .A(_04130_ ), .B(fanout_net_32 ), .C1(fanout_net_27 ), .C2(\myreg.Reg[10][7] ), .ZN(_04131_ ) );
OR2_X1 _12063_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[8][7] ), .ZN(_04132_ ) );
OAI211_X1 _12064_ ( .A(_04132_ ), .B(_03785_ ), .C1(_03560_ ), .C2(\myreg.Reg[9][7] ), .ZN(_04133_ ) );
NAND3_X1 _12065_ ( .A1(_04131_ ), .A2(_03782_ ), .A3(_04133_ ), .ZN(_04134_ ) );
MUX2_X1 _12066_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_27 ), .Z(_04135_ ) );
MUX2_X1 _12067_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_27 ), .Z(_04136_ ) );
MUX2_X1 _12068_ ( .A(_04135_ ), .B(_04136_ ), .S(_03481_ ), .Z(_04137_ ) );
OAI211_X1 _12069_ ( .A(fanout_net_34 ), .B(_04134_ ), .C1(_04137_ ), .C2(_03490_ ), .ZN(_04138_ ) );
NOR2_X1 _12070_ ( .A1(_03896_ ), .A2(\myreg.Reg[3][7] ), .ZN(_04139_ ) );
OAI21_X1 _12071_ ( .A(fanout_net_32 ), .B1(fanout_net_27 ), .B2(\myreg.Reg[2][7] ), .ZN(_04140_ ) );
NOR2_X1 _12072_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[0][7] ), .ZN(_04141_ ) );
OAI21_X1 _12073_ ( .A(_03481_ ), .B1(_03896_ ), .B2(\myreg.Reg[1][7] ), .ZN(_04142_ ) );
OAI221_X1 _12074_ ( .A(_03489_ ), .B1(_04139_ ), .B2(_04140_ ), .C1(_04141_ ), .C2(_04142_ ), .ZN(_04143_ ) );
MUX2_X1 _12075_ ( .A(\myreg.Reg[6][7] ), .B(\myreg.Reg[7][7] ), .S(fanout_net_27 ), .Z(_04144_ ) );
MUX2_X1 _12076_ ( .A(\myreg.Reg[4][7] ), .B(\myreg.Reg[5][7] ), .S(fanout_net_27 ), .Z(_04145_ ) );
MUX2_X1 _12077_ ( .A(_04144_ ), .B(_04145_ ), .S(_03481_ ), .Z(_04146_ ) );
OAI211_X1 _12078_ ( .A(_03493_ ), .B(_04143_ ), .C1(_04146_ ), .C2(_03490_ ), .ZN(_04147_ ) );
OAI211_X4 _12079_ ( .A(_04138_ ), .B(_04147_ ), .C1(_03511_ ), .C2(_03497_ ), .ZN(_04148_ ) );
NAND2_X4 _12080_ ( .A1(_04129_ ), .A2(_04148_ ), .ZN(_04149_ ) );
AOI211_X1 _12081_ ( .A(_03378_ ), .B(_04128_ ), .C1(_04149_ ), .C2(_03362_ ), .ZN(_04150_ ) );
OR2_X1 _12082_ ( .A1(_04127_ ), .A2(_04150_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
OR3_X4 _12083_ ( .A1(_03510_ ), .A2(_03496_ ), .A3(\EX_LS_result_reg [6] ), .ZN(_04151_ ) );
OR2_X1 _12084_ ( .A1(_04005_ ), .A2(\myreg.Reg[1][6] ), .ZN(_04152_ ) );
OAI211_X1 _12085_ ( .A(_04152_ ), .B(_03481_ ), .C1(fanout_net_27 ), .C2(\myreg.Reg[0][6] ), .ZN(_04153_ ) );
OR2_X1 _12086_ ( .A1(_04005_ ), .A2(\myreg.Reg[3][6] ), .ZN(_04154_ ) );
OAI211_X1 _12087_ ( .A(_04154_ ), .B(fanout_net_32 ), .C1(fanout_net_27 ), .C2(\myreg.Reg[2][6] ), .ZN(_04155_ ) );
NAND3_X1 _12088_ ( .A1(_04153_ ), .A2(_04155_ ), .A3(_03489_ ), .ZN(_04156_ ) );
MUX2_X1 _12089_ ( .A(\myreg.Reg[6][6] ), .B(\myreg.Reg[7][6] ), .S(fanout_net_27 ), .Z(_04157_ ) );
MUX2_X1 _12090_ ( .A(\myreg.Reg[4][6] ), .B(\myreg.Reg[5][6] ), .S(fanout_net_27 ), .Z(_04158_ ) );
MUX2_X1 _12091_ ( .A(_04157_ ), .B(_04158_ ), .S(_03855_ ), .Z(_04159_ ) );
OAI211_X1 _12092_ ( .A(_03493_ ), .B(_04156_ ), .C1(_04159_ ), .C2(_03782_ ), .ZN(_04160_ ) );
OR2_X1 _12093_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[14][6] ), .ZN(_04161_ ) );
OAI211_X1 _12094_ ( .A(_04161_ ), .B(fanout_net_32 ), .C1(_03896_ ), .C2(\myreg.Reg[15][6] ), .ZN(_04162_ ) );
OR2_X1 _12095_ ( .A1(fanout_net_27 ), .A2(\myreg.Reg[12][6] ), .ZN(_04163_ ) );
OAI211_X1 _12096_ ( .A(_04163_ ), .B(_03855_ ), .C1(_03779_ ), .C2(\myreg.Reg[13][6] ), .ZN(_04164_ ) );
NAND3_X1 _12097_ ( .A1(_04162_ ), .A2(_04164_ ), .A3(fanout_net_33 ), .ZN(_04165_ ) );
MUX2_X1 _12098_ ( .A(\myreg.Reg[8][6] ), .B(\myreg.Reg[9][6] ), .S(fanout_net_27 ), .Z(_04166_ ) );
MUX2_X1 _12099_ ( .A(\myreg.Reg[10][6] ), .B(\myreg.Reg[11][6] ), .S(fanout_net_27 ), .Z(_04167_ ) );
MUX2_X1 _12100_ ( .A(_04166_ ), .B(_04167_ ), .S(fanout_net_32 ), .Z(_04168_ ) );
OAI211_X1 _12101_ ( .A(fanout_net_34 ), .B(_04165_ ), .C1(_04168_ ), .C2(fanout_net_33 ), .ZN(_04169_ ) );
OAI211_X4 _12102_ ( .A(_04160_ ), .B(_04169_ ), .C1(_03873_ ), .C2(_03874_ ), .ZN(_04170_ ) );
NAND2_X1 _12103_ ( .A1(_04151_ ), .A2(_04170_ ), .ZN(_04171_ ) );
INV_X1 _12104_ ( .A(_04171_ ), .ZN(_04172_ ) );
MUX2_X1 _12105_ ( .A(\ID_EX_pc [6] ), .B(_04172_ ), .S(_03361_ ), .Z(_04173_ ) );
NAND3_X1 _12106_ ( .A1(_04106_ ), .A2(_03251_ ), .A3(_04107_ ), .ZN(_04174_ ) );
OR2_X2 _12107_ ( .A1(_03645_ ), .A2(_03441_ ), .ZN(_04175_ ) );
NAND3_X1 _12108_ ( .A1(_03449_ ), .A2(\mepc [6] ), .A3(_03463_ ), .ZN(_04176_ ) );
NAND3_X1 _12109_ ( .A1(_03449_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_03452_ ), .ZN(_04177_ ) );
NAND4_X1 _12110_ ( .A1(_03768_ ), .A2(_03842_ ), .A3(\mycsreg.CSReg[0][6] ), .A4(_03691_ ), .ZN(_04178_ ) );
NAND4_X1 _12111_ ( .A1(_03652_ ), .A2(_03842_ ), .A3(\mtvec [6] ), .A4(_03595_ ), .ZN(_04179_ ) );
NAND4_X1 _12112_ ( .A1(_04176_ ), .A2(_04177_ ), .A3(_04178_ ), .A4(_04179_ ), .ZN(_04180_ ) );
OAI21_X1 _12113_ ( .A(_04174_ ), .B1(_04175_ ), .B2(_04180_ ), .ZN(_04181_ ) );
AOI22_X1 _12114_ ( .A1(_04181_ ), .A2(fanout_net_7 ), .B1(fanout_net_6 ), .B2(_01708_ ), .ZN(_04182_ ) );
OAI21_X1 _12115_ ( .A(_04182_ ), .B1(fanout_net_6 ), .B2(_01707_ ), .ZN(_04183_ ) );
OAI211_X1 _12116_ ( .A(_03474_ ), .B(_04174_ ), .C1(_04175_ ), .C2(_04180_ ), .ZN(_04184_ ) );
NAND2_X1 _12117_ ( .A1(_04183_ ), .A2(_04184_ ), .ZN(_04185_ ) );
MUX2_X1 _12118_ ( .A(_04173_ ), .B(_04185_ ), .S(_03551_ ), .Z(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
NAND3_X1 _12119_ ( .A1(_04106_ ), .A2(_03238_ ), .A3(_04107_ ), .ZN(_04186_ ) );
NAND3_X1 _12120_ ( .A1(_03765_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_03599_ ), .ZN(_04187_ ) );
NAND3_X1 _12121_ ( .A1(_03765_ ), .A2(\mepc [5] ), .A3(_03463_ ), .ZN(_04188_ ) );
NAND4_X1 _12122_ ( .A1(_03690_ ), .A2(_03685_ ), .A3(\mtvec [5] ), .A4(_04072_ ), .ZN(_04189_ ) );
NAND4_X1 _12123_ ( .A1(_03768_ ), .A2(_03685_ ), .A3(\mycsreg.CSReg[0][5] ), .A4(_03691_ ), .ZN(_04190_ ) );
NAND4_X1 _12124_ ( .A1(_04187_ ), .A2(_04188_ ), .A3(_04189_ ), .A4(_04190_ ), .ZN(_04191_ ) );
OAI211_X1 _12125_ ( .A(_03474_ ), .B(_04186_ ), .C1(_04175_ ), .C2(_04191_ ), .ZN(_04192_ ) );
INV_X1 _12126_ ( .A(_04192_ ), .ZN(_04193_ ) );
AND2_X1 _12127_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [5] ), .ZN(_04194_ ) );
OR2_X1 _12128_ ( .A1(_04193_ ), .A2(_04194_ ), .ZN(_04195_ ) );
AOI21_X1 _12129_ ( .A(_04195_ ), .B1(_02381_ ), .B2(_01657_ ), .ZN(_04196_ ) );
BUF_X2 _12130_ ( .A(_03423_ ), .Z(_04197_ ) );
BUF_X2 _12131_ ( .A(_03431_ ), .Z(_04198_ ) );
NOR3_X1 _12132_ ( .A1(_04197_ ), .A2(\EX_LS_result_csreg_mem [5] ), .A3(_04198_ ), .ZN(_04199_ ) );
BUF_X2 _12133_ ( .A(_03460_ ), .Z(_04200_ ) );
NAND4_X1 _12134_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [5] ), .A4(_04200_ ), .ZN(_04201_ ) );
AND4_X1 _12135_ ( .A1(_03443_ ), .A2(_04187_ ), .A3(_04188_ ), .A4(_04201_ ), .ZN(_04202_ ) );
AND3_X1 _12136_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_04200_ ), .ZN(_04203_ ) );
NOR2_X1 _12137_ ( .A1(_03939_ ), .A2(_04203_ ), .ZN(_04204_ ) );
AOI21_X1 _12138_ ( .A(_04199_ ), .B1(_04202_ ), .B2(_04204_ ), .ZN(_04205_ ) );
OAI21_X1 _12139_ ( .A(_03698_ ), .B1(_04205_ ), .B2(_02379_ ), .ZN(_04206_ ) );
OR3_X4 _12140_ ( .A1(_03510_ ), .A2(_03496_ ), .A3(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04207_ ) );
OR2_X1 _12141_ ( .A1(_04005_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04208_ ) );
OAI211_X1 _12142_ ( .A(_04208_ ), .B(_03481_ ), .C1(fanout_net_27 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04209_ ) );
OR2_X1 _12143_ ( .A1(_04005_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04210_ ) );
OAI211_X1 _12144_ ( .A(_04210_ ), .B(fanout_net_32 ), .C1(fanout_net_27 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04211_ ) );
NAND3_X1 _12145_ ( .A1(_04209_ ), .A2(_04211_ ), .A3(_03489_ ), .ZN(_04212_ ) );
MUX2_X1 _12146_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04213_ ) );
MUX2_X1 _12147_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04214_ ) );
MUX2_X1 _12148_ ( .A(_04213_ ), .B(_04214_ ), .S(_03855_ ), .Z(_04215_ ) );
OAI211_X1 _12149_ ( .A(_03493_ ), .B(_04212_ ), .C1(_04215_ ), .C2(_03782_ ), .ZN(_04216_ ) );
OR2_X1 _12150_ ( .A1(_04005_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04217_ ) );
OAI211_X1 _12151_ ( .A(_04217_ ), .B(_03855_ ), .C1(fanout_net_27 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04218_ ) );
NAND2_X1 _12152_ ( .A1(_01647_ ), .A2(fanout_net_27 ), .ZN(_04219_ ) );
OAI211_X1 _12153_ ( .A(_04219_ ), .B(fanout_net_32 ), .C1(fanout_net_27 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04220_ ) );
NAND3_X1 _12154_ ( .A1(_04218_ ), .A2(fanout_net_33 ), .A3(_04220_ ), .ZN(_04221_ ) );
MUX2_X1 _12155_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04222_ ) );
MUX2_X1 _12156_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_04223_ ) );
MUX2_X1 _12157_ ( .A(_04222_ ), .B(_04223_ ), .S(fanout_net_32 ), .Z(_04224_ ) );
OAI211_X1 _12158_ ( .A(fanout_net_34 ), .B(_04221_ ), .C1(_04224_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04225_ ) );
OAI211_X1 _12159_ ( .A(_04216_ ), .B(_04225_ ), .C1(_03873_ ), .C2(_03874_ ), .ZN(_04226_ ) );
NAND2_X1 _12160_ ( .A1(_04207_ ), .A2(_04226_ ), .ZN(_04227_ ) );
INV_X1 _12161_ ( .A(_04227_ ), .ZN(_04228_ ) );
MUX2_X1 _12162_ ( .A(_02342_ ), .B(_04228_ ), .S(_03370_ ), .Z(_04229_ ) );
OAI22_X1 _12163_ ( .A1(_04196_ ), .A2(_04206_ ), .B1(_03762_ ), .B2(_04229_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
NAND3_X1 _12164_ ( .A1(_04106_ ), .A2(_03239_ ), .A3(_04107_ ), .ZN(_04230_ ) );
NAND3_X1 _12165_ ( .A1(_03765_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_03599_ ), .ZN(_04231_ ) );
NAND3_X1 _12166_ ( .A1(_03449_ ), .A2(\mepc [4] ), .A3(_03463_ ), .ZN(_04232_ ) );
NAND4_X1 _12167_ ( .A1(_03768_ ), .A2(_03460_ ), .A3(\mycsreg.CSReg[0][4] ), .A4(_03691_ ), .ZN(_04233_ ) );
NAND4_X1 _12168_ ( .A1(_03690_ ), .A2(_03460_ ), .A3(\mtvec [4] ), .A4(_03691_ ), .ZN(_04234_ ) );
NAND4_X1 _12169_ ( .A1(_04231_ ), .A2(_04232_ ), .A3(_04233_ ), .A4(_04234_ ), .ZN(_04235_ ) );
OAI211_X1 _12170_ ( .A(_03474_ ), .B(_04230_ ), .C1(_04175_ ), .C2(_04235_ ), .ZN(_04236_ ) );
INV_X1 _12171_ ( .A(_04236_ ), .ZN(_04237_ ) );
AOI21_X1 _12172_ ( .A(_04237_ ), .B1(fanout_net_6 ), .B2(\ID_EX_imm [4] ), .ZN(_04238_ ) );
INV_X1 _12173_ ( .A(_03394_ ), .ZN(_04239_ ) );
OAI21_X1 _12174_ ( .A(_04238_ ), .B1(fanout_net_6 ), .B2(_04239_ ), .ZN(_04240_ ) );
NOR3_X1 _12175_ ( .A1(_04197_ ), .A2(\EX_LS_result_csreg_mem [4] ), .A3(_04198_ ), .ZN(_04241_ ) );
NAND4_X1 _12176_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [4] ), .A4(_04200_ ), .ZN(_04242_ ) );
AND4_X1 _12177_ ( .A1(_03443_ ), .A2(_04231_ ), .A3(_04232_ ), .A4(_04242_ ), .ZN(_04243_ ) );
AND3_X1 _12178_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_04200_ ), .ZN(_04244_ ) );
NOR2_X1 _12179_ ( .A1(_03939_ ), .A2(_04244_ ), .ZN(_04245_ ) );
AOI21_X1 _12180_ ( .A(_04241_ ), .B1(_04243_ ), .B2(_04245_ ), .ZN(_04246_ ) );
OAI211_X1 _12181_ ( .A(_04240_ ), .B(_03379_ ), .C1(_02379_ ), .C2(_04246_ ), .ZN(_04247_ ) );
BUF_X4 _12182_ ( .A(_03700_ ), .Z(_04248_ ) );
NAND4_X1 _12183_ ( .A1(_02343_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_04249_ ) );
OR3_X4 _12184_ ( .A1(_03511_ ), .A2(_03874_ ), .A3(\EX_LS_result_reg [4] ), .ZN(_04250_ ) );
OR2_X1 _12185_ ( .A1(_03779_ ), .A2(\myreg.Reg[5][4] ), .ZN(_04251_ ) );
OAI211_X1 _12186_ ( .A(_04251_ ), .B(_03785_ ), .C1(fanout_net_27 ), .C2(\myreg.Reg[4][4] ), .ZN(_04252_ ) );
OR2_X1 _12187_ ( .A1(_03559_ ), .A2(\myreg.Reg[7][4] ), .ZN(_04253_ ) );
OAI211_X1 _12188_ ( .A(_04253_ ), .B(fanout_net_32 ), .C1(fanout_net_27 ), .C2(\myreg.Reg[6][4] ), .ZN(_04254_ ) );
NAND3_X1 _12189_ ( .A1(_04252_ ), .A2(_04254_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04255_ ) );
MUX2_X1 _12190_ ( .A(\myreg.Reg[2][4] ), .B(\myreg.Reg[3][4] ), .S(fanout_net_27 ), .Z(_04256_ ) );
MUX2_X1 _12191_ ( .A(\myreg.Reg[0][4] ), .B(\myreg.Reg[1][4] ), .S(fanout_net_27 ), .Z(_04257_ ) );
MUX2_X1 _12192_ ( .A(_04256_ ), .B(_04257_ ), .S(_03785_ ), .Z(_04258_ ) );
OAI211_X1 _12193_ ( .A(_03494_ ), .B(_04255_ ), .C1(_04258_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04259_ ) );
NOR2_X1 _12194_ ( .A1(_03896_ ), .A2(\myreg.Reg[11][4] ), .ZN(_04260_ ) );
OAI21_X1 _12195_ ( .A(fanout_net_32 ), .B1(fanout_net_28 ), .B2(\myreg.Reg[10][4] ), .ZN(_04261_ ) );
NOR2_X1 _12196_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[8][4] ), .ZN(_04262_ ) );
OAI21_X1 _12197_ ( .A(_03481_ ), .B1(_03560_ ), .B2(\myreg.Reg[9][4] ), .ZN(_04263_ ) );
OAI221_X1 _12198_ ( .A(_03782_ ), .B1(_04260_ ), .B2(_04261_ ), .C1(_04262_ ), .C2(_04263_ ), .ZN(_04264_ ) );
MUX2_X1 _12199_ ( .A(\myreg.Reg[12][4] ), .B(\myreg.Reg[13][4] ), .S(fanout_net_28 ), .Z(_04265_ ) );
MUX2_X1 _12200_ ( .A(\myreg.Reg[14][4] ), .B(\myreg.Reg[15][4] ), .S(fanout_net_28 ), .Z(_04266_ ) );
MUX2_X1 _12201_ ( .A(_04265_ ), .B(_04266_ ), .S(fanout_net_32 ), .Z(_04267_ ) );
OAI211_X1 _12202_ ( .A(fanout_net_34 ), .B(_04264_ ), .C1(_04267_ ), .C2(_03490_ ), .ZN(_04268_ ) );
OAI211_X2 _12203_ ( .A(_04259_ ), .B(_04268_ ), .C1(_03511_ ), .C2(_03497_ ), .ZN(_04269_ ) );
NAND2_X4 _12204_ ( .A1(_04250_ ), .A2(_04269_ ), .ZN(_04270_ ) );
INV_X1 _12205_ ( .A(_04270_ ), .ZN(_04271_ ) );
OAI211_X1 _12206_ ( .A(_04248_ ), .B(_04249_ ), .C1(_04271_ ), .C2(_01367_ ), .ZN(_04272_ ) );
NAND2_X1 _12207_ ( .A1(_04247_ ), .A2(_04272_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
NAND3_X1 _12208_ ( .A1(_04065_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_03599_ ), .ZN(_04273_ ) );
NAND3_X1 _12209_ ( .A1(_03765_ ), .A2(\mepc [3] ), .A3(_03463_ ), .ZN(_04274_ ) );
NAND4_X1 _12210_ ( .A1(_03768_ ), .A2(_03685_ ), .A3(\mycsreg.CSReg[0][3] ), .A4(_04072_ ), .ZN(_04275_ ) );
NAND4_X1 _12211_ ( .A1(_03690_ ), .A2(_03685_ ), .A3(\mtvec [3] ), .A4(_04072_ ), .ZN(_04276_ ) );
NAND4_X1 _12212_ ( .A1(_04273_ ), .A2(_04274_ ), .A3(_04275_ ), .A4(_04276_ ), .ZN(_04277_ ) );
AOI211_X1 _12213_ ( .A(_03441_ ), .B(_04277_ ), .C1(_04107_ ), .C2(_04106_ ), .ZN(_04278_ ) );
AND3_X1 _12214_ ( .A1(_04106_ ), .A2(_03240_ ), .A3(_04107_ ), .ZN(_04279_ ) );
NOR2_X1 _12215_ ( .A1(_04278_ ), .A2(_04279_ ), .ZN(_04280_ ) );
INV_X1 _12216_ ( .A(_04279_ ), .ZN(_04281_ ) );
OAI211_X1 _12217_ ( .A(_03474_ ), .B(_04281_ ), .C1(_04175_ ), .C2(_04277_ ), .ZN(_04282_ ) );
INV_X1 _12218_ ( .A(_04282_ ), .ZN(_04283_ ) );
AND2_X1 _12219_ ( .A1(fanout_net_6 ), .A2(\ID_EX_imm [3] ), .ZN(_04284_ ) );
OR2_X1 _12220_ ( .A1(_04283_ ), .A2(_04284_ ), .ZN(_04285_ ) );
AOI21_X1 _12221_ ( .A(\ID_EX_typ [0] ), .B1(_01500_ ), .B2(_01520_ ), .ZN(_04286_ ) );
OAI221_X1 _12222_ ( .A(_03379_ ), .B1(_02379_ ), .B2(_04280_ ), .C1(_04285_ ), .C2(_04286_ ), .ZN(_04287_ ) );
NAND4_X1 _12223_ ( .A1(_02344_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_04288_ ) );
OR3_X2 _12224_ ( .A1(_03873_ ), .A2(_03874_ ), .A3(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04289_ ) );
OR2_X1 _12225_ ( .A1(_04005_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04290_ ) );
OAI211_X1 _12226_ ( .A(_04290_ ), .B(fanout_net_32 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04291_ ) );
OR2_X1 _12227_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04292_ ) );
OAI211_X1 _12228_ ( .A(_04292_ ), .B(_03855_ ), .C1(_03896_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04293_ ) );
NAND3_X1 _12229_ ( .A1(_04291_ ), .A2(_03489_ ), .A3(_04293_ ), .ZN(_04294_ ) );
MUX2_X1 _12230_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04295_ ) );
MUX2_X1 _12231_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04296_ ) );
MUX2_X1 _12232_ ( .A(_04295_ ), .B(_04296_ ), .S(_03855_ ), .Z(_04297_ ) );
OAI211_X1 _12233_ ( .A(_03493_ ), .B(_04294_ ), .C1(_04297_ ), .C2(_03782_ ), .ZN(_04298_ ) );
OR2_X1 _12234_ ( .A1(_04005_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04299_ ) );
OAI211_X1 _12235_ ( .A(_04299_ ), .B(_03481_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04300_ ) );
OR2_X1 _12236_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04301_ ) );
OAI211_X1 _12237_ ( .A(_04301_ ), .B(fanout_net_32 ), .C1(_03896_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04302_ ) );
NAND3_X1 _12238_ ( .A1(_04300_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04302_ ), .ZN(_04303_ ) );
MUX2_X1 _12239_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04304_ ) );
MUX2_X1 _12240_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04305_ ) );
MUX2_X1 _12241_ ( .A(_04304_ ), .B(_04305_ ), .S(fanout_net_32 ), .Z(_04306_ ) );
OAI211_X1 _12242_ ( .A(fanout_net_34 ), .B(_04303_ ), .C1(_04306_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04307_ ) );
OAI211_X1 _12243_ ( .A(_04298_ ), .B(_04307_ ), .C1(_03873_ ), .C2(_03874_ ), .ZN(_04308_ ) );
NAND2_X1 _12244_ ( .A1(_04289_ ), .A2(_04308_ ), .ZN(_04309_ ) );
OAI211_X1 _12245_ ( .A(_04248_ ), .B(_04288_ ), .C1(_04309_ ), .C2(_01367_ ), .ZN(_04310_ ) );
NAND2_X1 _12246_ ( .A1(_04287_ ), .A2(_04310_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
NAND4_X1 _12247_ ( .A1(_02345_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_04311_ ) );
OR3_X1 _12248_ ( .A1(_03509_ ), .A2(_01377_ ), .A3(\EX_LS_result_reg [2] ), .ZN(_04312_ ) );
OR2_X1 _12249_ ( .A1(_03558_ ), .A2(\myreg.Reg[1][2] ), .ZN(_04313_ ) );
OAI211_X1 _12250_ ( .A(_04313_ ), .B(_03480_ ), .C1(fanout_net_28 ), .C2(\myreg.Reg[0][2] ), .ZN(_04314_ ) );
OR2_X1 _12251_ ( .A1(_03557_ ), .A2(\myreg.Reg[3][2] ), .ZN(_04315_ ) );
OAI211_X1 _12252_ ( .A(_04315_ ), .B(fanout_net_32 ), .C1(fanout_net_28 ), .C2(\myreg.Reg[2][2] ), .ZN(_04316_ ) );
NAND3_X1 _12253_ ( .A1(_04314_ ), .A2(_04316_ ), .A3(_03488_ ), .ZN(_04317_ ) );
MUX2_X1 _12254_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_28 ), .Z(_04318_ ) );
MUX2_X1 _12255_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_28 ), .Z(_04319_ ) );
MUX2_X1 _12256_ ( .A(_04318_ ), .B(_04319_ ), .S(_03480_ ), .Z(_04320_ ) );
OAI211_X1 _12257_ ( .A(_03492_ ), .B(_04317_ ), .C1(_04320_ ), .C2(_03488_ ), .ZN(_04321_ ) );
OR2_X1 _12258_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[14][2] ), .ZN(_04322_ ) );
OAI211_X1 _12259_ ( .A(_04322_ ), .B(fanout_net_32 ), .C1(_04005_ ), .C2(\myreg.Reg[15][2] ), .ZN(_04323_ ) );
OR2_X1 _12260_ ( .A1(fanout_net_28 ), .A2(\myreg.Reg[12][2] ), .ZN(_04324_ ) );
OAI211_X1 _12261_ ( .A(_04324_ ), .B(_03480_ ), .C1(_04005_ ), .C2(\myreg.Reg[13][2] ), .ZN(_04325_ ) );
NAND3_X1 _12262_ ( .A1(_04323_ ), .A2(_04325_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04326_ ) );
MUX2_X1 _12263_ ( .A(\myreg.Reg[8][2] ), .B(\myreg.Reg[9][2] ), .S(fanout_net_28 ), .Z(_04327_ ) );
MUX2_X1 _12264_ ( .A(\myreg.Reg[10][2] ), .B(\myreg.Reg[11][2] ), .S(fanout_net_28 ), .Z(_04328_ ) );
MUX2_X1 _12265_ ( .A(_04327_ ), .B(_04328_ ), .S(fanout_net_32 ), .Z(_04329_ ) );
OAI211_X1 _12266_ ( .A(fanout_net_34 ), .B(_04326_ ), .C1(_04329_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04330_ ) );
OAI211_X4 _12267_ ( .A(_04321_ ), .B(_04330_ ), .C1(_03510_ ), .C2(_03496_ ), .ZN(_04331_ ) );
NAND2_X2 _12268_ ( .A1(_04312_ ), .A2(_04331_ ), .ZN(_04332_ ) );
INV_X1 _12269_ ( .A(_04332_ ), .ZN(_04333_ ) );
OAI211_X1 _12270_ ( .A(_03364_ ), .B(_04311_ ), .C1(_04333_ ), .C2(_01367_ ), .ZN(_04334_ ) );
AND3_X1 _12271_ ( .A1(_03592_ ), .A2(\mepc [2] ), .A3(_03462_ ), .ZN(_04335_ ) );
OR2_X1 _12272_ ( .A1(_03527_ ), .A2(_04335_ ), .ZN(_04336_ ) );
NAND3_X1 _12273_ ( .A1(_03765_ ), .A2(\mycsreg.CSReg[3][2] ), .A3(_03599_ ), .ZN(_04337_ ) );
NAND4_X1 _12274_ ( .A1(_03768_ ), .A2(_03685_ ), .A3(\mycsreg.CSReg[0][2] ), .A4(_03691_ ), .ZN(_04338_ ) );
NAND4_X1 _12275_ ( .A1(_03690_ ), .A2(_03685_ ), .A3(\mtvec [2] ), .A4(_03691_ ), .ZN(_04339_ ) );
NAND3_X1 _12276_ ( .A1(_04337_ ), .A2(_04338_ ), .A3(_04339_ ), .ZN(_04340_ ) );
OAI21_X1 _12277_ ( .A(_03646_ ), .B1(_04336_ ), .B2(_04340_ ), .ZN(_04341_ ) );
NAND4_X1 _12278_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_03096_ ), .A4(_03606_ ), .ZN(_04342_ ) );
AND2_X1 _12279_ ( .A1(_04341_ ), .A2(_04342_ ), .ZN(_04343_ ) );
OAI22_X1 _12280_ ( .A1(_04343_ ), .A2(_03548_ ), .B1(_01351_ ), .B2(_01548_ ), .ZN(_04344_ ) );
AOI21_X1 _12281_ ( .A(_04344_ ), .B1(_02381_ ), .B2(_01547_ ), .ZN(_04345_ ) );
INV_X1 _12282_ ( .A(_04343_ ), .ZN(_04346_ ) );
OAI21_X1 _12283_ ( .A(_03698_ ), .B1(_04346_ ), .B2(_02379_ ), .ZN(_04347_ ) );
OAI21_X1 _12284_ ( .A(_04334_ ), .B1(_04345_ ), .B2(_04347_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
INV_X1 _12285_ ( .A(_02214_ ), .ZN(_04348_ ) );
OR3_X1 _12286_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [29] ), .A3(_03432_ ), .ZN(_04349_ ) );
BUF_X4 _12287_ ( .A(_03449_ ), .Z(_04350_ ) );
NAND3_X1 _12288_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_04069_ ), .ZN(_04351_ ) );
NAND4_X1 _12289_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [29] ), .A4(_04071_ ), .ZN(_04352_ ) );
NAND3_X1 _12290_ ( .A1(_03443_ ), .A2(_04351_ ), .A3(_04352_ ), .ZN(_04353_ ) );
NAND3_X1 _12291_ ( .A1(_04065_ ), .A2(\mepc [29] ), .A3(_04066_ ), .ZN(_04354_ ) );
NAND3_X1 _12292_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_04071_ ), .ZN(_04355_ ) );
OAI211_X1 _12293_ ( .A(_04354_ ), .B(_04355_ ), .C1(_04197_ ), .C2(_04198_ ), .ZN(_04356_ ) );
OAI21_X1 _12294_ ( .A(_04349_ ), .B1(_04353_ ), .B2(_04356_ ), .ZN(_04357_ ) );
AOI22_X1 _12295_ ( .A1(_04348_ ), .A2(_01351_ ), .B1(fanout_net_7 ), .B2(_04357_ ), .ZN(_04358_ ) );
OAI211_X1 _12296_ ( .A(_04358_ ), .B(_03551_ ), .C1(_02381_ ), .C2(\ID_EX_imm [29] ), .ZN(_04359_ ) );
OR3_X1 _12297_ ( .A1(_04357_ ), .A2(_03700_ ), .A3(_03548_ ), .ZN(_04360_ ) );
AND3_X1 _12298_ ( .A1(_01366_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_typ [7] ), .ZN(_04361_ ) );
OR3_X1 _12299_ ( .A1(_03512_ ), .A2(_03498_ ), .A3(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04362_ ) );
OR2_X1 _12300_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04363_ ) );
OAI211_X1 _12301_ ( .A(_04363_ ), .B(_03573_ ), .C1(_03741_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04364_ ) );
NAND2_X1 _12302_ ( .A1(_02196_ ), .A2(fanout_net_28 ), .ZN(_04365_ ) );
OAI211_X1 _12303_ ( .A(_04365_ ), .B(fanout_net_32 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04366_ ) );
NAND3_X1 _12304_ ( .A1(_04364_ ), .A2(_04366_ ), .A3(_03519_ ), .ZN(_04367_ ) );
MUX2_X1 _12305_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04368_ ) );
MUX2_X1 _12306_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04369_ ) );
MUX2_X1 _12307_ ( .A(_04368_ ), .B(_04369_ ), .S(_03616_ ), .Z(_04370_ ) );
OAI211_X1 _12308_ ( .A(_03494_ ), .B(_04367_ ), .C1(_04370_ ), .C2(_03665_ ), .ZN(_04371_ ) );
OR2_X1 _12309_ ( .A1(_03561_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04372_ ) );
OAI211_X1 _12310_ ( .A(_04372_ ), .B(_03573_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04373_ ) );
OR2_X1 _12311_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04374_ ) );
OAI211_X1 _12312_ ( .A(_04374_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03617_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04375_ ) );
NAND3_X1 _12313_ ( .A1(_04373_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04375_ ), .ZN(_04376_ ) );
MUX2_X1 _12314_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04377_ ) );
MUX2_X1 _12315_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_04378_ ) );
MUX2_X1 _12316_ ( .A(_04377_ ), .B(_04378_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04379_ ) );
OAI211_X1 _12317_ ( .A(fanout_net_34 ), .B(_04376_ ), .C1(_04379_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04380_ ) );
OAI211_X1 _12318_ ( .A(_04371_ ), .B(_04380_ ), .C1(_03553_ ), .C2(_03554_ ), .ZN(_04381_ ) );
NAND2_X1 _12319_ ( .A1(_04362_ ), .A2(_04381_ ), .ZN(_04382_ ) );
AOI21_X1 _12320_ ( .A(_04361_ ), .B1(_04382_ ), .B2(_03362_ ), .ZN(_04383_ ) );
OAI211_X1 _12321_ ( .A(_04359_ ), .B(_04360_ ), .C1(_03552_ ), .C2(_04383_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
INV_X16 _12322_ ( .A(_01571_ ), .ZN(_04384_ ) );
OR3_X1 _12323_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_03432_ ), .ZN(_04385_ ) );
NAND4_X1 _12324_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [1] ), .A4(_04071_ ), .ZN(_04386_ ) );
NAND3_X1 _12325_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_04069_ ), .ZN(_04387_ ) );
NAND3_X1 _12326_ ( .A1(_04065_ ), .A2(\mepc [1] ), .A3(_04066_ ), .ZN(_04388_ ) );
NAND3_X1 _12327_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_04120_ ), .ZN(_04389_ ) );
NAND4_X1 _12328_ ( .A1(_04386_ ), .A2(_04387_ ), .A3(_04388_ ), .A4(_04389_ ), .ZN(_04390_ ) );
OAI21_X1 _12329_ ( .A(_04385_ ), .B1(_03939_ ), .B2(_04390_ ), .ZN(_04391_ ) );
AOI22_X1 _12330_ ( .A1(_04384_ ), .A2(_01351_ ), .B1(fanout_net_7 ), .B2(_04391_ ), .ZN(_04392_ ) );
OAI211_X1 _12331_ ( .A(_04392_ ), .B(_03551_ ), .C1(_02381_ ), .C2(\ID_EX_imm [1] ), .ZN(_04393_ ) );
INV_X1 _12332_ ( .A(_03939_ ), .ZN(_04394_ ) );
AND2_X1 _12333_ ( .A1(_04387_ ), .A2(_04388_ ), .ZN(_04395_ ) );
AND2_X1 _12334_ ( .A1(_04386_ ), .A2(_04389_ ), .ZN(_04396_ ) );
NAND3_X1 _12335_ ( .A1(_04394_ ), .A2(_04395_ ), .A3(_04396_ ), .ZN(_04397_ ) );
NAND4_X1 _12336_ ( .A1(_04397_ ), .A2(_04385_ ), .A3(_03378_ ), .A4(_03702_ ), .ZN(_04398_ ) );
OR3_X4 _12337_ ( .A1(_03509_ ), .A2(_01377_ ), .A3(\EX_LS_result_reg [1] ), .ZN(_04399_ ) );
OR2_X1 _12338_ ( .A1(_03557_ ), .A2(\myreg.Reg[1][1] ), .ZN(_04400_ ) );
OAI211_X1 _12339_ ( .A(_04400_ ), .B(_03480_ ), .C1(fanout_net_28 ), .C2(\myreg.Reg[0][1] ), .ZN(_04401_ ) );
OR2_X1 _12340_ ( .A1(_03557_ ), .A2(\myreg.Reg[3][1] ), .ZN(_04402_ ) );
OAI211_X1 _12341_ ( .A(_04402_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_29 ), .C2(\myreg.Reg[2][1] ), .ZN(_04403_ ) );
NAND3_X1 _12342_ ( .A1(_04401_ ), .A2(_04403_ ), .A3(_03488_ ), .ZN(_04404_ ) );
MUX2_X1 _12343_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(fanout_net_29 ), .Z(_04405_ ) );
MUX2_X1 _12344_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(fanout_net_29 ), .Z(_04406_ ) );
MUX2_X1 _12345_ ( .A(_04405_ ), .B(_04406_ ), .S(_03479_ ), .Z(_04407_ ) );
OAI211_X1 _12346_ ( .A(_03492_ ), .B(_04404_ ), .C1(_04407_ ), .C2(_03488_ ), .ZN(_04408_ ) );
OR2_X1 _12347_ ( .A1(_03557_ ), .A2(\myreg.Reg[15][1] ), .ZN(_04409_ ) );
OAI211_X1 _12348_ ( .A(_04409_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_29 ), .C2(\myreg.Reg[14][1] ), .ZN(_04410_ ) );
OR2_X1 _12349_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[12][1] ), .ZN(_04411_ ) );
OAI211_X1 _12350_ ( .A(_04411_ ), .B(_03480_ ), .C1(_03558_ ), .C2(\myreg.Reg[13][1] ), .ZN(_04412_ ) );
NAND3_X1 _12351_ ( .A1(_04410_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04412_ ), .ZN(_04413_ ) );
MUX2_X1 _12352_ ( .A(\myreg.Reg[8][1] ), .B(\myreg.Reg[9][1] ), .S(fanout_net_29 ), .Z(_04414_ ) );
MUX2_X1 _12353_ ( .A(\myreg.Reg[10][1] ), .B(\myreg.Reg[11][1] ), .S(fanout_net_29 ), .Z(_04415_ ) );
MUX2_X1 _12354_ ( .A(_04414_ ), .B(_04415_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04416_ ) );
OAI211_X1 _12355_ ( .A(fanout_net_34 ), .B(_04413_ ), .C1(_04416_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04417_ ) );
OAI211_X4 _12356_ ( .A(_04408_ ), .B(_04417_ ), .C1(_03509_ ), .C2(_01377_ ), .ZN(_04418_ ) );
NAND2_X4 _12357_ ( .A1(_04399_ ), .A2(_04418_ ), .ZN(_04419_ ) );
MUX2_X1 _12358_ ( .A(_02347_ ), .B(_04419_ ), .S(_03370_ ), .Z(_04420_ ) );
OAI211_X1 _12359_ ( .A(_04393_ ), .B(_04398_ ), .C1(_03552_ ), .C2(_04420_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
AND3_X1 _12360_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_04200_ ), .ZN(_04421_ ) );
NAND3_X1 _12361_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][0] ), .A3(_04069_ ), .ZN(_04422_ ) );
NAND3_X1 _12362_ ( .A1(_03688_ ), .A2(\mepc [0] ), .A3(_04120_ ), .ZN(_04423_ ) );
NAND4_X1 _12363_ ( .A1(_03690_ ), .A2(_04120_ ), .A3(\mtvec [0] ), .A4(_04072_ ), .ZN(_04424_ ) );
NAND4_X1 _12364_ ( .A1(_03878_ ), .A2(_04422_ ), .A3(_04423_ ), .A4(_04424_ ), .ZN(_04425_ ) );
OAI21_X1 _12365_ ( .A(_03646_ ), .B1(_04421_ ), .B2(_04425_ ), .ZN(_04426_ ) );
NAND4_X1 _12366_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_04077_ ), .A4(_03606_ ), .ZN(_04427_ ) );
AOI21_X1 _12367_ ( .A(_03700_ ), .B1(_04426_ ), .B2(_04427_ ), .ZN(_04428_ ) );
NAND2_X1 _12368_ ( .A1(_04428_ ), .A2(_03702_ ), .ZN(_04429_ ) );
NAND3_X1 _12369_ ( .A1(_01576_ ), .A2(_01595_ ), .A3(_02381_ ), .ZN(_04430_ ) );
NAND3_X1 _12370_ ( .A1(_04426_ ), .A2(fanout_net_7 ), .A3(_04427_ ), .ZN(_04431_ ) );
NAND2_X1 _12371_ ( .A1(_01575_ ), .A2(\ID_EX_typ [0] ), .ZN(_04432_ ) );
NAND4_X1 _12372_ ( .A1(_04430_ ), .A2(_04431_ ), .A3(_03378_ ), .A4(_04432_ ), .ZN(_04433_ ) );
OR3_X2 _12373_ ( .A1(_03509_ ), .A2(_01377_ ), .A3(\EX_LS_result_reg [0] ), .ZN(_04434_ ) );
OR2_X1 _12374_ ( .A1(_03557_ ), .A2(\myreg.Reg[3][0] ), .ZN(_04435_ ) );
OAI211_X1 _12375_ ( .A(_04435_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_29 ), .C2(\myreg.Reg[2][0] ), .ZN(_04436_ ) );
OR2_X1 _12376_ ( .A1(fanout_net_29 ), .A2(\myreg.Reg[0][0] ), .ZN(_04437_ ) );
OAI211_X1 _12377_ ( .A(_04437_ ), .B(_03479_ ), .C1(_03557_ ), .C2(\myreg.Reg[1][0] ), .ZN(_04438_ ) );
NAND3_X1 _12378_ ( .A1(_04436_ ), .A2(_03487_ ), .A3(_04438_ ), .ZN(_04439_ ) );
MUX2_X1 _12379_ ( .A(\myreg.Reg[6][0] ), .B(\myreg.Reg[7][0] ), .S(fanout_net_29 ), .Z(_04440_ ) );
MUX2_X1 _12380_ ( .A(\myreg.Reg[4][0] ), .B(\myreg.Reg[5][0] ), .S(fanout_net_29 ), .Z(_04441_ ) );
MUX2_X1 _12381_ ( .A(_04440_ ), .B(_04441_ ), .S(_03479_ ), .Z(_04442_ ) );
OAI211_X1 _12382_ ( .A(_03492_ ), .B(_04439_ ), .C1(_04442_ ), .C2(_03487_ ), .ZN(_04443_ ) );
OR2_X1 _12383_ ( .A1(_03557_ ), .A2(\myreg.Reg[15][0] ), .ZN(_04444_ ) );
OAI211_X1 _12384_ ( .A(_04444_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_29 ), .C2(\myreg.Reg[14][0] ), .ZN(_04445_ ) );
OR2_X1 _12385_ ( .A1(_03557_ ), .A2(\myreg.Reg[13][0] ), .ZN(_04446_ ) );
OAI211_X1 _12386_ ( .A(_04446_ ), .B(_03479_ ), .C1(fanout_net_29 ), .C2(\myreg.Reg[12][0] ), .ZN(_04447_ ) );
NAND3_X1 _12387_ ( .A1(_04445_ ), .A2(_04447_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04448_ ) );
MUX2_X1 _12388_ ( .A(\myreg.Reg[8][0] ), .B(\myreg.Reg[9][0] ), .S(fanout_net_29 ), .Z(_04449_ ) );
MUX2_X1 _12389_ ( .A(\myreg.Reg[10][0] ), .B(\myreg.Reg[11][0] ), .S(fanout_net_29 ), .Z(_04450_ ) );
MUX2_X1 _12390_ ( .A(_04449_ ), .B(_04450_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04451_ ) );
OAI211_X1 _12391_ ( .A(fanout_net_34 ), .B(_04448_ ), .C1(_04451_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04452_ ) );
OAI211_X1 _12392_ ( .A(_04443_ ), .B(_04452_ ), .C1(_03509_ ), .C2(_01377_ ), .ZN(_04453_ ) );
NAND2_X4 _12393_ ( .A1(_04434_ ), .A2(_04453_ ), .ZN(_04454_ ) );
MUX2_X1 _12394_ ( .A(_02348_ ), .B(_04454_ ), .S(_03590_ ), .Z(_04455_ ) );
OAI211_X1 _12395_ ( .A(_04429_ ), .B(_04433_ ), .C1(_04455_ ), .C2(_03762_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
OR3_X1 _12396_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_03432_ ), .ZN(_04456_ ) );
NAND3_X1 _12397_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_04069_ ), .ZN(_04457_ ) );
NAND4_X1 _12398_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [28] ), .A4(_04071_ ), .ZN(_04458_ ) );
NAND3_X1 _12399_ ( .A1(_03443_ ), .A2(_04457_ ), .A3(_04458_ ), .ZN(_04459_ ) );
NAND3_X1 _12400_ ( .A1(_04065_ ), .A2(\mepc [28] ), .A3(_04066_ ), .ZN(_04460_ ) );
NAND3_X1 _12401_ ( .A1(_03467_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_04071_ ), .ZN(_04461_ ) );
OAI211_X1 _12402_ ( .A(_04460_ ), .B(_04461_ ), .C1(_04197_ ), .C2(_04198_ ), .ZN(_04462_ ) );
OAI21_X1 _12403_ ( .A(_04456_ ), .B1(_04459_ ), .B2(_04462_ ), .ZN(_04463_ ) );
AOI22_X1 _12404_ ( .A1(_02308_ ), .A2(_01351_ ), .B1(fanout_net_7 ), .B2(_04463_ ), .ZN(_04464_ ) );
OAI211_X1 _12405_ ( .A(_04464_ ), .B(_03551_ ), .C1(_02381_ ), .C2(\ID_EX_imm [28] ), .ZN(_04465_ ) );
OR3_X1 _12406_ ( .A1(_04463_ ), .A2(_03700_ ), .A3(_03548_ ), .ZN(_04466_ ) );
AND3_X1 _12407_ ( .A1(_01366_ ), .A2(\ID_EX_pc [28] ), .A3(\ID_EX_typ [7] ), .ZN(_04467_ ) );
OR3_X1 _12408_ ( .A1(_03512_ ), .A2(_03498_ ), .A3(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .ZN(_04468_ ) );
OR2_X1 _12409_ ( .A1(_03561_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04469_ ) );
OAI211_X1 _12410_ ( .A(_04469_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_29 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04470_ ) );
OR2_X1 _12411_ ( .A1(fanout_net_29 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04471_ ) );
OAI211_X1 _12412_ ( .A(_04471_ ), .B(_03616_ ), .C1(_03617_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04472_ ) );
NAND3_X1 _12413_ ( .A1(_04470_ ), .A2(_03519_ ), .A3(_04472_ ), .ZN(_04473_ ) );
MUX2_X1 _12414_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04474_ ) );
MUX2_X1 _12415_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04475_ ) );
MUX2_X1 _12416_ ( .A(_04474_ ), .B(_04475_ ), .S(_03624_ ), .Z(_04476_ ) );
OAI211_X1 _12417_ ( .A(fanout_net_34 ), .B(_04473_ ), .C1(_04476_ ), .C2(_03665_ ), .ZN(_04477_ ) );
OR2_X1 _12418_ ( .A1(fanout_net_29 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04478_ ) );
OAI211_X1 _12419_ ( .A(_04478_ ), .B(_03624_ ), .C1(_03627_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04479_ ) );
NOR2_X1 _12420_ ( .A1(_03617_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04480_ ) );
OAI21_X1 _12421_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_29 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04481_ ) );
OAI211_X1 _12422_ ( .A(_04479_ ), .B(_03519_ ), .C1(_04480_ ), .C2(_04481_ ), .ZN(_04482_ ) );
MUX2_X1 _12423_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04483_ ) );
MUX2_X1 _12424_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04484_ ) );
MUX2_X1 _12425_ ( .A(_04483_ ), .B(_04484_ ), .S(_03624_ ), .Z(_04485_ ) );
OAI211_X1 _12426_ ( .A(_03494_ ), .B(_04482_ ), .C1(_04485_ ), .C2(_03665_ ), .ZN(_04486_ ) );
OAI211_X1 _12427_ ( .A(_04477_ ), .B(_04486_ ), .C1(_03553_ ), .C2(_03554_ ), .ZN(_04487_ ) );
NAND2_X1 _12428_ ( .A1(_04468_ ), .A2(_04487_ ), .ZN(_04488_ ) );
AOI21_X1 _12429_ ( .A(_04467_ ), .B1(_04488_ ), .B2(_03362_ ), .ZN(_04489_ ) );
OAI211_X1 _12430_ ( .A(_04465_ ), .B(_04466_ ), .C1(_03552_ ), .C2(_04489_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
INV_X1 _12431_ ( .A(_01472_ ), .ZN(_04490_ ) );
OR3_X1 _12432_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_03432_ ), .ZN(_04491_ ) );
NAND3_X1 _12433_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_04069_ ), .ZN(_04492_ ) );
NAND4_X1 _12434_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [27] ), .A4(_04071_ ), .ZN(_04493_ ) );
NAND3_X1 _12435_ ( .A1(_03443_ ), .A2(_04492_ ), .A3(_04493_ ), .ZN(_04494_ ) );
NAND3_X1 _12436_ ( .A1(_04065_ ), .A2(\mepc [27] ), .A3(_04066_ ), .ZN(_04495_ ) );
NAND3_X1 _12437_ ( .A1(_03467_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_04071_ ), .ZN(_04496_ ) );
OAI211_X1 _12438_ ( .A(_04495_ ), .B(_04496_ ), .C1(_04197_ ), .C2(_04198_ ), .ZN(_04497_ ) );
OAI21_X1 _12439_ ( .A(_04491_ ), .B1(_04494_ ), .B2(_04497_ ), .ZN(_04498_ ) );
AOI22_X1 _12440_ ( .A1(_04490_ ), .A2(_01351_ ), .B1(fanout_net_7 ), .B2(_04498_ ), .ZN(_04499_ ) );
OAI211_X1 _12441_ ( .A(_04499_ ), .B(_03551_ ), .C1(_02381_ ), .C2(\ID_EX_imm [27] ), .ZN(_04500_ ) );
OR3_X1 _12442_ ( .A1(_04498_ ), .A2(_03700_ ), .A3(_03548_ ), .ZN(_04501_ ) );
AND3_X1 _12443_ ( .A1(_01366_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_04502_ ) );
INV_X1 _12444_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04503_ ) );
OR3_X1 _12445_ ( .A1(_03553_ ), .A2(_03554_ ), .A3(_04503_ ), .ZN(_04504_ ) );
OR2_X1 _12446_ ( .A1(fanout_net_29 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04505_ ) );
OAI211_X1 _12447_ ( .A(_04505_ ), .B(_03663_ ), .C1(_03568_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04506_ ) );
OR2_X1 _12448_ ( .A1(fanout_net_29 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04507_ ) );
OAI211_X1 _12449_ ( .A(_04507_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03568_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04508_ ) );
NAND3_X1 _12450_ ( .A1(_04506_ ), .A2(_04508_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04509_ ) );
MUX2_X1 _12451_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04510_ ) );
MUX2_X1 _12452_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04511_ ) );
MUX2_X1 _12453_ ( .A(_04510_ ), .B(_04511_ ), .S(_03567_ ), .Z(_04512_ ) );
OAI211_X1 _12454_ ( .A(_03556_ ), .B(_04509_ ), .C1(_04512_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04513_ ) );
NOR2_X1 _12455_ ( .A1(_03741_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04514_ ) );
OAI21_X1 _12456_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_29 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04515_ ) );
NOR2_X1 _12457_ ( .A1(fanout_net_29 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04516_ ) );
OAI21_X1 _12458_ ( .A(_03567_ ), .B1(_03741_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04517_ ) );
OAI221_X1 _12459_ ( .A(_03565_ ), .B1(_04514_ ), .B2(_04515_ ), .C1(_04516_ ), .C2(_04517_ ), .ZN(_04518_ ) );
MUX2_X1 _12460_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_29 ), .Z(_04519_ ) );
MUX2_X1 _12461_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04520_ ) );
MUX2_X1 _12462_ ( .A(_04519_ ), .B(_04520_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04521_ ) );
OAI211_X1 _12463_ ( .A(fanout_net_34 ), .B(_04518_ ), .C1(_04521_ ), .C2(_03575_ ), .ZN(_04522_ ) );
OAI211_X1 _12464_ ( .A(_04513_ ), .B(_04522_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_04523_ ) );
NAND2_X1 _12465_ ( .A1(_04504_ ), .A2(_04523_ ), .ZN(_04524_ ) );
AOI21_X1 _12466_ ( .A(_04502_ ), .B1(_04524_ ), .B2(_03362_ ), .ZN(_04525_ ) );
OAI211_X1 _12467_ ( .A(_04500_ ), .B(_04501_ ), .C1(_03762_ ), .C2(_04525_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
OR3_X1 _12468_ ( .A1(_04197_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_04198_ ), .ZN(_04526_ ) );
NAND4_X1 _12469_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [26] ), .A4(_04120_ ), .ZN(_04527_ ) );
NAND3_X1 _12470_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_04069_ ), .ZN(_04528_ ) );
NAND3_X1 _12471_ ( .A1(_04350_ ), .A2(\mepc [26] ), .A3(_04066_ ), .ZN(_04529_ ) );
NAND3_X1 _12472_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_04120_ ), .ZN(_04530_ ) );
NAND4_X1 _12473_ ( .A1(_04527_ ), .A2(_04528_ ), .A3(_04529_ ), .A4(_04530_ ), .ZN(_04531_ ) );
OAI21_X1 _12474_ ( .A(_04526_ ), .B1(_03939_ ), .B2(_04531_ ), .ZN(_04532_ ) );
AOI22_X1 _12475_ ( .A1(_04532_ ), .A2(fanout_net_7 ), .B1(\ID_EX_typ [0] ), .B2(_02183_ ), .ZN(_04533_ ) );
OAI211_X1 _12476_ ( .A(_03698_ ), .B(_04533_ ), .C1(_02182_ ), .C2(\ID_EX_typ [0] ), .ZN(_04534_ ) );
OR3_X1 _12477_ ( .A1(_04532_ ), .A2(_03356_ ), .A3(_03548_ ), .ZN(_04535_ ) );
AND3_X1 _12478_ ( .A1(_01366_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_04536_ ) );
OR2_X1 _12479_ ( .A1(_03627_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04537_ ) );
OAI211_X1 _12480_ ( .A(_04537_ ), .B(_03663_ ), .C1(fanout_net_30 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04538_ ) );
NAND2_X1 _12481_ ( .A1(_02164_ ), .A2(fanout_net_30 ), .ZN(_04539_ ) );
OAI211_X1 _12482_ ( .A(_04539_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_30 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04540_ ) );
NAND3_X1 _12483_ ( .A1(_04538_ ), .A2(_03665_ ), .A3(_04540_ ), .ZN(_04541_ ) );
MUX2_X1 _12484_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04542_ ) );
MUX2_X1 _12485_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04543_ ) );
MUX2_X1 _12486_ ( .A(_04542_ ), .B(_04543_ ), .S(_03663_ ), .Z(_04544_ ) );
OAI211_X1 _12487_ ( .A(fanout_net_34 ), .B(_04541_ ), .C1(_04544_ ), .C2(_03575_ ), .ZN(_04545_ ) );
MUX2_X1 _12488_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04546_ ) );
AND2_X1 _12489_ ( .A1(_04546_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_04547_ ) );
MUX2_X1 _12490_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04548_ ) );
AOI211_X1 _12491_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_04547_ ), .C1(_03663_ ), .C2(_04548_ ), .ZN(_04549_ ) );
MUX2_X1 _12492_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04550_ ) );
MUX2_X1 _12493_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04551_ ) );
MUX2_X1 _12494_ ( .A(_04550_ ), .B(_04551_ ), .S(_03616_ ), .Z(_04552_ ) );
OAI21_X1 _12495_ ( .A(_03556_ ), .B1(_04552_ ), .B2(_03665_ ), .ZN(_04553_ ) );
OAI221_X1 _12496_ ( .A(_04545_ ), .B1(_04549_ ), .B2(_04553_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_04554_ ) );
NOR2_X1 _12497_ ( .A1(_03511_ ), .A2(_03497_ ), .ZN(_04555_ ) );
NAND2_X1 _12498_ ( .A1(_04555_ ), .A2(\EX_LS_result_reg [26] ), .ZN(_04556_ ) );
NAND2_X1 _12499_ ( .A1(_04554_ ), .A2(_04556_ ), .ZN(_04557_ ) );
AOI21_X1 _12500_ ( .A(_04536_ ), .B1(_04557_ ), .B2(_03362_ ), .ZN(_04558_ ) );
OAI211_X1 _12501_ ( .A(_04534_ ), .B(_04535_ ), .C1(_04558_ ), .C2(_03762_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND3_X1 _12502_ ( .A1(_03592_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_03452_ ), .ZN(_04559_ ) );
NAND4_X1 _12503_ ( .A1(_03652_ ), .A2(_03842_ ), .A3(\mtvec [25] ), .A4(_03595_ ), .ZN(_04560_ ) );
AND2_X1 _12504_ ( .A1(_04559_ ), .A2(_04560_ ), .ZN(_04561_ ) );
NAND3_X1 _12505_ ( .A1(_03592_ ), .A2(\mepc [25] ), .A3(_03462_ ), .ZN(_04562_ ) );
NAND4_X1 _12506_ ( .A1(_03594_ ), .A2(_03842_ ), .A3(\mycsreg.CSReg[0][25] ), .A4(_03595_ ), .ZN(_04563_ ) );
AND2_X1 _12507_ ( .A1(_04562_ ), .A2(_04563_ ), .ZN(_04564_ ) );
AOI22_X1 _12508_ ( .A1(_04107_ ), .A2(_04106_ ), .B1(_04561_ ), .B2(_04564_ ), .ZN(_04565_ ) );
AND3_X1 _12509_ ( .A1(_04106_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_04107_ ), .ZN(_04566_ ) );
NOR2_X1 _12510_ ( .A1(_04565_ ), .A2(_04566_ ), .ZN(_04567_ ) );
NOR2_X1 _12511_ ( .A1(_04567_ ), .A2(_03547_ ), .ZN(_04568_ ) );
NAND3_X1 _12512_ ( .A1(_02138_ ), .A2(_01351_ ), .A3(_02157_ ), .ZN(_04569_ ) );
AOI22_X1 _12513_ ( .A1(_04567_ ), .A2(fanout_net_7 ), .B1(\ID_EX_typ [0] ), .B2(_02185_ ), .ZN(_04570_ ) );
AOI211_X1 _12514_ ( .A(_03357_ ), .B(_04568_ ), .C1(_04569_ ), .C2(_04570_ ), .ZN(_04571_ ) );
INV_X1 _12515_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04572_ ) );
OR3_X4 _12516_ ( .A1(_03512_ ), .A2(_03498_ ), .A3(_04572_ ), .ZN(_04573_ ) );
OR2_X1 _12517_ ( .A1(_03561_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04574_ ) );
OAI211_X1 _12518_ ( .A(_04574_ ), .B(_03616_ ), .C1(fanout_net_30 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04575_ ) );
OR2_X1 _12519_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04576_ ) );
OAI211_X1 _12520_ ( .A(_04576_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03617_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04577_ ) );
NAND3_X1 _12521_ ( .A1(_04575_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04577_ ), .ZN(_04578_ ) );
MUX2_X1 _12522_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04579_ ) );
MUX2_X1 _12523_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04580_ ) );
MUX2_X1 _12524_ ( .A(_04579_ ), .B(_04580_ ), .S(_03624_ ), .Z(_04581_ ) );
OAI211_X1 _12525_ ( .A(_03494_ ), .B(_04578_ ), .C1(_04581_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04582_ ) );
NOR2_X1 _12526_ ( .A1(_03627_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04583_ ) );
OAI21_X1 _12527_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_30 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04584_ ) );
NOR2_X1 _12528_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04585_ ) );
OAI21_X1 _12529_ ( .A(_03624_ ), .B1(_03617_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04586_ ) );
OAI221_X1 _12530_ ( .A(_03519_ ), .B1(_04583_ ), .B2(_04584_ ), .C1(_04585_ ), .C2(_04586_ ), .ZN(_04587_ ) );
MUX2_X1 _12531_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04588_ ) );
MUX2_X1 _12532_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04589_ ) );
MUX2_X1 _12533_ ( .A(_04588_ ), .B(_04589_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04590_ ) );
OAI211_X1 _12534_ ( .A(fanout_net_34 ), .B(_04587_ ), .C1(_04590_ ), .C2(_03665_ ), .ZN(_04591_ ) );
OAI211_X1 _12535_ ( .A(_04582_ ), .B(_04591_ ), .C1(_03553_ ), .C2(_03554_ ), .ZN(_04592_ ) );
NAND2_X1 _12536_ ( .A1(_04573_ ), .A2(_04592_ ), .ZN(_04593_ ) );
INV_X1 _12537_ ( .A(_04593_ ), .ZN(_04594_ ) );
MUX2_X1 _12538_ ( .A(_02351_ ), .B(_04594_ ), .S(_03362_ ), .Z(_04595_ ) );
AOI21_X1 _12539_ ( .A(_04571_ ), .B1(_04595_ ), .B2(_03358_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND4_X1 _12540_ ( .A1(_03690_ ), .A2(_04200_ ), .A3(\mtvec [24] ), .A4(_04072_ ), .ZN(_04596_ ) );
NAND3_X1 _12541_ ( .A1(_03443_ ), .A2(_03878_ ), .A3(_04596_ ), .ZN(_04597_ ) );
NAND3_X1 _12542_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_04069_ ), .ZN(_04598_ ) );
NAND3_X1 _12543_ ( .A1(_04350_ ), .A2(\mepc [24] ), .A3(_04066_ ), .ZN(_04599_ ) );
NAND4_X1 _12544_ ( .A1(_03768_ ), .A2(_04120_ ), .A3(\mycsreg.CSReg[0][24] ), .A4(_04072_ ), .ZN(_04600_ ) );
NAND3_X1 _12545_ ( .A1(_04598_ ), .A2(_04599_ ), .A3(_04600_ ), .ZN(_04601_ ) );
OAI21_X1 _12546_ ( .A(_03646_ ), .B1(_04597_ ), .B2(_04601_ ), .ZN(_04602_ ) );
NAND4_X1 _12547_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_04077_ ), .A4(_03606_ ), .ZN(_04603_ ) );
AOI21_X1 _12548_ ( .A(_03700_ ), .B1(_04602_ ), .B2(_04603_ ), .ZN(_04604_ ) );
NAND2_X1 _12549_ ( .A1(_04604_ ), .A2(_03702_ ), .ZN(_04605_ ) );
NAND3_X1 _12550_ ( .A1(_01475_ ), .A2(_02381_ ), .A3(_01495_ ), .ZN(_04606_ ) );
NAND3_X1 _12551_ ( .A1(_04602_ ), .A2(fanout_net_7 ), .A3(_04603_ ), .ZN(_04607_ ) );
NAND2_X1 _12552_ ( .A1(_01497_ ), .A2(\ID_EX_typ [0] ), .ZN(_04608_ ) );
NAND4_X1 _12553_ ( .A1(_04606_ ), .A2(_03698_ ), .A3(_04607_ ), .A4(_04608_ ), .ZN(_04609_ ) );
AND3_X1 _12554_ ( .A1(_01366_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_typ [7] ), .ZN(_04610_ ) );
OR2_X1 _12555_ ( .A1(_03562_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04611_ ) );
OAI211_X1 _12556_ ( .A(_04611_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_30 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04612_ ) );
OR2_X1 _12557_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04613_ ) );
OAI211_X1 _12558_ ( .A(_04613_ ), .B(_03567_ ), .C1(_03568_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04614_ ) );
NAND3_X1 _12559_ ( .A1(_04612_ ), .A2(_03565_ ), .A3(_04614_ ), .ZN(_04615_ ) );
MUX2_X1 _12560_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04616_ ) );
MUX2_X1 _12561_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04617_ ) );
MUX2_X1 _12562_ ( .A(_04616_ ), .B(_04617_ ), .S(_03573_ ), .Z(_04618_ ) );
OAI211_X1 _12563_ ( .A(fanout_net_34 ), .B(_04615_ ), .C1(_04618_ ), .C2(_03575_ ), .ZN(_04619_ ) );
NOR2_X1 _12564_ ( .A1(_03617_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04620_ ) );
OAI21_X1 _12565_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_30 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04621_ ) );
NOR2_X1 _12566_ ( .A1(fanout_net_30 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04622_ ) );
OAI21_X1 _12567_ ( .A(_03573_ ), .B1(_03741_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04623_ ) );
OAI221_X1 _12568_ ( .A(_03519_ ), .B1(_04620_ ), .B2(_04621_ ), .C1(_04622_ ), .C2(_04623_ ), .ZN(_04624_ ) );
MUX2_X1 _12569_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04625_ ) );
MUX2_X1 _12570_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_30 ), .Z(_04626_ ) );
MUX2_X1 _12571_ ( .A(_04625_ ), .B(_04626_ ), .S(_03573_ ), .Z(_04627_ ) );
OAI211_X1 _12572_ ( .A(_03556_ ), .B(_04624_ ), .C1(_04627_ ), .C2(_03575_ ), .ZN(_04628_ ) );
AOI21_X1 _12573_ ( .A(_04555_ ), .B1(_04619_ ), .B2(_04628_ ), .ZN(_04629_ ) );
NOR3_X1 _12574_ ( .A1(_03586_ ), .A2(_03587_ ), .A3(\EX_LS_result_reg [24] ), .ZN(_04630_ ) );
NOR2_X1 _12575_ ( .A1(_04629_ ), .A2(_04630_ ), .ZN(_04631_ ) );
AOI21_X1 _12576_ ( .A(_04610_ ), .B1(_04631_ ), .B2(_03362_ ), .ZN(_04632_ ) );
OAI211_X1 _12577_ ( .A(_04605_ ), .B(_04609_ ), .C1(_04632_ ), .C2(_03762_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _12578_ ( .A1(_04197_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_04198_ ), .ZN(_04633_ ) );
NAND3_X1 _12579_ ( .A1(_04350_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_04069_ ), .ZN(_04634_ ) );
NAND4_X1 _12580_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [23] ), .A4(_04120_ ), .ZN(_04635_ ) );
NAND3_X1 _12581_ ( .A1(_04065_ ), .A2(\mepc [23] ), .A3(_04066_ ), .ZN(_04636_ ) );
NAND3_X1 _12582_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_04120_ ), .ZN(_04637_ ) );
AND4_X1 _12583_ ( .A1(_04634_ ), .A2(_04635_ ), .A3(_04636_ ), .A4(_04637_ ), .ZN(_04638_ ) );
AOI21_X1 _12584_ ( .A(_04633_ ), .B1(_04638_ ), .B2(_04394_ ), .ZN(_04639_ ) );
AOI21_X1 _12585_ ( .A(\ID_EX_typ [0] ), .B1(_02022_ ), .B2(_02041_ ), .ZN(_04640_ ) );
AND2_X1 _12586_ ( .A1(\ID_EX_typ [0] ), .A2(\ID_EX_imm [23] ), .ZN(_04641_ ) );
OAI221_X1 _12587_ ( .A(_03378_ ), .B1(_02379_ ), .B2(_04639_ ), .C1(_04640_ ), .C2(_04641_ ), .ZN(_04642_ ) );
AND2_X1 _12588_ ( .A1(_04634_ ), .A2(_04636_ ), .ZN(_04643_ ) );
AND2_X1 _12589_ ( .A1(_04635_ ), .A2(_04637_ ), .ZN(_04644_ ) );
NAND3_X1 _12590_ ( .A1(_04394_ ), .A2(_04643_ ), .A3(_04644_ ), .ZN(_04645_ ) );
OR3_X1 _12591_ ( .A1(_04197_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_04198_ ), .ZN(_04646_ ) );
NAND4_X1 _12592_ ( .A1(_04645_ ), .A2(_04646_ ), .A3(_03378_ ), .A4(_03702_ ), .ZN(_04647_ ) );
OR3_X1 _12593_ ( .A1(_03553_ ), .A2(_03554_ ), .A3(\EX_LS_result_reg [23] ), .ZN(_04648_ ) );
OR2_X1 _12594_ ( .A1(_03627_ ), .A2(\myreg.Reg[9][23] ), .ZN(_04649_ ) );
OAI211_X1 _12595_ ( .A(_04649_ ), .B(_03663_ ), .C1(fanout_net_30 ), .C2(\myreg.Reg[8][23] ), .ZN(_04650_ ) );
OR2_X1 _12596_ ( .A1(_03627_ ), .A2(\myreg.Reg[11][23] ), .ZN(_04651_ ) );
OAI211_X1 _12597_ ( .A(_04651_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_30 ), .C2(\myreg.Reg[10][23] ), .ZN(_04652_ ) );
NAND3_X1 _12598_ ( .A1(_04650_ ), .A2(_04652_ ), .A3(_03665_ ), .ZN(_04653_ ) );
MUX2_X1 _12599_ ( .A(\myreg.Reg[14][23] ), .B(\myreg.Reg[15][23] ), .S(fanout_net_30 ), .Z(_04654_ ) );
MUX2_X1 _12600_ ( .A(\myreg.Reg[12][23] ), .B(\myreg.Reg[13][23] ), .S(fanout_net_30 ), .Z(_04655_ ) );
MUX2_X1 _12601_ ( .A(_04654_ ), .B(_04655_ ), .S(_03567_ ), .Z(_04656_ ) );
OAI211_X1 _12602_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04653_ ), .C1(_04656_ ), .C2(_03575_ ), .ZN(_04657_ ) );
NOR2_X1 _12603_ ( .A1(_03568_ ), .A2(\myreg.Reg[3][23] ), .ZN(_04658_ ) );
OAI21_X1 _12604_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myreg.Reg[2][23] ), .ZN(_04659_ ) );
NOR2_X1 _12605_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[0][23] ), .ZN(_04660_ ) );
OAI21_X1 _12606_ ( .A(_03567_ ), .B1(_03568_ ), .B2(\myreg.Reg[1][23] ), .ZN(_04661_ ) );
OAI221_X1 _12607_ ( .A(_03565_ ), .B1(_04658_ ), .B2(_04659_ ), .C1(_04660_ ), .C2(_04661_ ), .ZN(_04662_ ) );
MUX2_X1 _12608_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04663_ ) );
MUX2_X1 _12609_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04664_ ) );
MUX2_X1 _12610_ ( .A(_04663_ ), .B(_04664_ ), .S(_03567_ ), .Z(_04665_ ) );
OAI211_X1 _12611_ ( .A(_03556_ ), .B(_04662_ ), .C1(_04665_ ), .C2(_03575_ ), .ZN(_04666_ ) );
OAI211_X1 _12612_ ( .A(_04657_ ), .B(_04666_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_04667_ ) );
NAND2_X1 _12613_ ( .A1(_04648_ ), .A2(_04667_ ), .ZN(_04668_ ) );
MUX2_X1 _12614_ ( .A(_02353_ ), .B(_04668_ ), .S(_03590_ ), .Z(_04669_ ) );
OAI211_X1 _12615_ ( .A(_04642_ ), .B(_04647_ ), .C1(_04669_ ), .C2(_03762_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _12616_ ( .A1(_03765_ ), .A2(\mepc [22] ), .A3(_04066_ ), .ZN(_04670_ ) );
NAND3_X1 _12617_ ( .A1(_03592_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_03452_ ), .ZN(_04671_ ) );
NAND4_X1 _12618_ ( .A1(_03594_ ), .A2(_03530_ ), .A3(\mycsreg.CSReg[0][22] ), .A4(_03595_ ), .ZN(_04672_ ) );
NAND4_X1 _12619_ ( .A1(_03652_ ), .A2(_03530_ ), .A3(\mtvec [22] ), .A4(_03650_ ), .ZN(_04673_ ) );
AND3_X1 _12620_ ( .A1(_04671_ ), .A2(_04672_ ), .A3(_04673_ ), .ZN(_04674_ ) );
NAND3_X1 _12621_ ( .A1(_03528_ ), .A2(_04670_ ), .A3(_04674_ ), .ZN(_04675_ ) );
OAI21_X1 _12622_ ( .A(_04675_ ), .B1(_03538_ ), .B2(_03542_ ), .ZN(_04676_ ) );
NAND4_X1 _12623_ ( .A1(_03605_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_03096_ ), .A4(_03606_ ), .ZN(_04677_ ) );
AND2_X1 _12624_ ( .A1(_04676_ ), .A2(_04677_ ), .ZN(_04678_ ) );
INV_X1 _12625_ ( .A(_04678_ ), .ZN(_04679_ ) );
OAI22_X1 _12626_ ( .A1(_04678_ ), .A2(_03548_ ), .B1(_01351_ ), .B2(_02065_ ), .ZN(_04680_ ) );
AOI21_X1 _12627_ ( .A(\ID_EX_typ [0] ), .B1(_02044_ ), .B2(_02063_ ), .ZN(_04681_ ) );
OAI221_X1 _12628_ ( .A(_03379_ ), .B1(_02379_ ), .B2(_04679_ ), .C1(_04680_ ), .C2(_04681_ ), .ZN(_04682_ ) );
NAND4_X1 _12629_ ( .A1(_02354_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_04683_ ) );
OR3_X1 _12630_ ( .A1(_03512_ ), .A2(_03498_ ), .A3(\EX_LS_result_reg [22] ), .ZN(_04684_ ) );
OR2_X1 _12631_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[0][22] ), .ZN(_04685_ ) );
OAI211_X1 _12632_ ( .A(_04685_ ), .B(_03573_ ), .C1(_03741_ ), .C2(\myreg.Reg[1][22] ), .ZN(_04686_ ) );
OR2_X1 _12633_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[2][22] ), .ZN(_04687_ ) );
OAI211_X1 _12634_ ( .A(_04687_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03741_ ), .C2(\myreg.Reg[3][22] ), .ZN(_04688_ ) );
NAND3_X1 _12635_ ( .A1(_04686_ ), .A2(_04688_ ), .A3(_03519_ ), .ZN(_04689_ ) );
MUX2_X1 _12636_ ( .A(\myreg.Reg[6][22] ), .B(\myreg.Reg[7][22] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04690_ ) );
MUX2_X1 _12637_ ( .A(\myreg.Reg[4][22] ), .B(\myreg.Reg[5][22] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04691_ ) );
MUX2_X1 _12638_ ( .A(_04690_ ), .B(_04691_ ), .S(_03616_ ), .Z(_04692_ ) );
OAI211_X1 _12639_ ( .A(_03556_ ), .B(_04689_ ), .C1(_04692_ ), .C2(_03665_ ), .ZN(_04693_ ) );
OR2_X1 _12640_ ( .A1(_03561_ ), .A2(\myreg.Reg[15][22] ), .ZN(_04694_ ) );
OAI211_X1 _12641_ ( .A(_04694_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[14][22] ), .ZN(_04695_ ) );
OR2_X1 _12642_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[12][22] ), .ZN(_04696_ ) );
OAI211_X1 _12643_ ( .A(_04696_ ), .B(_03616_ ), .C1(_03617_ ), .C2(\myreg.Reg[13][22] ), .ZN(_04697_ ) );
NAND3_X1 _12644_ ( .A1(_04695_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04697_ ), .ZN(_04698_ ) );
MUX2_X1 _12645_ ( .A(\myreg.Reg[8][22] ), .B(\myreg.Reg[9][22] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04699_ ) );
MUX2_X1 _12646_ ( .A(\myreg.Reg[10][22] ), .B(\myreg.Reg[11][22] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04700_ ) );
MUX2_X1 _12647_ ( .A(_04699_ ), .B(_04700_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04701_ ) );
OAI211_X1 _12648_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04698_ ), .C1(_04701_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04702_ ) );
OAI211_X1 _12649_ ( .A(_04693_ ), .B(_04702_ ), .C1(_03586_ ), .C2(_03587_ ), .ZN(_04703_ ) );
NAND2_X1 _12650_ ( .A1(_04684_ ), .A2(_04703_ ), .ZN(_04704_ ) );
INV_X1 _12651_ ( .A(_04704_ ), .ZN(_04705_ ) );
OAI211_X1 _12652_ ( .A(_04248_ ), .B(_04683_ ), .C1(_04705_ ), .C2(_01367_ ), .ZN(_04706_ ) );
NAND2_X1 _12653_ ( .A1(_04682_ ), .A2(_04706_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
INV_X1 _12654_ ( .A(_02267_ ), .ZN(_04707_ ) );
OR3_X1 _12655_ ( .A1(_03424_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_03432_ ), .ZN(_04708_ ) );
NAND4_X1 _12656_ ( .A1(_03457_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [31] ), .A4(_04071_ ), .ZN(_04709_ ) );
NAND3_X1 _12657_ ( .A1(_04065_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_04069_ ), .ZN(_04710_ ) );
NAND3_X1 _12658_ ( .A1(_04065_ ), .A2(\mepc [31] ), .A3(_04066_ ), .ZN(_04711_ ) );
NAND3_X1 _12659_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04071_ ), .ZN(_04712_ ) );
NAND4_X1 _12660_ ( .A1(_04709_ ), .A2(_04710_ ), .A3(_04711_ ), .A4(_04712_ ), .ZN(_04713_ ) );
OAI21_X1 _12661_ ( .A(_04708_ ), .B1(_03939_ ), .B2(_04713_ ), .ZN(_04714_ ) );
AOI22_X1 _12662_ ( .A1(_04707_ ), .A2(_01351_ ), .B1(fanout_net_7 ), .B2(_04714_ ), .ZN(_04715_ ) );
OAI211_X1 _12663_ ( .A(_04715_ ), .B(_03551_ ), .C1(_02381_ ), .C2(\ID_EX_imm [31] ), .ZN(_04716_ ) );
AND2_X1 _12664_ ( .A1(_04710_ ), .A2(_04711_ ), .ZN(_04717_ ) );
AND2_X1 _12665_ ( .A1(_04709_ ), .A2(_04712_ ), .ZN(_04718_ ) );
NAND3_X1 _12666_ ( .A1(_04394_ ), .A2(_04717_ ), .A3(_04718_ ), .ZN(_04719_ ) );
NAND4_X1 _12667_ ( .A1(_04719_ ), .A2(_04708_ ), .A3(_03378_ ), .A4(_03702_ ), .ZN(_04720_ ) );
AND3_X1 _12668_ ( .A1(_01366_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_04721_ ) );
OR2_X1 _12669_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04722_ ) );
OAI211_X1 _12670_ ( .A(_04722_ ), .B(_03624_ ), .C1(_03627_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04723_ ) );
OR2_X1 _12671_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04724_ ) );
OAI211_X1 _12672_ ( .A(_04724_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_03627_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04725_ ) );
NAND3_X1 _12673_ ( .A1(_04723_ ), .A2(_04725_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04726_ ) );
MUX2_X1 _12674_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04727_ ) );
MUX2_X1 _12675_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04728_ ) );
MUX2_X1 _12676_ ( .A(_04727_ ), .B(_04728_ ), .S(_03624_ ), .Z(_04729_ ) );
OAI211_X1 _12677_ ( .A(_03494_ ), .B(_04726_ ), .C1(_04729_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04730_ ) );
NOR2_X1 _12678_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04731_ ) );
OAI21_X1 _12679_ ( .A(_03482_ ), .B1(_03561_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04732_ ) );
MUX2_X1 _12680_ ( .A(_02258_ ), .B(_02259_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04733_ ) );
OAI221_X1 _12681_ ( .A(_03490_ ), .B1(_04731_ ), .B2(_04732_ ), .C1(_04733_ ), .C2(_03616_ ), .ZN(_04734_ ) );
MUX2_X1 _12682_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04735_ ) );
MUX2_X1 _12683_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_04736_ ) );
MUX2_X1 _12684_ ( .A(_04735_ ), .B(_04736_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04737_ ) );
OAI211_X1 _12685_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_04734_ ), .C1(_04737_ ), .C2(_03565_ ), .ZN(_04738_ ) );
AOI21_X1 _12686_ ( .A(_04555_ ), .B1(_04730_ ), .B2(_04738_ ), .ZN(_04739_ ) );
AND2_X1 _12687_ ( .A1(_04555_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04740_ ) );
NOR2_X1 _12688_ ( .A1(_04739_ ), .A2(_04740_ ), .ZN(_04741_ ) );
AOI21_X1 _12689_ ( .A(_04721_ ), .B1(_04741_ ), .B2(_03362_ ), .ZN(_04742_ ) );
OAI211_X1 _12690_ ( .A(_04716_ ), .B(_04720_ ), .C1(_03762_ ), .C2(_04742_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
INV_X1 _12691_ ( .A(_03470_ ), .ZN(_04743_ ) );
AND2_X1 _12692_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_04744_ ) );
AND2_X1 _12693_ ( .A1(_04744_ ), .A2(\ID_EX_pc [4] ), .ZN(_04745_ ) );
AND2_X1 _12694_ ( .A1(_04745_ ), .A2(\ID_EX_pc [5] ), .ZN(_04746_ ) );
AND2_X1 _12695_ ( .A1(_04746_ ), .A2(\ID_EX_pc [6] ), .ZN(_04747_ ) );
AND2_X1 _12696_ ( .A1(_04747_ ), .A2(\ID_EX_pc [7] ), .ZN(_04748_ ) );
AND2_X1 _12697_ ( .A1(_04748_ ), .A2(\ID_EX_pc [8] ), .ZN(_04749_ ) );
AND2_X1 _12698_ ( .A1(_04749_ ), .A2(\ID_EX_pc [9] ), .ZN(_04750_ ) );
AND4_X1 _12699_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_04751_ ) );
AND2_X1 _12700_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_04752_ ) );
AND4_X2 _12701_ ( .A1(\ID_EX_pc [13] ), .A2(_04751_ ), .A3(\ID_EX_pc [12] ), .A4(_04752_ ), .ZN(_04753_ ) );
AND2_X1 _12702_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_04754_ ) );
NAND3_X1 _12703_ ( .A1(_04750_ ), .A2(_04753_ ), .A3(_04754_ ), .ZN(_04755_ ) );
NOR2_X1 _12704_ ( .A1(_04755_ ), .A2(_02327_ ), .ZN(_04756_ ) );
XNOR2_X1 _12705_ ( .A(_04756_ ), .B(_02326_ ), .ZN(_04757_ ) );
AND2_X2 _12706_ ( .A1(_01360_ ), .A2(_01355_ ), .ZN(_04758_ ) );
BUF_X4 _12707_ ( .A(_04758_ ), .Z(_04759_ ) );
AND2_X1 _12708_ ( .A1(_03876_ ), .A2(_03850_ ), .ZN(_04760_ ) );
NOR2_X1 _12709_ ( .A1(_03876_ ), .A2(_03850_ ), .ZN(_04761_ ) );
NOR2_X2 _12710_ ( .A1(_04760_ ), .A2(_04761_ ), .ZN(_04762_ ) );
INV_X1 _12711_ ( .A(_01808_ ), .ZN(_04763_ ) );
XNOR2_X1 _12712_ ( .A(_04763_ ), .B(_03913_ ), .ZN(_04764_ ) );
AND2_X1 _12713_ ( .A1(_04762_ ), .A2(_04764_ ), .ZN(_04765_ ) );
INV_X1 _12714_ ( .A(_01760_ ), .ZN(_04766_ ) );
XNOR2_X2 _12715_ ( .A(_04766_ ), .B(_03802_ ), .ZN(_04767_ ) );
XNOR2_X2 _12716_ ( .A(_03814_ ), .B(_03838_ ), .ZN(_04768_ ) );
AND3_X2 _12717_ ( .A1(_04765_ ), .A2(_04767_ ), .A3(_04768_ ), .ZN(_04769_ ) );
INV_X1 _12718_ ( .A(_04769_ ), .ZN(_04770_ ) );
NAND2_X1 _12719_ ( .A1(_01861_ ), .A2(_01881_ ), .ZN(_04771_ ) );
INV_X1 _12720_ ( .A(_04771_ ), .ZN(_04772_ ) );
XNOR2_X2 _12721_ ( .A(_04772_ ), .B(_03986_ ), .ZN(_04773_ ) );
INV_X1 _12722_ ( .A(_01905_ ), .ZN(_04774_ ) );
XNOR2_X2 _12723_ ( .A(_04774_ ), .B(_04025_ ), .ZN(_04775_ ) );
AND2_X2 _12724_ ( .A1(_04773_ ), .A2(_04775_ ), .ZN(_04776_ ) );
INV_X1 _12725_ ( .A(_01854_ ), .ZN(_04777_ ) );
XNOR2_X2 _12726_ ( .A(_04777_ ), .B(_04061_ ), .ZN(_04778_ ) );
INV_X1 _12727_ ( .A(_01832_ ), .ZN(_04779_ ) );
XNOR2_X2 _12728_ ( .A(_04779_ ), .B(_04104_ ), .ZN(_04780_ ) );
AND3_X1 _12729_ ( .A1(_04776_ ), .A2(_04778_ ), .A3(_04780_ ), .ZN(_04781_ ) );
INV_X1 _12730_ ( .A(_04781_ ), .ZN(_04782_ ) );
XNOR2_X2 _12731_ ( .A(_04384_ ), .B(_04419_ ), .ZN(_04783_ ) );
OAI21_X2 _12732_ ( .A(_04783_ ), .B1(_03359_ ), .B2(_04454_ ), .ZN(_04784_ ) );
NAND2_X1 _12733_ ( .A1(_04419_ ), .A2(_01571_ ), .ZN(_04785_ ) );
AND2_X4 _12734_ ( .A1(_04784_ ), .A2(_04785_ ), .ZN(_04786_ ) );
INV_X1 _12735_ ( .A(_01547_ ), .ZN(_04787_ ) );
XNOR2_X1 _12736_ ( .A(_04787_ ), .B(_04332_ ), .ZN(_04788_ ) );
INV_X2 _12737_ ( .A(_04788_ ), .ZN(_04789_ ) );
OR2_X4 _12738_ ( .A1(_04786_ ), .A2(_04789_ ), .ZN(_04790_ ) );
AND2_X1 _12739_ ( .A1(_04332_ ), .A2(_01547_ ), .ZN(_04791_ ) );
INV_X1 _12740_ ( .A(_04791_ ), .ZN(_04792_ ) );
AOI22_X4 _12741_ ( .A1(_04790_ ), .A2(_04792_ ), .B1(_01601_ ), .B2(_04309_ ), .ZN(_04793_ ) );
NOR2_X1 _12742_ ( .A1(_01601_ ), .A2(_04309_ ), .ZN(_04794_ ) );
OR2_X2 _12743_ ( .A1(_04793_ ), .A2(_04794_ ), .ZN(_04795_ ) );
AND2_X4 _12744_ ( .A1(_01684_ ), .A2(_04149_ ), .ZN(_04796_ ) );
NOR2_X2 _12745_ ( .A1(_01684_ ), .A2(_04149_ ), .ZN(_04797_ ) );
NOR2_X2 _12746_ ( .A1(_04796_ ), .A2(_04797_ ), .ZN(_04798_ ) );
INV_X4 _12747_ ( .A(_01707_ ), .ZN(_04799_ ) );
XNOR2_X1 _12748_ ( .A(_04799_ ), .B(_04171_ ), .ZN(_04800_ ) );
XNOR2_X2 _12749_ ( .A(_04239_ ), .B(_04270_ ), .ZN(_04801_ ) );
XNOR2_X1 _12750_ ( .A(_04227_ ), .B(_01657_ ), .ZN(_04802_ ) );
AND2_X1 _12751_ ( .A1(_04801_ ), .A2(_04802_ ), .ZN(_04803_ ) );
NAND4_X4 _12752_ ( .A1(_04795_ ), .A2(_04798_ ), .A3(_04800_ ), .A4(_04803_ ), .ZN(_04804_ ) );
AND2_X4 _12753_ ( .A1(_04270_ ), .A2(_03394_ ), .ZN(_04805_ ) );
AND2_X4 _12754_ ( .A1(_04802_ ), .A2(_04805_ ), .ZN(_04806_ ) );
AOI21_X4 _12755_ ( .A(_04806_ ), .B1(_01657_ ), .B2(_04228_ ), .ZN(_04807_ ) );
INV_X1 _12756_ ( .A(_04798_ ), .ZN(_04808_ ) );
INV_X1 _12757_ ( .A(_04800_ ), .ZN(_04809_ ) );
NOR3_X2 _12758_ ( .A1(_04807_ ), .A2(_04808_ ), .A3(_04809_ ), .ZN(_04810_ ) );
NAND2_X1 _12759_ ( .A1(_04171_ ), .A2(_01707_ ), .ZN(_04811_ ) );
NOR3_X1 _12760_ ( .A1(_04796_ ), .A2(_04797_ ), .A3(_04811_ ), .ZN(_04812_ ) );
NOR3_X1 _12761_ ( .A1(_04810_ ), .A2(_04796_ ), .A3(_04812_ ), .ZN(_04813_ ) );
AOI211_X2 _12762_ ( .A(_04770_ ), .B(_04782_ ), .C1(_04804_ ), .C2(_04813_ ), .ZN(_04814_ ) );
AND2_X1 _12763_ ( .A1(_03802_ ), .A2(_01760_ ), .ZN(_04815_ ) );
NAND2_X1 _12764_ ( .A1(_04061_ ), .A2(_01854_ ), .ZN(_04816_ ) );
INV_X2 _12765_ ( .A(_04778_ ), .ZN(_04817_ ) );
NAND2_X2 _12766_ ( .A1(_04104_ ), .A2(_01832_ ), .ZN(_04818_ ) );
OAI21_X2 _12767_ ( .A(_04816_ ), .B1(_04817_ ), .B2(_04818_ ), .ZN(_04819_ ) );
AND2_X4 _12768_ ( .A1(_04819_ ), .A2(_04776_ ), .ZN(_04820_ ) );
AND2_X1 _12769_ ( .A1(_03986_ ), .A2(_04771_ ), .ZN(_04821_ ) );
AND2_X1 _12770_ ( .A1(_04025_ ), .A2(_01905_ ), .ZN(_04822_ ) );
AND2_X1 _12771_ ( .A1(_04773_ ), .A2(_04822_ ), .ZN(_04823_ ) );
NOR3_X4 _12772_ ( .A1(_04820_ ), .A2(_04821_ ), .A3(_04823_ ), .ZN(_04824_ ) );
NOR2_X1 _12773_ ( .A1(_04824_ ), .A2(_04770_ ), .ZN(_04825_ ) );
AND2_X1 _12774_ ( .A1(_03838_ ), .A2(_01738_ ), .ZN(_04826_ ) );
AND2_X1 _12775_ ( .A1(_04767_ ), .A2(_04826_ ), .ZN(_04827_ ) );
INV_X1 _12776_ ( .A(_04760_ ), .ZN(_04828_ ) );
NAND2_X1 _12777_ ( .A1(_03913_ ), .A2(_01808_ ), .ZN(_04829_ ) );
AOI21_X1 _12778_ ( .A(_04761_ ), .B1(_04828_ ), .B2(_04829_ ), .ZN(_04830_ ) );
AND3_X1 _12779_ ( .A1(_04830_ ), .A2(_04767_ ), .A3(_04768_ ), .ZN(_04831_ ) );
OR4_X4 _12780_ ( .A1(_04815_ ), .A2(_04825_ ), .A3(_04827_ ), .A4(_04831_ ), .ZN(_04832_ ) );
NOR2_X2 _12781_ ( .A1(_04814_ ), .A2(_04832_ ), .ZN(_04833_ ) );
INV_X2 _12782_ ( .A(_04833_ ), .ZN(_04834_ ) );
NAND2_X1 _12783_ ( .A1(_01974_ ), .A2(_01994_ ), .ZN(_04835_ ) );
INV_X1 _12784_ ( .A(_04835_ ), .ZN(_04836_ ) );
XNOR2_X1 _12785_ ( .A(_04836_ ), .B(_03638_ ), .ZN(_04837_ ) );
XNOR2_X1 _12786_ ( .A(_02123_ ), .B(_03683_ ), .ZN(_04838_ ) );
AND2_X1 _12787_ ( .A1(_04837_ ), .A2(_04838_ ), .ZN(_04839_ ) );
INV_X1 _12788_ ( .A(_01969_ ), .ZN(_04840_ ) );
XNOR2_X1 _12789_ ( .A(_04840_ ), .B(_03760_ ), .ZN(_04841_ ) );
INV_X1 _12790_ ( .A(_01945_ ), .ZN(_04842_ ) );
XNOR2_X1 _12791_ ( .A(_04842_ ), .B(_03724_ ), .ZN(_04843_ ) );
NAND4_X4 _12792_ ( .A1(_04834_ ), .A2(_04839_ ), .A3(_04841_ ), .A4(_04843_ ), .ZN(_04844_ ) );
AND2_X1 _12793_ ( .A1(_03683_ ), .A2(_02018_ ), .ZN(_04845_ ) );
AND2_X1 _12794_ ( .A1(_04837_ ), .A2(_04845_ ), .ZN(_04846_ ) );
AOI21_X1 _12795_ ( .A(_04846_ ), .B1(_04835_ ), .B2(_03638_ ), .ZN(_04847_ ) );
AND2_X1 _12796_ ( .A1(_03724_ ), .A2(_01945_ ), .ZN(_04848_ ) );
NOR2_X1 _12797_ ( .A1(_03724_ ), .A2(_01945_ ), .ZN(_04849_ ) );
INV_X1 _12798_ ( .A(_03760_ ), .ZN(_04850_ ) );
NOR4_X4 _12799_ ( .A1(_04848_ ), .A2(_04849_ ), .A3(_04840_ ), .A4(_04850_ ), .ZN(_04851_ ) );
OAI211_X1 _12800_ ( .A(_04837_ ), .B(_04838_ ), .C1(_04851_ ), .C2(_04848_ ), .ZN(_04852_ ) );
AND2_X1 _12801_ ( .A1(_04847_ ), .A2(_04852_ ), .ZN(_04853_ ) );
NAND2_X4 _12802_ ( .A1(_04844_ ), .A2(_04853_ ), .ZN(_04854_ ) );
INV_X1 _12803_ ( .A(_02088_ ), .ZN(_04855_ ) );
XNOR2_X1 _12804_ ( .A(_04855_ ), .B(_03589_ ), .ZN(_04856_ ) );
NAND2_X1 _12805_ ( .A1(_04854_ ), .A2(_04856_ ), .ZN(_04857_ ) );
XNOR2_X1 _12806_ ( .A(_03524_ ), .B(_03472_ ), .ZN(_04858_ ) );
INV_X1 _12807_ ( .A(_04858_ ), .ZN(_04859_ ) );
NAND2_X1 _12808_ ( .A1(_03589_ ), .A2(_02088_ ), .ZN(_04860_ ) );
AND3_X1 _12809_ ( .A1(_04857_ ), .A2(_04859_ ), .A3(_04860_ ), .ZN(_04861_ ) );
AOI21_X1 _12810_ ( .A(_04859_ ), .B1(_04857_ ), .B2(_04860_ ), .ZN(_04862_ ) );
NOR2_X1 _12811_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .ZN(_04863_ ) );
AND3_X1 _12812_ ( .A1(_04863_ ), .A2(\ID_EX_typ [3] ), .A3(_02378_ ), .ZN(_04864_ ) );
AND2_X1 _12813_ ( .A1(_04864_ ), .A2(_02376_ ), .ZN(_04865_ ) );
INV_X1 _12814_ ( .A(_04865_ ), .ZN(_04866_ ) );
BUF_X2 _12815_ ( .A(_04866_ ), .Z(_04867_ ) );
NOR3_X1 _12816_ ( .A1(_04861_ ), .A2(_04862_ ), .A3(_04867_ ), .ZN(_04868_ ) );
XOR2_X1 _12817_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_04869_ ) );
XOR2_X1 _12818_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_04870_ ) );
AND2_X1 _12819_ ( .A1(_04869_ ), .A2(_04870_ ), .ZN(_04871_ ) );
AND2_X1 _12820_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_imm [13] ), .ZN(_04872_ ) );
NOR2_X1 _12821_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_imm [13] ), .ZN(_04873_ ) );
NOR2_X1 _12822_ ( .A1(_04872_ ), .A2(_04873_ ), .ZN(_04874_ ) );
XOR2_X1 _12823_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_04875_ ) );
AND3_X1 _12824_ ( .A1(_04871_ ), .A2(_04874_ ), .A3(_04875_ ), .ZN(_04876_ ) );
XOR2_X1 _12825_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_04877_ ) );
AND2_X1 _12826_ ( .A1(\ID_EX_pc [9] ), .A2(\ID_EX_imm [9] ), .ZN(_04878_ ) );
NOR2_X1 _12827_ ( .A1(\ID_EX_pc [9] ), .A2(\ID_EX_imm [9] ), .ZN(_04879_ ) );
NOR2_X1 _12828_ ( .A1(_04878_ ), .A2(_04879_ ), .ZN(_04880_ ) );
AND2_X1 _12829_ ( .A1(_04877_ ), .A2(_04880_ ), .ZN(_04881_ ) );
XOR2_X1 _12830_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_04882_ ) );
XOR2_X1 _12831_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_04883_ ) );
AND3_X1 _12832_ ( .A1(_04881_ ), .A2(_04882_ ), .A3(_04883_ ), .ZN(_04884_ ) );
XOR2_X1 _12833_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_04885_ ) );
INV_X1 _12834_ ( .A(_04885_ ), .ZN(_04886_ ) );
XOR2_X1 _12835_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_04887_ ) );
AND2_X1 _12836_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_04888_ ) );
AND2_X1 _12837_ ( .A1(_04887_ ), .A2(_04888_ ), .ZN(_04889_ ) );
AOI21_X1 _12838_ ( .A(_04889_ ), .B1(\ID_EX_pc [1] ), .B2(\ID_EX_imm [1] ), .ZN(_04890_ ) );
XOR2_X1 _12839_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_04891_ ) );
INV_X1 _12840_ ( .A(_04891_ ), .ZN(_04892_ ) );
AND2_X1 _12841_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_04893_ ) );
NOR2_X1 _12842_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_04894_ ) );
NOR2_X1 _12843_ ( .A1(_04893_ ), .A2(_04894_ ), .ZN(_04895_ ) );
INV_X1 _12844_ ( .A(_04895_ ), .ZN(_04896_ ) );
OR3_X1 _12845_ ( .A1(_04890_ ), .A2(_04892_ ), .A3(_04896_ ), .ZN(_04897_ ) );
AND2_X1 _12846_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_04898_ ) );
AOI21_X1 _12847_ ( .A(_04893_ ), .B1(_04895_ ), .B2(_04898_ ), .ZN(_04899_ ) );
AOI21_X1 _12848_ ( .A(_04886_ ), .B1(_04897_ ), .B2(_04899_ ), .ZN(_04900_ ) );
AND2_X1 _12849_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_04901_ ) );
AND2_X1 _12850_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_04902_ ) );
NOR3_X1 _12851_ ( .A1(_04900_ ), .A2(_04901_ ), .A3(_04902_ ), .ZN(_04903_ ) );
NOR2_X1 _12852_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_04904_ ) );
NOR2_X1 _12853_ ( .A1(_04903_ ), .A2(_04904_ ), .ZN(_04905_ ) );
XOR2_X1 _12854_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_04906_ ) );
AND2_X1 _12855_ ( .A1(_04905_ ), .A2(_04906_ ), .ZN(_04907_ ) );
AND2_X1 _12856_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_04908_ ) );
NOR2_X1 _12857_ ( .A1(_04907_ ), .A2(_04908_ ), .ZN(_04909_ ) );
NOR2_X1 _12858_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04910_ ) );
NOR2_X1 _12859_ ( .A1(_04909_ ), .A2(_04910_ ), .ZN(_04911_ ) );
AND2_X1 _12860_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04912_ ) );
OAI211_X1 _12861_ ( .A(_04876_ ), .B(_04884_ ), .C1(_04911_ ), .C2(_04912_ ), .ZN(_04913_ ) );
AND2_X1 _12862_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04914_ ) );
NAND2_X1 _12863_ ( .A1(_04869_ ), .A2(_04914_ ), .ZN(_04915_ ) );
OAI21_X1 _12864_ ( .A(_04915_ ), .B1(_02332_ ), .B2(_01761_ ), .ZN(_04916_ ) );
AND2_X1 _12865_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_04917_ ) );
NOR2_X1 _12866_ ( .A1(_04917_ ), .A2(_04872_ ), .ZN(_04918_ ) );
NOR2_X1 _12867_ ( .A1(_04918_ ), .A2(_04873_ ), .ZN(_04919_ ) );
AND2_X1 _12868_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_04920_ ) );
AND2_X1 _12869_ ( .A1(_04882_ ), .A2(_04920_ ), .ZN(_04921_ ) );
AOI21_X1 _12870_ ( .A(_04921_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_04922_ ) );
AND2_X1 _12871_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_04923_ ) );
AND2_X1 _12872_ ( .A1(_04880_ ), .A2(_04923_ ), .ZN(_04924_ ) );
OAI211_X1 _12873_ ( .A(_04882_ ), .B(_04883_ ), .C1(_04924_ ), .C2(_04878_ ), .ZN(_04925_ ) );
AND2_X1 _12874_ ( .A1(_04922_ ), .A2(_04925_ ), .ZN(_04926_ ) );
INV_X1 _12875_ ( .A(_04926_ ), .ZN(_04927_ ) );
AOI221_X4 _12876_ ( .A(_04916_ ), .B1(_04871_ ), .B2(_04919_ ), .C1(_04927_ ), .C2(_04876_ ), .ZN(_04928_ ) );
NAND2_X1 _12877_ ( .A1(_04913_ ), .A2(_04928_ ), .ZN(_04929_ ) );
XOR2_X1 _12878_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_04930_ ) );
XOR2_X1 _12879_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_04931_ ) );
AND2_X1 _12880_ ( .A1(_04930_ ), .A2(_04931_ ), .ZN(_04932_ ) );
XOR2_X1 _12881_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_04933_ ) );
XOR2_X1 _12882_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_04934_ ) );
AND2_X1 _12883_ ( .A1(_04933_ ), .A2(_04934_ ), .ZN(_04935_ ) );
NAND3_X1 _12884_ ( .A1(_04929_ ), .A2(_04932_ ), .A3(_04935_ ), .ZN(_04936_ ) );
AND2_X1 _12885_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_04937_ ) );
AND2_X1 _12886_ ( .A1(_04934_ ), .A2(_04937_ ), .ZN(_04938_ ) );
AOI21_X1 _12887_ ( .A(_04938_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_04939_ ) );
INV_X1 _12888_ ( .A(_04939_ ), .ZN(_04940_ ) );
AND2_X1 _12889_ ( .A1(_04940_ ), .A2(_04932_ ), .ZN(_04941_ ) );
AND2_X1 _12890_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_imm [19] ), .ZN(_04942_ ) );
AOI211_X1 _12891_ ( .A(_02329_ ), .B(_02019_ ), .C1(_02328_ ), .C2(_01975_ ), .ZN(_04943_ ) );
NOR3_X1 _12892_ ( .A1(_04941_ ), .A2(_04942_ ), .A3(_04943_ ), .ZN(_04944_ ) );
AND2_X1 _12893_ ( .A1(_04936_ ), .A2(_04944_ ), .ZN(_04945_ ) );
XOR2_X1 _12894_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_04946_ ) );
INV_X1 _12895_ ( .A(_04946_ ), .ZN(_04947_ ) );
NOR2_X1 _12896_ ( .A1(_04945_ ), .A2(_04947_ ), .ZN(_04948_ ) );
AND2_X1 _12897_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_04949_ ) );
XOR2_X1 _12898_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_04950_ ) );
NOR3_X1 _12899_ ( .A1(_04948_ ), .A2(_04949_ ), .A3(_04950_ ), .ZN(_04951_ ) );
NOR3_X1 _12900_ ( .A1(_02376_ ), .A2(\ID_EX_typ [1] ), .A3(\ID_EX_typ [0] ), .ZN(_04952_ ) );
AND2_X1 _12901_ ( .A1(\ID_EX_typ [3] ), .A2(fanout_net_7 ), .ZN(_04953_ ) );
AND2_X2 _12902_ ( .A1(_04952_ ), .A2(_04953_ ), .ZN(_04954_ ) );
INV_X1 _12903_ ( .A(_04954_ ), .ZN(_04955_ ) );
AND2_X1 _12904_ ( .A1(_04950_ ), .A2(_04949_ ), .ZN(_04956_ ) );
NOR3_X1 _12905_ ( .A1(_04951_ ), .A2(_04955_ ), .A3(_04956_ ), .ZN(_04957_ ) );
INV_X1 _12906_ ( .A(_04950_ ), .ZN(_04958_ ) );
OR3_X1 _12907_ ( .A1(_04945_ ), .A2(_04947_ ), .A3(_04958_ ), .ZN(_04959_ ) );
NAND2_X1 _12908_ ( .A1(_04957_ ), .A2(_04959_ ), .ZN(_04960_ ) );
NOR3_X1 _12909_ ( .A1(_02377_ ), .A2(_02378_ ), .A3(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ), .ZN(_04961_ ) );
BUF_X4 _12910_ ( .A(_04961_ ), .Z(_04962_ ) );
NOR2_X1 _12911_ ( .A1(_02380_ ), .A2(\ID_EX_typ [0] ), .ZN(_04963_ ) );
BUF_X4 _12912_ ( .A(_04963_ ), .Z(_04964_ ) );
NAND3_X1 _12913_ ( .A1(_04962_ ), .A2(\ID_EX_imm [21] ), .A3(_04964_ ), .ZN(_04965_ ) );
NAND2_X1 _12914_ ( .A1(_04960_ ), .A2(_04965_ ), .ZN(_04966_ ) );
OAI21_X1 _12915_ ( .A(_04759_ ), .B1(_04868_ ), .B2(_04966_ ), .ZN(_04967_ ) );
AND2_X1 _12916_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .ZN(_04968_ ) );
AND2_X2 _12917_ ( .A1(_04968_ ), .A2(fanout_net_7 ), .ZN(_04969_ ) );
INV_X1 _12918_ ( .A(_04969_ ), .ZN(_04970_ ) );
NAND2_X2 _12919_ ( .A1(_04454_ ), .A2(_02374_ ), .ZN(_04971_ ) );
NAND2_X1 _12920_ ( .A1(_01575_ ), .A2(fanout_net_8 ), .ZN(_04972_ ) );
NAND2_X4 _12921_ ( .A1(_04971_ ), .A2(_04972_ ), .ZN(_04973_ ) );
NAND3_X1 _12922_ ( .A1(_04399_ ), .A2(_04418_ ), .A3(_02373_ ), .ZN(_04974_ ) );
NAND2_X1 _12923_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [1] ), .ZN(_04975_ ) );
AND2_X2 _12924_ ( .A1(_04974_ ), .A2(_04975_ ), .ZN(_04976_ ) );
AND2_X4 _12925_ ( .A1(_04973_ ), .A2(_04976_ ), .ZN(_04977_ ) );
NAND3_X1 _12926_ ( .A1(_04312_ ), .A2(_04331_ ), .A3(_02374_ ), .ZN(_04978_ ) );
NAND2_X1 _12927_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [2] ), .ZN(_04979_ ) );
AND2_X1 _12928_ ( .A1(_04978_ ), .A2(_04979_ ), .ZN(_04980_ ) );
BUF_X4 _12929_ ( .A(_04980_ ), .Z(_04981_ ) );
AND2_X4 _12930_ ( .A1(_04977_ ), .A2(_04981_ ), .ZN(_04982_ ) );
NAND3_X1 _12931_ ( .A1(_04289_ ), .A2(_02374_ ), .A3(_04308_ ), .ZN(_04983_ ) );
NAND2_X1 _12932_ ( .A1(fanout_net_8 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_04984_ ) );
AND2_X4 _12933_ ( .A1(_04983_ ), .A2(_04984_ ), .ZN(_04985_ ) );
INV_X4 _12934_ ( .A(_04985_ ), .ZN(_04986_ ) );
AND2_X4 _12935_ ( .A1(_04982_ ), .A2(_04986_ ), .ZN(_04987_ ) );
NAND3_X1 _12936_ ( .A1(_04250_ ), .A2(_04269_ ), .A3(_02375_ ), .ZN(_04988_ ) );
NAND2_X1 _12937_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [4] ), .ZN(_04989_ ) );
AND2_X2 _12938_ ( .A1(_04988_ ), .A2(_04989_ ), .ZN(_04990_ ) );
AND2_X4 _12939_ ( .A1(_04987_ ), .A2(_04990_ ), .ZN(_04991_ ) );
NAND2_X1 _12940_ ( .A1(_04227_ ), .A2(_02374_ ), .ZN(_04992_ ) );
NAND2_X1 _12941_ ( .A1(_01660_ ), .A2(fanout_net_8 ), .ZN(_04993_ ) );
NAND2_X4 _12942_ ( .A1(_04992_ ), .A2(_04993_ ), .ZN(_04994_ ) );
INV_X1 _12943_ ( .A(_04994_ ), .ZN(_04995_ ) );
NOR2_X4 _12944_ ( .A1(_04991_ ), .A2(_04995_ ), .ZN(_04996_ ) );
NAND3_X1 _12945_ ( .A1(_04129_ ), .A2(_02374_ ), .A3(_04148_ ), .ZN(_04997_ ) );
NAND2_X1 _12946_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [7] ), .ZN(_04998_ ) );
AND2_X2 _12947_ ( .A1(_04997_ ), .A2(_04998_ ), .ZN(_04999_ ) );
NAND3_X1 _12948_ ( .A1(_04151_ ), .A2(_04170_ ), .A3(_02374_ ), .ZN(_05000_ ) );
NAND2_X1 _12949_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [6] ), .ZN(_05001_ ) );
AND2_X2 _12950_ ( .A1(_05000_ ), .A2(_05001_ ), .ZN(_05002_ ) );
AND2_X1 _12951_ ( .A1(_04999_ ), .A2(_05002_ ), .ZN(_05003_ ) );
INV_X1 _12952_ ( .A(_05003_ ), .ZN(_05004_ ) );
NOR2_X4 _12953_ ( .A1(_04996_ ), .A2(_05004_ ), .ZN(_05005_ ) );
NAND3_X1 _12954_ ( .A1(_04041_ ), .A2(_02375_ ), .A3(_04060_ ), .ZN(_05006_ ) );
NAND2_X1 _12955_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [9] ), .ZN(_05007_ ) );
AND2_X2 _12956_ ( .A1(_05006_ ), .A2(_05007_ ), .ZN(_05008_ ) );
NAND3_X1 _12957_ ( .A1(_04084_ ), .A2(_04103_ ), .A3(_02375_ ), .ZN(_05009_ ) );
NAND2_X1 _12958_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [8] ), .ZN(_05010_ ) );
AND2_X2 _12959_ ( .A1(_05009_ ), .A2(_05010_ ), .ZN(_05011_ ) );
NOR3_X1 _12960_ ( .A1(_05005_ ), .A2(_05008_ ), .A3(_05011_ ), .ZN(_05012_ ) );
AND2_X1 _12961_ ( .A1(_05008_ ), .A2(_05011_ ), .ZN(_05013_ ) );
AND2_X4 _12962_ ( .A1(_05005_ ), .A2(_05013_ ), .ZN(_05014_ ) );
OR2_X4 _12963_ ( .A1(_05012_ ), .A2(_05014_ ), .ZN(_05015_ ) );
INV_X1 _12964_ ( .A(_05005_ ), .ZN(_05016_ ) );
OR4_X1 _12965_ ( .A1(_04999_ ), .A2(_04991_ ), .A3(_05002_ ), .A4(_04995_ ), .ZN(_05017_ ) );
AOI21_X1 _12966_ ( .A(_04707_ ), .B1(_05016_ ), .B2(_05017_ ), .ZN(_05018_ ) );
AND2_X4 _12967_ ( .A1(_05015_ ), .A2(_05018_ ), .ZN(_05019_ ) );
NAND3_X1 _12968_ ( .A1(_03966_ ), .A2(_02374_ ), .A3(_03985_ ), .ZN(_05020_ ) );
NAND2_X1 _12969_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [11] ), .ZN(_05021_ ) );
AND2_X1 _12970_ ( .A1(_05020_ ), .A2(_05021_ ), .ZN(_05022_ ) );
NAND3_X1 _12971_ ( .A1(_04004_ ), .A2(_04024_ ), .A3(_02375_ ), .ZN(_05023_ ) );
NAND2_X1 _12972_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [10] ), .ZN(_05024_ ) );
AND2_X1 _12973_ ( .A1(_05023_ ), .A2(_05024_ ), .ZN(_05025_ ) );
BUF_X2 _12974_ ( .A(_02375_ ), .Z(_05026_ ) );
NAND3_X1 _12975_ ( .A1(_03661_ ), .A2(_03682_ ), .A3(_05026_ ), .ZN(_05027_ ) );
NAND2_X1 _12976_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [18] ), .ZN(_05028_ ) );
AND2_X1 _12977_ ( .A1(_05027_ ), .A2(_05028_ ), .ZN(_05029_ ) );
NAND3_X1 _12978_ ( .A1(_03704_ ), .A2(_05026_ ), .A3(_03723_ ), .ZN(_05030_ ) );
NAND2_X1 _12979_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [17] ), .ZN(_05031_ ) );
AND2_X4 _12980_ ( .A1(_05030_ ), .A2(_05031_ ), .ZN(_05032_ ) );
NAND3_X1 _12981_ ( .A1(_03739_ ), .A2(_03759_ ), .A3(_05026_ ), .ZN(_05033_ ) );
NAND2_X1 _12982_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [16] ), .ZN(_05034_ ) );
AND2_X1 _12983_ ( .A1(_05033_ ), .A2(_05034_ ), .ZN(_05035_ ) );
NAND3_X1 _12984_ ( .A1(_04554_ ), .A2(_04556_ ), .A3(_02376_ ), .ZN(_05036_ ) );
NAND2_X1 _12985_ ( .A1(_02183_ ), .A2(fanout_net_8 ), .ZN(_05037_ ) );
NAND2_X1 _12986_ ( .A1(_05036_ ), .A2(_05037_ ), .ZN(_05038_ ) );
AND4_X1 _12987_ ( .A1(_05029_ ), .A2(_05032_ ), .A3(_05035_ ), .A4(_05038_ ), .ZN(_05039_ ) );
OAI21_X1 _12988_ ( .A(_05026_ ), .B1(_04629_ ), .B2(_04630_ ), .ZN(_05040_ ) );
NAND2_X1 _12989_ ( .A1(_01497_ ), .A2(fanout_net_8 ), .ZN(_05041_ ) );
NAND2_X1 _12990_ ( .A1(_05040_ ), .A2(_05041_ ), .ZN(_05042_ ) );
NAND3_X1 _12991_ ( .A1(_04504_ ), .A2(_05026_ ), .A3(_04523_ ), .ZN(_05043_ ) );
NAND2_X1 _12992_ ( .A1(_01473_ ), .A2(fanout_net_8 ), .ZN(_05044_ ) );
NAND2_X1 _12993_ ( .A1(_05043_ ), .A2(_05044_ ), .ZN(_05045_ ) );
NAND3_X1 _12994_ ( .A1(_04684_ ), .A2(_04703_ ), .A3(_05026_ ), .ZN(_05046_ ) );
NAND2_X1 _12995_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [22] ), .ZN(_05047_ ) );
AND2_X2 _12996_ ( .A1(_05046_ ), .A2(_05047_ ), .ZN(_05048_ ) );
NAND3_X1 _12997_ ( .A1(_04573_ ), .A2(_02375_ ), .A3(_04592_ ), .ZN(_05049_ ) );
NAND2_X1 _12998_ ( .A1(_02185_ ), .A2(fanout_net_8 ), .ZN(_05050_ ) );
NAND2_X2 _12999_ ( .A1(_05049_ ), .A2(_05050_ ), .ZN(_05051_ ) );
NAND4_X1 _13000_ ( .A1(_05042_ ), .A2(_05045_ ), .A3(_05048_ ), .A4(_05051_ ), .ZN(_05052_ ) );
NAND2_X1 _13001_ ( .A1(_03935_ ), .A2(_02376_ ), .ZN(_05053_ ) );
OR2_X1 _13002_ ( .A1(_05026_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05054_ ) );
NAND2_X1 _13003_ ( .A1(_05053_ ), .A2(_05054_ ), .ZN(_05055_ ) );
NAND2_X1 _13004_ ( .A1(_04488_ ), .A2(_02376_ ), .ZN(_05056_ ) );
OR2_X1 _13005_ ( .A1(_05026_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05057_ ) );
NAND2_X1 _13006_ ( .A1(_05056_ ), .A2(_05057_ ), .ZN(_05058_ ) );
NAND2_X1 _13007_ ( .A1(_04382_ ), .A2(_02376_ ), .ZN(_05059_ ) );
NAND2_X1 _13008_ ( .A1(_02242_ ), .A2(fanout_net_8 ), .ZN(_05060_ ) );
NAND2_X1 _13009_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [23] ), .ZN(_05061_ ) );
NAND3_X1 _13010_ ( .A1(_04648_ ), .A2(_02376_ ), .A3(_04667_ ), .ZN(_05062_ ) );
NAND4_X1 _13011_ ( .A1(_05059_ ), .A2(_05060_ ), .A3(_05061_ ), .A4(_05062_ ), .ZN(_05063_ ) );
NOR4_X1 _13012_ ( .A1(_05052_ ), .A2(_05055_ ), .A3(_05058_ ), .A4(_05063_ ), .ZN(_05064_ ) );
NAND2_X1 _13013_ ( .A1(_03524_ ), .A2(_02376_ ), .ZN(_05065_ ) );
NAND2_X1 _13014_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [21] ), .ZN(_05066_ ) );
AND2_X2 _13015_ ( .A1(_05065_ ), .A2(_05066_ ), .ZN(_05067_ ) );
NAND2_X1 _13016_ ( .A1(_04741_ ), .A2(_05026_ ), .ZN(_05068_ ) );
NAND2_X1 _13017_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [31] ), .ZN(_05069_ ) );
AND2_X1 _13018_ ( .A1(_05068_ ), .A2(_05069_ ), .ZN(_05070_ ) );
NAND3_X1 _13019_ ( .A1(_03555_ ), .A2(_03588_ ), .A3(_05026_ ), .ZN(_05071_ ) );
NAND2_X1 _13020_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [20] ), .ZN(_05072_ ) );
AND2_X2 _13021_ ( .A1(_05071_ ), .A2(_05072_ ), .ZN(_05073_ ) );
NAND3_X1 _13022_ ( .A1(_03614_ ), .A2(_02375_ ), .A3(_03637_ ), .ZN(_05074_ ) );
NAND2_X1 _13023_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [19] ), .ZN(_05075_ ) );
AND2_X1 _13024_ ( .A1(_05074_ ), .A2(_05075_ ), .ZN(_05076_ ) );
AND4_X1 _13025_ ( .A1(_05067_ ), .A2(_05070_ ), .A3(_05073_ ), .A4(_05076_ ), .ZN(_05077_ ) );
NAND2_X1 _13026_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [15] ), .ZN(_05078_ ) );
NAND3_X2 _13027_ ( .A1(_03778_ ), .A2(_02375_ ), .A3(_03801_ ), .ZN(_05079_ ) );
NAND3_X1 _13028_ ( .A1(_03818_ ), .A2(_03837_ ), .A3(_02375_ ), .ZN(_05080_ ) );
NAND2_X1 _13029_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [14] ), .ZN(_05081_ ) );
AND4_X1 _13030_ ( .A1(_05078_ ), .A2(_05079_ ), .A3(_05080_ ), .A4(_05081_ ), .ZN(_05082_ ) );
NAND3_X2 _13031_ ( .A1(_03853_ ), .A2(_02374_ ), .A3(_03875_ ), .ZN(_05083_ ) );
NAND2_X1 _13032_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [13] ), .ZN(_05084_ ) );
AND2_X4 _13033_ ( .A1(_05083_ ), .A2(_05084_ ), .ZN(_05085_ ) );
NAND3_X1 _13034_ ( .A1(_03892_ ), .A2(_03912_ ), .A3(_02374_ ), .ZN(_05086_ ) );
NAND2_X1 _13035_ ( .A1(\ID_EX_typ [4] ), .A2(\ID_EX_imm [12] ), .ZN(_05087_ ) );
AND2_X2 _13036_ ( .A1(_05086_ ), .A2(_05087_ ), .ZN(_05088_ ) );
AND3_X1 _13037_ ( .A1(_05082_ ), .A2(_05085_ ), .A3(_05088_ ), .ZN(_05089_ ) );
AND4_X1 _13038_ ( .A1(_05039_ ), .A2(_05064_ ), .A3(_05077_ ), .A4(_05089_ ), .ZN(_05090_ ) );
NAND4_X1 _13039_ ( .A1(_05014_ ), .A2(_05022_ ), .A3(_05025_ ), .A4(_05090_ ), .ZN(_05091_ ) );
NOR4_X1 _13040_ ( .A1(_05042_ ), .A2(_05032_ ), .A3(_05038_ ), .A4(_05051_ ), .ZN(_05092_ ) );
INV_X1 _13041_ ( .A(_05045_ ), .ZN(_05093_ ) );
INV_X1 _13042_ ( .A(_05048_ ), .ZN(_05094_ ) );
AOI22_X1 _13043_ ( .A1(_05059_ ), .A2(_05060_ ), .B1(_05061_ ), .B2(_05062_ ), .ZN(_05095_ ) );
NAND4_X1 _13044_ ( .A1(_05092_ ), .A2(_05093_ ), .A3(_05094_ ), .A4(_05095_ ), .ZN(_05096_ ) );
AOI22_X1 _13045_ ( .A1(_05021_ ), .A2(_05020_ ), .B1(_05023_ ), .B2(_05024_ ), .ZN(_05097_ ) );
NAND3_X1 _13046_ ( .A1(_05058_ ), .A2(_05055_ ), .A3(_05097_ ), .ZN(_05098_ ) );
AND2_X2 _13047_ ( .A1(_05079_ ), .A2(_05078_ ), .ZN(_05099_ ) );
AND2_X4 _13048_ ( .A1(_05080_ ), .A2(_05081_ ), .ZN(_05100_ ) );
OR4_X1 _13049_ ( .A1(_05099_ ), .A2(_05100_ ), .A3(_05085_ ), .A4(_05088_ ), .ZN(_05101_ ) );
NOR3_X1 _13050_ ( .A1(_05096_ ), .A2(_05098_ ), .A3(_05101_ ), .ZN(_05102_ ) );
AOI22_X1 _13051_ ( .A1(_05068_ ), .A2(_05069_ ), .B1(_05075_ ), .B2(_05074_ ), .ZN(_05103_ ) );
NOR4_X1 _13052_ ( .A1(_05067_ ), .A2(_05073_ ), .A3(_05029_ ), .A4(_05035_ ), .ZN(_05104_ ) );
NAND3_X1 _13053_ ( .A1(_05102_ ), .A2(_05103_ ), .A3(_05104_ ), .ZN(_05105_ ) );
OAI21_X2 _13054_ ( .A(_05091_ ), .B1(_05014_ ), .B2(_05105_ ), .ZN(_05106_ ) );
AND2_X4 _13055_ ( .A1(_05019_ ), .A2(_05106_ ), .ZN(_05107_ ) );
BUF_X8 _13056_ ( .A(_05107_ ), .Z(_05108_ ) );
INV_X8 _13057_ ( .A(_05108_ ), .ZN(_05109_ ) );
BUF_X4 _13058_ ( .A(_04973_ ), .Z(_05110_ ) );
BUF_X2 _13059_ ( .A(_04976_ ), .Z(_05111_ ) );
XOR2_X1 _13060_ ( .A(_05110_ ), .B(_05111_ ), .Z(_05112_ ) );
BUF_X4 _13061_ ( .A(_04981_ ), .Z(_05113_ ) );
AND2_X1 _13062_ ( .A1(_05112_ ), .A2(_05113_ ), .ZN(_05114_ ) );
XNOR2_X1 _13063_ ( .A(_04982_ ), .B(_04985_ ), .ZN(_05115_ ) );
BUF_X2 _13064_ ( .A(_05115_ ), .Z(_05116_ ) );
NOR3_X1 _13065_ ( .A1(_05109_ ), .A2(_05114_ ), .A3(_05116_ ), .ZN(_05117_ ) );
XNOR2_X1 _13066_ ( .A(_04987_ ), .B(_04990_ ), .ZN(_05118_ ) );
BUF_X2 _13067_ ( .A(_05118_ ), .Z(_05119_ ) );
XNOR2_X1 _13068_ ( .A(_04991_ ), .B(_04994_ ), .ZN(_05120_ ) );
AND2_X1 _13069_ ( .A1(_05107_ ), .A2(_05120_ ), .ZN(_05121_ ) );
BUF_X4 _13070_ ( .A(_05121_ ), .Z(_05122_ ) );
NOR2_X1 _13071_ ( .A1(_05118_ ), .A2(_04994_ ), .ZN(_05123_ ) );
OAI22_X1 _13072_ ( .A1(_05117_ ), .A2(_05119_ ), .B1(_05122_ ), .B2(_05123_ ), .ZN(_05124_ ) );
INV_X2 _13073_ ( .A(_04981_ ), .ZN(_05125_ ) );
NAND2_X1 _13074_ ( .A1(_04973_ ), .A2(_04348_ ), .ZN(_05126_ ) );
BUF_X2 _13075_ ( .A(_04976_ ), .Z(_05127_ ) );
CLKBUF_X2 _13076_ ( .A(_04971_ ), .Z(_05128_ ) );
BUF_X2 _13077_ ( .A(_05128_ ), .Z(_05129_ ) );
CLKBUF_X2 _13078_ ( .A(_04972_ ), .Z(_05130_ ) );
BUF_X2 _13079_ ( .A(_05130_ ), .Z(_05131_ ) );
NAND3_X1 _13080_ ( .A1(_05129_ ), .A2(_01446_ ), .A3(_05131_ ), .ZN(_05132_ ) );
NAND3_X1 _13081_ ( .A1(_05126_ ), .A2(_05127_ ), .A3(_05132_ ), .ZN(_05133_ ) );
INV_X2 _13082_ ( .A(_04976_ ), .ZN(_05134_ ) );
NAND3_X1 _13083_ ( .A1(_05134_ ), .A2(_02268_ ), .A3(_04973_ ), .ZN(_05135_ ) );
AOI21_X1 _13084_ ( .A(_05125_ ), .B1(_05133_ ), .B2(_05135_ ), .ZN(_05136_ ) );
INV_X1 _13085_ ( .A(_02182_ ), .ZN(_05137_ ) );
AND3_X1 _13086_ ( .A1(_05128_ ), .A2(_05137_ ), .A3(_05130_ ), .ZN(_05138_ ) );
AOI21_X1 _13087_ ( .A(_02158_ ), .B1(_05128_ ), .B2(_05130_ ), .ZN(_05139_ ) );
NOR3_X1 _13088_ ( .A1(_05138_ ), .A2(_05134_ ), .A3(_05139_ ), .ZN(_05140_ ) );
AND3_X1 _13089_ ( .A1(_05128_ ), .A2(_02308_ ), .A3(_05130_ ), .ZN(_05141_ ) );
BUF_X2 _13090_ ( .A(_04971_ ), .Z(_05142_ ) );
BUF_X2 _13091_ ( .A(_04972_ ), .Z(_05143_ ) );
AOI21_X1 _13092_ ( .A(_01472_ ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_05144_ ) );
NOR3_X1 _13093_ ( .A1(_05141_ ), .A2(_05144_ ), .A3(_04976_ ), .ZN(_05145_ ) );
OAI21_X1 _13094_ ( .A(_05125_ ), .B1(_05140_ ), .B2(_05145_ ), .ZN(_05146_ ) );
INV_X1 _13095_ ( .A(_02064_ ), .ZN(_05147_ ) );
AND3_X1 _13096_ ( .A1(_05128_ ), .A2(_05147_ ), .A3(_05130_ ), .ZN(_05148_ ) );
AOI21_X1 _13097_ ( .A(_03472_ ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_05149_ ) );
OAI21_X1 _13098_ ( .A(_05127_ ), .B1(_05148_ ), .B2(_05149_ ), .ZN(_05150_ ) );
INV_X1 _13099_ ( .A(_01496_ ), .ZN(_05151_ ) );
AND3_X1 _13100_ ( .A1(_05128_ ), .A2(_05151_ ), .A3(_05130_ ), .ZN(_05152_ ) );
AOI21_X1 _13101_ ( .A(_02042_ ), .B1(_05128_ ), .B2(_05130_ ), .ZN(_05153_ ) );
OAI21_X1 _13102_ ( .A(_05134_ ), .B1(_05152_ ), .B2(_05153_ ), .ZN(_05154_ ) );
NAND3_X1 _13103_ ( .A1(_05150_ ), .A2(_05154_ ), .A3(_04981_ ), .ZN(_05155_ ) );
NAND2_X1 _13104_ ( .A1(_05146_ ), .A2(_05155_ ), .ZN(_05156_ ) );
MUX2_X1 _13105_ ( .A(_05136_ ), .B(_05156_ ), .S(_04986_ ), .Z(_05157_ ) );
BUF_X2 _13106_ ( .A(_04990_ ), .Z(_05158_ ) );
BUF_X2 _13107_ ( .A(_05158_ ), .Z(_05159_ ) );
NAND2_X1 _13108_ ( .A1(_05157_ ), .A2(_05159_ ), .ZN(_05160_ ) );
AOI21_X1 _13109_ ( .A(_04970_ ), .B1(_05124_ ), .B2(_05160_ ), .ZN(_05161_ ) );
NOR2_X1 _13110_ ( .A1(_01349_ ), .A2(\ID_EX_typ [1] ), .ZN(_05162_ ) );
AND2_X1 _13111_ ( .A1(_05162_ ), .A2(fanout_net_7 ), .ZN(_05163_ ) );
INV_X1 _13112_ ( .A(_05163_ ), .ZN(_05164_ ) );
BUF_X2 _13113_ ( .A(_05158_ ), .Z(_05165_ ) );
AND3_X1 _13114_ ( .A1(_05129_ ), .A2(_04779_ ), .A3(_05131_ ), .ZN(_05166_ ) );
BUF_X2 _13115_ ( .A(_05134_ ), .Z(_05167_ ) );
BUF_X2 _13116_ ( .A(_05167_ ), .Z(_05168_ ) );
CLKBUF_X2 _13117_ ( .A(_05128_ ), .Z(_05169_ ) );
CLKBUF_X2 _13118_ ( .A(_05130_ ), .Z(_05170_ ) );
AOI21_X1 _13119_ ( .A(_01854_ ), .B1(_05169_ ), .B2(_05170_ ), .ZN(_05171_ ) );
NOR3_X1 _13120_ ( .A1(_05166_ ), .A2(_05168_ ), .A3(_05171_ ), .ZN(_05172_ ) );
BUF_X2 _13121_ ( .A(_04971_ ), .Z(_05173_ ) );
BUF_X2 _13122_ ( .A(_04972_ ), .Z(_05174_ ) );
AND3_X1 _13123_ ( .A1(_05173_ ), .A2(_04799_ ), .A3(_05174_ ), .ZN(_05175_ ) );
AOI21_X1 _13124_ ( .A(_01684_ ), .B1(_05129_ ), .B2(_05131_ ), .ZN(_05176_ ) );
BUF_X2 _13125_ ( .A(_05111_ ), .Z(_05177_ ) );
NOR3_X1 _13126_ ( .A1(_05175_ ), .A2(_05176_ ), .A3(_05177_ ), .ZN(_05178_ ) );
NOR2_X1 _13127_ ( .A1(_05172_ ), .A2(_05178_ ), .ZN(_05179_ ) );
BUF_X4 _13128_ ( .A(_05113_ ), .Z(_05180_ ) );
NOR2_X1 _13129_ ( .A1(_05179_ ), .A2(_05180_ ), .ZN(_05181_ ) );
BUF_X4 _13130_ ( .A(_05125_ ), .Z(_05182_ ) );
AND3_X1 _13131_ ( .A1(_05129_ ), .A2(_04774_ ), .A3(_05131_ ), .ZN(_05183_ ) );
BUF_X2 _13132_ ( .A(_05127_ ), .Z(_05184_ ) );
AOI21_X1 _13133_ ( .A(_04771_ ), .B1(_05169_ ), .B2(_05170_ ), .ZN(_05185_ ) );
OR3_X1 _13134_ ( .A1(_05183_ ), .A2(_05184_ ), .A3(_05185_ ), .ZN(_05186_ ) );
AOI21_X1 _13135_ ( .A(_03850_ ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_05187_ ) );
INV_X1 _13136_ ( .A(_05187_ ), .ZN(_05188_ ) );
BUF_X4 _13137_ ( .A(_05110_ ), .Z(_05189_ ) );
OAI211_X1 _13138_ ( .A(_05188_ ), .B(_05177_ ), .C1(_01808_ ), .C2(_05189_ ), .ZN(_05190_ ) );
AOI21_X1 _13139_ ( .A(_05182_ ), .B1(_05186_ ), .B2(_05190_ ), .ZN(_05191_ ) );
NOR2_X1 _13140_ ( .A1(_05181_ ), .A2(_05191_ ), .ZN(_05192_ ) );
BUF_X2 _13141_ ( .A(_04986_ ), .Z(_05193_ ) );
BUF_X4 _13142_ ( .A(_05193_ ), .Z(_05194_ ) );
NOR2_X1 _13143_ ( .A1(_05192_ ), .A2(_05194_ ), .ZN(_05195_ ) );
AND3_X1 _13144_ ( .A1(_05128_ ), .A2(_04855_ ), .A3(_05130_ ), .ZN(_05196_ ) );
BUF_X4 _13145_ ( .A(_05134_ ), .Z(_05197_ ) );
NOR3_X1 _13146_ ( .A1(_05196_ ), .A2(_05197_ ), .A3(_05149_ ), .ZN(_05198_ ) );
AND3_X1 _13147_ ( .A1(_05128_ ), .A2(_02123_ ), .A3(_05130_ ), .ZN(_05199_ ) );
AOI21_X1 _13148_ ( .A(_04835_ ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_05200_ ) );
NOR3_X1 _13149_ ( .A1(_05199_ ), .A2(_05200_ ), .A3(_05184_ ), .ZN(_05201_ ) );
BUF_X4 _13150_ ( .A(_05125_ ), .Z(_05202_ ) );
OR3_X1 _13151_ ( .A1(_05198_ ), .A2(_05201_ ), .A3(_05202_ ), .ZN(_05203_ ) );
AOI21_X1 _13152_ ( .A(_01760_ ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_05204_ ) );
INV_X1 _13153_ ( .A(_05204_ ), .ZN(_05205_ ) );
OAI211_X1 _13154_ ( .A(_05205_ ), .B(_05168_ ), .C1(_01738_ ), .C2(_05189_ ), .ZN(_05206_ ) );
AOI21_X1 _13155_ ( .A(_01945_ ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_05207_ ) );
INV_X1 _13156_ ( .A(_05207_ ), .ZN(_05208_ ) );
OAI211_X1 _13157_ ( .A(_05208_ ), .B(_05177_ ), .C1(_01969_ ), .C2(_05189_ ), .ZN(_05209_ ) );
NAND3_X1 _13158_ ( .A1(_05206_ ), .A2(_05209_ ), .A3(_05182_ ), .ZN(_05210_ ) );
AND3_X1 _13159_ ( .A1(_05203_ ), .A2(_05193_ ), .A3(_05210_ ), .ZN(_05211_ ) );
OAI21_X1 _13160_ ( .A(_05165_ ), .B1(_05195_ ), .B2(_05211_ ), .ZN(_05212_ ) );
BUF_X2 _13161_ ( .A(_05111_ ), .Z(_05213_ ) );
BUF_X2 _13162_ ( .A(_05129_ ), .Z(_05214_ ) );
BUF_X2 _13163_ ( .A(_05131_ ), .Z(_05215_ ) );
AND3_X1 _13164_ ( .A1(_05214_ ), .A2(_04239_ ), .A3(_05215_ ), .ZN(_05216_ ) );
AOI21_X1 _13165_ ( .A(_01657_ ), .B1(_05129_ ), .B2(_05131_ ), .ZN(_05217_ ) );
OAI21_X1 _13166_ ( .A(_05213_ ), .B1(_05216_ ), .B2(_05217_ ), .ZN(_05218_ ) );
BUF_X4 _13167_ ( .A(_05197_ ), .Z(_05219_ ) );
AND3_X1 _13168_ ( .A1(_05214_ ), .A2(_04787_ ), .A3(_05215_ ), .ZN(_05220_ ) );
AOI21_X1 _13169_ ( .A(_01521_ ), .B1(_05214_ ), .B2(_05215_ ), .ZN(_05221_ ) );
OAI21_X1 _13170_ ( .A(_05219_ ), .B1(_05220_ ), .B2(_05221_ ), .ZN(_05222_ ) );
NAND2_X1 _13171_ ( .A1(_05218_ ), .A2(_05222_ ), .ZN(_05223_ ) );
NAND2_X1 _13172_ ( .A1(_05223_ ), .A2(_05180_ ), .ZN(_05224_ ) );
INV_X1 _13173_ ( .A(_03359_ ), .ZN(_05225_ ) );
AND3_X1 _13174_ ( .A1(_04971_ ), .A2(_05225_ ), .A3(_04972_ ), .ZN(_05226_ ) );
AOI21_X1 _13175_ ( .A(_01571_ ), .B1(_05214_ ), .B2(_05215_ ), .ZN(_05227_ ) );
NOR3_X1 _13176_ ( .A1(_05226_ ), .A2(_05168_ ), .A3(_05227_ ), .ZN(_05228_ ) );
BUF_X4 _13177_ ( .A(_05113_ ), .Z(_05229_ ) );
OR2_X1 _13178_ ( .A1(_05228_ ), .A2(_05229_ ), .ZN(_05230_ ) );
INV_X1 _13179_ ( .A(_04990_ ), .ZN(_05231_ ) );
BUF_X4 _13180_ ( .A(_05231_ ), .Z(_05232_ ) );
NAND4_X1 _13181_ ( .A1(_05224_ ), .A2(_05230_ ), .A3(_05194_ ), .A4(_05232_ ), .ZN(_05233_ ) );
AOI21_X1 _13182_ ( .A(_05164_ ), .B1(_05212_ ), .B2(_05233_ ), .ZN(_05234_ ) );
AND2_X2 _13183_ ( .A1(_04963_ ), .A2(fanout_net_7 ), .ZN(_05235_ ) );
AND3_X1 _13184_ ( .A1(_05157_ ), .A2(_05165_ ), .A3(_05235_ ), .ZN(_05236_ ) );
OR3_X1 _13185_ ( .A1(_05161_ ), .A2(_05234_ ), .A3(_05236_ ), .ZN(_05237_ ) );
OAI21_X1 _13186_ ( .A(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .B1(\ID_EX_typ [1] ), .B2(\ID_EX_typ [0] ), .ZN(_05238_ ) );
AND2_X2 _13187_ ( .A1(_05238_ ), .A2(_02379_ ), .ZN(_05239_ ) );
INV_X1 _13188_ ( .A(_05239_ ), .ZN(_05240_ ) );
XNOR2_X1 _13189_ ( .A(_05073_ ), .B(_02088_ ), .ZN(_05241_ ) );
INV_X1 _13190_ ( .A(_05241_ ), .ZN(_05242_ ) );
XNOR2_X2 _13191_ ( .A(_05085_ ), .B(_03850_ ), .ZN(_05243_ ) );
XNOR2_X2 _13192_ ( .A(_05088_ ), .B(_01808_ ), .ZN(_05244_ ) );
AND2_X1 _13193_ ( .A1(_05243_ ), .A2(_05244_ ), .ZN(_05245_ ) );
XNOR2_X2 _13194_ ( .A(_05099_ ), .B(_01760_ ), .ZN(_05246_ ) );
XNOR2_X1 _13195_ ( .A(_05100_ ), .B(_01738_ ), .ZN(_05247_ ) );
AND3_X4 _13196_ ( .A1(_05245_ ), .A2(_05246_ ), .A3(_05247_ ), .ZN(_05248_ ) );
INV_X1 _13197_ ( .A(_05248_ ), .ZN(_05249_ ) );
NOR2_X1 _13198_ ( .A1(_05022_ ), .A2(_04772_ ), .ZN(_05250_ ) );
NAND3_X1 _13199_ ( .A1(_05020_ ), .A2(_04772_ ), .A3(_05021_ ), .ZN(_05251_ ) );
NOR2_X1 _13200_ ( .A1(_05025_ ), .A2(_04774_ ), .ZN(_05252_ ) );
AOI21_X1 _13201_ ( .A(_05250_ ), .B1(_05251_ ), .B2(_05252_ ), .ZN(_05253_ ) );
XNOR2_X2 _13202_ ( .A(_05022_ ), .B(_04771_ ), .ZN(_05254_ ) );
XNOR2_X1 _13203_ ( .A(_05025_ ), .B(_01905_ ), .ZN(_05255_ ) );
AND2_X1 _13204_ ( .A1(_05254_ ), .A2(_05255_ ), .ZN(_05256_ ) );
NOR2_X1 _13205_ ( .A1(_05008_ ), .A2(_04777_ ), .ZN(_05257_ ) );
XNOR2_X1 _13206_ ( .A(_05008_ ), .B(_01854_ ), .ZN(_05258_ ) );
NOR2_X1 _13207_ ( .A1(_05011_ ), .A2(_04779_ ), .ZN(_05259_ ) );
AND2_X1 _13208_ ( .A1(_05258_ ), .A2(_05259_ ), .ZN(_05260_ ) );
OAI21_X1 _13209_ ( .A(_05256_ ), .B1(_05257_ ), .B2(_05260_ ), .ZN(_05261_ ) );
AOI21_X1 _13210_ ( .A(_05249_ ), .B1(_05253_ ), .B2(_05261_ ), .ZN(_05262_ ) );
NOR2_X1 _13211_ ( .A1(_05099_ ), .A2(_04766_ ), .ZN(_05263_ ) );
NOR2_X1 _13212_ ( .A1(_05088_ ), .A2(_04763_ ), .ZN(_05264_ ) );
AND2_X2 _13213_ ( .A1(_05243_ ), .A2(_05264_ ), .ZN(_05265_ ) );
INV_X1 _13214_ ( .A(_05085_ ), .ZN(_05266_ ) );
AOI21_X2 _13215_ ( .A(_05265_ ), .B1(_03850_ ), .B2(_05266_ ), .ZN(_05267_ ) );
INV_X1 _13216_ ( .A(_05246_ ), .ZN(_05268_ ) );
INV_X2 _13217_ ( .A(_05247_ ), .ZN(_05269_ ) );
NOR3_X1 _13218_ ( .A1(_05267_ ), .A2(_05268_ ), .A3(_05269_ ), .ZN(_05270_ ) );
NOR2_X1 _13219_ ( .A1(_05100_ ), .A2(_03814_ ), .ZN(_05271_ ) );
INV_X1 _13220_ ( .A(_05271_ ), .ZN(_05272_ ) );
AND3_X1 _13221_ ( .A1(_05079_ ), .A2(_04766_ ), .A3(_05078_ ), .ZN(_05273_ ) );
NOR3_X1 _13222_ ( .A1(_05272_ ), .A2(_05263_ ), .A3(_05273_ ), .ZN(_05274_ ) );
NOR4_X4 _13223_ ( .A1(_05262_ ), .A2(_05263_ ), .A3(_05270_ ), .A4(_05274_ ), .ZN(_05275_ ) );
XNOR2_X1 _13224_ ( .A(_05011_ ), .B(_01832_ ), .ZN(_05276_ ) );
AND2_X1 _13225_ ( .A1(_05258_ ), .A2(_05276_ ), .ZN(_05277_ ) );
AND2_X1 _13226_ ( .A1(_05256_ ), .A2(_05277_ ), .ZN(_05278_ ) );
NOR2_X1 _13227_ ( .A1(_04981_ ), .A2(_04787_ ), .ZN(_05279_ ) );
INV_X1 _13228_ ( .A(_05279_ ), .ZN(_05280_ ) );
AND3_X1 _13229_ ( .A1(_04974_ ), .A2(_04384_ ), .A3(_04975_ ), .ZN(_05281_ ) );
AOI21_X1 _13230_ ( .A(_04384_ ), .B1(_04975_ ), .B2(_04974_ ), .ZN(_05282_ ) );
NOR2_X2 _13231_ ( .A1(_05281_ ), .A2(_05282_ ), .ZN(_05283_ ) );
NOR2_X4 _13232_ ( .A1(_04973_ ), .A2(_05225_ ), .ZN(_05284_ ) );
AND2_X1 _13233_ ( .A1(_05283_ ), .A2(_05284_ ), .ZN(_05285_ ) );
NOR2_X2 _13234_ ( .A1(_05285_ ), .A2(_05282_ ), .ZN(_05286_ ) );
XNOR2_X1 _13235_ ( .A(_04981_ ), .B(_01547_ ), .ZN(_05287_ ) );
INV_X1 _13236_ ( .A(_05287_ ), .ZN(_05288_ ) );
OAI221_X1 _13237_ ( .A(_05280_ ), .B1(_01601_ ), .B2(_04986_ ), .C1(_05286_ ), .C2(_05288_ ), .ZN(_05289_ ) );
NOR2_X1 _13238_ ( .A1(_04985_ ), .A2(_01521_ ), .ZN(_05290_ ) );
INV_X1 _13239_ ( .A(_05290_ ), .ZN(_05291_ ) );
XNOR2_X1 _13240_ ( .A(_04999_ ), .B(_01684_ ), .ZN(_05292_ ) );
INV_X1 _13241_ ( .A(_01657_ ), .ZN(_05293_ ) );
XNOR2_X1 _13242_ ( .A(_04994_ ), .B(_05293_ ), .ZN(_05294_ ) );
XNOR2_X2 _13243_ ( .A(_05002_ ), .B(_01707_ ), .ZN(_05295_ ) );
XNOR2_X1 _13244_ ( .A(_04990_ ), .B(_03394_ ), .ZN(_05296_ ) );
AND4_X1 _13245_ ( .A1(_05292_ ), .A2(_05294_ ), .A3(_05295_ ), .A4(_05296_ ), .ZN(_05297_ ) );
AND3_X2 _13246_ ( .A1(_05289_ ), .A2(_05291_ ), .A3(_05297_ ), .ZN(_05298_ ) );
NOR2_X1 _13247_ ( .A1(_05002_ ), .A2(_04799_ ), .ZN(_05299_ ) );
NAND2_X1 _13248_ ( .A1(_05292_ ), .A2(_05299_ ), .ZN(_05300_ ) );
AND2_X1 _13249_ ( .A1(_05292_ ), .A2(_05295_ ), .ZN(_05301_ ) );
INV_X1 _13250_ ( .A(_05301_ ), .ZN(_05302_ ) );
AND2_X1 _13251_ ( .A1(_04994_ ), .A2(_01657_ ), .ZN(_05303_ ) );
NOR2_X1 _13252_ ( .A1(_04990_ ), .A2(_04239_ ), .ZN(_05304_ ) );
AOI21_X2 _13253_ ( .A(_05303_ ), .B1(_05294_ ), .B2(_05304_ ), .ZN(_05305_ ) );
OAI221_X2 _13254_ ( .A(_05300_ ), .B1(_04116_ ), .B2(_04999_ ), .C1(_05302_ ), .C2(_05305_ ), .ZN(_05306_ ) );
OAI211_X2 _13255_ ( .A(_05248_ ), .B(_05278_ ), .C1(_05298_ ), .C2(_05306_ ), .ZN(_05307_ ) );
AND2_X2 _13256_ ( .A1(_05275_ ), .A2(_05307_ ), .ZN(_05308_ ) );
XNOR2_X1 _13257_ ( .A(_05076_ ), .B(_04835_ ), .ZN(_05309_ ) );
XNOR2_X1 _13258_ ( .A(_05029_ ), .B(_02018_ ), .ZN(_05310_ ) );
AND2_X1 _13259_ ( .A1(_05309_ ), .A2(_05310_ ), .ZN(_05311_ ) );
XNOR2_X1 _13260_ ( .A(_05032_ ), .B(_01945_ ), .ZN(_05312_ ) );
XNOR2_X1 _13261_ ( .A(_05035_ ), .B(_01969_ ), .ZN(_05313_ ) );
AND2_X1 _13262_ ( .A1(_05312_ ), .A2(_05313_ ), .ZN(_05314_ ) );
NAND2_X1 _13263_ ( .A1(_05311_ ), .A2(_05314_ ), .ZN(_05315_ ) );
OR2_X4 _13264_ ( .A1(_05308_ ), .A2(_05315_ ), .ZN(_05316_ ) );
NOR2_X1 _13265_ ( .A1(_05032_ ), .A2(_04842_ ), .ZN(_05317_ ) );
NOR2_X1 _13266_ ( .A1(_05035_ ), .A2(_04840_ ), .ZN(_05318_ ) );
AOI21_X1 _13267_ ( .A(_05317_ ), .B1(_05312_ ), .B2(_05318_ ), .ZN(_05319_ ) );
INV_X1 _13268_ ( .A(_05319_ ), .ZN(_05320_ ) );
NAND2_X1 _13269_ ( .A1(_05320_ ), .A2(_05311_ ), .ZN(_05321_ ) );
OR2_X1 _13270_ ( .A1(_05076_ ), .A2(_04836_ ), .ZN(_05322_ ) );
NAND3_X1 _13271_ ( .A1(_05074_ ), .A2(_04836_ ), .A3(_05075_ ), .ZN(_05323_ ) );
NOR2_X1 _13272_ ( .A1(_05029_ ), .A2(_02123_ ), .ZN(_05324_ ) );
NAND3_X1 _13273_ ( .A1(_05322_ ), .A2(_05323_ ), .A3(_05324_ ), .ZN(_05325_ ) );
AND3_X1 _13274_ ( .A1(_05321_ ), .A2(_05322_ ), .A3(_05325_ ), .ZN(_05326_ ) );
AOI21_X1 _13275_ ( .A(_05242_ ), .B1(_05316_ ), .B2(_05326_ ), .ZN(_05327_ ) );
XNOR2_X1 _13276_ ( .A(_05067_ ), .B(_03472_ ), .ZN(_05328_ ) );
INV_X1 _13277_ ( .A(_05328_ ), .ZN(_05329_ ) );
NOR2_X1 _13278_ ( .A1(_05073_ ), .A2(_04855_ ), .ZN(_05330_ ) );
OR3_X1 _13279_ ( .A1(_05327_ ), .A2(_05329_ ), .A3(_05330_ ), .ZN(_05331_ ) );
OAI21_X1 _13280_ ( .A(_05329_ ), .B1(_05327_ ), .B2(_05330_ ), .ZN(_05332_ ) );
AOI21_X1 _13281_ ( .A(_05240_ ), .B1(_05331_ ), .B2(_05332_ ), .ZN(_05333_ ) );
AND2_X1 _13282_ ( .A1(_04968_ ), .A2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .ZN(_05334_ ) );
BUF_X2 _13283_ ( .A(_05334_ ), .Z(_05335_ ) );
AND2_X1 _13284_ ( .A1(_05328_ ), .A2(_05335_ ), .ZN(_05336_ ) );
INV_X1 _13285_ ( .A(_03472_ ), .ZN(_05337_ ) );
AND2_X1 _13286_ ( .A1(_05162_ ), .A2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .ZN(_05338_ ) );
INV_X1 _13287_ ( .A(_05338_ ), .ZN(_05339_ ) );
BUF_X2 _13288_ ( .A(_05339_ ), .Z(_05340_ ) );
NOR3_X1 _13289_ ( .A1(_05067_ ), .A2(_05337_ ), .A3(_05340_ ), .ZN(_05341_ ) );
AND2_X1 _13290_ ( .A1(_04963_ ), .A2(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ), .ZN(_05342_ ) );
INV_X1 _13291_ ( .A(_05342_ ), .ZN(_05343_ ) );
BUF_X4 _13292_ ( .A(_05343_ ), .Z(_05344_ ) );
AOI21_X1 _13293_ ( .A(_05344_ ), .B1(_05067_ ), .B2(_05337_ ), .ZN(_05345_ ) );
OR3_X1 _13294_ ( .A1(_05336_ ), .A2(_05341_ ), .A3(_05345_ ), .ZN(_05346_ ) );
NOR3_X1 _13295_ ( .A1(_05237_ ), .A2(_05333_ ), .A3(_05346_ ), .ZN(_05347_ ) );
AND2_X1 _13296_ ( .A1(_04961_ ), .A2(_04963_ ), .ZN(_05348_ ) );
NOR3_X1 _13297_ ( .A1(_04865_ ), .A2(_05348_ ), .A3(_04954_ ), .ZN(_05349_ ) );
NOR2_X1 _13298_ ( .A1(_02377_ ), .A2(\ID_EX_typ [2] ), .ZN(_05350_ ) );
NAND3_X1 _13299_ ( .A1(_05162_ ), .A2(_05350_ ), .A3(_02376_ ), .ZN(_05351_ ) );
NAND4_X1 _13300_ ( .A1(_04863_ ), .A2(\ID_EX_typ [4] ), .A3(\ID_EX_typ [3] ), .A4(_02378_ ), .ZN(_05352_ ) );
AND2_X1 _13301_ ( .A1(_05351_ ), .A2(_05352_ ), .ZN(_05353_ ) );
AND2_X1 _13302_ ( .A1(_05349_ ), .A2(_05353_ ), .ZN(_05354_ ) );
INV_X1 _13303_ ( .A(_04758_ ), .ZN(_05355_ ) );
NOR2_X1 _13304_ ( .A1(_05354_ ), .A2(_05355_ ), .ZN(_05356_ ) );
BUF_X4 _13305_ ( .A(_05356_ ), .Z(_05357_ ) );
OAI21_X1 _13306_ ( .A(_04967_ ), .B1(_05347_ ), .B2(_05357_ ), .ZN(_05358_ ) );
INV_X1 _13307_ ( .A(_01361_ ), .ZN(_05359_ ) );
BUF_X4 _13308_ ( .A(_05359_ ), .Z(_05360_ ) );
MUX2_X1 _13309_ ( .A(_04757_ ), .B(_05358_ ), .S(_05360_ ), .Z(_05361_ ) );
MUX2_X1 _13310_ ( .A(_04743_ ), .B(_05361_ ), .S(_03390_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
CLKBUF_X2 _13311_ ( .A(_03356_ ), .Z(_05362_ ) );
OR2_X1 _13312_ ( .A1(_03545_ ), .A2(_05362_ ), .ZN(_05363_ ) );
INV_X1 _13313_ ( .A(_05356_ ), .ZN(_05364_ ) );
BUF_X2 _13314_ ( .A(_05364_ ), .Z(_05365_ ) );
BUF_X4 _13315_ ( .A(_04969_ ), .Z(_05366_ ) );
INV_X1 _13316_ ( .A(_05116_ ), .ZN(_05367_ ) );
BUF_X2 _13317_ ( .A(_05367_ ), .Z(_05368_ ) );
BUF_X4 _13318_ ( .A(_05229_ ), .Z(_05369_ ) );
BUF_X4 _13319_ ( .A(_05369_ ), .Z(_05370_ ) );
INV_X1 _13320_ ( .A(_04973_ ), .ZN(_05371_ ) );
BUF_X4 _13321_ ( .A(_05219_ ), .Z(_05372_ ) );
OAI21_X1 _13322_ ( .A(_05370_ ), .B1(_05371_ ), .B2(_05372_ ), .ZN(_05373_ ) );
AND3_X1 _13323_ ( .A1(_05108_ ), .A2(_05368_ ), .A3(_05373_ ), .ZN(_05374_ ) );
INV_X1 _13324_ ( .A(_05374_ ), .ZN(_05375_ ) );
INV_X1 _13325_ ( .A(_05118_ ), .ZN(_05376_ ) );
INV_X1 _13326_ ( .A(_05123_ ), .ZN(_05377_ ) );
INV_X1 _13327_ ( .A(_05122_ ), .ZN(_05378_ ) );
AOI22_X1 _13328_ ( .A1(_05375_ ), .A2(_05376_ ), .B1(_05377_ ), .B2(_05378_ ), .ZN(_05379_ ) );
BUF_X4 _13329_ ( .A(_05232_ ), .Z(_05380_ ) );
BUF_X4 _13330_ ( .A(_05380_ ), .Z(_05381_ ) );
AND3_X1 _13331_ ( .A1(_05142_ ), .A2(_05337_ ), .A3(_05143_ ), .ZN(_05382_ ) );
AOI21_X1 _13332_ ( .A(_02088_ ), .B1(_05142_ ), .B2(_05143_ ), .ZN(_05383_ ) );
NOR3_X1 _13333_ ( .A1(_05382_ ), .A2(_05167_ ), .A3(_05383_ ), .ZN(_05384_ ) );
INV_X1 _13334_ ( .A(_02042_ ), .ZN(_05385_ ) );
AND3_X1 _13335_ ( .A1(_05169_ ), .A2(_05385_ ), .A3(_05170_ ), .ZN(_05386_ ) );
AOI21_X1 _13336_ ( .A(_02064_ ), .B1(_05173_ ), .B2(_05174_ ), .ZN(_05387_ ) );
NOR3_X1 _13337_ ( .A1(_05386_ ), .A2(_05387_ ), .A3(_05111_ ), .ZN(_05388_ ) );
NOR2_X1 _13338_ ( .A1(_05384_ ), .A2(_05388_ ), .ZN(_05389_ ) );
NAND2_X1 _13339_ ( .A1(_05389_ ), .A2(_05369_ ), .ZN(_05390_ ) );
INV_X1 _13340_ ( .A(_02158_ ), .ZN(_05391_ ) );
AND3_X1 _13341_ ( .A1(_05142_ ), .A2(_05391_ ), .A3(_05143_ ), .ZN(_05392_ ) );
AOI21_X1 _13342_ ( .A(_01496_ ), .B1(_05173_ ), .B2(_05174_ ), .ZN(_05393_ ) );
OAI21_X1 _13343_ ( .A(_05184_ ), .B1(_05392_ ), .B2(_05393_ ), .ZN(_05394_ ) );
AND3_X1 _13344_ ( .A1(_05173_ ), .A2(_04490_ ), .A3(_05174_ ), .ZN(_05395_ ) );
AOI21_X1 _13345_ ( .A(_02182_ ), .B1(_05173_ ), .B2(_05174_ ), .ZN(_05396_ ) );
OAI21_X1 _13346_ ( .A(_05197_ ), .B1(_05395_ ), .B2(_05396_ ), .ZN(_05397_ ) );
NAND2_X1 _13347_ ( .A1(_05394_ ), .A2(_05397_ ), .ZN(_05398_ ) );
BUF_X4 _13348_ ( .A(_05202_ ), .Z(_05399_ ) );
NAND2_X1 _13349_ ( .A1(_05398_ ), .A2(_05399_ ), .ZN(_05400_ ) );
NAND3_X1 _13350_ ( .A1(_05390_ ), .A2(_05194_ ), .A3(_05400_ ), .ZN(_05401_ ) );
AND3_X1 _13351_ ( .A1(_05173_ ), .A2(_04348_ ), .A3(_05174_ ), .ZN(_05402_ ) );
AOI21_X1 _13352_ ( .A(_02236_ ), .B1(_05173_ ), .B2(_05174_ ), .ZN(_05403_ ) );
NOR2_X1 _13353_ ( .A1(_05402_ ), .A2(_05403_ ), .ZN(_05404_ ) );
AOI21_X1 _13354_ ( .A(_03949_ ), .B1(_05173_ ), .B2(_05174_ ), .ZN(_05405_ ) );
AOI21_X1 _13355_ ( .A(_05405_ ), .B1(_04707_ ), .B2(_05371_ ), .ZN(_05406_ ) );
MUX2_X1 _13356_ ( .A(_05404_ ), .B(_05406_ ), .S(_05167_ ), .Z(_05407_ ) );
BUF_X4 _13357_ ( .A(_04985_ ), .Z(_05408_ ) );
BUF_X4 _13358_ ( .A(_05408_ ), .Z(_05409_ ) );
NAND3_X1 _13359_ ( .A1(_05407_ ), .A2(_05409_ ), .A3(_05370_ ), .ZN(_05410_ ) );
AOI21_X1 _13360_ ( .A(_05381_ ), .B1(_05401_ ), .B2(_05410_ ), .ZN(_05411_ ) );
OAI21_X1 _13361_ ( .A(_05366_ ), .B1(_05379_ ), .B2(_05411_ ), .ZN(_05412_ ) );
BUF_X2 _13362_ ( .A(_05163_ ), .Z(_05413_ ) );
AND3_X1 _13363_ ( .A1(_04116_ ), .A2(_05169_ ), .A3(_05170_ ), .ZN(_05414_ ) );
BUF_X2 _13364_ ( .A(_05168_ ), .Z(_05415_ ) );
AOI21_X1 _13365_ ( .A(_01832_ ), .B1(_05214_ ), .B2(_05215_ ), .ZN(_05416_ ) );
NOR3_X1 _13366_ ( .A1(_05414_ ), .A2(_05415_ ), .A3(_05416_ ), .ZN(_05417_ ) );
AND3_X1 _13367_ ( .A1(_05293_ ), .A2(_05169_ ), .A3(_05170_ ), .ZN(_05418_ ) );
AOI21_X1 _13368_ ( .A(_01707_ ), .B1(_05214_ ), .B2(_05215_ ), .ZN(_05419_ ) );
BUF_X2 _13369_ ( .A(_05184_ ), .Z(_05420_ ) );
NOR3_X1 _13370_ ( .A1(_05418_ ), .A2(_05419_ ), .A3(_05420_ ), .ZN(_05421_ ) );
NOR2_X1 _13371_ ( .A1(_05417_ ), .A2(_05421_ ), .ZN(_05422_ ) );
BUF_X4 _13372_ ( .A(_05180_ ), .Z(_05423_ ) );
NOR2_X1 _13373_ ( .A1(_05422_ ), .A2(_05423_ ), .ZN(_05424_ ) );
BUF_X2 _13374_ ( .A(_05193_ ), .Z(_05425_ ) );
BUF_X2 _13375_ ( .A(_05425_ ), .Z(_05426_ ) );
BUF_X2 _13376_ ( .A(_05426_ ), .Z(_05427_ ) );
BUF_X4 _13377_ ( .A(_05182_ ), .Z(_05428_ ) );
AND3_X1 _13378_ ( .A1(_05169_ ), .A2(_04772_ ), .A3(_05170_ ), .ZN(_05429_ ) );
AOI21_X1 _13379_ ( .A(_01808_ ), .B1(_05169_ ), .B2(_05170_ ), .ZN(_05430_ ) );
OR3_X1 _13380_ ( .A1(_05429_ ), .A2(_05219_ ), .A3(_05430_ ), .ZN(_05431_ ) );
AND3_X1 _13381_ ( .A1(_05169_ ), .A2(_04777_ ), .A3(_05170_ ), .ZN(_05432_ ) );
AOI21_X1 _13382_ ( .A(_01905_ ), .B1(_05214_ ), .B2(_05215_ ), .ZN(_05433_ ) );
OR3_X1 _13383_ ( .A1(_05432_ ), .A2(_05433_ ), .A3(_05213_ ), .ZN(_05434_ ) );
AOI21_X1 _13384_ ( .A(_05428_ ), .B1(_05431_ ), .B2(_05434_ ), .ZN(_05435_ ) );
NOR3_X1 _13385_ ( .A1(_05424_ ), .A2(_05427_ ), .A3(_05435_ ), .ZN(_05436_ ) );
NOR2_X1 _13386_ ( .A1(_05110_ ), .A2(_03850_ ), .ZN(_05437_ ) );
AOI21_X1 _13387_ ( .A(_01738_ ), .B1(_05129_ ), .B2(_05131_ ), .ZN(_05438_ ) );
OR3_X1 _13388_ ( .A1(_05437_ ), .A2(_05420_ ), .A3(_05438_ ), .ZN(_05439_ ) );
AND3_X1 _13389_ ( .A1(_05129_ ), .A2(_04766_ ), .A3(_05131_ ), .ZN(_05440_ ) );
AOI21_X1 _13390_ ( .A(_01969_ ), .B1(_05129_ ), .B2(_05131_ ), .ZN(_05441_ ) );
OR3_X1 _13391_ ( .A1(_05440_ ), .A2(_05415_ ), .A3(_05441_ ), .ZN(_05442_ ) );
AOI21_X1 _13392_ ( .A(_05370_ ), .B1(_05439_ ), .B2(_05442_ ), .ZN(_05443_ ) );
BUF_X2 _13393_ ( .A(_05213_ ), .Z(_05444_ ) );
AND3_X1 _13394_ ( .A1(_05142_ ), .A2(_04836_ ), .A3(_05143_ ), .ZN(_05445_ ) );
OAI21_X1 _13395_ ( .A(_05444_ ), .B1(_05445_ ), .B2(_05383_ ), .ZN(_05446_ ) );
AND3_X1 _13396_ ( .A1(_05173_ ), .A2(_04842_ ), .A3(_05174_ ), .ZN(_05447_ ) );
AOI21_X1 _13397_ ( .A(_02018_ ), .B1(_05173_ ), .B2(_05174_ ), .ZN(_05448_ ) );
OAI21_X1 _13398_ ( .A(_05415_ ), .B1(_05447_ ), .B2(_05448_ ), .ZN(_05449_ ) );
AND3_X1 _13399_ ( .A1(_05446_ ), .A2(_05449_ ), .A3(_05423_ ), .ZN(_05450_ ) );
BUF_X2 _13400_ ( .A(_05408_ ), .Z(_05451_ ) );
BUF_X2 _13401_ ( .A(_05451_ ), .Z(_05452_ ) );
NOR3_X1 _13402_ ( .A1(_05443_ ), .A2(_05450_ ), .A3(_05452_ ), .ZN(_05453_ ) );
NOR3_X1 _13403_ ( .A1(_05436_ ), .A2(_05381_ ), .A3(_05453_ ), .ZN(_05454_ ) );
AND2_X1 _13404_ ( .A1(_04977_ ), .A2(_03359_ ), .ZN(_05455_ ) );
INV_X1 _13405_ ( .A(_05455_ ), .ZN(_05456_ ) );
AND2_X1 _13406_ ( .A1(_05110_ ), .A2(_04787_ ), .ZN(_05457_ ) );
AND3_X1 _13407_ ( .A1(_05169_ ), .A2(_04384_ ), .A3(_05170_ ), .ZN(_05458_ ) );
OAI21_X1 _13408_ ( .A(_05219_ ), .B1(_05457_ ), .B2(_05458_ ), .ZN(_05459_ ) );
AND3_X1 _13409_ ( .A1(_05169_ ), .A2(_01601_ ), .A3(_05170_ ), .ZN(_05460_ ) );
AOI21_X1 _13410_ ( .A(_03394_ ), .B1(_05214_ ), .B2(_05215_ ), .ZN(_05461_ ) );
OAI21_X1 _13411_ ( .A(_05420_ ), .B1(_05460_ ), .B2(_05461_ ), .ZN(_05462_ ) );
NAND2_X1 _13412_ ( .A1(_05459_ ), .A2(_05462_ ), .ZN(_05463_ ) );
MUX2_X1 _13413_ ( .A(_05456_ ), .B(_05463_ ), .S(_05369_ ), .Z(_05464_ ) );
BUF_X4 _13414_ ( .A(_05409_ ), .Z(_05465_ ) );
BUF_X4 _13415_ ( .A(_05465_ ), .Z(_05466_ ) );
BUF_X2 _13416_ ( .A(_05159_ ), .Z(_05467_ ) );
NOR3_X1 _13417_ ( .A1(_05464_ ), .A2(_05466_ ), .A3(_05467_ ), .ZN(_05468_ ) );
OAI21_X1 _13418_ ( .A(_05413_ ), .B1(_05454_ ), .B2(_05468_ ), .ZN(_05469_ ) );
BUF_X4 _13419_ ( .A(_05344_ ), .Z(_05470_ ) );
AOI21_X1 _13420_ ( .A(_05470_ ), .B1(_05073_ ), .B2(_04855_ ), .ZN(_05471_ ) );
BUF_X2 _13421_ ( .A(_05335_ ), .Z(_05472_ ) );
AOI21_X1 _13422_ ( .A(_05471_ ), .B1(_05241_ ), .B2(_05472_ ), .ZN(_05473_ ) );
BUF_X2 _13423_ ( .A(_05235_ ), .Z(_05474_ ) );
BUF_X4 _13424_ ( .A(_05338_ ), .Z(_05475_ ) );
BUF_X4 _13425_ ( .A(_05475_ ), .Z(_05476_ ) );
AOI22_X1 _13426_ ( .A1(_05411_ ), .A2(_05474_ ), .B1(_05330_ ), .B2(_05476_ ), .ZN(_05477_ ) );
NAND4_X1 _13427_ ( .A1(_05412_ ), .A2(_05469_ ), .A3(_05473_ ), .A4(_05477_ ), .ZN(_05478_ ) );
BUF_X4 _13428_ ( .A(_05239_ ), .Z(_05479_ ) );
AND2_X4 _13429_ ( .A1(_05316_ ), .A2(_05326_ ), .ZN(_05480_ ) );
OAI21_X1 _13430_ ( .A(_05479_ ), .B1(_05480_ ), .B2(_05242_ ), .ZN(_05481_ ) );
AOI21_X1 _13431_ ( .A(_05481_ ), .B1(_05480_ ), .B2(_05242_ ), .ZN(_05482_ ) );
OAI21_X1 _13432_ ( .A(_05365_ ), .B1(_05478_ ), .B2(_05482_ ), .ZN(_05483_ ) );
CLKBUF_X2 _13433_ ( .A(_05359_ ), .Z(_05484_ ) );
AOI21_X1 _13434_ ( .A(_04867_ ), .B1(_04854_ ), .B2(_04856_ ), .ZN(_05485_ ) );
OAI21_X1 _13435_ ( .A(_05485_ ), .B1(_04856_ ), .B2(_04854_ ), .ZN(_05486_ ) );
BUF_X2 _13436_ ( .A(_04955_ ), .Z(_05487_ ) );
AND3_X1 _13437_ ( .A1(_04936_ ), .A2(_04944_ ), .A3(_04947_ ), .ZN(_05488_ ) );
OR3_X1 _13438_ ( .A1(_04948_ ), .A2(_05487_ ), .A3(_05488_ ), .ZN(_05489_ ) );
NAND2_X1 _13439_ ( .A1(_05486_ ), .A2(_05489_ ), .ZN(_05490_ ) );
BUF_X2 _13440_ ( .A(_04962_ ), .Z(_05491_ ) );
BUF_X2 _13441_ ( .A(_04964_ ), .Z(_05492_ ) );
AND3_X1 _13442_ ( .A1(_05491_ ), .A2(\ID_EX_imm [20] ), .A3(_05492_ ), .ZN(_05493_ ) );
OAI21_X1 _13443_ ( .A(_04759_ ), .B1(_05490_ ), .B2(_05493_ ), .ZN(_05494_ ) );
AND3_X1 _13444_ ( .A1(_05483_ ), .A2(_05484_ ), .A3(_05494_ ), .ZN(_05495_ ) );
NAND2_X1 _13445_ ( .A1(_04755_ ), .A2(\ID_EX_pc [20] ), .ZN(_05496_ ) );
BUF_X4 _13446_ ( .A(_01361_ ), .Z(_05497_ ) );
BUF_X2 _13447_ ( .A(_04750_ ), .Z(_05498_ ) );
NAND4_X1 _13448_ ( .A1(_05498_ ), .A2(_02327_ ), .A3(_04753_ ), .A4(_04754_ ), .ZN(_05499_ ) );
NAND3_X1 _13449_ ( .A1(_05496_ ), .A2(_05497_ ), .A3(_05499_ ), .ZN(_05500_ ) );
NAND2_X1 _13450_ ( .A1(_05500_ ), .A2(_03407_ ), .ZN(_05501_ ) );
OAI21_X1 _13451_ ( .A(_05363_ ), .B1(_05495_ ), .B2(_05501_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OR3_X1 _13452_ ( .A1(_04197_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_04198_ ), .ZN(_05502_ ) );
NOR2_X1 _13453_ ( .A1(_03527_ ), .A2(_03601_ ), .ZN(_05503_ ) );
NAND4_X1 _13454_ ( .A1(_04119_ ), .A2(\ID_EX_csr [2] ), .A3(\mtvec [19] ), .A4(_04200_ ), .ZN(_05504_ ) );
NAND3_X1 _13455_ ( .A1(_05503_ ), .A2(_03593_ ), .A3(_05504_ ), .ZN(_05505_ ) );
NAND3_X1 _13456_ ( .A1(_04122_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_04200_ ), .ZN(_05506_ ) );
OAI21_X1 _13457_ ( .A(_05506_ ), .B1(_04197_ ), .B2(_04198_ ), .ZN(_05507_ ) );
OAI211_X1 _13458_ ( .A(_05502_ ), .B(_03698_ ), .C1(_05505_ ), .C2(_05507_ ), .ZN(_05508_ ) );
BUF_X4 _13459_ ( .A(_05355_ ), .Z(_05509_ ) );
AND3_X1 _13460_ ( .A1(_04834_ ), .A2(_04841_ ), .A3(_04843_ ), .ZN(_05510_ ) );
OR3_X1 _13461_ ( .A1(_05510_ ), .A2(_04848_ ), .A3(_04851_ ), .ZN(_05511_ ) );
AOI21_X1 _13462_ ( .A(_04845_ ), .B1(_05511_ ), .B2(_04838_ ), .ZN(_05512_ ) );
XNOR2_X1 _13463_ ( .A(_05512_ ), .B(_04837_ ), .ZN(_05513_ ) );
BUF_X2 _13464_ ( .A(_04865_ ), .Z(_05514_ ) );
BUF_X2 _13465_ ( .A(_05514_ ), .Z(_05515_ ) );
NAND2_X1 _13466_ ( .A1(_05513_ ), .A2(_05515_ ), .ZN(_05516_ ) );
AOI21_X1 _13467_ ( .A(_04940_ ), .B1(_04929_ ), .B2(_04935_ ), .ZN(_05517_ ) );
INV_X1 _13468_ ( .A(_04930_ ), .ZN(_05518_ ) );
OR2_X1 _13469_ ( .A1(_05517_ ), .A2(_05518_ ), .ZN(_05519_ ) );
OAI21_X1 _13470_ ( .A(_05519_ ), .B1(_02329_ ), .B2(_02019_ ), .ZN(_05520_ ) );
AOI21_X1 _13471_ ( .A(_05487_ ), .B1(_05520_ ), .B2(_04931_ ), .ZN(_05521_ ) );
OAI21_X1 _13472_ ( .A(_05521_ ), .B1(_04931_ ), .B2(_05520_ ), .ZN(_05522_ ) );
AND2_X1 _13473_ ( .A1(_05516_ ), .A2(_05522_ ), .ZN(_05523_ ) );
BUF_X4 _13474_ ( .A(_04962_ ), .Z(_05524_ ) );
BUF_X4 _13475_ ( .A(_04964_ ), .Z(_05525_ ) );
NAND3_X1 _13476_ ( .A1(_05524_ ), .A2(\ID_EX_imm [19] ), .A3(_05525_ ), .ZN(_05526_ ) );
AOI21_X1 _13477_ ( .A(_05509_ ), .B1(_05523_ ), .B2(_05526_ ), .ZN(_05527_ ) );
BUF_X4 _13478_ ( .A(_05357_ ), .Z(_05528_ ) );
AND3_X1 _13479_ ( .A1(_05214_ ), .A2(_03814_ ), .A3(_05215_ ), .ZN(_05529_ ) );
OAI21_X1 _13480_ ( .A(_05444_ ), .B1(_05529_ ), .B2(_05204_ ), .ZN(_05530_ ) );
AND3_X1 _13481_ ( .A1(_05129_ ), .A2(_04763_ ), .A3(_05131_ ), .ZN(_05531_ ) );
OAI21_X1 _13482_ ( .A(_05415_ ), .B1(_05531_ ), .B2(_05187_ ), .ZN(_05532_ ) );
NAND3_X1 _13483_ ( .A1(_05530_ ), .A2(_05532_ ), .A3(_05428_ ), .ZN(_05533_ ) );
OAI21_X1 _13484_ ( .A(_05444_ ), .B1(_05199_ ), .B2(_05200_ ), .ZN(_05534_ ) );
AND3_X1 _13485_ ( .A1(_05214_ ), .A2(_04840_ ), .A3(_05215_ ), .ZN(_05535_ ) );
OAI21_X1 _13486_ ( .A(_05415_ ), .B1(_05535_ ), .B2(_05207_ ), .ZN(_05536_ ) );
NAND3_X1 _13487_ ( .A1(_05534_ ), .A2(_05536_ ), .A3(_05423_ ), .ZN(_05537_ ) );
AND3_X1 _13488_ ( .A1(_05533_ ), .A2(_05537_ ), .A3(_05426_ ), .ZN(_05538_ ) );
NOR3_X1 _13489_ ( .A1(_05175_ ), .A2(_05219_ ), .A3(_05176_ ), .ZN(_05539_ ) );
NOR3_X1 _13490_ ( .A1(_05216_ ), .A2(_05217_ ), .A3(_05213_ ), .ZN(_05540_ ) );
NOR2_X1 _13491_ ( .A1(_05539_ ), .A2(_05540_ ), .ZN(_05541_ ) );
NAND2_X1 _13492_ ( .A1(_05541_ ), .A2(_05428_ ), .ZN(_05542_ ) );
NOR3_X1 _13493_ ( .A1(_05183_ ), .A2(_05219_ ), .A3(_05185_ ), .ZN(_05543_ ) );
NOR3_X1 _13494_ ( .A1(_05166_ ), .A2(_05171_ ), .A3(_05213_ ), .ZN(_05544_ ) );
NOR2_X1 _13495_ ( .A1(_05543_ ), .A2(_05544_ ), .ZN(_05545_ ) );
NAND2_X1 _13496_ ( .A1(_05545_ ), .A2(_05423_ ), .ZN(_05546_ ) );
NAND2_X1 _13497_ ( .A1(_05542_ ), .A2(_05546_ ), .ZN(_05547_ ) );
AOI211_X1 _13498_ ( .A(_05380_ ), .B(_05538_ ), .C1(_05547_ ), .C2(_05466_ ), .ZN(_05548_ ) );
OAI21_X1 _13499_ ( .A(_05213_ ), .B1(_05220_ ), .B2(_05221_ ), .ZN(_05549_ ) );
NOR2_X1 _13500_ ( .A1(_05226_ ), .A2(_05227_ ), .ZN(_05550_ ) );
OAI21_X1 _13501_ ( .A(_05549_ ), .B1(_05550_ ), .B2(_05420_ ), .ZN(_05551_ ) );
BUF_X4 _13502_ ( .A(_05399_ ), .Z(_05552_ ) );
BUF_X2 _13503_ ( .A(_05165_ ), .Z(_05553_ ) );
NOR4_X1 _13504_ ( .A1(_05551_ ), .A2(_05466_ ), .A3(_05552_ ), .A4(_05553_ ), .ZN(_05554_ ) );
OAI21_X1 _13505_ ( .A(_05413_ ), .B1(_05548_ ), .B2(_05554_ ), .ZN(_05555_ ) );
AND2_X4 _13506_ ( .A1(_05122_ ), .A2(_05118_ ), .ZN(_05556_ ) );
NAND2_X1 _13507_ ( .A1(_05110_ ), .A2(_02214_ ), .ZN(_05557_ ) );
OAI211_X1 _13508_ ( .A(_05557_ ), .B(_05168_ ), .C1(_01446_ ), .C2(_05189_ ), .ZN(_05558_ ) );
OAI21_X1 _13509_ ( .A(_05177_ ), .B1(_05141_ ), .B2(_05144_ ), .ZN(_05559_ ) );
NAND3_X1 _13510_ ( .A1(_05558_ ), .A2(_05559_ ), .A3(_05229_ ), .ZN(_05560_ ) );
NAND4_X1 _13511_ ( .A1(_05202_ ), .A2(_02268_ ), .A3(_05213_ ), .A4(_05189_ ), .ZN(_05561_ ) );
NAND2_X1 _13512_ ( .A1(_05560_ ), .A2(_05561_ ), .ZN(_05562_ ) );
NAND2_X1 _13513_ ( .A1(_05562_ ), .A2(_05408_ ), .ZN(_05563_ ) );
NOR3_X1 _13514_ ( .A1(_05138_ ), .A2(_05139_ ), .A3(_05184_ ), .ZN(_05564_ ) );
NOR3_X1 _13515_ ( .A1(_05152_ ), .A2(_05167_ ), .A3(_05153_ ), .ZN(_05565_ ) );
OR3_X1 _13516_ ( .A1(_05564_ ), .A2(_05565_ ), .A3(_05113_ ), .ZN(_05566_ ) );
NOR3_X1 _13517_ ( .A1(_05196_ ), .A2(_05197_ ), .A3(_05200_ ), .ZN(_05567_ ) );
NOR3_X1 _13518_ ( .A1(_05148_ ), .A2(_05149_ ), .A3(_05184_ ), .ZN(_05568_ ) );
NOR2_X1 _13519_ ( .A1(_05567_ ), .A2(_05568_ ), .ZN(_05569_ ) );
NAND2_X1 _13520_ ( .A1(_05569_ ), .A2(_05180_ ), .ZN(_05570_ ) );
NAND2_X1 _13521_ ( .A1(_05566_ ), .A2(_05570_ ), .ZN(_05571_ ) );
OAI21_X1 _13522_ ( .A(_05563_ ), .B1(_05571_ ), .B2(_05409_ ), .ZN(_05572_ ) );
AND2_X1 _13523_ ( .A1(_05572_ ), .A2(_05165_ ), .ZN(_05573_ ) );
XNOR2_X1 _13524_ ( .A(_04977_ ), .B(_05113_ ), .ZN(_05574_ ) );
AND4_X1 _13525_ ( .A1(_05368_ ), .A2(_05108_ ), .A3(_05574_ ), .A4(_05120_ ), .ZN(_05575_ ) );
OR3_X1 _13526_ ( .A1(_05556_ ), .A2(_05573_ ), .A3(_05575_ ), .ZN(_05576_ ) );
AOI22_X1 _13527_ ( .A1(_05576_ ), .A2(_05366_ ), .B1(_05474_ ), .B2(_05573_ ), .ZN(_05577_ ) );
NAND3_X1 _13528_ ( .A1(_05322_ ), .A2(_05323_ ), .A3(_05472_ ), .ZN(_05578_ ) );
NOR3_X1 _13529_ ( .A1(_05076_ ), .A2(_04836_ ), .A3(_05340_ ), .ZN(_05579_ ) );
BUF_X4 _13530_ ( .A(_05342_ ), .Z(_05580_ ) );
AOI21_X1 _13531_ ( .A(_05579_ ), .B1(_05323_ ), .B2(_05580_ ), .ZN(_05581_ ) );
AND4_X1 _13532_ ( .A1(_05555_ ), .A2(_05577_ ), .A3(_05578_ ), .A4(_05581_ ), .ZN(_05582_ ) );
INV_X1 _13533_ ( .A(_05312_ ), .ZN(_05583_ ) );
INV_X1 _13534_ ( .A(_05313_ ), .ZN(_05584_ ) );
AOI211_X1 _13535_ ( .A(_05583_ ), .B(_05584_ ), .C1(_05275_ ), .C2(_05307_ ), .ZN(_05585_ ) );
NOR2_X1 _13536_ ( .A1(_05585_ ), .A2(_05320_ ), .ZN(_05586_ ) );
INV_X1 _13537_ ( .A(_05310_ ), .ZN(_05587_ ) );
NOR2_X1 _13538_ ( .A1(_05586_ ), .A2(_05587_ ), .ZN(_05588_ ) );
OR3_X1 _13539_ ( .A1(_05588_ ), .A2(_05309_ ), .A3(_05324_ ), .ZN(_05589_ ) );
OAI21_X1 _13540_ ( .A(_05309_ ), .B1(_05588_ ), .B2(_05324_ ), .ZN(_05590_ ) );
NAND3_X1 _13541_ ( .A1(_05589_ ), .A2(_05479_ ), .A3(_05590_ ), .ZN(_05591_ ) );
AOI21_X1 _13542_ ( .A(_05528_ ), .B1(_05582_ ), .B2(_05591_ ), .ZN(_05592_ ) );
NOR3_X1 _13543_ ( .A1(_05527_ ), .A2(_01362_ ), .A3(_05592_ ), .ZN(_05593_ ) );
NAND3_X1 _13544_ ( .A1(_05498_ ), .A2(\ID_EX_pc [18] ), .A3(_04753_ ), .ZN(_05594_ ) );
NAND2_X1 _13545_ ( .A1(_05594_ ), .A2(\ID_EX_pc [19] ), .ZN(_05595_ ) );
NAND4_X1 _13546_ ( .A1(_05498_ ), .A2(_02328_ ), .A3(\ID_EX_pc [18] ), .A4(_04753_ ), .ZN(_05596_ ) );
NAND3_X1 _13547_ ( .A1(_05595_ ), .A2(_05497_ ), .A3(_05596_ ), .ZN(_05597_ ) );
NAND2_X1 _13548_ ( .A1(_05597_ ), .A2(_03407_ ), .ZN(_05598_ ) );
OAI21_X1 _13549_ ( .A(_05508_ ), .B1(_05593_ ), .B2(_05598_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
INV_X1 _13550_ ( .A(_03657_ ), .ZN(_05599_ ) );
AND2_X2 _13551_ ( .A1(_04750_ ), .A2(_04753_ ), .ZN(_05600_ ) );
XNOR2_X1 _13552_ ( .A(_05600_ ), .B(_02329_ ), .ZN(_05601_ ) );
AOI21_X1 _13553_ ( .A(_04866_ ), .B1(_05511_ ), .B2(_04838_ ), .ZN(_05602_ ) );
OAI21_X1 _13554_ ( .A(_05602_ ), .B1(_04838_ ), .B2(_05511_ ), .ZN(_05603_ ) );
NAND2_X1 _13555_ ( .A1(_05517_ ), .A2(_05518_ ), .ZN(_05604_ ) );
NAND3_X1 _13556_ ( .A1(_05519_ ), .A2(_04954_ ), .A3(_05604_ ), .ZN(_05605_ ) );
NAND2_X1 _13557_ ( .A1(_05603_ ), .A2(_05605_ ), .ZN(_05606_ ) );
AND3_X1 _13558_ ( .A1(_04961_ ), .A2(\ID_EX_imm [18] ), .A3(_04963_ ), .ZN(_05607_ ) );
OAI21_X1 _13559_ ( .A(_04759_ ), .B1(_05606_ ), .B2(_05607_ ), .ZN(_05608_ ) );
NAND3_X1 _13560_ ( .A1(_05019_ ), .A2(_05106_ ), .A3(_05574_ ), .ZN(_05609_ ) );
NOR2_X1 _13561_ ( .A1(_05167_ ), .A2(_05110_ ), .ZN(_05610_ ) );
NOR3_X1 _13562_ ( .A1(_05609_ ), .A2(_05610_ ), .A3(_05116_ ), .ZN(_05611_ ) );
OAI22_X1 _13563_ ( .A1(_05122_ ), .A2(_05123_ ), .B1(_05611_ ), .B2(_05119_ ), .ZN(_05612_ ) );
OR3_X1 _13564_ ( .A1(_05445_ ), .A2(_05134_ ), .A3(_05448_ ), .ZN(_05613_ ) );
OR3_X1 _13565_ ( .A1(_05382_ ), .A2(_05383_ ), .A3(_05127_ ), .ZN(_05614_ ) );
AOI21_X1 _13566_ ( .A(_05125_ ), .B1(_05613_ ), .B2(_05614_ ), .ZN(_05615_ ) );
OR3_X1 _13567_ ( .A1(_05392_ ), .A2(_05393_ ), .A3(_05127_ ), .ZN(_05616_ ) );
INV_X1 _13568_ ( .A(_05387_ ), .ZN(_05617_ ) );
OAI211_X1 _13569_ ( .A(_05617_ ), .B(_05111_ ), .C1(_02042_ ), .C2(_05110_ ), .ZN(_05618_ ) );
AOI21_X1 _13570_ ( .A(_05113_ ), .B1(_05616_ ), .B2(_05618_ ), .ZN(_05619_ ) );
OR2_X1 _13571_ ( .A1(_05615_ ), .A2(_05619_ ), .ZN(_05620_ ) );
NOR3_X1 _13572_ ( .A1(_05395_ ), .A2(_05134_ ), .A3(_05396_ ), .ZN(_05621_ ) );
NOR3_X1 _13573_ ( .A1(_05402_ ), .A2(_05403_ ), .A3(_05127_ ), .ZN(_05622_ ) );
NOR2_X1 _13574_ ( .A1(_05621_ ), .A2(_05622_ ), .ZN(_05623_ ) );
NAND2_X1 _13575_ ( .A1(_05623_ ), .A2(_05113_ ), .ZN(_05624_ ) );
AND2_X1 _13576_ ( .A1(_05406_ ), .A2(_05111_ ), .ZN(_05625_ ) );
OAI21_X1 _13577_ ( .A(_05624_ ), .B1(_05113_ ), .B2(_05625_ ), .ZN(_05626_ ) );
INV_X1 _13578_ ( .A(_05626_ ), .ZN(_05627_ ) );
MUX2_X1 _13579_ ( .A(_05620_ ), .B(_05627_ ), .S(_05408_ ), .Z(_05628_ ) );
NAND2_X1 _13580_ ( .A1(_05628_ ), .A2(_05165_ ), .ZN(_05629_ ) );
AOI21_X1 _13581_ ( .A(_04970_ ), .B1(_05612_ ), .B2(_05629_ ), .ZN(_05630_ ) );
OAI21_X1 _13582_ ( .A(_05239_ ), .B1(_05586_ ), .B2(_05587_ ), .ZN(_05631_ ) );
AOI21_X1 _13583_ ( .A(_05631_ ), .B1(_05587_ ), .B2(_05586_ ), .ZN(_05632_ ) );
INV_X1 _13584_ ( .A(_05029_ ), .ZN(_05633_ ) );
NAND3_X1 _13585_ ( .A1(_05633_ ), .A2(_02018_ ), .A3(_05475_ ), .ZN(_05634_ ) );
INV_X1 _13586_ ( .A(_05235_ ), .ZN(_05635_ ) );
OAI21_X1 _13587_ ( .A(_05634_ ), .B1(_05629_ ), .B2(_05635_ ), .ZN(_05636_ ) );
OAI21_X1 _13588_ ( .A(_05184_ ), .B1(_05457_ ), .B2(_05458_ ), .ZN(_05637_ ) );
OAI21_X1 _13589_ ( .A(_05197_ ), .B1(_05371_ ), .B2(_05225_ ), .ZN(_05638_ ) );
AND3_X1 _13590_ ( .A1(_05637_ ), .A2(_05229_ ), .A3(_05638_ ), .ZN(_05639_ ) );
AND2_X1 _13591_ ( .A1(_05639_ ), .A2(_05193_ ), .ZN(_05640_ ) );
OAI21_X1 _13592_ ( .A(_05163_ ), .B1(_05640_ ), .B2(_05158_ ), .ZN(_05641_ ) );
OAI21_X1 _13593_ ( .A(_05197_ ), .B1(_05414_ ), .B2(_05416_ ), .ZN(_05642_ ) );
OAI21_X1 _13594_ ( .A(_05177_ ), .B1(_05432_ ), .B2(_05433_ ), .ZN(_05643_ ) );
NAND2_X1 _13595_ ( .A1(_05642_ ), .A2(_05643_ ), .ZN(_05644_ ) );
NAND2_X1 _13596_ ( .A1(_05644_ ), .A2(_05180_ ), .ZN(_05645_ ) );
OAI21_X1 _13597_ ( .A(_05177_ ), .B1(_05418_ ), .B2(_05419_ ), .ZN(_05646_ ) );
OAI21_X1 _13598_ ( .A(_05197_ ), .B1(_05460_ ), .B2(_05461_ ), .ZN(_05647_ ) );
NAND2_X1 _13599_ ( .A1(_05646_ ), .A2(_05647_ ), .ZN(_05648_ ) );
NAND2_X1 _13600_ ( .A1(_05648_ ), .A2(_05182_ ), .ZN(_05649_ ) );
NAND2_X1 _13601_ ( .A1(_05645_ ), .A2(_05649_ ), .ZN(_05650_ ) );
OR3_X1 _13602_ ( .A1(_05447_ ), .A2(_05167_ ), .A3(_05448_ ), .ZN(_05651_ ) );
OR3_X1 _13603_ ( .A1(_05440_ ), .A2(_05441_ ), .A3(_05111_ ), .ZN(_05652_ ) );
NAND3_X1 _13604_ ( .A1(_05651_ ), .A2(_05652_ ), .A3(_05229_ ), .ZN(_05653_ ) );
OR3_X1 _13605_ ( .A1(_05437_ ), .A2(_05167_ ), .A3(_05438_ ), .ZN(_05654_ ) );
OR3_X1 _13606_ ( .A1(_05429_ ), .A2(_05430_ ), .A3(_05111_ ), .ZN(_05655_ ) );
NAND3_X1 _13607_ ( .A1(_05654_ ), .A2(_05202_ ), .A3(_05655_ ), .ZN(_05656_ ) );
NAND2_X1 _13608_ ( .A1(_05653_ ), .A2(_05656_ ), .ZN(_05657_ ) );
MUX2_X1 _13609_ ( .A(_05650_ ), .B(_05657_ ), .S(_05193_ ), .Z(_05658_ ) );
AOI21_X1 _13610_ ( .A(_05641_ ), .B1(_05658_ ), .B2(_05159_ ), .ZN(_05659_ ) );
OAI21_X1 _13611_ ( .A(_05342_ ), .B1(_05633_ ), .B2(_02018_ ), .ZN(_05660_ ) );
INV_X1 _13612_ ( .A(_05334_ ), .ZN(_05661_ ) );
BUF_X4 _13613_ ( .A(_05661_ ), .Z(_05662_ ) );
OAI21_X1 _13614_ ( .A(_05660_ ), .B1(_05587_ ), .B2(_05662_ ), .ZN(_05663_ ) );
OR3_X1 _13615_ ( .A1(_05636_ ), .A2(_05659_ ), .A3(_05663_ ), .ZN(_05664_ ) );
NOR3_X1 _13616_ ( .A1(_05630_ ), .A2(_05632_ ), .A3(_05664_ ), .ZN(_05665_ ) );
OAI21_X1 _13617_ ( .A(_05608_ ), .B1(_05357_ ), .B2(_05665_ ), .ZN(_05666_ ) );
MUX2_X1 _13618_ ( .A(_05601_ ), .B(_05666_ ), .S(_05360_ ), .Z(_05667_ ) );
MUX2_X1 _13619_ ( .A(_05599_ ), .B(_05667_ ), .S(_03390_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
INV_X1 _13620_ ( .A(_03701_ ), .ZN(_05668_ ) );
INV_X1 _13621_ ( .A(_01360_ ), .ZN(_05669_ ) );
AND2_X1 _13622_ ( .A1(_04929_ ), .A2(_04933_ ), .ZN(_05670_ ) );
OR3_X1 _13623_ ( .A1(_05670_ ), .A2(_04934_ ), .A3(_04937_ ), .ZN(_05671_ ) );
BUF_X4 _13624_ ( .A(_04954_ ), .Z(_05672_ ) );
OAI21_X1 _13625_ ( .A(_04934_ ), .B1(_05670_ ), .B2(_04937_ ), .ZN(_05673_ ) );
NAND3_X1 _13626_ ( .A1(_05671_ ), .A2(_05672_ ), .A3(_05673_ ), .ZN(_05674_ ) );
NAND3_X1 _13627_ ( .A1(_04962_ ), .A2(\ID_EX_imm [17] ), .A3(_04964_ ), .ZN(_05675_ ) );
NAND2_X1 _13628_ ( .A1(_05674_ ), .A2(_05675_ ), .ZN(_05676_ ) );
AND2_X1 _13629_ ( .A1(_04834_ ), .A2(_04841_ ), .ZN(_05677_ ) );
AND2_X1 _13630_ ( .A1(_03760_ ), .A2(_01969_ ), .ZN(_05678_ ) );
NOR3_X1 _13631_ ( .A1(_05677_ ), .A2(_05678_ ), .A3(_04843_ ), .ZN(_05679_ ) );
NOR2_X1 _13632_ ( .A1(_05679_ ), .A2(_04867_ ), .ZN(_05680_ ) );
OAI21_X1 _13633_ ( .A(_04843_ ), .B1(_05677_ ), .B2(_05678_ ), .ZN(_05681_ ) );
AOI21_X1 _13634_ ( .A(_05676_ ), .B1(_05680_ ), .B2(_05681_ ), .ZN(_05682_ ) );
AOI21_X1 _13635_ ( .A(_05669_ ), .B1(_05682_ ), .B2(_01355_ ), .ZN(_05683_ ) );
OR3_X1 _13636_ ( .A1(_05609_ ), .A2(_05112_ ), .A3(_05116_ ), .ZN(_05684_ ) );
AOI22_X1 _13637_ ( .A1(_05378_ ), .A2(_05377_ ), .B1(_05684_ ), .B2(_05376_ ), .ZN(_05685_ ) );
OR3_X1 _13638_ ( .A1(_05140_ ), .A2(_05145_ ), .A3(_05202_ ), .ZN(_05686_ ) );
NAND3_X1 _13639_ ( .A1(_05133_ ), .A2(_05182_ ), .A3(_05135_ ), .ZN(_05687_ ) );
NAND3_X1 _13640_ ( .A1(_05686_ ), .A2(_05465_ ), .A3(_05687_ ), .ZN(_05688_ ) );
NAND3_X1 _13641_ ( .A1(_05150_ ), .A2(_05154_ ), .A3(_05202_ ), .ZN(_05689_ ) );
OAI21_X1 _13642_ ( .A(_05127_ ), .B1(_05199_ ), .B2(_05207_ ), .ZN(_05690_ ) );
OAI21_X1 _13643_ ( .A(_05134_ ), .B1(_05196_ ), .B2(_05200_ ), .ZN(_05691_ ) );
NAND3_X1 _13644_ ( .A1(_05690_ ), .A2(_05691_ ), .A3(_05229_ ), .ZN(_05692_ ) );
AND2_X1 _13645_ ( .A1(_05689_ ), .A2(_05692_ ), .ZN(_05693_ ) );
OAI21_X1 _13646_ ( .A(_05688_ ), .B1(_05452_ ), .B2(_05693_ ), .ZN(_05694_ ) );
AND2_X1 _13647_ ( .A1(_05694_ ), .A2(_05467_ ), .ZN(_05695_ ) );
OAI21_X1 _13648_ ( .A(_05366_ ), .B1(_05685_ ), .B2(_05695_ ), .ZN(_05696_ ) );
NAND2_X1 _13649_ ( .A1(_05179_ ), .A2(_05423_ ), .ZN(_05697_ ) );
NAND2_X1 _13650_ ( .A1(_05223_ ), .A2(_05428_ ), .ZN(_05698_ ) );
NAND3_X1 _13651_ ( .A1(_05697_ ), .A2(_05466_ ), .A3(_05698_ ), .ZN(_05699_ ) );
BUF_X2 _13652_ ( .A(_05370_ ), .Z(_05700_ ) );
AOI21_X1 _13653_ ( .A(_05700_ ), .B1(_05186_ ), .B2(_05190_ ), .ZN(_05701_ ) );
AOI21_X1 _13654_ ( .A(_05552_ ), .B1(_05206_ ), .B2(_05209_ ), .ZN(_05702_ ) );
OAI21_X1 _13655_ ( .A(_05427_ ), .B1(_05701_ ), .B2(_05702_ ), .ZN(_05703_ ) );
AOI21_X1 _13656_ ( .A(_05381_ ), .B1(_05699_ ), .B2(_05703_ ), .ZN(_05704_ ) );
AND4_X1 _13657_ ( .A1(_05427_ ), .A2(_05228_ ), .A3(_05700_ ), .A4(_05380_ ), .ZN(_05705_ ) );
OAI21_X1 _13658_ ( .A(_05413_ ), .B1(_05704_ ), .B2(_05705_ ), .ZN(_05706_ ) );
NAND3_X1 _13659_ ( .A1(_05694_ ), .A2(_05467_ ), .A3(_05474_ ), .ZN(_05707_ ) );
NAND3_X1 _13660_ ( .A1(_05696_ ), .A2(_05706_ ), .A3(_05707_ ), .ZN(_05708_ ) );
BUF_X2 _13661_ ( .A(_05240_ ), .Z(_05709_ ) );
AOI21_X1 _13662_ ( .A(_05584_ ), .B1(_05275_ ), .B2(_05307_ ), .ZN(_05710_ ) );
OR3_X1 _13663_ ( .A1(_05710_ ), .A2(_05583_ ), .A3(_05318_ ), .ZN(_05711_ ) );
OAI21_X1 _13664_ ( .A(_05583_ ), .B1(_05710_ ), .B2(_05318_ ), .ZN(_05712_ ) );
AOI21_X1 _13665_ ( .A(_05709_ ), .B1(_05711_ ), .B2(_05712_ ), .ZN(_05713_ ) );
AND2_X1 _13666_ ( .A1(_05312_ ), .A2(_05472_ ), .ZN(_05714_ ) );
AOI21_X1 _13667_ ( .A(_05470_ ), .B1(_05032_ ), .B2(_04842_ ), .ZN(_05715_ ) );
NOR3_X1 _13668_ ( .A1(_05032_ ), .A2(_04842_ ), .A3(_05340_ ), .ZN(_05716_ ) );
OR3_X1 _13669_ ( .A1(_05714_ ), .A2(_05715_ ), .A3(_05716_ ), .ZN(_05717_ ) );
OR3_X1 _13670_ ( .A1(_05708_ ), .A2(_05713_ ), .A3(_05717_ ), .ZN(_05718_ ) );
AOI21_X1 _13671_ ( .A(_05683_ ), .B1(_05718_ ), .B2(_05365_ ), .ZN(_05719_ ) );
AND3_X1 _13672_ ( .A1(_04752_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_05720_ ) );
AND2_X1 _13673_ ( .A1(_05498_ ), .A2(_05720_ ), .ZN(_05721_ ) );
NAND3_X1 _13674_ ( .A1(_05721_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05722_ ) );
NOR2_X1 _13675_ ( .A1(_05722_ ), .A2(_02331_ ), .ZN(_05723_ ) );
XNOR2_X1 _13676_ ( .A(_05723_ ), .B(_02330_ ), .ZN(_05724_ ) );
BUF_X4 _13677_ ( .A(_05360_ ), .Z(_05725_ ) );
OAI21_X1 _13678_ ( .A(_04248_ ), .B1(_05724_ ), .B2(_05725_ ), .ZN(_05726_ ) );
OAI21_X1 _13679_ ( .A(_05668_ ), .B1(_05719_ ), .B2(_05726_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
INV_X1 _13680_ ( .A(_03734_ ), .ZN(_05727_ ) );
INV_X1 _13681_ ( .A(_05120_ ), .ZN(_05728_ ) );
INV_X1 _13682_ ( .A(_04987_ ), .ZN(_05729_ ) );
AOI211_X1 _13683_ ( .A(_05728_ ), .B(_05109_ ), .C1(_05553_ ), .C2(_05729_ ), .ZN(_05730_ ) );
NAND2_X1 _13684_ ( .A1(_05407_ ), .A2(_05202_ ), .ZN(_05731_ ) );
OAI21_X1 _13685_ ( .A(_05731_ ), .B1(_05182_ ), .B2(_05398_ ), .ZN(_05732_ ) );
NOR2_X1 _13686_ ( .A1(_05389_ ), .A2(_05229_ ), .ZN(_05733_ ) );
OR3_X1 _13687_ ( .A1(_05447_ ), .A2(_05167_ ), .A3(_05441_ ), .ZN(_05734_ ) );
OR3_X1 _13688_ ( .A1(_05445_ ), .A2(_05448_ ), .A3(_05127_ ), .ZN(_05735_ ) );
AOI21_X1 _13689_ ( .A(_05125_ ), .B1(_05734_ ), .B2(_05735_ ), .ZN(_05736_ ) );
NOR2_X1 _13690_ ( .A1(_05733_ ), .A2(_05736_ ), .ZN(_05737_ ) );
INV_X1 _13691_ ( .A(_05737_ ), .ZN(_05738_ ) );
MUX2_X1 _13692_ ( .A(_05732_ ), .B(_05738_ ), .S(_05193_ ), .Z(_05739_ ) );
AND2_X1 _13693_ ( .A1(_05739_ ), .A2(_05159_ ), .ZN(_05740_ ) );
OAI21_X1 _13694_ ( .A(_05366_ ), .B1(_05730_ ), .B2(_05740_ ), .ZN(_05741_ ) );
NAND3_X1 _13695_ ( .A1(_05739_ ), .A2(_05467_ ), .A3(_05474_ ), .ZN(_05742_ ) );
NAND2_X1 _13696_ ( .A1(_05463_ ), .A2(_05552_ ), .ZN(_05743_ ) );
BUF_X2 _13697_ ( .A(_05369_ ), .Z(_05744_ ) );
NAND2_X1 _13698_ ( .A1(_05422_ ), .A2(_05744_ ), .ZN(_05745_ ) );
NAND3_X1 _13699_ ( .A1(_05743_ ), .A2(_05745_ ), .A3(_05465_ ), .ZN(_05746_ ) );
BUF_X2 _13700_ ( .A(_05159_ ), .Z(_05747_ ) );
NAND3_X1 _13701_ ( .A1(_05439_ ), .A2(_05442_ ), .A3(_05744_ ), .ZN(_05748_ ) );
NAND3_X1 _13702_ ( .A1(_05431_ ), .A2(_05434_ ), .A3(_05552_ ), .ZN(_05749_ ) );
NAND3_X1 _13703_ ( .A1(_05748_ ), .A2(_05749_ ), .A3(_05426_ ), .ZN(_05750_ ) );
AND3_X1 _13704_ ( .A1(_05746_ ), .A2(_05747_ ), .A3(_05750_ ), .ZN(_05751_ ) );
AND3_X1 _13705_ ( .A1(_04977_ ), .A2(_03359_ ), .A3(_05370_ ), .ZN(_05752_ ) );
AND2_X1 _13706_ ( .A1(_05752_ ), .A2(_05426_ ), .ZN(_05753_ ) );
OAI21_X1 _13707_ ( .A(_05413_ ), .B1(_05753_ ), .B2(_05747_ ), .ZN(_05754_ ) );
OAI211_X1 _13708_ ( .A(_05741_ ), .B(_05742_ ), .C1(_05751_ ), .C2(_05754_ ), .ZN(_05755_ ) );
AND3_X1 _13709_ ( .A1(_05275_ ), .A2(_05307_ ), .A3(_05584_ ), .ZN(_05756_ ) );
NOR3_X1 _13710_ ( .A1(_05756_ ), .A2(_05710_ ), .A3(_05240_ ), .ZN(_05757_ ) );
NAND3_X1 _13711_ ( .A1(_05033_ ), .A2(_04840_ ), .A3(_05034_ ), .ZN(_05758_ ) );
AOI22_X1 _13712_ ( .A1(_05318_ ), .A2(_05475_ ), .B1(_05758_ ), .B2(_05580_ ), .ZN(_05759_ ) );
OAI21_X1 _13713_ ( .A(_05759_ ), .B1(_05584_ ), .B2(_05662_ ), .ZN(_05760_ ) );
OR3_X1 _13714_ ( .A1(_05755_ ), .A2(_05757_ ), .A3(_05760_ ), .ZN(_05761_ ) );
AND2_X1 _13715_ ( .A1(_05761_ ), .A2(_05365_ ), .ZN(_05762_ ) );
AOI21_X1 _13716_ ( .A(_04867_ ), .B1(_04834_ ), .B2(_04841_ ), .ZN(_05763_ ) );
OAI21_X1 _13717_ ( .A(_05763_ ), .B1(_04834_ ), .B2(_04841_ ), .ZN(_05764_ ) );
AOI21_X1 _13718_ ( .A(_04955_ ), .B1(_04929_ ), .B2(_04933_ ), .ZN(_05765_ ) );
OAI21_X1 _13719_ ( .A(_05765_ ), .B1(_04929_ ), .B2(_04933_ ), .ZN(_05766_ ) );
NAND3_X1 _13720_ ( .A1(_05491_ ), .A2(\ID_EX_imm [16] ), .A3(_05492_ ), .ZN(_05767_ ) );
AND2_X1 _13721_ ( .A1(_05766_ ), .A2(_05767_ ), .ZN(_05768_ ) );
AOI21_X1 _13722_ ( .A(_05509_ ), .B1(_05764_ ), .B2(_05768_ ), .ZN(_05769_ ) );
NOR3_X1 _13723_ ( .A1(_05762_ ), .A2(_01362_ ), .A3(_05769_ ), .ZN(_05770_ ) );
XNOR2_X1 _13724_ ( .A(_05722_ ), .B(\ID_EX_pc [16] ), .ZN(_05771_ ) );
OAI21_X1 _13725_ ( .A(_04248_ ), .B1(_05771_ ), .B2(_05725_ ), .ZN(_05772_ ) );
OAI21_X1 _13726_ ( .A(_05727_ ), .B1(_05770_ ), .B2(_05772_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OR2_X1 _13727_ ( .A1(_03774_ ), .A2(_05362_ ), .ZN(_05773_ ) );
INV_X1 _13728_ ( .A(_04762_ ), .ZN(_05774_ ) );
INV_X1 _13729_ ( .A(_04764_ ), .ZN(_05775_ ) );
AND2_X1 _13730_ ( .A1(_04804_ ), .A2(_04813_ ), .ZN(_05776_ ) );
OR2_X1 _13731_ ( .A1(_05776_ ), .A2(_04782_ ), .ZN(_05777_ ) );
AOI211_X1 _13732_ ( .A(_05774_ ), .B(_05775_ ), .C1(_05777_ ), .C2(_04824_ ), .ZN(_05778_ ) );
OAI21_X1 _13733_ ( .A(_04768_ ), .B1(_05778_ ), .B2(_04830_ ), .ZN(_05779_ ) );
INV_X1 _13734_ ( .A(_04826_ ), .ZN(_05780_ ) );
AND2_X1 _13735_ ( .A1(_05779_ ), .A2(_05780_ ), .ZN(_05781_ ) );
XNOR2_X1 _13736_ ( .A(_05781_ ), .B(_04767_ ), .ZN(_05782_ ) );
NAND2_X1 _13737_ ( .A1(_05782_ ), .A2(_05514_ ), .ZN(_05783_ ) );
NOR2_X1 _13738_ ( .A1(_04911_ ), .A2(_04912_ ), .ZN(_05784_ ) );
INV_X1 _13739_ ( .A(_05784_ ), .ZN(_05785_ ) );
AND2_X1 _13740_ ( .A1(_05785_ ), .A2(_04884_ ), .ZN(_05786_ ) );
NOR2_X1 _13741_ ( .A1(_05786_ ), .A2(_04927_ ), .ZN(_05787_ ) );
INV_X1 _13742_ ( .A(_04875_ ), .ZN(_05788_ ) );
NOR2_X1 _13743_ ( .A1(_05787_ ), .A2(_05788_ ), .ZN(_05789_ ) );
INV_X1 _13744_ ( .A(_05789_ ), .ZN(_05790_ ) );
AOI21_X1 _13745_ ( .A(_04873_ ), .B1(_05790_ ), .B2(_04918_ ), .ZN(_05791_ ) );
AND2_X1 _13746_ ( .A1(_05791_ ), .A2(_04870_ ), .ZN(_05792_ ) );
OR3_X1 _13747_ ( .A1(_05792_ ), .A2(_04869_ ), .A3(_04914_ ), .ZN(_05793_ ) );
OAI21_X1 _13748_ ( .A(_04869_ ), .B1(_05792_ ), .B2(_04914_ ), .ZN(_05794_ ) );
NAND3_X1 _13749_ ( .A1(_05793_ ), .A2(_05672_ ), .A3(_05794_ ), .ZN(_05795_ ) );
NAND3_X1 _13750_ ( .A1(_05491_ ), .A2(\ID_EX_imm [15] ), .A3(_05492_ ), .ZN(_05796_ ) );
AND3_X1 _13751_ ( .A1(_05783_ ), .A2(_05795_ ), .A3(_05796_ ), .ZN(_05797_ ) );
AOI21_X1 _13752_ ( .A(_05669_ ), .B1(_05797_ ), .B2(_01355_ ), .ZN(_05798_ ) );
BUF_X4 _13753_ ( .A(_04970_ ), .Z(_05799_ ) );
INV_X1 _13754_ ( .A(_05556_ ), .ZN(_05800_ ) );
NOR3_X1 _13755_ ( .A1(_05535_ ), .A2(_05219_ ), .A3(_05204_ ), .ZN(_05801_ ) );
NOR3_X1 _13756_ ( .A1(_05199_ ), .A2(_05207_ ), .A3(_05213_ ), .ZN(_05802_ ) );
OAI21_X1 _13757_ ( .A(_05370_ ), .B1(_05801_ ), .B2(_05802_ ), .ZN(_05803_ ) );
BUF_X2 _13758_ ( .A(_05194_ ), .Z(_05804_ ) );
OAI211_X1 _13759_ ( .A(_05803_ ), .B(_05804_ ), .C1(_05569_ ), .C2(_05700_ ), .ZN(_05805_ ) );
OAI21_X1 _13760_ ( .A(_05229_ ), .B1(_05565_ ), .B2(_05564_ ), .ZN(_05806_ ) );
NAND3_X1 _13761_ ( .A1(_05558_ ), .A2(_05559_ ), .A3(_05202_ ), .ZN(_05807_ ) );
NAND2_X1 _13762_ ( .A1(_05806_ ), .A2(_05807_ ), .ZN(_05808_ ) );
OAI211_X1 _13763_ ( .A(_05805_ ), .B(_05747_ ), .C1(_05427_ ), .C2(_05808_ ), .ZN(_05809_ ) );
NAND4_X1 _13764_ ( .A1(_04982_ ), .A2(_02268_ ), .A3(_05427_ ), .A4(_05381_ ), .ZN(_05810_ ) );
AND2_X1 _13765_ ( .A1(_05809_ ), .A2(_05810_ ), .ZN(_05811_ ) );
AOI21_X1 _13766_ ( .A(_05799_ ), .B1(_05800_ ), .B2(_05811_ ), .ZN(_05812_ ) );
BUF_X2 _13767_ ( .A(_05635_ ), .Z(_05813_ ) );
AOI21_X1 _13768_ ( .A(_05813_ ), .B1(_05809_ ), .B2(_05810_ ), .ZN(_05814_ ) );
OAI21_X1 _13769_ ( .A(_05423_ ), .B1(_05539_ ), .B2(_05540_ ), .ZN(_05815_ ) );
OAI211_X1 _13770_ ( .A(_05815_ ), .B(_05465_ ), .C1(_05744_ ), .C2(_05551_ ), .ZN(_05816_ ) );
OAI21_X1 _13771_ ( .A(_05428_ ), .B1(_05543_ ), .B2(_05544_ ), .ZN(_05817_ ) );
BUF_X2 _13772_ ( .A(_05425_ ), .Z(_05818_ ) );
NAND2_X1 _13773_ ( .A1(_05530_ ), .A2(_05532_ ), .ZN(_05819_ ) );
OAI211_X1 _13774_ ( .A(_05817_ ), .B(_05818_ ), .C1(_05552_ ), .C2(_05819_ ), .ZN(_05820_ ) );
AND2_X1 _13775_ ( .A1(_05158_ ), .A2(_05163_ ), .ZN(_05821_ ) );
BUF_X2 _13776_ ( .A(_05821_ ), .Z(_05822_ ) );
NAND3_X1 _13777_ ( .A1(_05816_ ), .A2(_05820_ ), .A3(_05822_ ), .ZN(_05823_ ) );
OAI221_X1 _13778_ ( .A(_05823_ ), .B1(_05273_ ), .B2(_05470_ ), .C1(_05268_ ), .C2(_05662_ ), .ZN(_05824_ ) );
NOR3_X1 _13779_ ( .A1(_05812_ ), .A2(_05814_ ), .A3(_05824_ ), .ZN(_05825_ ) );
OAI21_X1 _13780_ ( .A(_05278_ ), .B1(_05298_ ), .B2(_05306_ ), .ZN(_05826_ ) );
AND2_X1 _13781_ ( .A1(_05261_ ), .A2(_05253_ ), .ZN(_05827_ ) );
AND2_X1 _13782_ ( .A1(_05826_ ), .A2(_05827_ ), .ZN(_05828_ ) );
INV_X1 _13783_ ( .A(_05828_ ), .ZN(_05829_ ) );
NAND2_X1 _13784_ ( .A1(_05829_ ), .A2(_05245_ ), .ZN(_05830_ ) );
AOI21_X1 _13785_ ( .A(_05269_ ), .B1(_05830_ ), .B2(_05267_ ), .ZN(_05831_ ) );
INV_X1 _13786_ ( .A(_05831_ ), .ZN(_05832_ ) );
AOI21_X1 _13787_ ( .A(_05246_ ), .B1(_05832_ ), .B2(_05272_ ), .ZN(_05833_ ) );
NOR3_X1 _13788_ ( .A1(_05831_ ), .A2(_05268_ ), .A3(_05271_ ), .ZN(_05834_ ) );
OAI21_X1 _13789_ ( .A(_05479_ ), .B1(_05833_ ), .B2(_05834_ ), .ZN(_05835_ ) );
OR3_X1 _13790_ ( .A1(_05099_ ), .A2(_04766_ ), .A3(_05340_ ), .ZN(_05836_ ) );
NAND3_X1 _13791_ ( .A1(_05825_ ), .A2(_05835_ ), .A3(_05836_ ), .ZN(_05837_ ) );
AOI21_X1 _13792_ ( .A(_05798_ ), .B1(_05365_ ), .B2(_05837_ ), .ZN(_05838_ ) );
NAND3_X1 _13793_ ( .A1(_05498_ ), .A2(\ID_EX_pc [14] ), .A3(_05720_ ), .ZN(_05839_ ) );
NAND2_X1 _13794_ ( .A1(_05839_ ), .A2(\ID_EX_pc [15] ), .ZN(_05840_ ) );
NAND4_X1 _13795_ ( .A1(_05498_ ), .A2(_02332_ ), .A3(\ID_EX_pc [14] ), .A4(_05720_ ), .ZN(_05841_ ) );
NAND3_X1 _13796_ ( .A1(_05840_ ), .A2(_05497_ ), .A3(_05841_ ), .ZN(_05842_ ) );
NAND2_X1 _13797_ ( .A1(_05842_ ), .A2(_03407_ ), .ZN(_05843_ ) );
OAI21_X1 _13798_ ( .A(_05773_ ), .B1(_05838_ ), .B2(_05843_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
INV_X1 _13799_ ( .A(_03813_ ), .ZN(_05844_ ) );
XNOR2_X1 _13800_ ( .A(_05721_ ), .B(_02333_ ), .ZN(_05845_ ) );
OR3_X1 _13801_ ( .A1(_05778_ ), .A2(_04768_ ), .A3(_04830_ ), .ZN(_05846_ ) );
AND3_X1 _13802_ ( .A1(_05846_ ), .A2(_05514_ ), .A3(_05779_ ), .ZN(_05847_ ) );
AOI21_X1 _13803_ ( .A(_04955_ ), .B1(_05791_ ), .B2(_04870_ ), .ZN(_05848_ ) );
OAI21_X1 _13804_ ( .A(_05848_ ), .B1(_04870_ ), .B2(_05791_ ), .ZN(_05849_ ) );
NAND3_X1 _13805_ ( .A1(_04962_ ), .A2(\ID_EX_imm [14] ), .A3(_04964_ ), .ZN(_05850_ ) );
NAND2_X1 _13806_ ( .A1(_05849_ ), .A2(_05850_ ), .ZN(_05851_ ) );
OAI21_X1 _13807_ ( .A(_04759_ ), .B1(_05847_ ), .B2(_05851_ ), .ZN(_05852_ ) );
NAND3_X1 _13808_ ( .A1(_05830_ ), .A2(_05269_ ), .A3(_05267_ ), .ZN(_05853_ ) );
AND3_X1 _13809_ ( .A1(_05832_ ), .A2(_05239_ ), .A3(_05853_ ), .ZN(_05854_ ) );
AOI21_X1 _13810_ ( .A(_05113_ ), .B1(_05613_ ), .B2(_05614_ ), .ZN(_05855_ ) );
OR3_X1 _13811_ ( .A1(_05440_ ), .A2(_05134_ ), .A3(_05438_ ), .ZN(_05856_ ) );
OR3_X1 _13812_ ( .A1(_05447_ ), .A2(_05441_ ), .A3(_05127_ ), .ZN(_05857_ ) );
AOI21_X1 _13813_ ( .A(_05125_ ), .B1(_05856_ ), .B2(_05857_ ), .ZN(_05858_ ) );
NOR3_X1 _13814_ ( .A1(_05855_ ), .A2(_05858_ ), .A3(_04985_ ), .ZN(_05859_ ) );
NOR2_X1 _13815_ ( .A1(_05623_ ), .A2(_05113_ ), .ZN(_05860_ ) );
AOI21_X1 _13816_ ( .A(_05125_ ), .B1(_05616_ ), .B2(_05618_ ), .ZN(_05861_ ) );
NOR2_X1 _13817_ ( .A1(_05860_ ), .A2(_05861_ ), .ZN(_05862_ ) );
AOI211_X1 _13818_ ( .A(_05231_ ), .B(_05859_ ), .C1(_05409_ ), .C2(_05862_ ), .ZN(_05863_ ) );
AND3_X1 _13819_ ( .A1(_05406_ ), .A2(_04981_ ), .A3(_05184_ ), .ZN(_05864_ ) );
AND3_X1 _13820_ ( .A1(_05864_ ), .A2(_05193_ ), .A3(_05231_ ), .ZN(_05865_ ) );
NOR2_X1 _13821_ ( .A1(_05863_ ), .A2(_05865_ ), .ZN(_05866_ ) );
NOR2_X1 _13822_ ( .A1(_05866_ ), .A2(_05635_ ), .ZN(_05867_ ) );
INV_X1 _13823_ ( .A(_05821_ ), .ZN(_05868_ ) );
NAND2_X1 _13824_ ( .A1(_05637_ ), .A2(_05638_ ), .ZN(_05869_ ) );
NAND2_X1 _13825_ ( .A1(_05869_ ), .A2(_05399_ ), .ZN(_05870_ ) );
NAND2_X1 _13826_ ( .A1(_05648_ ), .A2(_05369_ ), .ZN(_05871_ ) );
NAND3_X1 _13827_ ( .A1(_05870_ ), .A2(_05409_ ), .A3(_05871_ ), .ZN(_05872_ ) );
NAND3_X1 _13828_ ( .A1(_05654_ ), .A2(_05369_ ), .A3(_05655_ ), .ZN(_05873_ ) );
NAND2_X1 _13829_ ( .A1(_05644_ ), .A2(_05399_ ), .ZN(_05874_ ) );
NAND3_X1 _13830_ ( .A1(_05873_ ), .A2(_05425_ ), .A3(_05874_ ), .ZN(_05875_ ) );
AOI21_X1 _13831_ ( .A(_05868_ ), .B1(_05872_ ), .B2(_05875_ ), .ZN(_05876_ ) );
OAI22_X1 _13832_ ( .A1(_05269_ ), .A2(_05661_ ), .B1(_05272_ ), .B2(_05339_ ), .ZN(_05877_ ) );
OR4_X1 _13833_ ( .A1(_05854_ ), .A2(_05867_ ), .A3(_05876_ ), .A4(_05877_ ), .ZN(_05878_ ) );
AND2_X1 _13834_ ( .A1(_05610_ ), .A2(_04981_ ), .ZN(_05879_ ) );
AND2_X1 _13835_ ( .A1(_05115_ ), .A2(_05879_ ), .ZN(_05880_ ) );
INV_X1 _13836_ ( .A(_05880_ ), .ZN(_05881_ ) );
NAND4_X1 _13837_ ( .A1(_05108_ ), .A2(_05119_ ), .A3(_05120_ ), .A4(_05881_ ), .ZN(_05882_ ) );
AOI21_X1 _13838_ ( .A(_04970_ ), .B1(_05882_ ), .B2(_05866_ ), .ZN(_05883_ ) );
AOI21_X1 _13839_ ( .A(_05470_ ), .B1(_05100_ ), .B2(_03814_ ), .ZN(_05884_ ) );
NOR3_X1 _13840_ ( .A1(_05878_ ), .A2(_05883_ ), .A3(_05884_ ), .ZN(_05885_ ) );
OAI21_X1 _13841_ ( .A(_05852_ ), .B1(_05885_ ), .B2(_05357_ ), .ZN(_05886_ ) );
MUX2_X1 _13842_ ( .A(_05845_ ), .B(_05886_ ), .S(_05360_ ), .Z(_05887_ ) );
MUX2_X1 _13843_ ( .A(_05844_ ), .B(_05887_ ), .S(_03390_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
OR2_X1 _13844_ ( .A1(_03848_ ), .A2(_05362_ ), .ZN(_05888_ ) );
NAND2_X1 _13845_ ( .A1(_05243_ ), .A2(_05472_ ), .ZN(_05889_ ) );
AND2_X1 _13846_ ( .A1(_05690_ ), .A2(_05691_ ), .ZN(_05890_ ) );
OAI211_X1 _13847_ ( .A(_05205_ ), .B(_05134_ ), .C1(_01969_ ), .C2(_05110_ ), .ZN(_05891_ ) );
OAI211_X1 _13848_ ( .A(_05188_ ), .B(_05127_ ), .C1(_01738_ ), .C2(_05110_ ), .ZN(_05892_ ) );
NAND2_X1 _13849_ ( .A1(_05891_ ), .A2(_05892_ ), .ZN(_05893_ ) );
MUX2_X1 _13850_ ( .A(_05890_ ), .B(_05893_ ), .S(_04981_ ), .Z(_05894_ ) );
OR2_X1 _13851_ ( .A1(_05894_ ), .A2(_05408_ ), .ZN(_05895_ ) );
OAI211_X1 _13852_ ( .A(_05895_ ), .B(_05165_ ), .C1(_05818_ ), .C2(_05156_ ), .ZN(_05896_ ) );
NAND3_X1 _13853_ ( .A1(_05136_ ), .A2(_05818_ ), .A3(_05232_ ), .ZN(_05897_ ) );
AOI21_X1 _13854_ ( .A(_05813_ ), .B1(_05896_ ), .B2(_05897_ ), .ZN(_05898_ ) );
AND2_X1 _13855_ ( .A1(_05114_ ), .A2(_05193_ ), .ZN(_05899_ ) );
OR4_X4 _13856_ ( .A1(_05376_ ), .A2(_05109_ ), .A3(_05728_ ), .A4(_05899_ ), .ZN(_05900_ ) );
AND2_X1 _13857_ ( .A1(_05896_ ), .A2(_05897_ ), .ZN(_05901_ ) );
AOI21_X1 _13858_ ( .A(_04970_ ), .B1(_05900_ ), .B2(_05901_ ), .ZN(_05902_ ) );
NAND3_X1 _13859_ ( .A1(_05224_ ), .A2(_05230_ ), .A3(_05452_ ), .ZN(_05903_ ) );
OAI21_X1 _13860_ ( .A(_05903_ ), .B1(_05192_ ), .B2(_05466_ ), .ZN(_05904_ ) );
AOI211_X1 _13861_ ( .A(_05898_ ), .B(_05902_ ), .C1(_05822_ ), .C2(_05904_ ), .ZN(_05905_ ) );
OAI21_X1 _13862_ ( .A(_05580_ ), .B1(_05266_ ), .B2(_03850_ ), .ZN(_05906_ ) );
NAND3_X1 _13863_ ( .A1(_05266_ ), .A2(_03850_ ), .A3(_05476_ ), .ZN(_05907_ ) );
AND4_X1 _13864_ ( .A1(_05889_ ), .A2(_05905_ ), .A3(_05906_ ), .A4(_05907_ ), .ZN(_05908_ ) );
INV_X1 _13865_ ( .A(_05244_ ), .ZN(_05909_ ) );
AOI21_X1 _13866_ ( .A(_05909_ ), .B1(_05826_ ), .B2(_05827_ ), .ZN(_05910_ ) );
NOR2_X1 _13867_ ( .A1(_05910_ ), .A2(_05264_ ), .ZN(_05911_ ) );
XNOR2_X1 _13868_ ( .A(_05911_ ), .B(_05243_ ), .ZN(_05912_ ) );
NAND2_X1 _13869_ ( .A1(_05912_ ), .A2(_05479_ ), .ZN(_05913_ ) );
AOI21_X1 _13870_ ( .A(_05528_ ), .B1(_05908_ ), .B2(_05913_ ), .ZN(_05914_ ) );
AND2_X1 _13871_ ( .A1(_05777_ ), .A2(_04824_ ), .ZN(_05915_ ) );
OR2_X1 _13872_ ( .A1(_05915_ ), .A2(_05775_ ), .ZN(_05916_ ) );
AND3_X1 _13873_ ( .A1(_05916_ ), .A2(_04829_ ), .A3(_05774_ ), .ZN(_05917_ ) );
AOI21_X1 _13874_ ( .A(_05774_ ), .B1(_05916_ ), .B2(_04829_ ), .ZN(_05918_ ) );
OR3_X1 _13875_ ( .A1(_05917_ ), .A2(_05918_ ), .A3(_04867_ ), .ZN(_05919_ ) );
OR3_X1 _13876_ ( .A1(_05789_ ), .A2(_04917_ ), .A3(_04874_ ), .ZN(_05920_ ) );
OAI21_X1 _13877_ ( .A(_04874_ ), .B1(_05789_ ), .B2(_04917_ ), .ZN(_05921_ ) );
NAND3_X1 _13878_ ( .A1(_05920_ ), .A2(_05672_ ), .A3(_05921_ ), .ZN(_05922_ ) );
NAND3_X1 _13879_ ( .A1(_05491_ ), .A2(\ID_EX_imm [13] ), .A3(_05492_ ), .ZN(_05923_ ) );
AND2_X1 _13880_ ( .A1(_05922_ ), .A2(_05923_ ), .ZN(_05924_ ) );
AOI21_X1 _13881_ ( .A(_05509_ ), .B1(_05919_ ), .B2(_05924_ ), .ZN(_05925_ ) );
NOR3_X1 _13882_ ( .A1(_05914_ ), .A2(_05925_ ), .A3(_01362_ ), .ZN(_05926_ ) );
NAND4_X1 _13883_ ( .A1(_05498_ ), .A2(_02334_ ), .A3(\ID_EX_pc [12] ), .A4(_04752_ ), .ZN(_05927_ ) );
NAND3_X1 _13884_ ( .A1(_04749_ ), .A2(\ID_EX_pc [9] ), .A3(_04752_ ), .ZN(_05928_ ) );
OAI21_X1 _13885_ ( .A(\ID_EX_pc [13] ), .B1(_05928_ ), .B2(_02335_ ), .ZN(_05929_ ) );
NAND3_X1 _13886_ ( .A1(_05927_ ), .A2(_05497_ ), .A3(_05929_ ), .ZN(_05930_ ) );
NAND2_X1 _13887_ ( .A1(_05930_ ), .A2(_03407_ ), .ZN(_05931_ ) );
OAI21_X1 _13888_ ( .A(_05888_ ), .B1(_05926_ ), .B2(_05931_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
INV_X1 _13889_ ( .A(_03890_ ), .ZN(_05932_ ) );
OAI211_X1 _13890_ ( .A(_05122_ ), .B(_05119_ ), .C1(_05466_ ), .C2(_05373_ ), .ZN(_05933_ ) );
AOI21_X1 _13891_ ( .A(_05804_ ), .B1(_05390_ ), .B2(_05400_ ), .ZN(_05934_ ) );
OR3_X1 _13892_ ( .A1(_05437_ ), .A2(_05197_ ), .A3(_05430_ ), .ZN(_05935_ ) );
OR3_X1 _13893_ ( .A1(_05440_ ), .A2(_05438_ ), .A3(_05184_ ), .ZN(_05936_ ) );
NAND3_X1 _13894_ ( .A1(_05935_ ), .A2(_05180_ ), .A3(_05936_ ), .ZN(_05937_ ) );
NAND3_X1 _13895_ ( .A1(_05734_ ), .A2(_05735_ ), .A3(_05182_ ), .ZN(_05938_ ) );
AOI21_X1 _13896_ ( .A(_05452_ ), .B1(_05937_ ), .B2(_05938_ ), .ZN(_05939_ ) );
NOR3_X1 _13897_ ( .A1(_05934_ ), .A2(_05939_ ), .A3(_05381_ ), .ZN(_05940_ ) );
AND4_X1 _13898_ ( .A1(_05427_ ), .A2(_05407_ ), .A3(_05700_ ), .A4(_05380_ ), .ZN(_05941_ ) );
NOR2_X1 _13899_ ( .A1(_05940_ ), .A2(_05941_ ), .ZN(_05942_ ) );
AOI21_X1 _13900_ ( .A(_05799_ ), .B1(_05933_ ), .B2(_05942_ ), .ZN(_05943_ ) );
NOR2_X1 _13901_ ( .A1(_05910_ ), .A2(_05709_ ), .ZN(_05944_ ) );
OAI21_X1 _13902_ ( .A(_05944_ ), .B1(_05244_ ), .B2(_05829_ ), .ZN(_05945_ ) );
OAI21_X1 _13903_ ( .A(_05474_ ), .B1(_05940_ ), .B2(_05941_ ), .ZN(_05946_ ) );
INV_X1 _13904_ ( .A(_05088_ ), .ZN(_05947_ ) );
NAND3_X1 _13905_ ( .A1(_05947_ ), .A2(_01808_ ), .A3(_05476_ ), .ZN(_05948_ ) );
AOI21_X1 _13906_ ( .A(_05344_ ), .B1(_05088_ ), .B2(_04763_ ), .ZN(_05949_ ) );
OAI21_X1 _13907_ ( .A(_05818_ ), .B1(_05424_ ), .B2(_05435_ ), .ZN(_05950_ ) );
OAI21_X1 _13908_ ( .A(_05950_ ), .B1(_05464_ ), .B2(_05426_ ), .ZN(_05951_ ) );
AOI221_X4 _13909_ ( .A(_05949_ ), .B1(_05244_ ), .B2(_05335_ ), .C1(_05951_ ), .C2(_05822_ ), .ZN(_05952_ ) );
NAND4_X1 _13910_ ( .A1(_05945_ ), .A2(_05946_ ), .A3(_05948_ ), .A4(_05952_ ), .ZN(_05953_ ) );
OAI21_X1 _13911_ ( .A(_05365_ ), .B1(_05943_ ), .B2(_05953_ ), .ZN(_05954_ ) );
NAND3_X1 _13912_ ( .A1(_05777_ ), .A2(_05775_ ), .A3(_04824_ ), .ZN(_05955_ ) );
AND3_X1 _13913_ ( .A1(_05916_ ), .A2(_05515_ ), .A3(_05955_ ), .ZN(_05956_ ) );
OR3_X1 _13914_ ( .A1(_05786_ ), .A2(_04875_ ), .A3(_04927_ ), .ZN(_05957_ ) );
NAND3_X1 _13915_ ( .A1(_05790_ ), .A2(_05672_ ), .A3(_05957_ ), .ZN(_05958_ ) );
NAND3_X1 _13916_ ( .A1(_05524_ ), .A2(\ID_EX_imm [12] ), .A3(_05525_ ), .ZN(_05959_ ) );
NAND2_X1 _13917_ ( .A1(_05958_ ), .A2(_05959_ ), .ZN(_05960_ ) );
OAI21_X1 _13918_ ( .A(_04759_ ), .B1(_05956_ ), .B2(_05960_ ), .ZN(_05961_ ) );
AND3_X1 _13919_ ( .A1(_05954_ ), .A2(_05484_ ), .A3(_05961_ ), .ZN(_05962_ ) );
XNOR2_X1 _13920_ ( .A(_05928_ ), .B(\ID_EX_pc [12] ), .ZN(_05963_ ) );
OAI21_X1 _13921_ ( .A(_04248_ ), .B1(_05963_ ), .B2(_05725_ ), .ZN(_05964_ ) );
OAI21_X1 _13922_ ( .A(_05932_ ), .B1(_05962_ ), .B2(_05964_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
INV_X1 _13923_ ( .A(_03947_ ), .ZN(_05965_ ) );
AND3_X1 _13924_ ( .A1(_04750_ ), .A2(\ID_EX_pc [11] ), .A3(\ID_EX_pc [10] ), .ZN(_05966_ ) );
AND3_X1 _13925_ ( .A1(_05966_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_05967_ ) );
AND3_X1 _13926_ ( .A1(_05967_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05968_ ) );
AND3_X1 _13927_ ( .A1(_05968_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_05969_ ) );
AND3_X1 _13928_ ( .A1(_05969_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_05970_ ) );
AND3_X1 _13929_ ( .A1(_05970_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05971_ ) );
AND3_X1 _13930_ ( .A1(_05971_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_05972_ ) );
AND3_X1 _13931_ ( .A1(_05972_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_05973_ ) );
AND3_X1 _13932_ ( .A1(_05973_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_05974_ ) );
AND3_X1 _13933_ ( .A1(_05974_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_05975_ ) );
XNOR2_X1 _13934_ ( .A(_05975_ ), .B(_02325_ ), .ZN(_05976_ ) );
XOR2_X1 _13935_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_05977_ ) );
INV_X1 _13936_ ( .A(_05977_ ), .ZN(_05978_ ) );
XOR2_X1 _13937_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_05979_ ) );
XOR2_X1 _13938_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_05980_ ) );
AND2_X1 _13939_ ( .A1(_05979_ ), .A2(_05980_ ), .ZN(_05981_ ) );
INV_X1 _13940_ ( .A(_05981_ ), .ZN(_05982_ ) );
NOR4_X1 _13941_ ( .A1(_04945_ ), .A2(_04947_ ), .A3(_04958_ ), .A4(_05982_ ), .ZN(_05983_ ) );
AND2_X1 _13942_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_05984_ ) );
AND2_X1 _13943_ ( .A1(_05979_ ), .A2(_05984_ ), .ZN(_05985_ ) );
AOI21_X1 _13944_ ( .A(_05985_ ), .B1(\ID_EX_pc [23] ), .B2(\ID_EX_imm [23] ), .ZN(_05986_ ) );
AOI21_X1 _13945_ ( .A(_04956_ ), .B1(\ID_EX_pc [21] ), .B2(\ID_EX_imm [21] ), .ZN(_05987_ ) );
OAI21_X1 _13946_ ( .A(_05986_ ), .B1(_05987_ ), .B2(_05982_ ), .ZN(_05988_ ) );
OR2_X1 _13947_ ( .A1(_05983_ ), .A2(_05988_ ), .ZN(_05989_ ) );
XOR2_X1 _13948_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_05990_ ) );
AND2_X1 _13949_ ( .A1(_05989_ ), .A2(_05990_ ), .ZN(_05991_ ) );
AND2_X1 _13950_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_05992_ ) );
AND2_X1 _13951_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_05993_ ) );
OR3_X1 _13952_ ( .A1(_05991_ ), .A2(_05992_ ), .A3(_05993_ ), .ZN(_05994_ ) );
XOR2_X1 _13953_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_05995_ ) );
XOR2_X1 _13954_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_05996_ ) );
NOR2_X1 _13955_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_05997_ ) );
INV_X1 _13956_ ( .A(_05997_ ), .ZN(_05998_ ) );
NAND4_X1 _13957_ ( .A1(_05994_ ), .A2(_05995_ ), .A3(_05996_ ), .A4(_05998_ ), .ZN(_05999_ ) );
AND2_X1 _13958_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_06000_ ) );
AND2_X1 _13959_ ( .A1(_05995_ ), .A2(_06000_ ), .ZN(_06001_ ) );
AOI21_X1 _13960_ ( .A(_06001_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_06002_ ) );
AOI21_X1 _13961_ ( .A(_05978_ ), .B1(_05999_ ), .B2(_06002_ ), .ZN(_06003_ ) );
AND2_X1 _13962_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_06004_ ) );
OAI22_X1 _13963_ ( .A1(_06003_ ), .A2(_06004_ ), .B1(\ID_EX_pc [29] ), .B2(\ID_EX_imm [29] ), .ZN(_06005_ ) );
INV_X1 _13964_ ( .A(\ID_EX_imm [29] ), .ZN(_06006_ ) );
OAI21_X1 _13965_ ( .A(_06005_ ), .B1(_02336_ ), .B2(_06006_ ), .ZN(_06007_ ) );
XOR2_X1 _13966_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_06008_ ) );
AOI21_X1 _13967_ ( .A(_04955_ ), .B1(_06007_ ), .B2(_06008_ ), .ZN(_06009_ ) );
OAI21_X1 _13968_ ( .A(_06009_ ), .B1(_06008_ ), .B2(_06007_ ), .ZN(_06010_ ) );
NAND3_X1 _13969_ ( .A1(_04962_ ), .A2(\ID_EX_imm [30] ), .A3(_04964_ ), .ZN(_06011_ ) );
NAND2_X1 _13970_ ( .A1(_06010_ ), .A2(_06011_ ), .ZN(_06012_ ) );
XNOR2_X1 _13971_ ( .A(_04488_ ), .B(_02236_ ), .ZN(_06013_ ) );
XNOR2_X1 _13972_ ( .A(_04382_ ), .B(_02214_ ), .ZN(_06014_ ) );
XNOR2_X1 _13973_ ( .A(_04524_ ), .B(_01472_ ), .ZN(_06015_ ) );
INV_X1 _13974_ ( .A(_06015_ ), .ZN(_06016_ ) );
XNOR2_X1 _13975_ ( .A(_04557_ ), .B(_02182_ ), .ZN(_06017_ ) );
INV_X1 _13976_ ( .A(_06017_ ), .ZN(_06018_ ) );
XNOR2_X1 _13977_ ( .A(_05385_ ), .B(_04668_ ), .ZN(_06019_ ) );
XNOR2_X1 _13978_ ( .A(_05147_ ), .B(_04704_ ), .ZN(_06020_ ) );
AND2_X1 _13979_ ( .A1(_06019_ ), .A2(_06020_ ), .ZN(_06021_ ) );
NAND4_X4 _13980_ ( .A1(_04854_ ), .A2(_04858_ ), .A3(_04856_ ), .A4(_06021_ ), .ZN(_06022_ ) );
AND3_X1 _13981_ ( .A1(_04858_ ), .A2(_02088_ ), .A3(_03589_ ), .ZN(_06023_ ) );
NOR2_X1 _13982_ ( .A1(_03524_ ), .A2(_05337_ ), .ZN(_06024_ ) );
OAI21_X1 _13983_ ( .A(_06021_ ), .B1(_06023_ ), .B2(_06024_ ), .ZN(_06025_ ) );
AND2_X1 _13984_ ( .A1(_04668_ ), .A2(_02042_ ), .ZN(_06026_ ) );
INV_X1 _13985_ ( .A(_06026_ ), .ZN(_06027_ ) );
AND2_X1 _13986_ ( .A1(_04704_ ), .A2(_02064_ ), .ZN(_06028_ ) );
NAND2_X1 _13987_ ( .A1(_06019_ ), .A2(_06028_ ), .ZN(_06029_ ) );
AND3_X1 _13988_ ( .A1(_06025_ ), .A2(_06027_ ), .A3(_06029_ ), .ZN(_06030_ ) );
NAND2_X4 _13989_ ( .A1(_06022_ ), .A2(_06030_ ), .ZN(_06031_ ) );
XNOR2_X1 _13990_ ( .A(_04593_ ), .B(_02158_ ), .ZN(_06032_ ) );
XNOR2_X1 _13991_ ( .A(_04631_ ), .B(_01496_ ), .ZN(_06033_ ) );
NAND3_X4 _13992_ ( .A1(_06031_ ), .A2(_06032_ ), .A3(_06033_ ), .ZN(_06034_ ) );
NOR2_X1 _13993_ ( .A1(_04631_ ), .A2(_05151_ ), .ZN(_06035_ ) );
AND2_X1 _13994_ ( .A1(_06032_ ), .A2(_06035_ ), .ZN(_06036_ ) );
AOI21_X1 _13995_ ( .A(_06036_ ), .B1(_02158_ ), .B2(_04594_ ), .ZN(_06037_ ) );
AOI211_X2 _13996_ ( .A(_06016_ ), .B(_06018_ ), .C1(_06034_ ), .C2(_06037_ ), .ZN(_06038_ ) );
NOR2_X1 _13997_ ( .A1(_04557_ ), .A2(_05137_ ), .ZN(_06039_ ) );
NAND2_X1 _13998_ ( .A1(_06015_ ), .A2(_06039_ ), .ZN(_06040_ ) );
OAI21_X1 _13999_ ( .A(_06040_ ), .B1(_04490_ ), .B2(_04524_ ), .ZN(_06041_ ) );
OAI211_X1 _14000_ ( .A(_06013_ ), .B(_06014_ ), .C1(_06038_ ), .C2(_06041_ ), .ZN(_06042_ ) );
NAND3_X1 _14001_ ( .A1(_02214_ ), .A2(_04362_ ), .A3(_04381_ ), .ZN(_06043_ ) );
NAND4_X1 _14002_ ( .A1(_06014_ ), .A2(_02236_ ), .A3(_04487_ ), .A4(_04468_ ), .ZN(_06044_ ) );
AND3_X2 _14003_ ( .A1(_06042_ ), .A2(_06043_ ), .A3(_06044_ ), .ZN(_06045_ ) );
XNOR2_X1 _14004_ ( .A(_03935_ ), .B(_01446_ ), .ZN(_06046_ ) );
OR2_X4 _14005_ ( .A1(_06045_ ), .A2(_06046_ ), .ZN(_06047_ ) );
AOI21_X1 _14006_ ( .A(_04866_ ), .B1(_06045_ ), .B2(_06046_ ), .ZN(_06048_ ) );
AND2_X4 _14007_ ( .A1(_06047_ ), .A2(_06048_ ), .ZN(_06049_ ) );
OAI21_X4 _14008_ ( .A(_04758_ ), .B1(_06012_ ), .B2(_06049_ ), .ZN(_06050_ ) );
AND4_X1 _14009_ ( .A1(_05019_ ), .A2(_05106_ ), .A3(_05123_ ), .A4(_05881_ ), .ZN(_06051_ ) );
AND3_X1 _14010_ ( .A1(_05864_ ), .A2(_04986_ ), .A3(_04990_ ), .ZN(_06052_ ) );
OR2_X1 _14011_ ( .A1(_06051_ ), .A2(_06052_ ), .ZN(_06053_ ) );
OAI21_X1 _14012_ ( .A(_04969_ ), .B1(_05556_ ), .B2(_06053_ ), .ZN(_06054_ ) );
AOI21_X1 _14013_ ( .A(_05159_ ), .B1(_05872_ ), .B2(_05875_ ), .ZN(_06055_ ) );
OR3_X1 _14014_ ( .A1(_05402_ ), .A2(_05219_ ), .A3(_05405_ ), .ZN(_06056_ ) );
NOR2_X1 _14015_ ( .A1(_05395_ ), .A2(_05403_ ), .ZN(_06057_ ) );
INV_X1 _14016_ ( .A(_06057_ ), .ZN(_06058_ ) );
OAI211_X1 _14017_ ( .A(_06056_ ), .B(_05423_ ), .C1(_05444_ ), .C2(_06058_ ), .ZN(_06059_ ) );
OR3_X1 _14018_ ( .A1(_05392_ ), .A2(_05168_ ), .A3(_05396_ ), .ZN(_06060_ ) );
OR3_X1 _14019_ ( .A1(_05386_ ), .A2(_05393_ ), .A3(_05177_ ), .ZN(_06061_ ) );
NAND3_X1 _14020_ ( .A1(_06060_ ), .A2(_06061_ ), .A3(_05428_ ), .ZN(_06062_ ) );
NAND3_X1 _14021_ ( .A1(_06059_ ), .A2(_05194_ ), .A3(_06062_ ), .ZN(_06063_ ) );
NAND3_X1 _14022_ ( .A1(_05651_ ), .A2(_05652_ ), .A3(_05399_ ), .ZN(_06064_ ) );
OAI21_X1 _14023_ ( .A(_05177_ ), .B1(_05382_ ), .B2(_05387_ ), .ZN(_06065_ ) );
OAI21_X1 _14024_ ( .A(_05168_ ), .B1(_05445_ ), .B2(_05383_ ), .ZN(_06066_ ) );
NAND2_X1 _14025_ ( .A1(_06065_ ), .A2(_06066_ ), .ZN(_06067_ ) );
NAND2_X1 _14026_ ( .A1(_06067_ ), .A2(_05369_ ), .ZN(_06068_ ) );
NAND3_X1 _14027_ ( .A1(_06064_ ), .A2(_06068_ ), .A3(_05451_ ), .ZN(_06069_ ) );
AOI21_X1 _14028_ ( .A(_05232_ ), .B1(_06063_ ), .B2(_06069_ ), .ZN(_06070_ ) );
OAI21_X1 _14029_ ( .A(_05413_ ), .B1(_06055_ ), .B2(_06070_ ), .ZN(_06071_ ) );
OAI21_X1 _14030_ ( .A(_05580_ ), .B1(_05055_ ), .B2(_03949_ ), .ZN(_06072_ ) );
AND2_X1 _14031_ ( .A1(_06052_ ), .A2(_05235_ ), .ZN(_06073_ ) );
AOI21_X1 _14032_ ( .A(_01446_ ), .B1(_05053_ ), .B2(_05054_ ), .ZN(_06074_ ) );
AND3_X1 _14033_ ( .A1(_05053_ ), .A2(_01446_ ), .A3(_05054_ ), .ZN(_06075_ ) );
NOR2_X1 _14034_ ( .A1(_06075_ ), .A2(_06074_ ), .ZN(_06076_ ) );
AOI221_X4 _14035_ ( .A(_06073_ ), .B1(_05475_ ), .B2(_06074_ ), .C1(_05334_ ), .C2(_06076_ ), .ZN(_06077_ ) );
NAND4_X1 _14036_ ( .A1(_06054_ ), .A2(_06071_ ), .A3(_06072_ ), .A4(_06077_ ), .ZN(_06078_ ) );
XNOR2_X1 _14037_ ( .A(_05058_ ), .B(_02308_ ), .ZN(_06079_ ) );
NAND2_X1 _14038_ ( .A1(_05059_ ), .A2(_05060_ ), .ZN(_06080_ ) );
XNOR2_X1 _14039_ ( .A(_06080_ ), .B(_04348_ ), .ZN(_06081_ ) );
NAND2_X1 _14040_ ( .A1(_06079_ ), .A2(_06081_ ), .ZN(_06082_ ) );
INV_X2 _14041_ ( .A(_05480_ ), .ZN(_06083_ ) );
AND2_X1 _14042_ ( .A1(_05062_ ), .A2(_05061_ ), .ZN(_06084_ ) );
XNOR2_X1 _14043_ ( .A(_06084_ ), .B(_02042_ ), .ZN(_06085_ ) );
XNOR2_X1 _14044_ ( .A(_05048_ ), .B(_02064_ ), .ZN(_06086_ ) );
AND2_X1 _14045_ ( .A1(_06085_ ), .A2(_06086_ ), .ZN(_06087_ ) );
AND2_X1 _14046_ ( .A1(_05328_ ), .A2(_05241_ ), .ZN(_06088_ ) );
NAND3_X2 _14047_ ( .A1(_06083_ ), .A2(_06087_ ), .A3(_06088_ ), .ZN(_06089_ ) );
NAND2_X1 _14048_ ( .A1(_05328_ ), .A2(_05330_ ), .ZN(_06090_ ) );
OAI21_X1 _14049_ ( .A(_06090_ ), .B1(_05337_ ), .B2(_05067_ ), .ZN(_06091_ ) );
NAND2_X1 _14050_ ( .A1(_06091_ ), .A2(_06087_ ), .ZN(_06092_ ) );
OR2_X1 _14051_ ( .A1(_06084_ ), .A2(_05385_ ), .ZN(_06093_ ) );
NAND3_X1 _14052_ ( .A1(_06085_ ), .A2(_02064_ ), .A3(_05094_ ), .ZN(_06094_ ) );
AND3_X1 _14053_ ( .A1(_06092_ ), .A2(_06093_ ), .A3(_06094_ ), .ZN(_06095_ ) );
AND2_X2 _14054_ ( .A1(_06089_ ), .A2(_06095_ ), .ZN(_06096_ ) );
INV_X2 _14055_ ( .A(_06096_ ), .ZN(_06097_ ) );
XNOR2_X1 _14056_ ( .A(_05045_ ), .B(_01472_ ), .ZN(_06098_ ) );
NOR2_X1 _14057_ ( .A1(_05038_ ), .A2(_05137_ ), .ZN(_06099_ ) );
AOI21_X1 _14058_ ( .A(_02182_ ), .B1(_05036_ ), .B2(_05037_ ), .ZN(_06100_ ) );
NOR2_X1 _14059_ ( .A1(_06099_ ), .A2(_06100_ ), .ZN(_06101_ ) );
XNOR2_X1 _14060_ ( .A(_05051_ ), .B(_02158_ ), .ZN(_06102_ ) );
INV_X1 _14061_ ( .A(_06102_ ), .ZN(_06103_ ) );
NOR2_X1 _14062_ ( .A1(_05042_ ), .A2(_05151_ ), .ZN(_06104_ ) );
AOI21_X1 _14063_ ( .A(_01496_ ), .B1(_05040_ ), .B2(_05041_ ), .ZN(_06105_ ) );
NOR3_X1 _14064_ ( .A1(_06103_ ), .A2(_06104_ ), .A3(_06105_ ), .ZN(_06106_ ) );
NAND4_X4 _14065_ ( .A1(_06097_ ), .A2(_06098_ ), .A3(_06101_ ), .A4(_06106_ ), .ZN(_06107_ ) );
AND2_X1 _14066_ ( .A1(_06099_ ), .A2(_06098_ ), .ZN(_06108_ ) );
NOR2_X1 _14067_ ( .A1(_05051_ ), .A2(_05391_ ), .ZN(_06109_ ) );
AND2_X1 _14068_ ( .A1(_05051_ ), .A2(_05391_ ), .ZN(_06110_ ) );
INV_X1 _14069_ ( .A(_06110_ ), .ZN(_06111_ ) );
AOI21_X1 _14070_ ( .A(_06109_ ), .B1(_06111_ ), .B2(_06104_ ), .ZN(_06112_ ) );
INV_X1 _14071_ ( .A(_06098_ ), .ZN(_06113_ ) );
INV_X1 _14072_ ( .A(_06101_ ), .ZN(_06114_ ) );
NOR3_X1 _14073_ ( .A1(_06112_ ), .A2(_06113_ ), .A3(_06114_ ), .ZN(_06115_ ) );
AOI211_X1 _14074_ ( .A(_06108_ ), .B(_06115_ ), .C1(_01472_ ), .C2(_05093_ ), .ZN(_06116_ ) );
AOI21_X2 _14075_ ( .A(_06082_ ), .B1(_06107_ ), .B2(_06116_ ), .ZN(_06117_ ) );
AND2_X1 _14076_ ( .A1(_05058_ ), .A2(_02236_ ), .ZN(_06118_ ) );
NAND2_X1 _14077_ ( .A1(_06118_ ), .A2(_06081_ ), .ZN(_06119_ ) );
AND2_X1 _14078_ ( .A1(_06080_ ), .A2(_02214_ ), .ZN(_06120_ ) );
INV_X1 _14079_ ( .A(_06120_ ), .ZN(_06121_ ) );
NAND2_X1 _14080_ ( .A1(_06119_ ), .A2(_06121_ ), .ZN(_06122_ ) );
NOR2_X2 _14081_ ( .A1(_06117_ ), .A2(_06122_ ), .ZN(_06123_ ) );
XNOR2_X2 _14082_ ( .A(_06123_ ), .B(_06076_ ), .ZN(_06124_ ) );
AOI21_X2 _14083_ ( .A(_06078_ ), .B1(_06124_ ), .B2(_05239_ ), .ZN(_06125_ ) );
OAI21_X2 _14084_ ( .A(_06050_ ), .B1(_06125_ ), .B2(_05357_ ), .ZN(_06126_ ) );
MUX2_X2 _14085_ ( .A(_05976_ ), .B(_06126_ ), .S(_05360_ ), .Z(_06127_ ) );
MUX2_X2 _14086_ ( .A(_05965_ ), .B(_06127_ ), .S(_03390_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
OR2_X1 _14087_ ( .A1(_03962_ ), .A2(_05362_ ), .ZN(_06128_ ) );
INV_X1 _14088_ ( .A(_04780_ ), .ZN(_06129_ ) );
AOI211_X1 _14089_ ( .A(_04817_ ), .B(_06129_ ), .C1(_04804_ ), .C2(_04813_ ), .ZN(_06130_ ) );
OAI21_X1 _14090_ ( .A(_04775_ ), .B1(_06130_ ), .B2(_04819_ ), .ZN(_06131_ ) );
INV_X1 _14091_ ( .A(_04822_ ), .ZN(_06132_ ) );
AND2_X1 _14092_ ( .A1(_06131_ ), .A2(_06132_ ), .ZN(_06133_ ) );
XNOR2_X1 _14093_ ( .A(_06133_ ), .B(_04773_ ), .ZN(_06134_ ) );
AND2_X1 _14094_ ( .A1(_06134_ ), .A2(_05515_ ), .ZN(_06135_ ) );
INV_X1 _14095_ ( .A(_04883_ ), .ZN(_06136_ ) );
OAI21_X1 _14096_ ( .A(_04881_ ), .B1(_04911_ ), .B2(_04912_ ), .ZN(_06137_ ) );
INV_X1 _14097_ ( .A(_04879_ ), .ZN(_06138_ ) );
AOI21_X1 _14098_ ( .A(_04878_ ), .B1(_06138_ ), .B2(_04923_ ), .ZN(_06139_ ) );
AOI21_X1 _14099_ ( .A(_06136_ ), .B1(_06137_ ), .B2(_06139_ ), .ZN(_06140_ ) );
OR3_X1 _14100_ ( .A1(_06140_ ), .A2(_04920_ ), .A3(_04882_ ), .ZN(_06141_ ) );
OAI21_X1 _14101_ ( .A(_04882_ ), .B1(_06140_ ), .B2(_04920_ ), .ZN(_06142_ ) );
NAND3_X1 _14102_ ( .A1(_06141_ ), .A2(_05672_ ), .A3(_06142_ ), .ZN(_06143_ ) );
NAND3_X1 _14103_ ( .A1(_05524_ ), .A2(\ID_EX_imm [11] ), .A3(_05525_ ), .ZN(_06144_ ) );
NAND2_X1 _14104_ ( .A1(_06143_ ), .A2(_06144_ ), .ZN(_06145_ ) );
OAI21_X1 _14105_ ( .A(_04759_ ), .B1(_06135_ ), .B2(_06145_ ), .ZN(_06146_ ) );
AND2_X2 _14106_ ( .A1(_05120_ ), .A2(_05118_ ), .ZN(_06147_ ) );
OAI211_X1 _14107_ ( .A(_05108_ ), .B(_06147_ ), .C1(_05368_ ), .C2(_05574_ ), .ZN(_06148_ ) );
AOI21_X1 _14108_ ( .A(_05804_ ), .B1(_05566_ ), .B2(_05570_ ), .ZN(_06149_ ) );
OAI21_X1 _14109_ ( .A(_05399_ ), .B1(_05801_ ), .B2(_05802_ ), .ZN(_06150_ ) );
OAI21_X1 _14110_ ( .A(_05420_ ), .B1(_05531_ ), .B2(_05185_ ), .ZN(_06151_ ) );
OAI21_X1 _14111_ ( .A(_05415_ ), .B1(_05529_ ), .B2(_05187_ ), .ZN(_06152_ ) );
NAND3_X1 _14112_ ( .A1(_06151_ ), .A2(_06152_ ), .A3(_05369_ ), .ZN(_06153_ ) );
AND3_X1 _14113_ ( .A1(_06150_ ), .A2(_05804_ ), .A3(_06153_ ), .ZN(_06154_ ) );
OAI21_X1 _14114_ ( .A(_05467_ ), .B1(_06149_ ), .B2(_06154_ ), .ZN(_06155_ ) );
AOI21_X1 _14115_ ( .A(_05451_ ), .B1(_05560_ ), .B2(_05561_ ), .ZN(_06156_ ) );
OR2_X1 _14116_ ( .A1(_06156_ ), .A2(_05747_ ), .ZN(_06157_ ) );
NAND2_X1 _14117_ ( .A1(_06155_ ), .A2(_06157_ ), .ZN(_06158_ ) );
AOI21_X1 _14118_ ( .A(_05799_ ), .B1(_06148_ ), .B2(_06158_ ), .ZN(_06159_ ) );
INV_X1 _14119_ ( .A(_05255_ ), .ZN(_06160_ ) );
OAI21_X1 _14120_ ( .A(_05277_ ), .B1(_05298_ ), .B2(_05306_ ), .ZN(_06161_ ) );
AOI21_X1 _14121_ ( .A(_05257_ ), .B1(_05258_ ), .B2(_05259_ ), .ZN(_06162_ ) );
AOI21_X1 _14122_ ( .A(_06160_ ), .B1(_06161_ ), .B2(_06162_ ), .ZN(_06163_ ) );
OR3_X1 _14123_ ( .A1(_06163_ ), .A2(_05252_ ), .A3(_05254_ ), .ZN(_06164_ ) );
OAI21_X1 _14124_ ( .A(_05254_ ), .B1(_06163_ ), .B2(_05252_ ), .ZN(_06165_ ) );
NAND3_X1 _14125_ ( .A1(_06164_ ), .A2(_05479_ ), .A3(_06165_ ), .ZN(_06166_ ) );
NAND3_X1 _14126_ ( .A1(_06155_ ), .A2(_05474_ ), .A3(_06157_ ), .ZN(_06167_ ) );
NAND2_X1 _14127_ ( .A1(_05251_ ), .A2(_05580_ ), .ZN(_06168_ ) );
NAND3_X1 _14128_ ( .A1(_05542_ ), .A2(_05546_ ), .A3(_05194_ ), .ZN(_06169_ ) );
OR3_X1 _14129_ ( .A1(_05551_ ), .A2(_05425_ ), .A3(_05399_ ), .ZN(_06170_ ) );
AOI21_X1 _14130_ ( .A(_05868_ ), .B1(_06169_ ), .B2(_06170_ ), .ZN(_06171_ ) );
AOI221_X4 _14131_ ( .A(_06171_ ), .B1(_05250_ ), .B2(_05475_ ), .C1(_05254_ ), .C2(_05335_ ), .ZN(_06172_ ) );
NAND4_X1 _14132_ ( .A1(_06166_ ), .A2(_06167_ ), .A3(_06168_ ), .A4(_06172_ ), .ZN(_06173_ ) );
OAI21_X1 _14133_ ( .A(_05364_ ), .B1(_06159_ ), .B2(_06173_ ), .ZN(_06174_ ) );
AND3_X1 _14134_ ( .A1(_06146_ ), .A2(_05484_ ), .A3(_06174_ ), .ZN(_06175_ ) );
AOI21_X1 _14135_ ( .A(_02337_ ), .B1(_05498_ ), .B2(\ID_EX_pc [10] ), .ZN(_06176_ ) );
AND4_X1 _14136_ ( .A1(_02337_ ), .A2(_04749_ ), .A3(\ID_EX_pc [10] ), .A4(\ID_EX_pc [9] ), .ZN(_06177_ ) );
OR3_X1 _14137_ ( .A1(_06176_ ), .A2(_05360_ ), .A3(_06177_ ), .ZN(_06178_ ) );
NAND2_X1 _14138_ ( .A1(_06178_ ), .A2(_03407_ ), .ZN(_06179_ ) );
OAI21_X1 _14139_ ( .A(_06128_ ), .B1(_06175_ ), .B2(_06179_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
AND2_X1 _14140_ ( .A1(_05108_ ), .A2(_05367_ ), .ZN(_06180_ ) );
NOR3_X1 _14141_ ( .A1(_05609_ ), .A2(_05610_ ), .A3(_05368_ ), .ZN(_06181_ ) );
OAI21_X1 _14142_ ( .A(_06147_ ), .B1(_06180_ ), .B2(_06181_ ), .ZN(_06182_ ) );
OR3_X1 _14143_ ( .A1(_05437_ ), .A2(_05213_ ), .A3(_05430_ ), .ZN(_06183_ ) );
OR3_X1 _14144_ ( .A1(_05429_ ), .A2(_05168_ ), .A3(_05433_ ), .ZN(_06184_ ) );
AOI21_X1 _14145_ ( .A(_05399_ ), .B1(_06183_ ), .B2(_06184_ ), .ZN(_06185_ ) );
AOI21_X1 _14146_ ( .A(_05180_ ), .B1(_05856_ ), .B2(_05857_ ), .ZN(_06186_ ) );
OR3_X1 _14147_ ( .A1(_06185_ ), .A2(_06186_ ), .A3(_05409_ ), .ZN(_06187_ ) );
OAI211_X1 _14148_ ( .A(_06187_ ), .B(_05159_ ), .C1(_05426_ ), .C2(_05620_ ), .ZN(_06188_ ) );
NAND3_X1 _14149_ ( .A1(_05627_ ), .A2(_05804_ ), .A3(_05380_ ), .ZN(_06189_ ) );
AND2_X1 _14150_ ( .A1(_06188_ ), .A2(_06189_ ), .ZN(_06190_ ) );
AOI21_X1 _14151_ ( .A(_05799_ ), .B1(_06182_ ), .B2(_06190_ ), .ZN(_06191_ ) );
AOI21_X1 _14152_ ( .A(_05813_ ), .B1(_06188_ ), .B2(_06189_ ), .ZN(_06192_ ) );
NAND3_X1 _14153_ ( .A1(_05645_ ), .A2(_05649_ ), .A3(_05818_ ), .ZN(_06193_ ) );
NAND4_X1 _14154_ ( .A1(_05637_ ), .A2(_05451_ ), .A3(_05370_ ), .A4(_05638_ ), .ZN(_06194_ ) );
AOI21_X1 _14155_ ( .A(_05868_ ), .B1(_06193_ ), .B2(_06194_ ), .ZN(_06195_ ) );
NOR3_X1 _14156_ ( .A1(_06191_ ), .A2(_06192_ ), .A3(_06195_ ), .ZN(_06196_ ) );
NAND2_X1 _14157_ ( .A1(_05255_ ), .A2(_05472_ ), .ZN(_06197_ ) );
INV_X1 _14158_ ( .A(_05025_ ), .ZN(_06198_ ) );
NAND3_X1 _14159_ ( .A1(_06198_ ), .A2(_01905_ ), .A3(_05475_ ), .ZN(_06199_ ) );
OAI21_X1 _14160_ ( .A(_05580_ ), .B1(_06198_ ), .B2(_01905_ ), .ZN(_06200_ ) );
AND3_X1 _14161_ ( .A1(_06197_ ), .A2(_06199_ ), .A3(_06200_ ), .ZN(_06201_ ) );
NAND2_X1 _14162_ ( .A1(_06196_ ), .A2(_06201_ ), .ZN(_06202_ ) );
AND3_X1 _14163_ ( .A1(_06161_ ), .A2(_06160_ ), .A3(_06162_ ), .ZN(_06203_ ) );
NOR3_X1 _14164_ ( .A1(_06203_ ), .A2(_06163_ ), .A3(_05709_ ), .ZN(_06204_ ) );
OAI21_X1 _14165_ ( .A(_05364_ ), .B1(_06202_ ), .B2(_06204_ ), .ZN(_06205_ ) );
OR3_X1 _14166_ ( .A1(_06130_ ), .A2(_04775_ ), .A3(_04819_ ), .ZN(_06206_ ) );
AND3_X1 _14167_ ( .A1(_06206_ ), .A2(_05515_ ), .A3(_06131_ ), .ZN(_06207_ ) );
AND3_X1 _14168_ ( .A1(_06137_ ), .A2(_06136_ ), .A3(_06139_ ), .ZN(_06208_ ) );
OR3_X1 _14169_ ( .A1(_06208_ ), .A2(_06140_ ), .A3(_04955_ ), .ZN(_06209_ ) );
NAND3_X1 _14170_ ( .A1(_05491_ ), .A2(\ID_EX_imm [10] ), .A3(_05492_ ), .ZN(_06210_ ) );
NAND2_X1 _14171_ ( .A1(_06209_ ), .A2(_06210_ ), .ZN(_06211_ ) );
OAI21_X1 _14172_ ( .A(_04759_ ), .B1(_06207_ ), .B2(_06211_ ), .ZN(_06212_ ) );
AND3_X1 _14173_ ( .A1(_06205_ ), .A2(_05484_ ), .A3(_06212_ ), .ZN(_06213_ ) );
XNOR2_X1 _14174_ ( .A(_05498_ ), .B(_02338_ ), .ZN(_06214_ ) );
OAI21_X1 _14175_ ( .A(_03364_ ), .B1(_06214_ ), .B2(_05725_ ), .ZN(_06215_ ) );
OAI22_X1 _14176_ ( .A1(_06213_ ), .A2(_06215_ ), .B1(_03358_ ), .B2(_03999_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
INV_X1 _14177_ ( .A(_04037_ ), .ZN(_06216_ ) );
XNOR2_X1 _14178_ ( .A(_04749_ ), .B(_02339_ ), .ZN(_06217_ ) );
OR2_X1 _14179_ ( .A1(_05776_ ), .A2(_06129_ ), .ZN(_06218_ ) );
AND2_X1 _14180_ ( .A1(_06218_ ), .A2(_04818_ ), .ZN(_06219_ ) );
OAI21_X1 _14181_ ( .A(_05514_ ), .B1(_06219_ ), .B2(_04817_ ), .ZN(_06220_ ) );
AOI21_X1 _14182_ ( .A(_06220_ ), .B1(_04817_ ), .B2(_06219_ ), .ZN(_06221_ ) );
AND2_X1 _14183_ ( .A1(_05785_ ), .A2(_04877_ ), .ZN(_06222_ ) );
OR3_X1 _14184_ ( .A1(_06222_ ), .A2(_04923_ ), .A3(_04880_ ), .ZN(_06223_ ) );
OAI21_X1 _14185_ ( .A(_04880_ ), .B1(_06222_ ), .B2(_04923_ ), .ZN(_06224_ ) );
AND3_X1 _14186_ ( .A1(_06223_ ), .A2(_04954_ ), .A3(_06224_ ), .ZN(_06225_ ) );
OR2_X1 _14187_ ( .A1(_06221_ ), .A2(_06225_ ), .ZN(_06226_ ) );
AND3_X1 _14188_ ( .A1(_04961_ ), .A2(\ID_EX_imm [9] ), .A3(_04963_ ), .ZN(_06227_ ) );
OAI21_X1 _14189_ ( .A(_04758_ ), .B1(_06226_ ), .B2(_06227_ ), .ZN(_06228_ ) );
NOR3_X1 _14190_ ( .A1(_05609_ ), .A2(_05112_ ), .A3(_05368_ ), .ZN(_06229_ ) );
OAI21_X1 _14191_ ( .A(_06147_ ), .B1(_06180_ ), .B2(_06229_ ), .ZN(_06230_ ) );
NAND3_X1 _14192_ ( .A1(_05689_ ), .A2(_05692_ ), .A3(_05408_ ), .ZN(_06231_ ) );
NAND2_X1 _14193_ ( .A1(_05893_ ), .A2(_05182_ ), .ZN(_06232_ ) );
OAI21_X1 _14194_ ( .A(_05111_ ), .B1(_05183_ ), .B2(_05171_ ), .ZN(_06233_ ) );
OAI21_X1 _14195_ ( .A(_05167_ ), .B1(_05531_ ), .B2(_05185_ ), .ZN(_06234_ ) );
NAND3_X1 _14196_ ( .A1(_06233_ ), .A2(_06234_ ), .A3(_05229_ ), .ZN(_06235_ ) );
NAND2_X1 _14197_ ( .A1(_06232_ ), .A2(_06235_ ), .ZN(_06236_ ) );
OAI211_X1 _14198_ ( .A(_05158_ ), .B(_06231_ ), .C1(_06236_ ), .C2(_05409_ ), .ZN(_06237_ ) );
NAND4_X1 _14199_ ( .A1(_05686_ ), .A2(_05425_ ), .A3(_05232_ ), .A4(_05687_ ), .ZN(_06238_ ) );
AND2_X1 _14200_ ( .A1(_06237_ ), .A2(_06238_ ), .ZN(_06239_ ) );
AOI21_X1 _14201_ ( .A(_04970_ ), .B1(_06230_ ), .B2(_06239_ ), .ZN(_06240_ ) );
AOI21_X1 _14202_ ( .A(_05635_ ), .B1(_06237_ ), .B2(_06238_ ), .ZN(_06241_ ) );
NAND3_X1 _14203_ ( .A1(_05697_ ), .A2(_05194_ ), .A3(_05698_ ), .ZN(_06242_ ) );
NAND4_X1 _14204_ ( .A1(_05550_ ), .A2(_05451_ ), .A3(_05370_ ), .A4(_05444_ ), .ZN(_06243_ ) );
AOI21_X1 _14205_ ( .A(_05868_ ), .B1(_06242_ ), .B2(_06243_ ), .ZN(_06244_ ) );
OR3_X1 _14206_ ( .A1(_06240_ ), .A2(_06241_ ), .A3(_06244_ ), .ZN(_06245_ ) );
OAI21_X1 _14207_ ( .A(_05276_ ), .B1(_05298_ ), .B2(_05306_ ), .ZN(_06246_ ) );
INV_X1 _14208_ ( .A(_05259_ ), .ZN(_06247_ ) );
INV_X1 _14209_ ( .A(_05258_ ), .ZN(_06248_ ) );
AND3_X1 _14210_ ( .A1(_06246_ ), .A2(_06247_ ), .A3(_06248_ ), .ZN(_06249_ ) );
AOI21_X1 _14211_ ( .A(_06248_ ), .B1(_06246_ ), .B2(_06247_ ), .ZN(_06250_ ) );
NOR3_X1 _14212_ ( .A1(_06249_ ), .A2(_06250_ ), .A3(_05240_ ), .ZN(_06251_ ) );
AND2_X1 _14213_ ( .A1(_05258_ ), .A2(_05335_ ), .ZN(_06252_ ) );
NOR3_X1 _14214_ ( .A1(_05008_ ), .A2(_04777_ ), .A3(_05340_ ), .ZN(_06253_ ) );
AOI21_X1 _14215_ ( .A(_05344_ ), .B1(_05008_ ), .B2(_04777_ ), .ZN(_06254_ ) );
OR3_X1 _14216_ ( .A1(_06252_ ), .A2(_06253_ ), .A3(_06254_ ), .ZN(_06255_ ) );
NOR3_X1 _14217_ ( .A1(_06245_ ), .A2(_06251_ ), .A3(_06255_ ), .ZN(_06256_ ) );
OAI21_X1 _14218_ ( .A(_06228_ ), .B1(_06256_ ), .B2(_05357_ ), .ZN(_06257_ ) );
MUX2_X1 _14219_ ( .A(_06217_ ), .B(_06257_ ), .S(_05360_ ), .Z(_06258_ ) );
MUX2_X1 _14220_ ( .A(_06216_ ), .B(_06258_ ), .S(_03390_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
INV_X1 _14221_ ( .A(_04082_ ), .ZN(_06259_ ) );
NOR2_X1 _14222_ ( .A1(_04982_ ), .A2(_05465_ ), .ZN(_06260_ ) );
INV_X1 _14223_ ( .A(_06260_ ), .ZN(_06261_ ) );
NAND4_X1 _14224_ ( .A1(_05108_ ), .A2(_05119_ ), .A3(_06261_ ), .A4(_05120_ ), .ZN(_06262_ ) );
NAND3_X1 _14225_ ( .A1(_05935_ ), .A2(_05182_ ), .A3(_05936_ ), .ZN(_06263_ ) );
OAI21_X1 _14226_ ( .A(_05177_ ), .B1(_05432_ ), .B2(_05416_ ), .ZN(_06264_ ) );
OAI21_X1 _14227_ ( .A(_05197_ ), .B1(_05429_ ), .B2(_05433_ ), .ZN(_06265_ ) );
NAND2_X1 _14228_ ( .A1(_06264_ ), .A2(_06265_ ), .ZN(_06266_ ) );
NAND2_X1 _14229_ ( .A1(_06266_ ), .A2(_05180_ ), .ZN(_06267_ ) );
AND3_X1 _14230_ ( .A1(_06263_ ), .A2(_05818_ ), .A3(_06267_ ), .ZN(_06268_ ) );
AOI211_X1 _14231_ ( .A(_05380_ ), .B(_06268_ ), .C1(_05738_ ), .C2(_05452_ ), .ZN(_06269_ ) );
AOI21_X1 _14232_ ( .A(_05553_ ), .B1(_05732_ ), .B2(_05804_ ), .ZN(_06270_ ) );
OR2_X1 _14233_ ( .A1(_06269_ ), .A2(_06270_ ), .ZN(_06271_ ) );
AOI21_X1 _14234_ ( .A(_05799_ ), .B1(_06262_ ), .B2(_06271_ ), .ZN(_06272_ ) );
OR3_X1 _14235_ ( .A1(_05298_ ), .A2(_05306_ ), .A3(_05276_ ), .ZN(_06273_ ) );
NAND3_X1 _14236_ ( .A1(_06273_ ), .A2(_05479_ ), .A3(_06246_ ), .ZN(_06274_ ) );
OR3_X1 _14237_ ( .A1(_06269_ ), .A2(_06270_ ), .A3(_05813_ ), .ZN(_06275_ ) );
INV_X1 _14238_ ( .A(_05011_ ), .ZN(_06276_ ) );
NAND3_X1 _14239_ ( .A1(_06276_ ), .A2(_01832_ ), .A3(_05476_ ), .ZN(_06277_ ) );
AOI21_X1 _14240_ ( .A(_05344_ ), .B1(_05011_ ), .B2(_04779_ ), .ZN(_06278_ ) );
NAND3_X1 _14241_ ( .A1(_05743_ ), .A2(_05745_ ), .A3(_05804_ ), .ZN(_06279_ ) );
NAND4_X1 _14242_ ( .A1(_04977_ ), .A2(_03359_ ), .A3(_05465_ ), .A4(_05700_ ), .ZN(_06280_ ) );
AOI21_X1 _14243_ ( .A(_05868_ ), .B1(_06279_ ), .B2(_06280_ ), .ZN(_06281_ ) );
AOI211_X1 _14244_ ( .A(_06278_ ), .B(_06281_ ), .C1(_05276_ ), .C2(_05472_ ), .ZN(_06282_ ) );
NAND4_X1 _14245_ ( .A1(_06274_ ), .A2(_06275_ ), .A3(_06277_ ), .A4(_06282_ ), .ZN(_06283_ ) );
OAI21_X1 _14246_ ( .A(_05365_ ), .B1(_06272_ ), .B2(_06283_ ), .ZN(_06284_ ) );
NAND3_X1 _14247_ ( .A1(_04804_ ), .A2(_04813_ ), .A3(_06129_ ), .ZN(_06285_ ) );
AND3_X1 _14248_ ( .A1(_06218_ ), .A2(_05515_ ), .A3(_06285_ ), .ZN(_06286_ ) );
AOI21_X1 _14249_ ( .A(_05487_ ), .B1(_05785_ ), .B2(_04877_ ), .ZN(_06287_ ) );
OAI21_X1 _14250_ ( .A(_06287_ ), .B1(_05785_ ), .B2(_04877_ ), .ZN(_06288_ ) );
NAND3_X1 _14251_ ( .A1(_05524_ ), .A2(\ID_EX_imm [8] ), .A3(_05525_ ), .ZN(_06289_ ) );
NAND2_X1 _14252_ ( .A1(_06288_ ), .A2(_06289_ ), .ZN(_06290_ ) );
OAI21_X1 _14253_ ( .A(_04759_ ), .B1(_06286_ ), .B2(_06290_ ), .ZN(_06291_ ) );
AND3_X1 _14254_ ( .A1(_06284_ ), .A2(_05484_ ), .A3(_06291_ ), .ZN(_06292_ ) );
XNOR2_X1 _14255_ ( .A(_04748_ ), .B(_02340_ ), .ZN(_06293_ ) );
OAI21_X1 _14256_ ( .A(_03364_ ), .B1(_06293_ ), .B2(_05725_ ), .ZN(_06294_ ) );
OAI21_X1 _14257_ ( .A(_06259_ ), .B1(_06292_ ), .B2(_06294_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
NAND2_X1 _14258_ ( .A1(_04114_ ), .A2(_03379_ ), .ZN(_06295_ ) );
XNOR2_X1 _14259_ ( .A(_04747_ ), .B(\ID_EX_pc [7] ), .ZN(_06296_ ) );
NOR2_X1 _14260_ ( .A1(_06296_ ), .A2(_05484_ ), .ZN(_06297_ ) );
OAI21_X1 _14261_ ( .A(_04803_ ), .B1(_04793_ ), .B2(_04794_ ), .ZN(_06298_ ) );
AND2_X1 _14262_ ( .A1(_06298_ ), .A2(_04807_ ), .ZN(_06299_ ) );
OR2_X1 _14263_ ( .A1(_06299_ ), .A2(_04809_ ), .ZN(_06300_ ) );
AND3_X1 _14264_ ( .A1(_06300_ ), .A2(_04811_ ), .A3(_04808_ ), .ZN(_06301_ ) );
AOI21_X1 _14265_ ( .A(_04808_ ), .B1(_06300_ ), .B2(_04811_ ), .ZN(_06302_ ) );
NOR3_X1 _14266_ ( .A1(_06301_ ), .A2(_06302_ ), .A3(_04867_ ), .ZN(_06303_ ) );
NOR2_X1 _14267_ ( .A1(_04912_ ), .A2(_04910_ ), .ZN(_06304_ ) );
OR3_X1 _14268_ ( .A1(_04907_ ), .A2(_04908_ ), .A3(_06304_ ), .ZN(_06305_ ) );
OAI21_X1 _14269_ ( .A(_06304_ ), .B1(_04907_ ), .B2(_04908_ ), .ZN(_06306_ ) );
NAND3_X1 _14270_ ( .A1(_06305_ ), .A2(_05672_ ), .A3(_06306_ ), .ZN(_06307_ ) );
NAND3_X1 _14271_ ( .A1(_05491_ ), .A2(\ID_EX_imm [7] ), .A3(_05492_ ), .ZN(_06308_ ) );
NAND2_X1 _14272_ ( .A1(_06307_ ), .A2(_06308_ ), .ZN(_06309_ ) );
OAI21_X1 _14273_ ( .A(_04759_ ), .B1(_06303_ ), .B2(_06309_ ), .ZN(_06310_ ) );
NAND3_X1 _14274_ ( .A1(_05122_ ), .A2(_05119_ ), .A3(_05368_ ), .ZN(_06311_ ) );
AND3_X1 _14275_ ( .A1(_04977_ ), .A2(_02268_ ), .A3(_05180_ ), .ZN(_06312_ ) );
MUX2_X1 _14276_ ( .A(_06312_ ), .B(_05808_ ), .S(_05425_ ), .Z(_06313_ ) );
NAND2_X1 _14277_ ( .A1(_06313_ ), .A2(_05380_ ), .ZN(_06314_ ) );
OR3_X1 _14278_ ( .A1(_05166_ ), .A2(_05176_ ), .A3(_05197_ ), .ZN(_06315_ ) );
OR3_X1 _14279_ ( .A1(_05183_ ), .A2(_05171_ ), .A3(_05184_ ), .ZN(_06316_ ) );
NAND2_X1 _14280_ ( .A1(_06315_ ), .A2(_06316_ ), .ZN(_06317_ ) );
NAND2_X1 _14281_ ( .A1(_06317_ ), .A2(_05744_ ), .ZN(_06318_ ) );
NAND3_X1 _14282_ ( .A1(_06151_ ), .A2(_06152_ ), .A3(_05428_ ), .ZN(_06319_ ) );
AOI21_X1 _14283_ ( .A(_05465_ ), .B1(_06318_ ), .B2(_06319_ ), .ZN(_06320_ ) );
OAI21_X1 _14284_ ( .A(_05428_ ), .B1(_05567_ ), .B2(_05568_ ), .ZN(_06321_ ) );
AOI21_X1 _14285_ ( .A(_05818_ ), .B1(_06321_ ), .B2(_05803_ ), .ZN(_06322_ ) );
OAI21_X1 _14286_ ( .A(_05553_ ), .B1(_06320_ ), .B2(_06322_ ), .ZN(_06323_ ) );
AND2_X1 _14287_ ( .A1(_06314_ ), .A2(_06323_ ), .ZN(_06324_ ) );
AOI21_X1 _14288_ ( .A(_05799_ ), .B1(_06311_ ), .B2(_06324_ ), .ZN(_06325_ ) );
INV_X1 _14289_ ( .A(_05292_ ), .ZN(_06326_ ) );
NAND4_X1 _14290_ ( .A1(_05289_ ), .A2(_05291_ ), .A3(_05296_ ), .A4(_05294_ ), .ZN(_06327_ ) );
NAND2_X1 _14291_ ( .A1(_06327_ ), .A2(_05305_ ), .ZN(_06328_ ) );
NAND2_X1 _14292_ ( .A1(_06328_ ), .A2(_05295_ ), .ZN(_06329_ ) );
INV_X1 _14293_ ( .A(_05299_ ), .ZN(_06330_ ) );
AOI21_X1 _14294_ ( .A(_06326_ ), .B1(_06329_ ), .B2(_06330_ ), .ZN(_06331_ ) );
AOI211_X1 _14295_ ( .A(_05299_ ), .B(_05292_ ), .C1(_06328_ ), .C2(_05295_ ), .ZN(_06332_ ) );
NOR3_X1 _14296_ ( .A1(_06331_ ), .A2(_06332_ ), .A3(_05709_ ), .ZN(_06333_ ) );
AOI21_X1 _14297_ ( .A(_05813_ ), .B1(_06314_ ), .B2(_06323_ ), .ZN(_06334_ ) );
AOI21_X1 _14298_ ( .A(_05470_ ), .B1(_04999_ ), .B2(_04116_ ), .ZN(_06335_ ) );
OAI211_X1 _14299_ ( .A(_05549_ ), .B(_05428_ ), .C1(_05550_ ), .C2(_05444_ ), .ZN(_06336_ ) );
AOI21_X1 _14300_ ( .A(_05451_ ), .B1(_05815_ ), .B2(_06336_ ), .ZN(_06337_ ) );
NAND2_X1 _14301_ ( .A1(_06337_ ), .A2(_05822_ ), .ZN(_06338_ ) );
OR3_X1 _14302_ ( .A1(_04116_ ), .A2(_04999_ ), .A3(_05339_ ), .ZN(_06339_ ) );
OAI211_X1 _14303_ ( .A(_06338_ ), .B(_06339_ ), .C1(_06326_ ), .C2(_05662_ ), .ZN(_06340_ ) );
OR3_X1 _14304_ ( .A1(_06334_ ), .A2(_06335_ ), .A3(_06340_ ), .ZN(_06341_ ) );
NOR3_X1 _14305_ ( .A1(_06325_ ), .A2(_06333_ ), .A3(_06341_ ), .ZN(_06342_ ) );
OAI21_X1 _14306_ ( .A(_06310_ ), .B1(_06342_ ), .B2(_05528_ ), .ZN(_06343_ ) );
AOI21_X1 _14307_ ( .A(_06297_ ), .B1(_06343_ ), .B2(_05725_ ), .ZN(_06344_ ) );
OAI21_X1 _14308_ ( .A(_06295_ ), .B1(_06344_ ), .B2(_03762_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
OAI211_X1 _14309_ ( .A(_03698_ ), .B(_04174_ ), .C1(_04175_ ), .C2(_04180_ ), .ZN(_06345_ ) );
NOR3_X1 _14310_ ( .A1(_05109_ ), .A2(_05116_ ), .A3(_05879_ ), .ZN(_06346_ ) );
NAND2_X1 _14311_ ( .A1(_06346_ ), .A2(_06147_ ), .ZN(_06347_ ) );
NAND4_X1 _14312_ ( .A1(_05406_ ), .A2(_04985_ ), .A3(_05229_ ), .A4(_05213_ ), .ZN(_06348_ ) );
OAI211_X1 _14313_ ( .A(_05381_ ), .B(_06348_ ), .C1(_05862_ ), .C2(_05466_ ), .ZN(_06349_ ) );
AOI21_X1 _14314_ ( .A(_05700_ ), .B1(_06183_ ), .B2(_06184_ ), .ZN(_06350_ ) );
OAI21_X1 _14315_ ( .A(_05444_ ), .B1(_05414_ ), .B2(_05419_ ), .ZN(_06351_ ) );
OAI21_X1 _14316_ ( .A(_05372_ ), .B1(_05432_ ), .B2(_05416_ ), .ZN(_06352_ ) );
AND3_X1 _14317_ ( .A1(_06351_ ), .A2(_06352_ ), .A3(_05744_ ), .ZN(_06353_ ) );
OAI21_X1 _14318_ ( .A(_05427_ ), .B1(_06350_ ), .B2(_06353_ ), .ZN(_06354_ ) );
OAI21_X1 _14319_ ( .A(_05466_ ), .B1(_05855_ ), .B2(_05858_ ), .ZN(_06355_ ) );
NAND3_X1 _14320_ ( .A1(_06354_ ), .A2(_05467_ ), .A3(_06355_ ), .ZN(_06356_ ) );
NAND2_X1 _14321_ ( .A1(_06349_ ), .A2(_06356_ ), .ZN(_06357_ ) );
AOI21_X1 _14322_ ( .A(_05799_ ), .B1(_06347_ ), .B2(_06357_ ), .ZN(_06358_ ) );
AOI21_X1 _14323_ ( .A(_05709_ ), .B1(_06328_ ), .B2(_05295_ ), .ZN(_06359_ ) );
OAI21_X1 _14324_ ( .A(_06359_ ), .B1(_05295_ ), .B2(_06328_ ), .ZN(_06360_ ) );
AND3_X1 _14325_ ( .A1(_05870_ ), .A2(_05425_ ), .A3(_05871_ ), .ZN(_06361_ ) );
AND2_X1 _14326_ ( .A1(_06361_ ), .A2(_05822_ ), .ZN(_06362_ ) );
NAND3_X1 _14327_ ( .A1(_05000_ ), .A2(_04799_ ), .A3(_05001_ ), .ZN(_06363_ ) );
AOI221_X4 _14328_ ( .A(_06362_ ), .B1(_06363_ ), .B2(_05342_ ), .C1(_05295_ ), .C2(_05335_ ), .ZN(_06364_ ) );
NAND3_X1 _14329_ ( .A1(_06349_ ), .A2(_05474_ ), .A3(_06356_ ), .ZN(_06365_ ) );
OR3_X1 _14330_ ( .A1(_05002_ ), .A2(_04799_ ), .A3(_05340_ ), .ZN(_06366_ ) );
NAND4_X1 _14331_ ( .A1(_06360_ ), .A2(_06364_ ), .A3(_06365_ ), .A4(_06366_ ), .ZN(_06367_ ) );
OAI21_X1 _14332_ ( .A(_05365_ ), .B1(_06358_ ), .B2(_06367_ ), .ZN(_06368_ ) );
NAND3_X1 _14333_ ( .A1(_06298_ ), .A2(_04809_ ), .A3(_04807_ ), .ZN(_06369_ ) );
AND3_X1 _14334_ ( .A1(_06300_ ), .A2(_05515_ ), .A3(_06369_ ), .ZN(_06370_ ) );
AOI21_X1 _14335_ ( .A(_05487_ ), .B1(_04905_ ), .B2(_04906_ ), .ZN(_06371_ ) );
OAI21_X1 _14336_ ( .A(_06371_ ), .B1(_04906_ ), .B2(_04905_ ), .ZN(_06372_ ) );
NAND3_X1 _14337_ ( .A1(_05491_ ), .A2(\ID_EX_imm [6] ), .A3(_05492_ ), .ZN(_06373_ ) );
NAND2_X1 _14338_ ( .A1(_06372_ ), .A2(_06373_ ), .ZN(_06374_ ) );
OAI21_X1 _14339_ ( .A(_04759_ ), .B1(_06370_ ), .B2(_06374_ ), .ZN(_06375_ ) );
AND3_X1 _14340_ ( .A1(_06368_ ), .A2(_05484_ ), .A3(_06375_ ), .ZN(_06376_ ) );
AOI21_X1 _14341_ ( .A(\ID_EX_pc [6] ), .B1(_04745_ ), .B2(\ID_EX_pc [5] ), .ZN(_06377_ ) );
OAI21_X1 _14342_ ( .A(_05497_ ), .B1(_04747_ ), .B2(_06377_ ), .ZN(_06378_ ) );
NAND2_X1 _14343_ ( .A1(_06378_ ), .A2(_03407_ ), .ZN(_06379_ ) );
OAI21_X1 _14344_ ( .A(_06345_ ), .B1(_06376_ ), .B2(_06379_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
XNOR2_X1 _14345_ ( .A(_04745_ ), .B(_02342_ ), .ZN(_06380_ ) );
AND2_X1 _14346_ ( .A1(_04795_ ), .A2(_04801_ ), .ZN(_06381_ ) );
OR3_X1 _14347_ ( .A1(_06381_ ), .A2(_04805_ ), .A3(_04802_ ), .ZN(_06382_ ) );
OAI21_X1 _14348_ ( .A(_04802_ ), .B1(_06381_ ), .B2(_04805_ ), .ZN(_06383_ ) );
AND3_X1 _14349_ ( .A1(_06382_ ), .A2(_05514_ ), .A3(_06383_ ), .ZN(_06384_ ) );
NOR2_X1 _14350_ ( .A1(_04901_ ), .A2(_04904_ ), .ZN(_06385_ ) );
OR3_X1 _14351_ ( .A1(_04900_ ), .A2(_04902_ ), .A3(_06385_ ), .ZN(_06386_ ) );
OAI21_X1 _14352_ ( .A(_06385_ ), .B1(_04900_ ), .B2(_04902_ ), .ZN(_06387_ ) );
NAND3_X1 _14353_ ( .A1(_06386_ ), .A2(_04954_ ), .A3(_06387_ ), .ZN(_06388_ ) );
NAND3_X1 _14354_ ( .A1(_04962_ ), .A2(\ID_EX_imm [5] ), .A3(_04964_ ), .ZN(_06389_ ) );
NAND2_X1 _14355_ ( .A1(_06388_ ), .A2(_06389_ ), .ZN(_06390_ ) );
OAI21_X1 _14356_ ( .A(_04758_ ), .B1(_06384_ ), .B2(_06390_ ), .ZN(_06391_ ) );
AND2_X1 _14357_ ( .A1(_05294_ ), .A2(_05334_ ), .ZN(_06392_ ) );
INV_X1 _14358_ ( .A(_06147_ ), .ZN(_06393_ ) );
NOR4_X4 _14359_ ( .A1(_05109_ ), .A2(_05114_ ), .A3(_05116_ ), .A4(_06393_ ), .ZN(_06394_ ) );
NAND2_X1 _14360_ ( .A1(_05157_ ), .A2(_05231_ ), .ZN(_06395_ ) );
NAND3_X1 _14361_ ( .A1(_06233_ ), .A2(_06234_ ), .A3(_05125_ ), .ZN(_06396_ ) );
NOR3_X1 _14362_ ( .A1(_05166_ ), .A2(_05176_ ), .A3(_05111_ ), .ZN(_06397_ ) );
NOR3_X1 _14363_ ( .A1(_05175_ ), .A2(_05167_ ), .A3(_05217_ ), .ZN(_06398_ ) );
NOR2_X1 _14364_ ( .A1(_06397_ ), .A2(_06398_ ), .ZN(_06399_ ) );
OAI211_X1 _14365_ ( .A(_06396_ ), .B(_04986_ ), .C1(_06399_ ), .C2(_05202_ ), .ZN(_06400_ ) );
OAI211_X1 _14366_ ( .A(_05158_ ), .B(_06400_ ), .C1(_05894_ ), .C2(_05193_ ), .ZN(_06401_ ) );
NAND2_X1 _14367_ ( .A1(_06395_ ), .A2(_06401_ ), .ZN(_06402_ ) );
OAI21_X2 _14368_ ( .A(_04969_ ), .B1(_06394_ ), .B2(_06402_ ), .ZN(_06403_ ) );
NAND2_X1 _14369_ ( .A1(_06402_ ), .A2(_05235_ ), .ZN(_06404_ ) );
NAND4_X1 _14370_ ( .A1(_05224_ ), .A2(_05230_ ), .A3(_05425_ ), .A4(_05158_ ), .ZN(_06405_ ) );
OAI211_X1 _14371_ ( .A(_06403_ ), .B(_06404_ ), .C1(_05164_ ), .C2(_06405_ ), .ZN(_06406_ ) );
AND3_X1 _14372_ ( .A1(_04994_ ), .A2(_01657_ ), .A3(_05475_ ), .ZN(_06407_ ) );
AOI21_X1 _14373_ ( .A(_05343_ ), .B1(_04995_ ), .B2(_05293_ ), .ZN(_06408_ ) );
OR4_X2 _14374_ ( .A1(_06392_ ), .A2(_06406_ ), .A3(_06407_ ), .A4(_06408_ ), .ZN(_06409_ ) );
NAND2_X1 _14375_ ( .A1(_05289_ ), .A2(_05291_ ), .ZN(_06410_ ) );
INV_X1 _14376_ ( .A(_05296_ ), .ZN(_06411_ ) );
NOR2_X1 _14377_ ( .A1(_06410_ ), .A2(_06411_ ), .ZN(_06412_ ) );
OR3_X1 _14378_ ( .A1(_06412_ ), .A2(_05304_ ), .A3(_05294_ ), .ZN(_06413_ ) );
OAI21_X1 _14379_ ( .A(_05294_ ), .B1(_06412_ ), .B2(_05304_ ), .ZN(_06414_ ) );
AND2_X1 _14380_ ( .A1(_06414_ ), .A2(_05239_ ), .ZN(_06415_ ) );
AOI21_X1 _14381_ ( .A(_06409_ ), .B1(_06413_ ), .B2(_06415_ ), .ZN(_06416_ ) );
OAI21_X1 _14382_ ( .A(_06391_ ), .B1(_06416_ ), .B2(_05357_ ), .ZN(_06417_ ) );
MUX2_X1 _14383_ ( .A(_06380_ ), .B(_06417_ ), .S(_05360_ ), .Z(_06418_ ) );
MUX2_X1 _14384_ ( .A(_04205_ ), .B(_06418_ ), .S(_03390_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
XNOR2_X1 _14385_ ( .A(_04744_ ), .B(_02343_ ), .ZN(_06419_ ) );
NOR3_X1 _14386_ ( .A1(_04793_ ), .A2(_04794_ ), .A3(_04801_ ), .ZN(_06420_ ) );
NOR3_X1 _14387_ ( .A1(_06381_ ), .A2(_06420_ ), .A3(_04866_ ), .ZN(_06421_ ) );
AND3_X1 _14388_ ( .A1(_04897_ ), .A2(_04899_ ), .A3(_04886_ ), .ZN(_06422_ ) );
NOR3_X1 _14389_ ( .A1(_06422_ ), .A2(_04900_ ), .A3(_04955_ ), .ZN(_06423_ ) );
OR2_X1 _14390_ ( .A1(_06421_ ), .A2(_06423_ ), .ZN(_06424_ ) );
AND3_X1 _14391_ ( .A1(_04961_ ), .A2(\ID_EX_imm [4] ), .A3(_04963_ ), .ZN(_06425_ ) );
OAI21_X1 _14392_ ( .A(_04758_ ), .B1(_06424_ ), .B2(_06425_ ), .ZN(_06426_ ) );
NAND4_X1 _14393_ ( .A1(_05108_ ), .A2(_05368_ ), .A3(_05373_ ), .A4(_06147_ ), .ZN(_06427_ ) );
AOI21_X1 _14394_ ( .A(_05425_ ), .B1(_05937_ ), .B2(_05938_ ), .ZN(_06428_ ) );
OAI21_X1 _14395_ ( .A(_05420_ ), .B1(_05418_ ), .B2(_05461_ ), .ZN(_06429_ ) );
OAI21_X1 _14396_ ( .A(_05219_ ), .B1(_05414_ ), .B2(_05419_ ), .ZN(_06430_ ) );
NAND2_X1 _14397_ ( .A1(_06429_ ), .A2(_06430_ ), .ZN(_06431_ ) );
MUX2_X1 _14398_ ( .A(_06266_ ), .B(_06431_ ), .S(_05369_ ), .Z(_06432_ ) );
AOI211_X1 _14399_ ( .A(_05232_ ), .B(_06428_ ), .C1(_05818_ ), .C2(_06432_ ), .ZN(_06433_ ) );
AOI21_X1 _14400_ ( .A(_05165_ ), .B1(_05401_ ), .B2(_05410_ ), .ZN(_06434_ ) );
NOR2_X1 _14401_ ( .A1(_06433_ ), .A2(_06434_ ), .ZN(_06435_ ) );
AOI21_X1 _14402_ ( .A(_05799_ ), .B1(_06427_ ), .B2(_06435_ ), .ZN(_06436_ ) );
NAND3_X1 _14403_ ( .A1(_05380_ ), .A2(_03394_ ), .A3(_05475_ ), .ZN(_06437_ ) );
XNOR2_X1 _14404_ ( .A(_06410_ ), .B(_06411_ ), .ZN(_06438_ ) );
OAI221_X1 _14405_ ( .A(_06437_ ), .B1(_05240_ ), .B2(_06438_ ), .C1(_06435_ ), .C2(_05813_ ), .ZN(_06439_ ) );
OR3_X1 _14406_ ( .A1(_05464_ ), .A2(_05451_ ), .A3(_05868_ ), .ZN(_06440_ ) );
OAI21_X1 _14407_ ( .A(_05580_ ), .B1(_05380_ ), .B2(_03394_ ), .ZN(_06441_ ) );
OAI211_X1 _14408_ ( .A(_06440_ ), .B(_06441_ ), .C1(_06411_ ), .C2(_05662_ ), .ZN(_06442_ ) );
NOR3_X1 _14409_ ( .A1(_06436_ ), .A2(_06439_ ), .A3(_06442_ ), .ZN(_06443_ ) );
OAI21_X1 _14410_ ( .A(_06426_ ), .B1(_06443_ ), .B2(_05357_ ), .ZN(_06444_ ) );
MUX2_X1 _14411_ ( .A(_06419_ ), .B(_06444_ ), .S(_05359_ ), .Z(_06445_ ) );
MUX2_X1 _14412_ ( .A(_04246_ ), .B(_06445_ ), .S(_03390_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
XOR2_X1 _14413_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .Z(_06446_ ) );
AND2_X1 _14414_ ( .A1(_04790_ ), .A2(_04792_ ), .ZN(_06447_ ) );
XNOR2_X1 _14415_ ( .A(_04309_ ), .B(_01521_ ), .ZN(_06448_ ) );
XNOR2_X1 _14416_ ( .A(_06447_ ), .B(_06448_ ), .ZN(_06449_ ) );
AND2_X1 _14417_ ( .A1(_06449_ ), .A2(_05514_ ), .ZN(_06450_ ) );
OR2_X1 _14418_ ( .A1(_04890_ ), .A2(_04892_ ), .ZN(_06451_ ) );
INV_X1 _14419_ ( .A(_04898_ ), .ZN(_06452_ ) );
AND3_X1 _14420_ ( .A1(_06451_ ), .A2(_06452_ ), .A3(_04896_ ), .ZN(_06453_ ) );
AOI21_X1 _14421_ ( .A(_04896_ ), .B1(_06451_ ), .B2(_06452_ ), .ZN(_06454_ ) );
OR3_X1 _14422_ ( .A1(_06453_ ), .A2(_06454_ ), .A3(_04955_ ), .ZN(_06455_ ) );
NAND3_X1 _14423_ ( .A1(_04962_ ), .A2(\ID_EX_imm [3] ), .A3(_04964_ ), .ZN(_06456_ ) );
NAND2_X1 _14424_ ( .A1(_06455_ ), .A2(_06456_ ), .ZN(_06457_ ) );
OAI21_X1 _14425_ ( .A(_04758_ ), .B1(_06450_ ), .B2(_06457_ ), .ZN(_06458_ ) );
AND4_X1 _14426_ ( .A1(_05119_ ), .A2(_05122_ ), .A3(_05368_ ), .A4(_05574_ ), .ZN(_06459_ ) );
NAND2_X1 _14427_ ( .A1(_05572_ ), .A2(_05232_ ), .ZN(_06460_ ) );
NAND3_X1 _14428_ ( .A1(_06150_ ), .A2(_05409_ ), .A3(_06153_ ), .ZN(_06461_ ) );
NOR2_X1 _14429_ ( .A1(_05216_ ), .A2(_05221_ ), .ZN(_06462_ ) );
NOR2_X1 _14430_ ( .A1(_05175_ ), .A2(_05217_ ), .ZN(_06463_ ) );
MUX2_X1 _14431_ ( .A(_06462_ ), .B(_06463_ ), .S(_05168_ ), .Z(_06464_ ) );
MUX2_X1 _14432_ ( .A(_06317_ ), .B(_06464_ ), .S(_05369_ ), .Z(_06465_ ) );
OAI211_X1 _14433_ ( .A(_05165_ ), .B(_06461_ ), .C1(_06465_ ), .C2(_05451_ ), .ZN(_06466_ ) );
NAND2_X1 _14434_ ( .A1(_06460_ ), .A2(_06466_ ), .ZN(_06467_ ) );
OAI21_X1 _14435_ ( .A(_04969_ ), .B1(_06459_ ), .B2(_06467_ ), .ZN(_06468_ ) );
XNOR2_X1 _14436_ ( .A(_04985_ ), .B(_01601_ ), .ZN(_06469_ ) );
NOR2_X1 _14437_ ( .A1(_05286_ ), .A2(_05288_ ), .ZN(_06470_ ) );
OAI21_X1 _14438_ ( .A(_06469_ ), .B1(_06470_ ), .B2(_05279_ ), .ZN(_06471_ ) );
INV_X1 _14439_ ( .A(_06469_ ), .ZN(_06472_ ) );
OAI211_X1 _14440_ ( .A(_05280_ ), .B(_06472_ ), .C1(_05286_ ), .C2(_05288_ ), .ZN(_06473_ ) );
NAND3_X1 _14441_ ( .A1(_06471_ ), .A2(_05239_ ), .A3(_06473_ ), .ZN(_06474_ ) );
AND3_X1 _14442_ ( .A1(_05451_ ), .A2(_01521_ ), .A3(_05475_ ), .ZN(_06475_ ) );
NOR4_X1 _14443_ ( .A1(_05551_ ), .A2(_05408_ ), .A3(_05399_ ), .A4(_05232_ ), .ZN(_06476_ ) );
NAND2_X1 _14444_ ( .A1(_06476_ ), .A2(_05413_ ), .ZN(_06477_ ) );
OAI221_X1 _14445_ ( .A(_06477_ ), .B1(_05290_ ), .B2(_05344_ ), .C1(_06472_ ), .C2(_05662_ ), .ZN(_06478_ ) );
AOI211_X1 _14446_ ( .A(_06475_ ), .B(_06478_ ), .C1(_06467_ ), .C2(_05235_ ), .ZN(_06479_ ) );
AND3_X1 _14447_ ( .A1(_06468_ ), .A2(_06474_ ), .A3(_06479_ ), .ZN(_06480_ ) );
OAI21_X1 _14448_ ( .A(_06458_ ), .B1(_06480_ ), .B2(_05357_ ), .ZN(_06481_ ) );
MUX2_X1 _14449_ ( .A(_06446_ ), .B(_06481_ ), .S(_05359_ ), .Z(_06482_ ) );
MUX2_X1 _14450_ ( .A(_04280_ ), .B(_06482_ ), .S(_05362_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
OR2_X1 _14451_ ( .A1(_04343_ ), .A2(_05362_ ), .ZN(_06483_ ) );
NAND3_X1 _14452_ ( .A1(_04784_ ), .A2(_04785_ ), .A3(_04789_ ), .ZN(_06484_ ) );
NAND3_X1 _14453_ ( .A1(_04790_ ), .A2(_05514_ ), .A3(_06484_ ), .ZN(_06485_ ) );
NAND2_X1 _14454_ ( .A1(_04890_ ), .A2(_04892_ ), .ZN(_06486_ ) );
NAND3_X1 _14455_ ( .A1(_06451_ ), .A2(_05672_ ), .A3(_06486_ ), .ZN(_06487_ ) );
NAND3_X1 _14456_ ( .A1(_05491_ ), .A2(\ID_EX_imm [2] ), .A3(_05492_ ), .ZN(_06488_ ) );
AND3_X1 _14457_ ( .A1(_06485_ ), .A2(_06487_ ), .A3(_06488_ ), .ZN(_06489_ ) );
AOI21_X1 _14458_ ( .A(_05669_ ), .B1(_06489_ ), .B2(_01355_ ), .ZN(_06490_ ) );
NAND2_X1 _14459_ ( .A1(_05628_ ), .A2(_05381_ ), .ZN(_06491_ ) );
OR3_X1 _14460_ ( .A1(_06185_ ), .A2(_06186_ ), .A3(_05194_ ), .ZN(_06492_ ) );
OAI21_X1 _14461_ ( .A(_05372_ ), .B1(_05418_ ), .B2(_05461_ ), .ZN(_06493_ ) );
NOR2_X1 _14462_ ( .A1(_05457_ ), .A2(_05460_ ), .ZN(_06494_ ) );
OAI211_X1 _14463_ ( .A(_05744_ ), .B(_06493_ ), .C1(_06494_ ), .C2(_05372_ ), .ZN(_06495_ ) );
NAND3_X1 _14464_ ( .A1(_06351_ ), .A2(_06352_ ), .A3(_05552_ ), .ZN(_06496_ ) );
NAND3_X1 _14465_ ( .A1(_06495_ ), .A2(_05426_ ), .A3(_06496_ ), .ZN(_06497_ ) );
NAND3_X1 _14466_ ( .A1(_06492_ ), .A2(_05747_ ), .A3(_06497_ ), .ZN(_06498_ ) );
AOI21_X1 _14467_ ( .A(_05813_ ), .B1(_06491_ ), .B2(_06498_ ), .ZN(_06499_ ) );
NOR2_X1 _14468_ ( .A1(_05609_ ), .A2(_05610_ ), .ZN(_06500_ ) );
NAND3_X1 _14469_ ( .A1(_06500_ ), .A2(_05368_ ), .A3(_06147_ ), .ZN(_06501_ ) );
AND2_X1 _14470_ ( .A1(_06491_ ), .A2(_06498_ ), .ZN(_06502_ ) );
AOI21_X1 _14471_ ( .A(_05799_ ), .B1(_06501_ ), .B2(_06502_ ), .ZN(_06503_ ) );
AOI211_X1 _14472_ ( .A(_06499_ ), .B(_06503_ ), .C1(_05640_ ), .C2(_05822_ ), .ZN(_06504_ ) );
AOI21_X1 _14473_ ( .A(_05709_ ), .B1(_05286_ ), .B2(_05288_ ), .ZN(_06505_ ) );
OAI21_X1 _14474_ ( .A(_06505_ ), .B1(_05286_ ), .B2(_05288_ ), .ZN(_06506_ ) );
AOI21_X1 _14475_ ( .A(_05470_ ), .B1(_05700_ ), .B2(_04787_ ), .ZN(_06507_ ) );
AOI221_X4 _14476_ ( .A(_06507_ ), .B1(_05279_ ), .B2(_05476_ ), .C1(_05287_ ), .C2(_05472_ ), .ZN(_06508_ ) );
NAND3_X1 _14477_ ( .A1(_06504_ ), .A2(_06506_ ), .A3(_06508_ ), .ZN(_06509_ ) );
AOI21_X1 _14478_ ( .A(_06490_ ), .B1(_06509_ ), .B2(_05365_ ), .ZN(_06510_ ) );
OAI21_X1 _14479_ ( .A(_03364_ ), .B1(_05725_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06511_ ) );
OAI21_X1 _14480_ ( .A(_06483_ ), .B1(_06510_ ), .B2(_06511_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
OR2_X1 _14481_ ( .A1(_04357_ ), .A2(_05362_ ), .ZN(_06512_ ) );
NOR2_X1 _14482_ ( .A1(_06003_ ), .A2(_06004_ ), .ZN(_06513_ ) );
XNOR2_X1 _14483_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .ZN(_06514_ ) );
AOI21_X1 _14484_ ( .A(_05487_ ), .B1(_06513_ ), .B2(_06514_ ), .ZN(_06515_ ) );
OAI21_X1 _14485_ ( .A(_06515_ ), .B1(_06513_ ), .B2(_06514_ ), .ZN(_06516_ ) );
NAND3_X1 _14486_ ( .A1(_05524_ ), .A2(\ID_EX_imm [29] ), .A3(_05525_ ), .ZN(_06517_ ) );
AND2_X1 _14487_ ( .A1(_06516_ ), .A2(_06517_ ), .ZN(_06518_ ) );
OR2_X1 _14488_ ( .A1(_02308_ ), .A2(_04488_ ), .ZN(_06519_ ) );
NOR2_X1 _14489_ ( .A1(_06038_ ), .A2(_06041_ ), .ZN(_06520_ ) );
INV_X1 _14490_ ( .A(_06013_ ), .ZN(_06521_ ) );
OAI21_X1 _14491_ ( .A(_06519_ ), .B1(_06520_ ), .B2(_06521_ ), .ZN(_06522_ ) );
AOI21_X1 _14492_ ( .A(_04867_ ), .B1(_06522_ ), .B2(_06014_ ), .ZN(_06523_ ) );
OAI21_X1 _14493_ ( .A(_06523_ ), .B1(_06014_ ), .B2(_06522_ ), .ZN(_06524_ ) );
AOI21_X1 _14494_ ( .A(_05509_ ), .B1(_06518_ ), .B2(_06524_ ), .ZN(_06525_ ) );
INV_X1 _14495_ ( .A(_06079_ ), .ZN(_06526_ ) );
AOI21_X1 _14496_ ( .A(_06526_ ), .B1(_06107_ ), .B2(_06116_ ), .ZN(_06527_ ) );
OR3_X1 _14497_ ( .A1(_06527_ ), .A2(_06081_ ), .A3(_06118_ ), .ZN(_06528_ ) );
OAI21_X1 _14498_ ( .A(_06081_ ), .B1(_06527_ ), .B2(_06118_ ), .ZN(_06529_ ) );
NAND3_X1 _14499_ ( .A1(_06528_ ), .A2(_05479_ ), .A3(_06529_ ), .ZN(_06530_ ) );
AND2_X1 _14500_ ( .A1(_05136_ ), .A2(_05193_ ), .ZN(_06531_ ) );
AOI22_X1 _14501_ ( .A1(_05122_ ), .A2(_05119_ ), .B1(_05747_ ), .B2(_06531_ ), .ZN(_06532_ ) );
OR3_X1 _14502_ ( .A1(_05109_ ), .A2(_05728_ ), .A3(_05899_ ), .ZN(_06533_ ) );
NAND2_X1 _14503_ ( .A1(_06532_ ), .A2(_06533_ ), .ZN(_06534_ ) );
NAND2_X1 _14504_ ( .A1(_06534_ ), .A2(_05366_ ), .ZN(_06535_ ) );
NAND3_X1 _14505_ ( .A1(_05203_ ), .A2(_05465_ ), .A3(_05210_ ), .ZN(_06536_ ) );
OR3_X1 _14506_ ( .A1(_05138_ ), .A2(_05144_ ), .A3(_05420_ ), .ZN(_06537_ ) );
OAI211_X1 _14507_ ( .A(_05126_ ), .B(_05444_ ), .C1(_02236_ ), .C2(_05189_ ), .ZN(_06538_ ) );
NAND3_X1 _14508_ ( .A1(_06537_ ), .A2(_05370_ ), .A3(_06538_ ), .ZN(_06539_ ) );
OAI21_X1 _14509_ ( .A(_05444_ ), .B1(_05152_ ), .B2(_05139_ ), .ZN(_06540_ ) );
OAI21_X1 _14510_ ( .A(_05372_ ), .B1(_05148_ ), .B2(_05153_ ), .ZN(_06541_ ) );
AND2_X1 _14511_ ( .A1(_06540_ ), .A2(_06541_ ), .ZN(_06542_ ) );
OAI211_X1 _14512_ ( .A(_06539_ ), .B(_05426_ ), .C1(_06542_ ), .C2(_05744_ ), .ZN(_06543_ ) );
NAND3_X1 _14513_ ( .A1(_06536_ ), .A2(_05553_ ), .A3(_06543_ ), .ZN(_06544_ ) );
AND2_X1 _14514_ ( .A1(_06544_ ), .A2(_05413_ ), .ZN(_06545_ ) );
OAI21_X1 _14515_ ( .A(_06545_ ), .B1(_05467_ ), .B2(_05904_ ), .ZN(_06546_ ) );
OAI21_X1 _14516_ ( .A(_05580_ ), .B1(_06080_ ), .B2(_02214_ ), .ZN(_06547_ ) );
AND3_X1 _14517_ ( .A1(_06531_ ), .A2(_05165_ ), .A3(_05235_ ), .ZN(_06548_ ) );
AOI221_X4 _14518_ ( .A(_06548_ ), .B1(_05475_ ), .B2(_06120_ ), .C1(_05335_ ), .C2(_06081_ ), .ZN(_06549_ ) );
AND4_X1 _14519_ ( .A1(_06535_ ), .A2(_06546_ ), .A3(_06547_ ), .A4(_06549_ ), .ZN(_06550_ ) );
AOI21_X1 _14520_ ( .A(_05528_ ), .B1(_06530_ ), .B2(_06550_ ), .ZN(_06551_ ) );
NOR3_X1 _14521_ ( .A1(_06525_ ), .A2(_06551_ ), .A3(_01362_ ), .ZN(_06552_ ) );
AND4_X1 _14522_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_06553_ ) );
AND4_X1 _14523_ ( .A1(\ID_EX_pc [21] ), .A2(_06553_ ), .A3(\ID_EX_pc [20] ), .A4(_04754_ ), .ZN(_06554_ ) );
AND2_X1 _14524_ ( .A1(_05600_ ), .A2(_06554_ ), .ZN(_06555_ ) );
AND3_X1 _14525_ ( .A1(_06555_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_06556_ ) );
NAND2_X1 _14526_ ( .A1(_06556_ ), .A2(\ID_EX_pc [28] ), .ZN(_06557_ ) );
NAND2_X1 _14527_ ( .A1(_06557_ ), .A2(\ID_EX_pc [29] ), .ZN(_06558_ ) );
NAND3_X1 _14528_ ( .A1(_06556_ ), .A2(_02336_ ), .A3(\ID_EX_pc [28] ), .ZN(_06559_ ) );
NAND3_X1 _14529_ ( .A1(_06558_ ), .A2(_05497_ ), .A3(_06559_ ), .ZN(_06560_ ) );
NAND2_X1 _14530_ ( .A1(_06560_ ), .A2(_03407_ ), .ZN(_06561_ ) );
OAI21_X1 _14531_ ( .A(_06512_ ), .B1(_06552_ ), .B2(_06561_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
NAND3_X1 _14532_ ( .A1(_04397_ ), .A2(_04385_ ), .A3(_03698_ ), .ZN(_06562_ ) );
OR3_X1 _14533_ ( .A1(_04783_ ), .A2(_03359_ ), .A3(_04454_ ), .ZN(_06563_ ) );
NAND3_X1 _14534_ ( .A1(_06563_ ), .A2(_05514_ ), .A3(_04784_ ), .ZN(_06564_ ) );
NOR2_X1 _14535_ ( .A1(_04889_ ), .A2(_04955_ ), .ZN(_06565_ ) );
OAI21_X1 _14536_ ( .A(_06565_ ), .B1(_04888_ ), .B2(_04887_ ), .ZN(_06566_ ) );
NAND3_X1 _14537_ ( .A1(_05491_ ), .A2(\ID_EX_imm [1] ), .A3(_05492_ ), .ZN(_06567_ ) );
AND3_X1 _14538_ ( .A1(_06564_ ), .A2(_06566_ ), .A3(_06567_ ), .ZN(_06568_ ) );
AOI21_X1 _14539_ ( .A(_05669_ ), .B1(_06568_ ), .B2(_01355_ ), .ZN(_06569_ ) );
NOR4_X1 _14540_ ( .A1(_05609_ ), .A2(_05112_ ), .A3(_05116_ ), .A4(_06393_ ), .ZN(_06570_ ) );
NOR3_X1 _14541_ ( .A1(_05220_ ), .A2(_05372_ ), .A3(_05227_ ), .ZN(_06571_ ) );
AOI211_X1 _14542_ ( .A(_05552_ ), .B(_06571_ ), .C1(_05372_ ), .C2(_06462_ ), .ZN(_06572_ ) );
NOR3_X1 _14543_ ( .A1(_06398_ ), .A2(_06397_ ), .A3(_05744_ ), .ZN(_06573_ ) );
OAI21_X1 _14544_ ( .A(_05804_ ), .B1(_06572_ ), .B2(_06573_ ), .ZN(_06574_ ) );
OAI211_X1 _14545_ ( .A(_06574_ ), .B(_05747_ ), .C1(_05427_ ), .C2(_06236_ ), .ZN(_06575_ ) );
NAND2_X1 _14546_ ( .A1(_05694_ ), .A2(_05381_ ), .ZN(_06576_ ) );
NAND2_X1 _14547_ ( .A1(_06575_ ), .A2(_06576_ ), .ZN(_06577_ ) );
OAI21_X1 _14548_ ( .A(_05366_ ), .B1(_06570_ ), .B2(_06577_ ), .ZN(_06578_ ) );
AOI21_X1 _14549_ ( .A(_05709_ ), .B1(_05283_ ), .B2(_05284_ ), .ZN(_06579_ ) );
OAI21_X1 _14550_ ( .A(_06579_ ), .B1(_05284_ ), .B2(_05283_ ), .ZN(_06580_ ) );
NAND2_X1 _14551_ ( .A1(_06577_ ), .A2(_05474_ ), .ZN(_06581_ ) );
AND3_X1 _14552_ ( .A1(_05550_ ), .A2(_05700_ ), .A3(_05444_ ), .ZN(_06582_ ) );
NAND3_X1 _14553_ ( .A1(_06582_ ), .A2(_05427_ ), .A3(_05822_ ), .ZN(_06583_ ) );
NAND2_X1 _14554_ ( .A1(_05282_ ), .A2(_05476_ ), .ZN(_06584_ ) );
NOR2_X1 _14555_ ( .A1(_05281_ ), .A2(_05470_ ), .ZN(_06585_ ) );
AOI21_X1 _14556_ ( .A(_06585_ ), .B1(_05283_ ), .B2(_05472_ ), .ZN(_06586_ ) );
AND4_X1 _14557_ ( .A1(_06581_ ), .A2(_06583_ ), .A3(_06584_ ), .A4(_06586_ ), .ZN(_06587_ ) );
NAND3_X1 _14558_ ( .A1(_06578_ ), .A2(_06580_ ), .A3(_06587_ ), .ZN(_06588_ ) );
AOI21_X1 _14559_ ( .A(_06569_ ), .B1(_06588_ ), .B2(_05365_ ), .ZN(_06589_ ) );
OAI21_X1 _14560_ ( .A(_03364_ ), .B1(_05725_ ), .B2(\ID_EX_pc [1] ), .ZN(_06590_ ) );
OAI21_X1 _14561_ ( .A(_06562_ ), .B1(_06589_ ), .B2(_06590_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
NOR2_X1 _14562_ ( .A1(_06079_ ), .A2(_06081_ ), .ZN(_06591_ ) );
AND3_X1 _14563_ ( .A1(_05068_ ), .A2(_02268_ ), .A3(_05069_ ), .ZN(_06592_ ) );
AOI21_X1 _14564_ ( .A(_02268_ ), .B1(_05068_ ), .B2(_05069_ ), .ZN(_06593_ ) );
NOR3_X1 _14565_ ( .A1(_06076_ ), .A2(_06592_ ), .A3(_06593_ ), .ZN(_06594_ ) );
AND2_X1 _14566_ ( .A1(_06591_ ), .A2(_06594_ ), .ZN(_06595_ ) );
NOR2_X1 _14567_ ( .A1(_06104_ ), .A2(_06105_ ), .ZN(_06596_ ) );
INV_X1 _14568_ ( .A(_06596_ ), .ZN(_06597_ ) );
NOR2_X1 _14569_ ( .A1(_06101_ ), .A2(_06098_ ), .ZN(_06598_ ) );
NAND3_X1 _14570_ ( .A1(_06597_ ), .A2(_06103_ ), .A3(_06598_ ), .ZN(_06599_ ) );
INV_X1 _14571_ ( .A(_06085_ ), .ZN(_06600_ ) );
INV_X1 _14572_ ( .A(_06086_ ), .ZN(_06601_ ) );
NAND3_X1 _14573_ ( .A1(_05242_ ), .A2(_06600_ ), .A3(_06601_ ), .ZN(_06602_ ) );
OR2_X1 _14574_ ( .A1(_05328_ ), .A2(_06602_ ), .ZN(_06603_ ) );
OR2_X1 _14575_ ( .A1(_05309_ ), .A2(_05310_ ), .ZN(_06604_ ) );
NOR4_X1 _14576_ ( .A1(_06603_ ), .A2(_05312_ ), .A3(_05313_ ), .A4(_06604_ ), .ZN(_06605_ ) );
NOR2_X1 _14577_ ( .A1(_05247_ ), .A2(_05246_ ), .ZN(_06606_ ) );
INV_X1 _14578_ ( .A(_06606_ ), .ZN(_06607_ ) );
NOR3_X1 _14579_ ( .A1(_06607_ ), .A2(_05244_ ), .A3(_05243_ ), .ZN(_06608_ ) );
OR3_X1 _14580_ ( .A1(_05254_ ), .A2(_05255_ ), .A3(_05276_ ), .ZN(_06609_ ) );
AND3_X1 _14581_ ( .A1(_06326_ ), .A2(_01707_ ), .A3(_05002_ ), .ZN(_06610_ ) );
OR3_X1 _14582_ ( .A1(_05294_ ), .A2(_04239_ ), .A3(_05231_ ), .ZN(_06611_ ) );
NAND3_X1 _14583_ ( .A1(_04992_ ), .A2(_01657_ ), .A3(_04993_ ), .ZN(_06612_ ) );
AOI211_X1 _14584_ ( .A(_05292_ ), .B(_05295_ ), .C1(_06611_ ), .C2(_06612_ ), .ZN(_06613_ ) );
AOI211_X1 _14585_ ( .A(_06610_ ), .B(_06613_ ), .C1(_01684_ ), .C2(_04999_ ), .ZN(_06614_ ) );
NOR4_X1 _14586_ ( .A1(_05292_ ), .A2(_05294_ ), .A3(_05295_ ), .A4(_05296_ ), .ZN(_06615_ ) );
NOR3_X1 _14587_ ( .A1(_06469_ ), .A2(_04787_ ), .A3(_05125_ ), .ZN(_06616_ ) );
AOI21_X1 _14588_ ( .A(_01601_ ), .B1(_04984_ ), .B2(_04983_ ), .ZN(_06617_ ) );
OR2_X1 _14589_ ( .A1(_06616_ ), .A2(_06617_ ), .ZN(_06618_ ) );
NAND3_X1 _14590_ ( .A1(_04974_ ), .A2(_01571_ ), .A3(_04975_ ), .ZN(_06619_ ) );
OAI21_X1 _14591_ ( .A(_06619_ ), .B1(_05283_ ), .B2(_05226_ ), .ZN(_06620_ ) );
AND3_X1 _14592_ ( .A1(_05288_ ), .A2(_06472_ ), .A3(_06620_ ), .ZN(_06621_ ) );
OAI21_X1 _14593_ ( .A(_06615_ ), .B1(_06618_ ), .B2(_06621_ ), .ZN(_06622_ ) );
AOI211_X1 _14594_ ( .A(_05258_ ), .B(_06609_ ), .C1(_06614_ ), .C2(_06622_ ), .ZN(_06623_ ) );
NOR2_X1 _14595_ ( .A1(_05255_ ), .A2(_05254_ ), .ZN(_06624_ ) );
NOR3_X1 _14596_ ( .A1(_05258_ ), .A2(_04779_ ), .A3(_06276_ ), .ZN(_06625_ ) );
AND3_X1 _14597_ ( .A1(_05006_ ), .A2(_01854_ ), .A3(_05007_ ), .ZN(_06626_ ) );
OAI21_X1 _14598_ ( .A(_06624_ ), .B1(_06625_ ), .B2(_06626_ ), .ZN(_06627_ ) );
OR3_X1 _14599_ ( .A1(_05254_ ), .A2(_04774_ ), .A3(_06198_ ), .ZN(_06628_ ) );
NAND3_X1 _14600_ ( .A1(_05020_ ), .A2(_04771_ ), .A3(_05021_ ), .ZN(_06629_ ) );
NAND3_X1 _14601_ ( .A1(_06627_ ), .A2(_06628_ ), .A3(_06629_ ), .ZN(_06630_ ) );
OAI21_X1 _14602_ ( .A(_06608_ ), .B1(_06623_ ), .B2(_06630_ ), .ZN(_06631_ ) );
NOR3_X1 _14603_ ( .A1(_05243_ ), .A2(_04763_ ), .A3(_05947_ ), .ZN(_06632_ ) );
AND3_X1 _14604_ ( .A1(_05083_ ), .A2(_03850_ ), .A3(_05084_ ), .ZN(_06633_ ) );
OAI21_X1 _14605_ ( .A(_06606_ ), .B1(_06632_ ), .B2(_06633_ ), .ZN(_06634_ ) );
NAND3_X1 _14606_ ( .A1(_05268_ ), .A2(_01738_ ), .A3(_05100_ ), .ZN(_06635_ ) );
NAND3_X1 _14607_ ( .A1(_06631_ ), .A2(_06634_ ), .A3(_06635_ ), .ZN(_06636_ ) );
AND3_X1 _14608_ ( .A1(_05079_ ), .A2(_01760_ ), .A3(_05078_ ), .ZN(_06637_ ) );
OAI21_X1 _14609_ ( .A(_06605_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06638_ ) );
NAND3_X1 _14610_ ( .A1(_05030_ ), .A2(_01945_ ), .A3(_05031_ ), .ZN(_06639_ ) );
NAND3_X1 _14611_ ( .A1(_05583_ ), .A2(_01969_ ), .A3(_05035_ ), .ZN(_06640_ ) );
AOI21_X1 _14612_ ( .A(_06604_ ), .B1(_06639_ ), .B2(_06640_ ), .ZN(_06641_ ) );
AOI21_X1 _14613_ ( .A(_06641_ ), .B1(_04835_ ), .B2(_05076_ ), .ZN(_06642_ ) );
OR3_X1 _14614_ ( .A1(_05309_ ), .A2(_02123_ ), .A3(_05633_ ), .ZN(_06643_ ) );
AOI21_X1 _14615_ ( .A(_06603_ ), .B1(_06642_ ), .B2(_06643_ ), .ZN(_06644_ ) );
AND3_X1 _14616_ ( .A1(_05329_ ), .A2(_02088_ ), .A3(_05073_ ), .ZN(_06645_ ) );
AOI21_X1 _14617_ ( .A(_06645_ ), .B1(_03472_ ), .B2(_05067_ ), .ZN(_06646_ ) );
NOR3_X1 _14618_ ( .A1(_06646_ ), .A2(_06085_ ), .A3(_06086_ ), .ZN(_06647_ ) );
AOI211_X1 _14619_ ( .A(_06644_ ), .B(_06647_ ), .C1(_02042_ ), .C2(_06084_ ), .ZN(_06648_ ) );
AND2_X1 _14620_ ( .A1(_06638_ ), .A2(_06648_ ), .ZN(_06649_ ) );
NAND3_X1 _14621_ ( .A1(_06600_ ), .A2(_02064_ ), .A3(_05048_ ), .ZN(_06650_ ) );
AOI21_X1 _14622_ ( .A(_06599_ ), .B1(_06649_ ), .B2(_06650_ ), .ZN(_06651_ ) );
AND3_X1 _14623_ ( .A1(_06103_ ), .A2(_01496_ ), .A3(_05042_ ), .ZN(_06652_ ) );
AOI21_X1 _14624_ ( .A(_05391_ ), .B1(_05049_ ), .B2(_05050_ ), .ZN(_06653_ ) );
OAI21_X1 _14625_ ( .A(_06598_ ), .B1(_06652_ ), .B2(_06653_ ), .ZN(_06654_ ) );
NAND3_X1 _14626_ ( .A1(_06113_ ), .A2(_02182_ ), .A3(_05038_ ), .ZN(_06655_ ) );
NAND2_X1 _14627_ ( .A1(_05045_ ), .A2(_01472_ ), .ZN(_06656_ ) );
NAND3_X1 _14628_ ( .A1(_06654_ ), .A2(_06655_ ), .A3(_06656_ ), .ZN(_06657_ ) );
OAI21_X1 _14629_ ( .A(_06595_ ), .B1(_06651_ ), .B2(_06657_ ), .ZN(_06658_ ) );
OR3_X1 _14630_ ( .A1(_06081_ ), .A2(_05058_ ), .A3(_02308_ ), .ZN(_06659_ ) );
OAI21_X1 _14631_ ( .A(_06659_ ), .B1(_04348_ ), .B2(_06080_ ), .ZN(_06660_ ) );
NAND2_X1 _14632_ ( .A1(_06660_ ), .A2(_06594_ ), .ZN(_06661_ ) );
NAND3_X1 _14633_ ( .A1(_02380_ ), .A2(_01349_ ), .A3(\ID_EX_typ [2] ), .ZN(_06662_ ) );
NOR2_X1 _14634_ ( .A1(_06592_ ), .A2(_06593_ ), .ZN(_06663_ ) );
AND3_X1 _14635_ ( .A1(_03949_ ), .A2(_05053_ ), .A3(_05054_ ), .ZN(_06664_ ) );
AOI211_X1 _14636_ ( .A(_06592_ ), .B(_06662_ ), .C1(_06663_ ), .C2(_06664_ ), .ZN(_06665_ ) );
AND3_X1 _14637_ ( .A1(_06658_ ), .A2(_06661_ ), .A3(_06665_ ), .ZN(_06666_ ) );
NAND4_X1 _14638_ ( .A1(_05019_ ), .A2(_04994_ ), .A3(_04991_ ), .A4(_05106_ ), .ZN(_06667_ ) );
NOR2_X1 _14639_ ( .A1(_05739_ ), .A2(_05159_ ), .ZN(_06668_ ) );
AND3_X1 _14640_ ( .A1(_06263_ ), .A2(_05408_ ), .A3(_06267_ ), .ZN(_06669_ ) );
AOI21_X1 _14641_ ( .A(_05180_ ), .B1(_06429_ ), .B2(_06430_ ), .ZN(_06670_ ) );
AND2_X1 _14642_ ( .A1(_05110_ ), .A2(_05225_ ), .ZN(_06671_ ) );
NOR3_X1 _14643_ ( .A1(_06671_ ), .A2(_05458_ ), .A3(_05219_ ), .ZN(_06672_ ) );
AOI21_X1 _14644_ ( .A(_06672_ ), .B1(_05415_ ), .B2(_06494_ ), .ZN(_06673_ ) );
AOI21_X1 _14645_ ( .A(_06670_ ), .B1(_05423_ ), .B2(_06673_ ), .ZN(_06674_ ) );
AOI211_X1 _14646_ ( .A(_05232_ ), .B(_06669_ ), .C1(_06674_ ), .C2(_05194_ ), .ZN(_06675_ ) );
OR2_X1 _14647_ ( .A1(_06668_ ), .A2(_06675_ ), .ZN(_06676_ ) );
AOI21_X1 _14648_ ( .A(_04970_ ), .B1(_06667_ ), .B2(_06676_ ), .ZN(_06677_ ) );
NOR3_X1 _14649_ ( .A1(_06668_ ), .A2(_05813_ ), .A3(_06675_ ), .ZN(_06678_ ) );
AND3_X1 _14650_ ( .A1(_05752_ ), .A2(_05804_ ), .A3(_05822_ ), .ZN(_06679_ ) );
NOR4_X1 _14651_ ( .A1(_06666_ ), .A2(_06677_ ), .A3(_06678_ ), .A4(_06679_ ), .ZN(_06680_ ) );
OR3_X1 _14652_ ( .A1(_06671_ ), .A2(_05284_ ), .A3(_05240_ ), .ZN(_06681_ ) );
AOI21_X1 _14653_ ( .A(_05470_ ), .B1(_05189_ ), .B2(_05225_ ), .ZN(_06682_ ) );
NOR3_X1 _14654_ ( .A1(_06671_ ), .A2(_05284_ ), .A3(_05662_ ), .ZN(_06683_ ) );
AOI211_X1 _14655_ ( .A(_06682_ ), .B(_06683_ ), .C1(_05284_ ), .C2(_05476_ ), .ZN(_06684_ ) );
AND3_X1 _14656_ ( .A1(_06680_ ), .A2(_06681_ ), .A3(_06684_ ), .ZN(_06685_ ) );
OAI21_X1 _14657_ ( .A(_05484_ ), .B1(_06685_ ), .B2(_05528_ ), .ZN(_06686_ ) );
AND2_X1 _14658_ ( .A1(_06663_ ), .A2(_06664_ ), .ZN(_06687_ ) );
NOR3_X1 _14659_ ( .A1(_06687_ ), .A2(_05353_ ), .A3(_06593_ ), .ZN(_06688_ ) );
NAND3_X1 _14660_ ( .A1(_06658_ ), .A2(_06688_ ), .A3(_06661_ ), .ZN(_06689_ ) );
XNOR2_X1 _14661_ ( .A(_04454_ ), .B(_03359_ ), .ZN(_06690_ ) );
NAND2_X1 _14662_ ( .A1(_06690_ ), .A2(_05515_ ), .ZN(_06691_ ) );
AND2_X1 _14663_ ( .A1(_06689_ ), .A2(_06691_ ), .ZN(_06692_ ) );
NOR2_X1 _14664_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_06693_ ) );
NOR3_X1 _14665_ ( .A1(_05487_ ), .A2(_04888_ ), .A3(_06693_ ), .ZN(_06694_ ) );
AOI21_X1 _14666_ ( .A(_06694_ ), .B1(\ID_EX_imm [0] ), .B2(_05348_ ), .ZN(_06695_ ) );
AOI21_X1 _14667_ ( .A(_05509_ ), .B1(_06692_ ), .B2(_06695_ ), .ZN(_06696_ ) );
OAI221_X1 _14668_ ( .A(_04248_ ), .B1(\ID_EX_pc [0] ), .B2(_05484_ ), .C1(_06686_ ), .C2(_06696_ ), .ZN(_06697_ ) );
INV_X1 _14669_ ( .A(_04428_ ), .ZN(_06698_ ) );
NAND2_X1 _14670_ ( .A1(_06697_ ), .A2(_06698_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
OR2_X1 _14671_ ( .A1(_04463_ ), .A2(_05362_ ), .ZN(_06699_ ) );
AND3_X1 _14672_ ( .A1(_05999_ ), .A2(_06002_ ), .A3(_05978_ ), .ZN(_06700_ ) );
OR3_X1 _14673_ ( .A1(_06700_ ), .A2(_06003_ ), .A3(_05487_ ), .ZN(_06701_ ) );
NAND3_X1 _14674_ ( .A1(_05524_ ), .A2(\ID_EX_imm [28] ), .A3(_05525_ ), .ZN(_06702_ ) );
AND2_X1 _14675_ ( .A1(_06701_ ), .A2(_06702_ ), .ZN(_06703_ ) );
OAI21_X1 _14676_ ( .A(_05515_ ), .B1(_06520_ ), .B2(_06521_ ), .ZN(_06704_ ) );
NOR3_X1 _14677_ ( .A1(_06038_ ), .A2(_06041_ ), .A3(_06013_ ), .ZN(_06705_ ) );
OR2_X1 _14678_ ( .A1(_06704_ ), .A2(_06705_ ), .ZN(_06706_ ) );
AOI21_X1 _14679_ ( .A(_05509_ ), .B1(_06703_ ), .B2(_06706_ ), .ZN(_06707_ ) );
AND3_X1 _14680_ ( .A1(_06107_ ), .A2(_06116_ ), .A3(_06526_ ), .ZN(_06708_ ) );
OR3_X1 _14681_ ( .A1(_06708_ ), .A2(_06527_ ), .A3(_05709_ ), .ZN(_06709_ ) );
OAI211_X1 _14682_ ( .A(_05108_ ), .B(_05123_ ), .C1(_05452_ ), .C2(_05373_ ), .ZN(_06710_ ) );
NAND3_X1 _14683_ ( .A1(_05407_ ), .A2(_05818_ ), .A3(_05744_ ), .ZN(_06711_ ) );
OAI21_X1 _14684_ ( .A(_06710_ ), .B1(_05381_ ), .B2(_06711_ ), .ZN(_06712_ ) );
OAI21_X1 _14685_ ( .A(_05366_ ), .B1(_05556_ ), .B2(_06712_ ), .ZN(_06713_ ) );
OAI21_X1 _14686_ ( .A(_05465_ ), .B1(_05443_ ), .B2(_05450_ ), .ZN(_06714_ ) );
OR3_X1 _14687_ ( .A1(_05392_ ), .A2(_05396_ ), .A3(_05420_ ), .ZN(_06715_ ) );
OAI211_X1 _14688_ ( .A(_06715_ ), .B(_05370_ ), .C1(_06058_ ), .C2(_05372_ ), .ZN(_06716_ ) );
OR3_X1 _14689_ ( .A1(_05386_ ), .A2(_05415_ ), .A3(_05393_ ), .ZN(_06717_ ) );
OAI211_X1 _14690_ ( .A(_05617_ ), .B(_05372_ ), .C1(_03472_ ), .C2(_05189_ ), .ZN(_06718_ ) );
NAND2_X1 _14691_ ( .A1(_06717_ ), .A2(_06718_ ), .ZN(_06719_ ) );
OAI211_X1 _14692_ ( .A(_06716_ ), .B(_05818_ ), .C1(_05744_ ), .C2(_06719_ ), .ZN(_06720_ ) );
NAND3_X1 _14693_ ( .A1(_06714_ ), .A2(_06720_ ), .A3(_05553_ ), .ZN(_06721_ ) );
AND2_X1 _14694_ ( .A1(_06721_ ), .A2(_05413_ ), .ZN(_06722_ ) );
OAI21_X1 _14695_ ( .A(_06722_ ), .B1(_05467_ ), .B2(_05951_ ), .ZN(_06723_ ) );
NAND3_X1 _14696_ ( .A1(_05058_ ), .A2(_02236_ ), .A3(_05476_ ), .ZN(_06724_ ) );
OR3_X1 _14697_ ( .A1(_06711_ ), .A2(_05380_ ), .A3(_05813_ ), .ZN(_06725_ ) );
NAND2_X1 _14698_ ( .A1(_06079_ ), .A2(_05335_ ), .ZN(_06726_ ) );
OAI21_X1 _14699_ ( .A(_05580_ ), .B1(_05058_ ), .B2(_02236_ ), .ZN(_06727_ ) );
AND3_X1 _14700_ ( .A1(_06725_ ), .A2(_06726_ ), .A3(_06727_ ), .ZN(_06728_ ) );
AND4_X1 _14701_ ( .A1(_06713_ ), .A2(_06723_ ), .A3(_06724_ ), .A4(_06728_ ), .ZN(_06729_ ) );
AOI21_X1 _14702_ ( .A(_05528_ ), .B1(_06709_ ), .B2(_06729_ ), .ZN(_06730_ ) );
NOR3_X1 _14703_ ( .A1(_06707_ ), .A2(_01362_ ), .A3(_06730_ ), .ZN(_06731_ ) );
XNOR2_X1 _14704_ ( .A(_06556_ ), .B(_02346_ ), .ZN(_06732_ ) );
OAI21_X1 _14705_ ( .A(_03364_ ), .B1(_06732_ ), .B2(_05725_ ), .ZN(_06733_ ) );
OAI21_X1 _14706_ ( .A(_06699_ ), .B1(_06731_ ), .B2(_06733_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
OR2_X1 _14707_ ( .A1(_04498_ ), .A2(_05362_ ), .ZN(_06734_ ) );
AND2_X1 _14708_ ( .A1(_06034_ ), .A2(_06037_ ), .ZN(_06735_ ) );
OR2_X1 _14709_ ( .A1(_06735_ ), .A2(_06018_ ), .ZN(_06736_ ) );
INV_X1 _14710_ ( .A(_06039_ ), .ZN(_06737_ ) );
AND3_X1 _14711_ ( .A1(_06736_ ), .A2(_06737_ ), .A3(_06016_ ), .ZN(_06738_ ) );
AOI21_X1 _14712_ ( .A(_06016_ ), .B1(_06736_ ), .B2(_06737_ ), .ZN(_06739_ ) );
OR3_X1 _14713_ ( .A1(_06738_ ), .A2(_06739_ ), .A3(_04867_ ), .ZN(_06740_ ) );
NAND3_X1 _14714_ ( .A1(_05994_ ), .A2(_05996_ ), .A3(_05998_ ), .ZN(_06741_ ) );
OAI21_X1 _14715_ ( .A(_06741_ ), .B1(_02350_ ), .B2(_02183_ ), .ZN(_06742_ ) );
AOI21_X1 _14716_ ( .A(_05487_ ), .B1(_06742_ ), .B2(_05995_ ), .ZN(_06743_ ) );
OAI21_X1 _14717_ ( .A(_06743_ ), .B1(_05995_ ), .B2(_06742_ ), .ZN(_06744_ ) );
NAND3_X1 _14718_ ( .A1(_05524_ ), .A2(\ID_EX_imm [27] ), .A3(_05525_ ), .ZN(_06745_ ) );
AND2_X1 _14719_ ( .A1(_06744_ ), .A2(_06745_ ), .ZN(_06746_ ) );
AOI21_X1 _14720_ ( .A(_05509_ ), .B1(_06740_ ), .B2(_06746_ ), .ZN(_06747_ ) );
NAND2_X1 _14721_ ( .A1(_06097_ ), .A2(_06106_ ), .ZN(_06748_ ) );
AND2_X2 _14722_ ( .A1(_06748_ ), .A2(_06112_ ), .ZN(_06749_ ) );
OR2_X4 _14723_ ( .A1(_06749_ ), .A2(_06114_ ), .ZN(_06750_ ) );
INV_X1 _14724_ ( .A(_06099_ ), .ZN(_06751_ ) );
AND3_X4 _14725_ ( .A1(_06750_ ), .A2(_06113_ ), .A3(_06751_ ), .ZN(_06752_ ) );
AOI21_X1 _14726_ ( .A(_06113_ ), .B1(_06750_ ), .B2(_06751_ ), .ZN(_06753_ ) );
OR3_X2 _14727_ ( .A1(_06752_ ), .A2(_06753_ ), .A3(_05709_ ), .ZN(_06754_ ) );
NAND2_X1 _14728_ ( .A1(_06098_ ), .A2(_05472_ ), .ZN(_06755_ ) );
AOI22_X1 _14729_ ( .A1(_05122_ ), .A2(_05119_ ), .B1(_05553_ ), .B2(_06156_ ), .ZN(_06756_ ) );
OAI211_X1 _14730_ ( .A(_05108_ ), .B(_05123_ ), .C1(_05368_ ), .C2(_05574_ ), .ZN(_06757_ ) );
AOI21_X1 _14731_ ( .A(_04970_ ), .B1(_06756_ ), .B2(_06757_ ), .ZN(_06758_ ) );
OAI21_X1 _14732_ ( .A(_05420_ ), .B1(_05148_ ), .B2(_05153_ ), .ZN(_06759_ ) );
OAI21_X1 _14733_ ( .A(_05415_ ), .B1(_05196_ ), .B2(_05149_ ), .ZN(_06760_ ) );
AND2_X1 _14734_ ( .A1(_06759_ ), .A2(_06760_ ), .ZN(_06761_ ) );
OR3_X1 _14735_ ( .A1(_05138_ ), .A2(_05168_ ), .A3(_05144_ ), .ZN(_06762_ ) );
OR3_X1 _14736_ ( .A1(_05152_ ), .A2(_05139_ ), .A3(_05177_ ), .ZN(_06763_ ) );
NAND2_X1 _14737_ ( .A1(_06762_ ), .A2(_06763_ ), .ZN(_06764_ ) );
MUX2_X1 _14738_ ( .A(_06761_ ), .B(_06764_ ), .S(_05423_ ), .Z(_06765_ ) );
NOR2_X1 _14739_ ( .A1(_06765_ ), .A2(_05452_ ), .ZN(_06766_ ) );
AND3_X1 _14740_ ( .A1(_05533_ ), .A2(_05537_ ), .A3(_05451_ ), .ZN(_06767_ ) );
NOR3_X1 _14741_ ( .A1(_06766_ ), .A2(_05868_ ), .A3(_06767_ ), .ZN(_06768_ ) );
NOR2_X1 _14742_ ( .A1(_05158_ ), .A2(_05164_ ), .ZN(_06769_ ) );
INV_X1 _14743_ ( .A(_06769_ ), .ZN(_06770_ ) );
AOI21_X1 _14744_ ( .A(_06770_ ), .B1(_06169_ ), .B2(_06170_ ), .ZN(_06771_ ) );
AND3_X1 _14745_ ( .A1(_06156_ ), .A2(_05553_ ), .A3(_05235_ ), .ZN(_06772_ ) );
NOR4_X1 _14746_ ( .A1(_06758_ ), .A2(_06768_ ), .A3(_06771_ ), .A4(_06772_ ), .ZN(_06773_ ) );
OAI21_X1 _14747_ ( .A(_05580_ ), .B1(_05093_ ), .B2(_01472_ ), .ZN(_06774_ ) );
NAND3_X1 _14748_ ( .A1(_05093_ ), .A2(_01472_ ), .A3(_05476_ ), .ZN(_06775_ ) );
AND4_X1 _14749_ ( .A1(_06755_ ), .A2(_06773_ ), .A3(_06774_ ), .A4(_06775_ ), .ZN(_06776_ ) );
AOI21_X2 _14750_ ( .A(_05528_ ), .B1(_06754_ ), .B2(_06776_ ), .ZN(_06777_ ) );
NOR3_X1 _14751_ ( .A1(_06747_ ), .A2(_06777_ ), .A3(_01362_ ), .ZN(_06778_ ) );
NAND3_X1 _14752_ ( .A1(_05600_ ), .A2(\ID_EX_pc [26] ), .A3(_06554_ ), .ZN(_06779_ ) );
NAND2_X1 _14753_ ( .A1(_06779_ ), .A2(\ID_EX_pc [27] ), .ZN(_06780_ ) );
NAND4_X1 _14754_ ( .A1(_05600_ ), .A2(_02349_ ), .A3(\ID_EX_pc [26] ), .A4(_06554_ ), .ZN(_06781_ ) );
NAND3_X1 _14755_ ( .A1(_06780_ ), .A2(_05497_ ), .A3(_06781_ ), .ZN(_06782_ ) );
NAND2_X1 _14756_ ( .A1(_06782_ ), .A2(_03407_ ), .ZN(_06783_ ) );
OAI21_X1 _14757_ ( .A(_06734_ ), .B1(_06778_ ), .B2(_06783_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
OR2_X1 _14758_ ( .A1(_04532_ ), .A2(_03357_ ), .ZN(_06784_ ) );
AOI21_X1 _14759_ ( .A(_05182_ ), .B1(_06060_ ), .B2(_06061_ ), .ZN(_06785_ ) );
AND3_X1 _14760_ ( .A1(_06065_ ), .A2(_06066_ ), .A3(_05202_ ), .ZN(_06786_ ) );
OR3_X1 _14761_ ( .A1(_06785_ ), .A2(_06786_ ), .A3(_05408_ ), .ZN(_06787_ ) );
NAND2_X1 _14762_ ( .A1(_06787_ ), .A2(_05821_ ), .ZN(_06788_ ) );
AOI21_X1 _14763_ ( .A(_06788_ ), .B1(_05452_ ), .B2(_05657_ ), .ZN(_06789_ ) );
AOI21_X1 _14764_ ( .A(_06770_ ), .B1(_06193_ ), .B2(_06194_ ), .ZN(_06790_ ) );
OR2_X1 _14765_ ( .A1(_06789_ ), .A2(_06790_ ), .ZN(_06791_ ) );
INV_X1 _14766_ ( .A(_06180_ ), .ZN(_06792_ ) );
AND3_X1 _14767_ ( .A1(_05019_ ), .A2(_05106_ ), .A3(_05574_ ), .ZN(_06793_ ) );
OAI211_X1 _14768_ ( .A(_06793_ ), .B(_05116_ ), .C1(_05372_ ), .C2(_05189_ ), .ZN(_06794_ ) );
AOI21_X1 _14769_ ( .A(_05377_ ), .B1(_06792_ ), .B2(_06794_ ), .ZN(_06795_ ) );
NOR2_X1 _14770_ ( .A1(_05626_ ), .A2(_05409_ ), .ZN(_06796_ ) );
AND2_X1 _14771_ ( .A1(_06796_ ), .A2(_05158_ ), .ZN(_06797_ ) );
OR3_X1 _14772_ ( .A1(_06795_ ), .A2(_05556_ ), .A3(_06797_ ), .ZN(_06798_ ) );
XNOR2_X1 _14773_ ( .A(_06749_ ), .B(_06101_ ), .ZN(_06799_ ) );
AOI221_X4 _14774_ ( .A(_06791_ ), .B1(_05366_ ), .B2(_06798_ ), .C1(_06799_ ), .C2(_05239_ ), .ZN(_06800_ ) );
OAI22_X1 _14775_ ( .A1(_06114_ ), .A2(_05662_ ), .B1(_05344_ ), .B2(_06100_ ), .ZN(_06801_ ) );
AOI221_X4 _14776_ ( .A(_06801_ ), .B1(_05476_ ), .B2(_06099_ ), .C1(_06797_ ), .C2(_05474_ ), .ZN(_06802_ ) );
AOI21_X1 _14777_ ( .A(_05528_ ), .B1(_06800_ ), .B2(_06802_ ), .ZN(_06803_ ) );
NAND2_X1 _14778_ ( .A1(_06741_ ), .A2(_05672_ ), .ZN(_06804_ ) );
AOI21_X1 _14779_ ( .A(_05996_ ), .B1(_05994_ ), .B2(_05998_ ), .ZN(_06805_ ) );
OR2_X1 _14780_ ( .A1(_06804_ ), .A2(_06805_ ), .ZN(_06806_ ) );
NAND3_X1 _14781_ ( .A1(_05491_ ), .A2(\ID_EX_imm [26] ), .A3(_05492_ ), .ZN(_06807_ ) );
AND2_X1 _14782_ ( .A1(_06806_ ), .A2(_06807_ ), .ZN(_06808_ ) );
NAND3_X1 _14783_ ( .A1(_06034_ ), .A2(_06018_ ), .A3(_06037_ ), .ZN(_06809_ ) );
NAND3_X1 _14784_ ( .A1(_06736_ ), .A2(_05515_ ), .A3(_06809_ ), .ZN(_06810_ ) );
AOI21_X1 _14785_ ( .A(_05509_ ), .B1(_06808_ ), .B2(_06810_ ), .ZN(_06811_ ) );
NOR3_X1 _14786_ ( .A1(_06803_ ), .A2(_01362_ ), .A3(_06811_ ), .ZN(_06812_ ) );
AOI21_X1 _14787_ ( .A(_02350_ ), .B1(_05600_ ), .B2(_06554_ ), .ZN(_06813_ ) );
AND4_X1 _14788_ ( .A1(_02350_ ), .A2(_05498_ ), .A3(_04753_ ), .A4(_06554_ ), .ZN(_06814_ ) );
OR3_X1 _14789_ ( .A1(_06813_ ), .A2(_05360_ ), .A3(_06814_ ), .ZN(_06815_ ) );
NAND2_X1 _14790_ ( .A1(_06815_ ), .A2(_04248_ ), .ZN(_06816_ ) );
OAI21_X1 _14791_ ( .A(_06784_ ), .B1(_06812_ ), .B2(_06816_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
OAI21_X1 _14792_ ( .A(_03379_ ), .B1(_04565_ ), .B2(_04566_ ), .ZN(_06817_ ) );
AOI21_X1 _14793_ ( .A(_06035_ ), .B1(_06031_ ), .B2(_06033_ ), .ZN(_06818_ ) );
XNOR2_X1 _14794_ ( .A(_06818_ ), .B(_06032_ ), .ZN(_06819_ ) );
NAND2_X1 _14795_ ( .A1(_06819_ ), .A2(_05514_ ), .ZN(_06820_ ) );
NOR2_X1 _14796_ ( .A1(_05992_ ), .A2(_05997_ ), .ZN(_06821_ ) );
OR3_X1 _14797_ ( .A1(_05991_ ), .A2(_05993_ ), .A3(_06821_ ), .ZN(_06822_ ) );
OAI21_X1 _14798_ ( .A(_06821_ ), .B1(_05991_ ), .B2(_05993_ ), .ZN(_06823_ ) );
NAND3_X1 _14799_ ( .A1(_06822_ ), .A2(_05672_ ), .A3(_06823_ ), .ZN(_06824_ ) );
NAND3_X1 _14800_ ( .A1(_04962_ ), .A2(\ID_EX_imm [25] ), .A3(_04964_ ), .ZN(_06825_ ) );
AND3_X1 _14801_ ( .A1(_06820_ ), .A2(_06824_ ), .A3(_06825_ ), .ZN(_06826_ ) );
AOI21_X1 _14802_ ( .A(_05669_ ), .B1(_06826_ ), .B2(_01355_ ), .ZN(_06827_ ) );
AOI21_X1 _14803_ ( .A(_06597_ ), .B1(_06089_ ), .B2(_06095_ ), .ZN(_06828_ ) );
NOR2_X1 _14804_ ( .A1(_06828_ ), .A2(_06104_ ), .ZN(_06829_ ) );
XNOR2_X1 _14805_ ( .A(_06829_ ), .B(_06102_ ), .ZN(_06830_ ) );
NAND2_X1 _14806_ ( .A1(_06830_ ), .A2(_05479_ ), .ZN(_06831_ ) );
OR3_X1 _14807_ ( .A1(_05198_ ), .A2(_05201_ ), .A3(_05700_ ), .ZN(_06832_ ) );
OAI211_X1 _14808_ ( .A(_05427_ ), .B(_06832_ ), .C1(_06542_ ), .C2(_05552_ ), .ZN(_06833_ ) );
OAI21_X1 _14809_ ( .A(_05466_ ), .B1(_05701_ ), .B2(_05702_ ), .ZN(_06834_ ) );
AOI21_X1 _14810_ ( .A(_05868_ ), .B1(_06833_ ), .B2(_06834_ ), .ZN(_06835_ ) );
NOR3_X1 _14811_ ( .A1(_05051_ ), .A2(_05391_ ), .A3(_05340_ ), .ZN(_06836_ ) );
AOI21_X1 _14812_ ( .A(_06770_ ), .B1(_06242_ ), .B2(_06243_ ), .ZN(_06837_ ) );
NOR3_X1 _14813_ ( .A1(_06835_ ), .A2(_06836_ ), .A3(_06837_ ), .ZN(_06838_ ) );
OAI21_X1 _14814_ ( .A(_05123_ ), .B1(_06180_ ), .B2(_06229_ ), .ZN(_06839_ ) );
AND3_X1 _14815_ ( .A1(_05686_ ), .A2(_05426_ ), .A3(_05687_ ), .ZN(_06840_ ) );
AND2_X1 _14816_ ( .A1(_06840_ ), .A2(_05747_ ), .ZN(_06841_ ) );
AOI21_X1 _14817_ ( .A(_06841_ ), .B1(_05122_ ), .B2(_05119_ ), .ZN(_06842_ ) );
AOI21_X1 _14818_ ( .A(_05799_ ), .B1(_06839_ ), .B2(_06842_ ), .ZN(_06843_ ) );
NOR3_X1 _14819_ ( .A1(_06110_ ), .A2(_06109_ ), .A3(_05662_ ), .ZN(_06844_ ) );
AOI21_X1 _14820_ ( .A(_05470_ ), .B1(_05051_ ), .B2(_05391_ ), .ZN(_06845_ ) );
AND3_X1 _14821_ ( .A1(_06840_ ), .A2(_05467_ ), .A3(_05474_ ), .ZN(_06846_ ) );
NOR4_X1 _14822_ ( .A1(_06843_ ), .A2(_06844_ ), .A3(_06845_ ), .A4(_06846_ ), .ZN(_06847_ ) );
NAND3_X1 _14823_ ( .A1(_06831_ ), .A2(_06838_ ), .A3(_06847_ ), .ZN(_06848_ ) );
AOI21_X1 _14824_ ( .A(_06827_ ), .B1(_06848_ ), .B2(_05365_ ), .ZN(_06849_ ) );
AND3_X1 _14825_ ( .A1(_04754_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_06850_ ) );
AND2_X1 _14826_ ( .A1(_05600_ ), .A2(_06850_ ), .ZN(_06851_ ) );
AND3_X1 _14827_ ( .A1(_06851_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_06852_ ) );
NAND2_X1 _14828_ ( .A1(_06852_ ), .A2(\ID_EX_pc [24] ), .ZN(_06853_ ) );
NAND2_X1 _14829_ ( .A1(_06853_ ), .A2(\ID_EX_pc [25] ), .ZN(_06854_ ) );
NAND3_X1 _14830_ ( .A1(_06852_ ), .A2(_02351_ ), .A3(\ID_EX_pc [24] ), .ZN(_06855_ ) );
NAND3_X1 _14831_ ( .A1(_06854_ ), .A2(_05497_ ), .A3(_06855_ ), .ZN(_06856_ ) );
NAND2_X1 _14832_ ( .A1(_06856_ ), .A2(_04248_ ), .ZN(_06857_ ) );
OAI21_X1 _14833_ ( .A(_06817_ ), .B1(_06849_ ), .B2(_06857_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
INV_X1 _14834_ ( .A(_04604_ ), .ZN(_06858_ ) );
AOI21_X1 _14835_ ( .A(_04867_ ), .B1(_06031_ ), .B2(_06033_ ), .ZN(_06859_ ) );
OAI21_X1 _14836_ ( .A(_06859_ ), .B1(_06031_ ), .B2(_06033_ ), .ZN(_06860_ ) );
AOI21_X1 _14837_ ( .A(_05487_ ), .B1(_05989_ ), .B2(_05990_ ), .ZN(_06861_ ) );
OAI21_X1 _14838_ ( .A(_06861_ ), .B1(_05989_ ), .B2(_05990_ ), .ZN(_06862_ ) );
AND2_X1 _14839_ ( .A1(_06860_ ), .A2(_06862_ ), .ZN(_06863_ ) );
NAND3_X1 _14840_ ( .A1(_05524_ ), .A2(\ID_EX_imm [24] ), .A3(_05525_ ), .ZN(_06864_ ) );
AOI21_X1 _14841_ ( .A(_05509_ ), .B1(_06863_ ), .B2(_06864_ ), .ZN(_06865_ ) );
NAND4_X1 _14842_ ( .A1(_05019_ ), .A2(_06261_ ), .A3(_05106_ ), .A4(_05123_ ), .ZN(_06866_ ) );
NAND3_X1 _14843_ ( .A1(_05732_ ), .A2(_05804_ ), .A3(_05747_ ), .ZN(_06867_ ) );
NAND2_X1 _14844_ ( .A1(_06866_ ), .A2(_06867_ ), .ZN(_06868_ ) );
OAI21_X1 _14845_ ( .A(_05366_ ), .B1(_05556_ ), .B2(_06868_ ), .ZN(_06869_ ) );
NAND2_X1 _14846_ ( .A1(_06719_ ), .A2(_05700_ ), .ZN(_06870_ ) );
NAND3_X1 _14847_ ( .A1(_05446_ ), .A2(_05449_ ), .A3(_05552_ ), .ZN(_06871_ ) );
AOI21_X1 _14848_ ( .A(_05466_ ), .B1(_06870_ ), .B2(_06871_ ), .ZN(_06872_ ) );
AND3_X1 _14849_ ( .A1(_05748_ ), .A2(_05749_ ), .A3(_05452_ ), .ZN(_06873_ ) );
OAI21_X1 _14850_ ( .A(_05822_ ), .B1(_06872_ ), .B2(_06873_ ), .ZN(_06874_ ) );
NOR3_X1 _14851_ ( .A1(_06104_ ), .A2(_05662_ ), .A3(_06105_ ), .ZN(_06875_ ) );
AOI21_X1 _14852_ ( .A(_05344_ ), .B1(_05042_ ), .B2(_05151_ ), .ZN(_06876_ ) );
NOR3_X1 _14853_ ( .A1(_05042_ ), .A2(_05151_ ), .A3(_05340_ ), .ZN(_06877_ ) );
NOR3_X1 _14854_ ( .A1(_06875_ ), .A2(_06876_ ), .A3(_06877_ ), .ZN(_06878_ ) );
NOR2_X1 _14855_ ( .A1(_06867_ ), .A2(_05813_ ), .ZN(_06879_ ) );
AOI21_X1 _14856_ ( .A(_06770_ ), .B1(_06279_ ), .B2(_06280_ ), .ZN(_06880_ ) );
NOR2_X1 _14857_ ( .A1(_06879_ ), .A2(_06880_ ), .ZN(_06881_ ) );
AND4_X1 _14858_ ( .A1(_06869_ ), .A2(_06874_ ), .A3(_06878_ ), .A4(_06881_ ), .ZN(_06882_ ) );
NOR2_X1 _14859_ ( .A1(_06828_ ), .A2(_05709_ ), .ZN(_06883_ ) );
OAI21_X1 _14860_ ( .A(_06883_ ), .B1(_06097_ ), .B2(_06596_ ), .ZN(_06884_ ) );
AOI21_X1 _14861_ ( .A(_05528_ ), .B1(_06882_ ), .B2(_06884_ ), .ZN(_06885_ ) );
NOR3_X1 _14862_ ( .A1(_06865_ ), .A2(_01362_ ), .A3(_06885_ ), .ZN(_06886_ ) );
XNOR2_X1 _14863_ ( .A(_06852_ ), .B(_02352_ ), .ZN(_06887_ ) );
OAI21_X1 _14864_ ( .A(_03364_ ), .B1(_06887_ ), .B2(_05725_ ), .ZN(_06888_ ) );
OAI21_X1 _14865_ ( .A(_06858_ ), .B1(_06886_ ), .B2(_06888_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
NAND4_X1 _14866_ ( .A1(_03690_ ), .A2(_04200_ ), .A3(\mtvec [23] ), .A4(_04072_ ), .ZN(_06889_ ) );
AND2_X1 _14867_ ( .A1(_04634_ ), .A2(_06889_ ), .ZN(_06890_ ) );
NAND4_X1 _14868_ ( .A1(_03768_ ), .A2(_04200_ ), .A3(\mycsreg.CSReg[0][23] ), .A4(_04072_ ), .ZN(_06891_ ) );
AND2_X1 _14869_ ( .A1(_04636_ ), .A2(_06891_ ), .ZN(_06892_ ) );
AOI22_X1 _14870_ ( .A1(_04107_ ), .A2(_04106_ ), .B1(_06890_ ), .B2(_06892_ ), .ZN(_06893_ ) );
AND3_X1 _14871_ ( .A1(_04106_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_04107_ ), .ZN(_06894_ ) );
OAI21_X1 _14872_ ( .A(_03698_ ), .B1(_06893_ ), .B2(_06894_ ), .ZN(_06895_ ) );
OAI21_X1 _14873_ ( .A(_06020_ ), .B1(_04862_ ), .B2(_06024_ ), .ZN(_06896_ ) );
INV_X1 _14874_ ( .A(_06028_ ), .ZN(_06897_ ) );
AND2_X1 _14875_ ( .A1(_06896_ ), .A2(_06897_ ), .ZN(_06898_ ) );
XNOR2_X1 _14876_ ( .A(_06898_ ), .B(_06019_ ), .ZN(_06899_ ) );
NAND2_X1 _14877_ ( .A1(_06899_ ), .A2(_05515_ ), .ZN(_06900_ ) );
NAND2_X1 _14878_ ( .A1(_04959_ ), .A2(_05987_ ), .ZN(_06901_ ) );
AND2_X1 _14879_ ( .A1(_06901_ ), .A2(_05980_ ), .ZN(_06902_ ) );
OR3_X1 _14880_ ( .A1(_06902_ ), .A2(_05979_ ), .A3(_05984_ ), .ZN(_06903_ ) );
OAI21_X1 _14881_ ( .A(_05979_ ), .B1(_06902_ ), .B2(_05984_ ), .ZN(_06904_ ) );
NAND3_X1 _14882_ ( .A1(_06903_ ), .A2(_05672_ ), .A3(_06904_ ), .ZN(_06905_ ) );
AND2_X1 _14883_ ( .A1(_06900_ ), .A2(_06905_ ), .ZN(_06906_ ) );
NAND3_X1 _14884_ ( .A1(_05524_ ), .A2(\ID_EX_imm [23] ), .A3(_05525_ ), .ZN(_06907_ ) );
AOI21_X1 _14885_ ( .A(_05509_ ), .B1(_06906_ ), .B2(_06907_ ), .ZN(_06908_ ) );
AOI211_X1 _14886_ ( .A(_05728_ ), .B(_05109_ ), .C1(_05553_ ), .C2(_05116_ ), .ZN(_06909_ ) );
AND2_X1 _14887_ ( .A1(_06313_ ), .A2(_05159_ ), .ZN(_06910_ ) );
OAI21_X1 _14888_ ( .A(_04969_ ), .B1(_06909_ ), .B2(_06910_ ), .ZN(_06911_ ) );
NAND3_X1 _14889_ ( .A1(_06313_ ), .A2(_05747_ ), .A3(_05235_ ), .ZN(_06912_ ) );
NAND2_X1 _14890_ ( .A1(_06911_ ), .A2(_06912_ ), .ZN(_06913_ ) );
OAI21_X1 _14891_ ( .A(_05413_ ), .B1(_06337_ ), .B2(_05553_ ), .ZN(_06914_ ) );
OAI211_X1 _14892_ ( .A(_05817_ ), .B(_05465_ ), .C1(_05552_ ), .C2(_05819_ ), .ZN(_06915_ ) );
NAND3_X1 _14893_ ( .A1(_06759_ ), .A2(_06760_ ), .A3(_05423_ ), .ZN(_06916_ ) );
NAND3_X1 _14894_ ( .A1(_05534_ ), .A2(_05536_ ), .A3(_05428_ ), .ZN(_06917_ ) );
NAND2_X1 _14895_ ( .A1(_06916_ ), .A2(_06917_ ), .ZN(_06918_ ) );
OAI21_X1 _14896_ ( .A(_06915_ ), .B1(_05452_ ), .B2(_06918_ ), .ZN(_06919_ ) );
AOI21_X1 _14897_ ( .A(_06914_ ), .B1(_05467_ ), .B2(_06919_ ), .ZN(_06920_ ) );
OR2_X1 _14898_ ( .A1(_06913_ ), .A2(_06920_ ), .ZN(_06921_ ) );
AND2_X1 _14899_ ( .A1(_06085_ ), .A2(_05472_ ), .ZN(_06922_ ) );
NOR3_X1 _14900_ ( .A1(_06084_ ), .A2(_05385_ ), .A3(_05340_ ), .ZN(_06923_ ) );
AOI21_X1 _14901_ ( .A(_05470_ ), .B1(_06084_ ), .B2(_05385_ ), .ZN(_06924_ ) );
NOR4_X1 _14902_ ( .A1(_06921_ ), .A2(_06922_ ), .A3(_06923_ ), .A4(_06924_ ), .ZN(_06925_ ) );
AOI211_X1 _14903_ ( .A(_05329_ ), .B(_05242_ ), .C1(_05316_ ), .C2(_05326_ ), .ZN(_06926_ ) );
OAI21_X1 _14904_ ( .A(_06086_ ), .B1(_06926_ ), .B2(_06091_ ), .ZN(_06927_ ) );
OR2_X1 _14905_ ( .A1(_05048_ ), .A2(_05147_ ), .ZN(_06928_ ) );
AND3_X1 _14906_ ( .A1(_06927_ ), .A2(_06085_ ), .A3(_06928_ ), .ZN(_06929_ ) );
AOI21_X1 _14907_ ( .A(_06085_ ), .B1(_06927_ ), .B2(_06928_ ), .ZN(_06930_ ) );
OAI21_X1 _14908_ ( .A(_05479_ ), .B1(_06929_ ), .B2(_06930_ ), .ZN(_06931_ ) );
AOI21_X1 _14909_ ( .A(_05357_ ), .B1(_06925_ ), .B2(_06931_ ), .ZN(_06932_ ) );
NOR3_X1 _14910_ ( .A1(_06908_ ), .A2(_01362_ ), .A3(_06932_ ), .ZN(_06933_ ) );
NAND3_X1 _14911_ ( .A1(_05600_ ), .A2(\ID_EX_pc [22] ), .A3(_06850_ ), .ZN(_06934_ ) );
NAND2_X1 _14912_ ( .A1(_06934_ ), .A2(\ID_EX_pc [23] ), .ZN(_06935_ ) );
NAND4_X1 _14913_ ( .A1(_05600_ ), .A2(_02353_ ), .A3(\ID_EX_pc [22] ), .A4(_06850_ ), .ZN(_06936_ ) );
NAND3_X1 _14914_ ( .A1(_06935_ ), .A2(_05497_ ), .A3(_06936_ ), .ZN(_06937_ ) );
NAND2_X1 _14915_ ( .A1(_06937_ ), .A2(_04248_ ), .ZN(_06938_ ) );
OAI21_X1 _14916_ ( .A(_06895_ ), .B1(_06933_ ), .B2(_06938_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NOR4_X1 _14917_ ( .A1(_05109_ ), .A2(_05116_ ), .A3(_05377_ ), .A4(_05879_ ), .ZN(_06939_ ) );
OAI21_X1 _14918_ ( .A(_06348_ ), .B1(_05862_ ), .B2(_05408_ ), .ZN(_06940_ ) );
AND2_X1 _14919_ ( .A1(_06940_ ), .A2(_05158_ ), .ZN(_06941_ ) );
OR3_X4 _14920_ ( .A1(_05556_ ), .A2(_06939_ ), .A3(_06941_ ), .ZN(_06942_ ) );
AOI22_X1 _14921_ ( .A1(_06942_ ), .A2(_04969_ ), .B1(_05235_ ), .B2(_06941_ ), .ZN(_06943_ ) );
OAI21_X1 _14922_ ( .A(_05413_ ), .B1(_06361_ ), .B2(_05159_ ), .ZN(_06944_ ) );
NAND3_X1 _14923_ ( .A1(_05873_ ), .A2(_05409_ ), .A3(_05874_ ), .ZN(_06945_ ) );
NAND3_X1 _14924_ ( .A1(_06064_ ), .A2(_06068_ ), .A3(_05425_ ), .ZN(_06946_ ) );
AND3_X1 _14925_ ( .A1(_06945_ ), .A2(_06946_ ), .A3(_05165_ ), .ZN(_06947_ ) );
OR2_X1 _14926_ ( .A1(_06944_ ), .A2(_06947_ ), .ZN(_06948_ ) );
NAND2_X1 _14927_ ( .A1(_06943_ ), .A2(_06948_ ), .ZN(_06949_ ) );
AND2_X1 _14928_ ( .A1(_06086_ ), .A2(_05335_ ), .ZN(_06950_ ) );
NOR3_X1 _14929_ ( .A1(_05048_ ), .A2(_05147_ ), .A3(_05340_ ), .ZN(_06951_ ) );
AOI21_X1 _14930_ ( .A(_05344_ ), .B1(_05048_ ), .B2(_05147_ ), .ZN(_06952_ ) );
NOR4_X1 _14931_ ( .A1(_06949_ ), .A2(_06950_ ), .A3(_06951_ ), .A4(_06952_ ), .ZN(_06953_ ) );
OR3_X1 _14932_ ( .A1(_06926_ ), .A2(_06086_ ), .A3(_06091_ ), .ZN(_06954_ ) );
NAND3_X1 _14933_ ( .A1(_06954_ ), .A2(_05239_ ), .A3(_06927_ ), .ZN(_06955_ ) );
AOI21_X1 _14934_ ( .A(_05356_ ), .B1(_06953_ ), .B2(_06955_ ), .ZN(_06956_ ) );
OR3_X1 _14935_ ( .A1(_04862_ ), .A2(_06024_ ), .A3(_06020_ ), .ZN(_06957_ ) );
NAND3_X1 _14936_ ( .A1(_06957_ ), .A2(_05514_ ), .A3(_06896_ ), .ZN(_06958_ ) );
AOI21_X1 _14937_ ( .A(_04955_ ), .B1(_06901_ ), .B2(_05980_ ), .ZN(_06959_ ) );
OAI21_X1 _14938_ ( .A(_06959_ ), .B1(_05980_ ), .B2(_06901_ ), .ZN(_06960_ ) );
NAND3_X1 _14939_ ( .A1(_04962_ ), .A2(\ID_EX_imm [22] ), .A3(_04964_ ), .ZN(_06961_ ) );
AND2_X1 _14940_ ( .A1(_06960_ ), .A2(_06961_ ), .ZN(_06962_ ) );
AOI21_X1 _14941_ ( .A(_05355_ ), .B1(_06958_ ), .B2(_06962_ ), .ZN(_06963_ ) );
OAI21_X1 _14942_ ( .A(_05360_ ), .B1(_06956_ ), .B2(_06963_ ), .ZN(_06964_ ) );
XNOR2_X1 _14943_ ( .A(_06851_ ), .B(\ID_EX_pc [22] ), .ZN(_06965_ ) );
OAI21_X1 _14944_ ( .A(_06964_ ), .B1(_05484_ ), .B2(_06965_ ), .ZN(_06966_ ) );
MUX2_X1 _14945_ ( .A(_04679_ ), .B(_06966_ ), .S(_05362_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NAND3_X1 _14946_ ( .A1(_04719_ ), .A2(_04708_ ), .A3(_03698_ ), .ZN(_06967_ ) );
INV_X1 _14947_ ( .A(_06076_ ), .ZN(_06968_ ) );
NOR2_X1 _14948_ ( .A1(_06123_ ), .A2(_06968_ ), .ZN(_06969_ ) );
INV_X1 _14949_ ( .A(_06663_ ), .ZN(_06970_ ) );
OR3_X1 _14950_ ( .A1(_06969_ ), .A2(_06074_ ), .A3(_06970_ ), .ZN(_06971_ ) );
OAI21_X1 _14951_ ( .A(_06970_ ), .B1(_06969_ ), .B2(_06074_ ), .ZN(_06972_ ) );
NAND3_X1 _14952_ ( .A1(_06971_ ), .A2(_05479_ ), .A3(_06972_ ), .ZN(_06973_ ) );
NAND3_X1 _14953_ ( .A1(_05816_ ), .A2(_05820_ ), .A3(_06769_ ), .ZN(_06974_ ) );
OR3_X1 _14954_ ( .A1(_05070_ ), .A2(_04707_ ), .A3(_05339_ ), .ZN(_06975_ ) );
AOI21_X1 _14955_ ( .A(_05344_ ), .B1(_05070_ ), .B2(_04707_ ), .ZN(_06976_ ) );
AOI21_X1 _14956_ ( .A(_06976_ ), .B1(_06970_ ), .B2(_05335_ ), .ZN(_06977_ ) );
NAND3_X1 _14957_ ( .A1(_04982_ ), .A2(_02268_ ), .A3(_05194_ ), .ZN(_06978_ ) );
OR3_X1 _14958_ ( .A1(_06978_ ), .A2(_05232_ ), .A3(_05635_ ), .ZN(_06979_ ) );
NAND4_X1 _14959_ ( .A1(_06974_ ), .A2(_06975_ ), .A3(_06977_ ), .A4(_06979_ ), .ZN(_06980_ ) );
OAI211_X1 _14960_ ( .A(_05126_ ), .B(_05415_ ), .C1(_02236_ ), .C2(_05189_ ), .ZN(_06981_ ) );
OAI211_X1 _14961_ ( .A(_05420_ ), .B(_05132_ ), .C1(_05371_ ), .C2(_02268_ ), .ZN(_06982_ ) );
NAND2_X1 _14962_ ( .A1(_06981_ ), .A2(_06982_ ), .ZN(_06983_ ) );
MUX2_X1 _14963_ ( .A(_06983_ ), .B(_06764_ ), .S(_05399_ ), .Z(_06984_ ) );
MUX2_X1 _14964_ ( .A(_06918_ ), .B(_06984_ ), .S(_05426_ ), .Z(_06985_ ) );
OAI22_X1 _14965_ ( .A1(_05109_ ), .A2(_05728_ ), .B1(_05381_ ), .B2(_06978_ ), .ZN(_06986_ ) );
AOI221_X4 _14966_ ( .A(_06980_ ), .B1(_05822_ ), .B2(_06985_ ), .C1(_06986_ ), .C2(_05366_ ), .ZN(_06987_ ) );
AOI21_X1 _14967_ ( .A(_05528_ ), .B1(_06973_ ), .B2(_06987_ ), .ZN(_06988_ ) );
OAI21_X1 _14968_ ( .A(_06047_ ), .B1(_01446_ ), .B2(_03935_ ), .ZN(_06989_ ) );
XNOR2_X1 _14969_ ( .A(_04741_ ), .B(_02268_ ), .ZN(_06990_ ) );
AOI21_X1 _14970_ ( .A(_04867_ ), .B1(_06989_ ), .B2(_06990_ ), .ZN(_06991_ ) );
OAI21_X1 _14971_ ( .A(_06991_ ), .B1(_06989_ ), .B2(_06990_ ), .ZN(_06992_ ) );
NAND2_X1 _14972_ ( .A1(_06007_ ), .A2(_06008_ ), .ZN(_06993_ ) );
OAI21_X1 _14973_ ( .A(_06993_ ), .B1(_02325_ ), .B2(_01447_ ), .ZN(_06994_ ) );
XOR2_X1 _14974_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .Z(_06995_ ) );
OR2_X1 _14975_ ( .A1(_06994_ ), .A2(_06995_ ), .ZN(_06996_ ) );
AOI21_X1 _14976_ ( .A(_05487_ ), .B1(_06994_ ), .B2(_06995_ ), .ZN(_06997_ ) );
NAND2_X1 _14977_ ( .A1(_06996_ ), .A2(_06997_ ), .ZN(_06998_ ) );
NAND3_X1 _14978_ ( .A1(_05524_ ), .A2(\ID_EX_imm [31] ), .A3(_05525_ ), .ZN(_06999_ ) );
NAND4_X1 _14979_ ( .A1(_06992_ ), .A2(_01355_ ), .A3(_06998_ ), .A4(_06999_ ), .ZN(_07000_ ) );
AOI21_X1 _14980_ ( .A(_06988_ ), .B1(_07000_ ), .B2(_01360_ ), .ZN(_07001_ ) );
AND2_X1 _14981_ ( .A1(_05975_ ), .A2(\ID_EX_pc [30] ), .ZN(_07002_ ) );
OAI21_X1 _14982_ ( .A(_05497_ ), .B1(_07002_ ), .B2(_02324_ ), .ZN(_07003_ ) );
AND3_X1 _14983_ ( .A1(_05975_ ), .A2(_02324_ ), .A3(\ID_EX_pc [30] ), .ZN(_07004_ ) );
OAI21_X1 _14984_ ( .A(_03364_ ), .B1(_07003_ ), .B2(_07004_ ), .ZN(_07005_ ) );
OAI21_X1 _14985_ ( .A(_06967_ ), .B1(_07001_ ), .B2(_07005_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
NOR4_X1 _14986_ ( .A1(_01347_ ), .A2(fanout_net_4 ), .A3(EXU_valid_LSU ), .A4(excp_written ), .ZN(\myexu.state_$_OR__B_Y_$_ANDNOT__B_Y ) );
AOI21_X1 _14987_ ( .A(_01343_ ), .B1(_01344_ ), .B2(_01340_ ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _14988_ ( .A(IDU_ready_IFU ), .ZN(_07006_ ) );
NAND2_X1 _14989_ ( .A1(_07006_ ), .A2(IDU_valid_EXU ), .ZN(_07007_ ) );
OAI21_X1 _14990_ ( .A(_07007_ ), .B1(_02599_ ), .B2(_02592_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _14991_ ( .A1(_02591_ ), .A2(_02592_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _14992_ ( .A(_02525_ ), .ZN(_07008_ ) );
AND4_X1 _14993_ ( .A1(_02432_ ), .A2(_02434_ ), .A3(_02436_ ), .A4(_02439_ ), .ZN(_07009_ ) );
AND2_X1 _14994_ ( .A1(_02476_ ), .A2(_07009_ ), .ZN(_07010_ ) );
INV_X1 _14995_ ( .A(_07010_ ), .ZN(_07011_ ) );
AOI211_X1 _14996_ ( .A(_07006_ ), .B(_07008_ ), .C1(_02400_ ), .C2(_07011_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _14997_ ( .A1(_02591_ ), .A2(_02592_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14998_ ( .A1(_02591_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_02403_ ), .A4(_07008_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _14999_ ( .A1(_02916_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_02403_ ), .A4(_02524_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _15000_ ( .A(_03074_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _15001_ ( .A(_07007_ ), .B1(_07008_ ), .B2(_07006_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _15002_ ( .A1(_02525_ ), .A2(_07006_ ), .B1(_01217_ ), .B2(_01347_ ), .ZN(_07012_ ) );
INV_X1 _15003_ ( .A(loaduse_clear ), .ZN(_07013_ ) );
AOI221_X4 _15004_ ( .A(_07012_ ), .B1(\myidu.state [2] ), .B2(_07013_ ), .C1(_02591_ ), .C2(_03074_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
NAND3_X1 _15005_ ( .A1(_02450_ ), .A2(IDU_valid_EXU ), .A3(_03128_ ), .ZN(_07014_ ) );
NAND3_X1 _15006_ ( .A1(_02450_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_07015_ ) );
AOI21_X1 _15007_ ( .A(_02651_ ), .B1(_02641_ ), .B2(_02399_ ), .ZN(_07016_ ) );
OAI211_X1 _15008_ ( .A(_02586_ ), .B(_02552_ ), .C1(_02537_ ), .C2(_02545_ ), .ZN(_07017_ ) );
NOR4_X1 _15009_ ( .A1(_02564_ ), .A2(_02565_ ), .A3(_07017_ ), .A4(_02569_ ), .ZN(_07018_ ) );
AND2_X2 _15010_ ( .A1(_02576_ ), .A2(_02676_ ), .ZN(_07019_ ) );
AOI21_X1 _15011_ ( .A(_02659_ ), .B1(_07018_ ), .B2(_07019_ ), .ZN(_07020_ ) );
OR2_X1 _15012_ ( .A1(_07016_ ), .A2(_07020_ ), .ZN(_07021_ ) );
NAND3_X1 _15013_ ( .A1(_02741_ ), .A2(_02402_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_E ), .ZN(_07022_ ) );
OAI211_X1 _15014_ ( .A(_07014_ ), .B(_07015_ ), .C1(_07021_ ), .C2(_07022_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI221_X1 _15015_ ( .A(_02450_ ), .B1(EXU_valid_LSU ), .B2(_01347_ ), .C1(_02525_ ), .C2(_07006_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _15016_ ( .A(_02450_ ), .B(_02526_ ), .C1(_07016_ ), .C2(_07020_ ), .ZN(_07023_ ) );
NAND3_X1 _15017_ ( .A1(_02450_ ), .A2(\myidu.state [2] ), .A3(_07013_ ), .ZN(_07024_ ) );
NAND2_X1 _15018_ ( .A1(_07023_ ), .A2(_07024_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _15019_ ( .A1(_03072_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_07025_ ) );
NOR2_X1 _15020_ ( .A1(_03072_ ), .A2(IDU_ready_IFU ), .ZN(_07026_ ) );
OR2_X1 _15021_ ( .A1(_07026_ ), .A2(fanout_net_4 ), .ZN(_07027_ ) );
AOI211_X1 _15022_ ( .A(_07025_ ), .B(_07027_ ), .C1(_01201_ ), .C2(_03072_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
NAND3_X1 _15023_ ( .A1(_01201_ ), .A2(_03072_ ), .A3(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_07028_ ) );
NAND2_X1 _15024_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_07029_ ) );
NAND3_X1 _15025_ ( .A1(_07028_ ), .A2(_02524_ ), .A3(_07029_ ), .ZN(_07030_ ) );
NOR3_X1 _15026_ ( .A1(_01202_ ), .A2(_07027_ ), .A3(_07030_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__A_Y ) );
AND3_X1 _15027_ ( .A1(_03178_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_03179_ ), .ZN(_07031_ ) );
AOI21_X1 _15028_ ( .A(_07031_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B2(_03182_ ), .ZN(_07032_ ) );
MUX2_X1 _15029_ ( .A(\io_master_rdata [31] ), .B(_07032_ ), .S(_02360_ ), .Z(_07033_ ) );
AND2_X1 _15030_ ( .A1(_07033_ ), .A2(_01314_ ), .ZN(\myifu.data_in [31] ) );
OR2_X1 _15031_ ( .A1(_02361_ ), .A2(\io_master_rdata [30] ), .ZN(_07034_ ) );
BUF_X4 _15032_ ( .A(_01324_ ), .Z(_07035_ ) );
BUF_X4 _15033_ ( .A(_07035_ ), .Z(_07036_ ) );
BUF_X4 _15034_ ( .A(_01326_ ), .Z(_07037_ ) );
BUF_X4 _15035_ ( .A(_07037_ ), .Z(_07038_ ) );
BUF_X4 _15036_ ( .A(_02357_ ), .Z(_07039_ ) );
BUF_X4 _15037_ ( .A(_07039_ ), .Z(_07040_ ) );
MUX2_X1 _15038_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03182_ ), .Z(_07041_ ) );
NAND4_X1 _15039_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07041_ ), .ZN(_07042_ ) );
AND3_X1 _15040_ ( .A1(_07034_ ), .A2(_01314_ ), .A3(_07042_ ), .ZN(\myifu.data_in [30] ) );
OR2_X1 _15041_ ( .A1(_03201_ ), .A2(\io_master_rdata [21] ), .ZN(_07043_ ) );
MUX2_X1 _15042_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\io_master_araddr [2] ), .Z(_07044_ ) );
NAND4_X1 _15043_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07044_ ), .ZN(_07045_ ) );
AND3_X1 _15044_ ( .A1(_07043_ ), .A2(_01277_ ), .A3(_07045_ ), .ZN(\myifu.data_in [21] ) );
OR2_X1 _15045_ ( .A1(_02360_ ), .A2(\io_master_rdata [20] ), .ZN(_07046_ ) );
NAND2_X1 _15046_ ( .A1(_03182_ ), .A2(_00823_ ), .ZN(_07047_ ) );
BUF_X4 _15047_ ( .A(_03181_ ), .Z(_07048_ ) );
OAI211_X1 _15048_ ( .A(_03200_ ), .B(_07047_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_07048_ ), .ZN(_07049_ ) );
AND3_X1 _15049_ ( .A1(_07046_ ), .A2(_07049_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [20] ) );
OR2_X4 _15050_ ( .A1(_02360_ ), .A2(\io_master_rdata [19] ), .ZN(_07050_ ) );
MUX2_X1 _15051_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03180_ ), .Z(_07051_ ) );
NAND4_X1 _15052_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07051_ ), .ZN(_07052_ ) );
AND3_X1 _15053_ ( .A1(_07050_ ), .A2(_01277_ ), .A3(_07052_ ), .ZN(\myifu.data_in [19] ) );
OR2_X2 _15054_ ( .A1(_02360_ ), .A2(\io_master_rdata [18] ), .ZN(_07053_ ) );
NAND2_X1 _15055_ ( .A1(_03182_ ), .A2(_00833_ ), .ZN(_07054_ ) );
OAI211_X1 _15056_ ( .A(_03200_ ), .B(_07054_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_07048_ ), .ZN(_07055_ ) );
AND3_X1 _15057_ ( .A1(_07053_ ), .A2(_07055_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [18] ) );
NOR2_X4 _15058_ ( .A1(_02361_ ), .A2(\io_master_rdata [17] ), .ZN(_07056_ ) );
MUX2_X1 _15059_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03180_ ), .Z(_07057_ ) );
AND4_X1 _15060_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07057_ ), .ZN(_07058_ ) );
NOR3_X1 _15061_ ( .A1(_07056_ ), .A2(_01258_ ), .A3(_07058_ ), .ZN(\myifu.data_in [17] ) );
OR2_X2 _15062_ ( .A1(_02360_ ), .A2(\io_master_rdata [16] ), .ZN(_07059_ ) );
NAND2_X1 _15063_ ( .A1(_03182_ ), .A2(_00842_ ), .ZN(_07060_ ) );
OAI211_X1 _15064_ ( .A(_03200_ ), .B(_07060_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_07048_ ), .ZN(_07061_ ) );
AND3_X1 _15065_ ( .A1(_07059_ ), .A2(_07061_ ), .A3(_01314_ ), .ZN(\myifu.data_in [16] ) );
MUX2_X1 _15066_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03180_ ), .Z(_07062_ ) );
NAND4_X1 _15067_ ( .A1(_01324_ ), .A2(_01326_ ), .A3(_02357_ ), .A4(_07062_ ), .ZN(_07063_ ) );
OAI21_X2 _15068_ ( .A(_07063_ ), .B1(_02360_ ), .B2(\io_master_rdata [15] ), .ZN(_07064_ ) );
NOR2_X1 _15069_ ( .A1(_07064_ ), .A2(_03167_ ), .ZN(\myifu.data_in [15] ) );
OR2_X1 _15070_ ( .A1(_03201_ ), .A2(\io_master_rdata [14] ), .ZN(_07065_ ) );
MUX2_X1 _15071_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_07048_ ), .Z(_07066_ ) );
NAND4_X1 _15072_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07066_ ), .ZN(_07067_ ) );
AND3_X1 _15073_ ( .A1(_07065_ ), .A2(_01277_ ), .A3(_07067_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _15074_ ( .A1(_03202_ ), .A2(\io_master_rdata [13] ), .ZN(_07068_ ) );
MUX2_X1 _15075_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\io_master_araddr [2] ), .Z(_07069_ ) );
NAND4_X1 _15076_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07069_ ), .ZN(_07070_ ) );
AND3_X1 _15077_ ( .A1(_07068_ ), .A2(\io_master_arburst [0] ), .A3(_07070_ ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _15078_ ( .A1(_03201_ ), .A2(\io_master_rdata [12] ), .ZN(_07071_ ) );
NAND2_X1 _15079_ ( .A1(\io_master_araddr [2] ), .A2(_00857_ ), .ZN(_07072_ ) );
OAI211_X1 _15080_ ( .A(_03201_ ), .B(_07072_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_07073_ ) );
AND3_X1 _15081_ ( .A1(_07071_ ), .A2(_07073_ ), .A3(_01277_ ), .ZN(\myifu.data_in [12] ) );
MUX2_X1 _15082_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\io_master_araddr [2] ), .Z(_07074_ ) );
NAND4_X1 _15083_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07074_ ), .ZN(_07075_ ) );
OAI21_X1 _15084_ ( .A(_07075_ ), .B1(_03202_ ), .B2(\io_master_rdata [29] ), .ZN(_07076_ ) );
NOR2_X1 _15085_ ( .A1(_07076_ ), .A2(_01258_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _15086_ ( .A1(_03200_ ), .A2(\io_master_rdata [11] ), .ZN(_07077_ ) );
MUX2_X1 _15087_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03181_ ), .Z(_07078_ ) );
NAND4_X1 _15088_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07078_ ), .ZN(_07079_ ) );
AND3_X1 _15089_ ( .A1(_07077_ ), .A2(_01277_ ), .A3(_07079_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _15090_ ( .A1(_03201_ ), .A2(\io_master_rdata [10] ), .ZN(_07080_ ) );
MUX2_X1 _15091_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\io_master_araddr [2] ), .Z(_07081_ ) );
NAND4_X1 _15092_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07081_ ), .ZN(_07082_ ) );
AND3_X1 _15093_ ( .A1(_07080_ ), .A2(_01277_ ), .A3(_07082_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _15094_ ( .A1(_03201_ ), .A2(\io_master_rdata [9] ), .ZN(_07083_ ) );
MUX2_X1 _15095_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_07048_ ), .Z(_07084_ ) );
NAND4_X1 _15096_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07084_ ), .ZN(_07085_ ) );
AND3_X1 _15097_ ( .A1(_07083_ ), .A2(\io_master_arburst [0] ), .A3(_07085_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _15098_ ( .A1(_03201_ ), .A2(\io_master_rdata [8] ), .ZN(_07086_ ) );
NAND2_X1 _15099_ ( .A1(\io_master_araddr [2] ), .A2(_00872_ ), .ZN(_07087_ ) );
OAI211_X1 _15100_ ( .A(_03201_ ), .B(_07087_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_07088_ ) );
AND3_X1 _15101_ ( .A1(_07086_ ), .A2(_07088_ ), .A3(_01314_ ), .ZN(\myifu.data_in [8] ) );
MUX2_X1 _15102_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03182_ ), .Z(_07089_ ) );
NAND4_X1 _15103_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07089_ ), .ZN(_07090_ ) );
OAI21_X1 _15104_ ( .A(_07090_ ), .B1(_02361_ ), .B2(\io_master_rdata [7] ), .ZN(_07091_ ) );
NOR2_X1 _15105_ ( .A1(_07091_ ), .A2(_01258_ ), .ZN(\myifu.data_in [7] ) );
NAND2_X1 _15106_ ( .A1(_07048_ ), .A2(_00878_ ), .ZN(_07092_ ) );
OAI211_X1 _15107_ ( .A(_03200_ ), .B(_07092_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_07048_ ), .ZN(_07093_ ) );
OAI21_X1 _15108_ ( .A(_07093_ ), .B1(\io_master_rdata [6] ), .B2(_02361_ ), .ZN(_07094_ ) );
NOR2_X1 _15109_ ( .A1(_07094_ ), .A2(_01258_ ), .ZN(\myifu.data_in [6] ) );
MUX2_X1 _15110_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\io_master_araddr [2] ), .Z(_07095_ ) );
NAND4_X1 _15111_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07095_ ), .ZN(_07096_ ) );
OAI21_X1 _15112_ ( .A(_07096_ ), .B1(_03202_ ), .B2(\io_master_rdata [5] ), .ZN(_07097_ ) );
NOR2_X1 _15113_ ( .A1(_07097_ ), .A2(_03167_ ), .ZN(\myifu.data_in [5] ) );
NAND2_X1 _15114_ ( .A1(_03182_ ), .A2(_00886_ ), .ZN(_07098_ ) );
OAI211_X1 _15115_ ( .A(_03200_ ), .B(_07098_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_07048_ ), .ZN(_07099_ ) );
OAI21_X1 _15116_ ( .A(_07099_ ), .B1(\io_master_rdata [4] ), .B2(_02361_ ), .ZN(_07100_ ) );
NOR2_X1 _15117_ ( .A1(_07100_ ), .A2(_01258_ ), .ZN(\myifu.data_in [4] ) );
MUX2_X1 _15118_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03180_ ), .Z(_07101_ ) );
NAND4_X1 _15119_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07101_ ), .ZN(_07102_ ) );
OAI21_X1 _15120_ ( .A(_07102_ ), .B1(_02360_ ), .B2(\io_master_rdata [3] ), .ZN(_07103_ ) );
NOR2_X1 _15121_ ( .A1(_07103_ ), .A2(_03167_ ), .ZN(\myifu.data_in [3] ) );
NAND2_X1 _15122_ ( .A1(_03182_ ), .A2(_00892_ ), .ZN(_07104_ ) );
OAI211_X1 _15123_ ( .A(_03200_ ), .B(_07104_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_07048_ ), .ZN(_07105_ ) );
OAI21_X1 _15124_ ( .A(_07105_ ), .B1(\io_master_rdata [2] ), .B2(_03200_ ), .ZN(_07106_ ) );
NOR2_X1 _15125_ ( .A1(_07106_ ), .A2(_03167_ ), .ZN(\myifu.data_in [2] ) );
OR2_X1 _15126_ ( .A1(_02359_ ), .A2(\io_master_rdata [28] ), .ZN(_07107_ ) );
NAND2_X1 _15127_ ( .A1(_03181_ ), .A2(_00863_ ), .ZN(_07108_ ) );
OAI211_X2 _15128_ ( .A(_02360_ ), .B(_07108_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03181_ ), .ZN(_07109_ ) );
AND3_X1 _15129_ ( .A1(_07107_ ), .A2(_07109_ ), .A3(_01277_ ), .ZN(\myifu.data_in [28] ) );
MUX2_X1 _15130_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03181_ ), .Z(_07110_ ) );
NAND4_X1 _15131_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07110_ ), .ZN(_07111_ ) );
OAI21_X1 _15132_ ( .A(_07111_ ), .B1(_02361_ ), .B2(\io_master_rdata [1] ), .ZN(_07112_ ) );
NOR2_X1 _15133_ ( .A1(_07112_ ), .A2(_01258_ ), .ZN(\myifu.data_in [1] ) );
MUX2_X1 _15134_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .B(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .S(_03181_ ), .Z(_07113_ ) );
NAND4_X1 _15135_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07113_ ), .ZN(_07114_ ) );
OAI21_X1 _15136_ ( .A(_07114_ ), .B1(_02361_ ), .B2(\io_master_rdata [0] ), .ZN(_07115_ ) );
NOR2_X1 _15137_ ( .A1(_07115_ ), .A2(_03167_ ), .ZN(\myifu.data_in [0] ) );
OR2_X4 _15138_ ( .A1(_02360_ ), .A2(\io_master_rdata [27] ), .ZN(_07116_ ) );
MUX2_X1 _15139_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03180_ ), .Z(_07117_ ) );
NAND4_X1 _15140_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07117_ ), .ZN(_07118_ ) );
AND3_X1 _15141_ ( .A1(_07116_ ), .A2(\io_master_arburst [0] ), .A3(_07118_ ), .ZN(\myifu.data_in [27] ) );
OR2_X4 _15142_ ( .A1(_02359_ ), .A2(\io_master_rdata [26] ), .ZN(_07119_ ) );
MUX2_X1 _15143_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03180_ ), .Z(_07120_ ) );
NAND4_X1 _15144_ ( .A1(_01324_ ), .A2(_01326_ ), .A3(_02357_ ), .A4(_07120_ ), .ZN(_07121_ ) );
AND3_X1 _15145_ ( .A1(_07119_ ), .A2(_01277_ ), .A3(_07121_ ), .ZN(\myifu.data_in [26] ) );
OR2_X1 _15146_ ( .A1(_03201_ ), .A2(\io_master_rdata [25] ), .ZN(_07122_ ) );
MUX2_X1 _15147_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_07048_ ), .Z(_07123_ ) );
NAND4_X1 _15148_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07123_ ), .ZN(_07124_ ) );
AND3_X1 _15149_ ( .A1(_07122_ ), .A2(\io_master_arburst [0] ), .A3(_07124_ ), .ZN(\myifu.data_in [25] ) );
OR2_X4 _15150_ ( .A1(_02359_ ), .A2(\io_master_rdata [24] ), .ZN(_07125_ ) );
NAND2_X1 _15151_ ( .A1(_03181_ ), .A2(_00993_ ), .ZN(_07126_ ) );
OAI211_X1 _15152_ ( .A(_02359_ ), .B(_07126_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03181_ ), .ZN(_07127_ ) );
AND3_X1 _15153_ ( .A1(_07125_ ), .A2(_07127_ ), .A3(_01314_ ), .ZN(\myifu.data_in [24] ) );
MUX2_X1 _15154_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03182_ ), .Z(_07128_ ) );
NAND4_X1 _15155_ ( .A1(_07036_ ), .A2(_07038_ ), .A3(_07040_ ), .A4(_07128_ ), .ZN(_07129_ ) );
OAI21_X1 _15156_ ( .A(_07129_ ), .B1(_02361_ ), .B2(\io_master_rdata [23] ), .ZN(_07130_ ) );
NOR2_X1 _15157_ ( .A1(_07130_ ), .A2(_03167_ ), .ZN(\myifu.data_in [23] ) );
OR2_X1 _15158_ ( .A1(_03200_ ), .A2(\io_master_rdata [22] ), .ZN(_07131_ ) );
MUX2_X1 _15159_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03181_ ), .Z(_07132_ ) );
NAND4_X1 _15160_ ( .A1(_07035_ ), .A2(_07037_ ), .A3(_07039_ ), .A4(_07132_ ), .ZN(_07133_ ) );
AND3_X1 _15161_ ( .A1(_07131_ ), .A2(\io_master_arburst [0] ), .A3(_07133_ ), .ZN(\myifu.data_in [22] ) );
INV_X1 _15162_ ( .A(_03151_ ), .ZN(_07134_ ) );
OR2_X1 _15163_ ( .A1(_00210_ ), .A2(_07134_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
OR2_X1 _15164_ ( .A1(_00211_ ), .A2(_07134_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
OR2_X1 _15165_ ( .A1(_00212_ ), .A2(_07134_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND3_X1 _15166_ ( .A1(\IF_ID_pc [3] ), .A2(\IF_ID_pc [2] ), .A3(\myifu.myicache.valid_data_in ), .ZN(_07135_ ) );
NAND2_X1 _15167_ ( .A1(_07135_ ), .A2(_03151_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
INV_X1 _15168_ ( .A(_02676_ ), .ZN(_07136_ ) );
OAI21_X1 _15169_ ( .A(\IF_ID_inst [8] ), .B1(_02577_ ), .B2(_07136_ ), .ZN(_07137_ ) );
AOI21_X1 _15170_ ( .A(_02757_ ), .B1(_02408_ ), .B2(\IF_ID_inst [16] ), .ZN(_07138_ ) );
OAI211_X1 _15171_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B(_02566_ ), .C1(_02536_ ), .C2(_02555_ ), .ZN(_07139_ ) );
AND3_X1 _15172_ ( .A1(_02560_ ), .A2(_07139_ ), .A3(_02563_ ), .ZN(_07140_ ) );
NAND2_X1 _15173_ ( .A1(_07140_ ), .A2(_02711_ ), .ZN(_07141_ ) );
NOR4_X1 _15174_ ( .A1(_07141_ ), .A2(_02408_ ), .A3(_02636_ ), .A4(_02639_ ), .ZN(_07142_ ) );
NOR4_X1 _15175_ ( .A1(_02666_ ), .A2(_02702_ ), .A3(_02703_ ), .A4(_02470_ ), .ZN(_07143_ ) );
AND4_X1 _15176_ ( .A1(_02705_ ), .A2(_07019_ ), .A3(_02607_ ), .A4(_07143_ ), .ZN(_07144_ ) );
AND2_X1 _15177_ ( .A1(_07142_ ), .A2(_07144_ ), .ZN(_07145_ ) );
INV_X1 _15178_ ( .A(_02641_ ), .ZN(_07146_ ) );
NOR2_X1 _15179_ ( .A1(_07145_ ), .A2(_07146_ ), .ZN(_07147_ ) );
OAI211_X1 _15180_ ( .A(_07137_ ), .B(_07138_ ), .C1(_07147_ ), .C2(_02406_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
NOR2_X1 _15181_ ( .A1(_02640_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(_07148_ ) );
AND2_X1 _15182_ ( .A1(_02487_ ), .A2(\IF_ID_inst [31] ), .ZN(_07149_ ) );
AOI21_X1 _15183_ ( .A(_02401_ ), .B1(_07019_ ), .B2(_02705_ ), .ZN(_07150_ ) );
OR3_X1 _15184_ ( .A1(_07148_ ), .A2(_07149_ ), .A3(_07150_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
INV_X1 _15185_ ( .A(_07148_ ), .ZN(_07151_ ) );
OAI21_X1 _15186_ ( .A(\IF_ID_inst [31] ), .B1(_02577_ ), .B2(_07136_ ), .ZN(_07152_ ) );
AND2_X1 _15187_ ( .A1(_07151_ ), .A2(_07152_ ), .ZN(_07153_ ) );
BUF_X4 _15188_ ( .A(_07153_ ), .Z(_07154_ ) );
INV_X1 _15189_ ( .A(_07149_ ), .ZN(_07155_ ) );
BUF_X4 _15190_ ( .A(_07155_ ), .Z(_07156_ ) );
BUF_X4 _15191_ ( .A(_02705_ ), .Z(_07157_ ) );
OAI211_X1 _15192_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02405_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _15193_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02406_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _15194_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02409_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
OAI21_X1 _15195_ ( .A(\IF_ID_inst [19] ), .B1(_02487_ ), .B2(_02493_ ), .ZN(_07158_ ) );
BUF_X2 _15196_ ( .A(_02641_ ), .Z(_07159_ ) );
OAI211_X1 _15197_ ( .A(_07152_ ), .B(_07158_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI21_X1 _15198_ ( .A(\IF_ID_inst [18] ), .B1(_02487_ ), .B2(_02493_ ), .ZN(_07160_ ) );
OAI211_X1 _15199_ ( .A(_07152_ ), .B(_07160_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
NOR2_X1 _15200_ ( .A1(_02487_ ), .A2(_02493_ ), .ZN(_07161_ ) );
OAI221_X1 _15201_ ( .A(_07152_ ), .B1(_02595_ ), .B2(_07161_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI21_X1 _15202_ ( .A(\IF_ID_inst [16] ), .B1(_02487_ ), .B2(_02493_ ), .ZN(_07162_ ) );
OAI211_X1 _15203_ ( .A(_07152_ ), .B(_07162_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _15204_ ( .A(_07152_ ), .B1(_02624_ ), .B2(_07161_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _15205_ ( .A(_07152_ ), .B1(_02531_ ), .B2(_07161_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _15206_ ( .A(_07152_ ), .B1(_02392_ ), .B2(_07161_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _15207_ ( .A(_07152_ ), .B1(_02455_ ), .B2(_07161_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _15208_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02410_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
AOI21_X1 _15209_ ( .A(_02821_ ), .B1(_02577_ ), .B2(\IF_ID_inst [31] ), .ZN(_07163_ ) );
OAI221_X1 _15210_ ( .A(_07163_ ), .B1(_02473_ ), .B2(_02676_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
OAI221_X1 _15211_ ( .A(_02830_ ), .B1(_02405_ ), .B2(_07019_ ), .C1(_07159_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
OAI221_X1 _15212_ ( .A(_02834_ ), .B1(_02410_ ), .B2(_07019_ ), .C1(_02641_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
OAI221_X1 _15213_ ( .A(_02796_ ), .B1(_02411_ ), .B2(_07019_ ), .C1(_02641_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
OAI221_X1 _15214_ ( .A(_02790_ ), .B1(_02412_ ), .B2(_07019_ ), .C1(_02641_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
OAI221_X1 _15215_ ( .A(_02751_ ), .B1(_02413_ ), .B2(_07019_ ), .C1(_02641_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
OAI221_X1 _15216_ ( .A(_02781_ ), .B1(_02414_ ), .B2(_07019_ ), .C1(_02641_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _15217_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02411_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _15218_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02412_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _15219_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02413_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _15220_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02414_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _15221_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02415_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _15222_ ( .A(_07154_ ), .B(_07156_ ), .C1(_02416_ ), .C2(_07157_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _15223_ ( .A(_07153_ ), .B(_07155_ ), .C1(_02417_ ), .C2(_02705_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _15224_ ( .A(\IF_ID_inst [11] ), .B1(_02577_ ), .B2(_07136_ ), .ZN(_07164_ ) );
AOI21_X1 _15225_ ( .A(_02775_ ), .B1(_02408_ ), .B2(\IF_ID_inst [19] ), .ZN(_07165_ ) );
OAI211_X1 _15226_ ( .A(_07164_ ), .B(_07165_ ), .C1(_07147_ ), .C2(_02415_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _15227_ ( .A(\IF_ID_inst [10] ), .B1(_02577_ ), .B2(_07136_ ), .ZN(_07166_ ) );
AOI21_X1 _15228_ ( .A(_02768_ ), .B1(_02408_ ), .B2(\IF_ID_inst [18] ), .ZN(_07167_ ) );
OAI211_X1 _15229_ ( .A(_07166_ ), .B(_07167_ ), .C1(_07147_ ), .C2(_02416_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _15230_ ( .A(\IF_ID_inst [9] ), .B1(_02577_ ), .B2(_07136_ ), .ZN(_07168_ ) );
AND3_X1 _15231_ ( .A1(_02484_ ), .A2(\IF_ID_inst [22] ), .A3(_02466_ ), .ZN(_07169_ ) );
AOI221_X4 _15232_ ( .A(_07169_ ), .B1(\IF_ID_inst [17] ), .B2(_02408_ ), .C1(_07146_ ), .C2(\IF_ID_inst [22] ), .ZN(_07170_ ) );
INV_X1 _15233_ ( .A(_07145_ ), .ZN(_07171_ ) );
OAI211_X1 _15234_ ( .A(_07168_ ), .B(_07170_ ), .C1(_07171_ ), .C2(_02417_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OAI21_X1 _15235_ ( .A(\IF_ID_inst [7] ), .B1(_02459_ ), .B2(_02465_ ), .ZN(_07172_ ) );
OAI221_X1 _15236_ ( .A(_07172_ ), .B1(_02624_ ), .B2(_02400_ ), .C1(_07147_ ), .C2(_02409_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AOI21_X1 _15237_ ( .A(_01258_ ), .B1(_03220_ ), .B2(_03221_ ), .ZN(_07173_ ) );
INV_X1 _15238_ ( .A(_07173_ ), .ZN(_07174_ ) );
NOR2_X2 _15239_ ( .A1(_07174_ ), .A2(_03226_ ), .ZN(_07175_ ) );
INV_X1 _15240_ ( .A(_07175_ ), .ZN(_07176_ ) );
BUF_X4 _15241_ ( .A(_07176_ ), .Z(_07177_ ) );
AND3_X1 _15242_ ( .A1(_01248_ ), .A2(_01206_ ), .A3(_01276_ ), .ZN(_07178_ ) );
INV_X1 _15243_ ( .A(_03228_ ), .ZN(_07179_ ) );
NOR3_X1 _15244_ ( .A1(_07179_ ), .A2(\io_master_rid [1] ), .A3(_03229_ ), .ZN(_07180_ ) );
AND3_X1 _15245_ ( .A1(_01206_ ), .A2(io_master_rlast ), .A3(_07180_ ), .ZN(_07181_ ) );
NOR2_X1 _15246_ ( .A1(_07178_ ), .A2(_07181_ ), .ZN(_07182_ ) );
INV_X1 _15247_ ( .A(_07182_ ), .ZN(_07183_ ) );
INV_X1 _15248_ ( .A(_07180_ ), .ZN(_07184_ ) );
NOR4_X4 _15249_ ( .A1(_02361_ ), .A2(io_master_rlast ), .A3(_01258_ ), .A4(_07184_ ), .ZN(_07185_ ) );
OAI21_X2 _15250_ ( .A(_02498_ ), .B1(_07183_ ), .B2(_07185_ ), .ZN(_07186_ ) );
BUF_X4 _15251_ ( .A(_07186_ ), .Z(_07187_ ) );
BUF_X4 _15252_ ( .A(_07187_ ), .Z(_07188_ ) );
OAI21_X1 _15253_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07189_ ) );
NOR2_X2 _15254_ ( .A1(_07176_ ), .A2(_07186_ ), .ZN(_07190_ ) );
INV_X1 _15255_ ( .A(_07190_ ), .ZN(_07191_ ) );
BUF_X4 _15256_ ( .A(_07191_ ), .Z(_07192_ ) );
OAI211_X1 _15257_ ( .A(fanout_net_41 ), .B(_07189_ ), .C1(_07192_ ), .C2(\myifu.data_in [8] ), .ZN(_07193_ ) );
MUX2_X1 _15258_ ( .A(\myifu.myicache.data[0][8] ), .B(\myifu.myicache.data[1][8] ), .S(fanout_net_36 ), .Z(_07194_ ) );
MUX2_X1 _15259_ ( .A(\myifu.myicache.data[2][8] ), .B(\myifu.myicache.data[3][8] ), .S(fanout_net_37 ), .Z(_07195_ ) );
MUX2_X1 _15260_ ( .A(_07194_ ), .B(_07195_ ), .S(fanout_net_40 ), .Z(_07196_ ) );
NOR2_X1 _15261_ ( .A1(\myifu.state [1] ), .A2(fanout_net_41 ), .ZN(_07197_ ) );
BUF_X4 _15262_ ( .A(_07197_ ), .Z(_07198_ ) );
NAND2_X1 _15263_ ( .A1(_07196_ ), .A2(_07198_ ), .ZN(_07199_ ) );
NAND2_X1 _15264_ ( .A1(_07193_ ), .A2(_07199_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
OR4_X1 _15265_ ( .A1(_03226_ ), .A2(_07174_ ), .A3(_07186_ ), .A4(\myifu.data_in [31] ), .ZN(_07200_ ) );
OAI211_X1 _15266_ ( .A(_07200_ ), .B(fanout_net_41 ), .C1(_07190_ ), .C2(_02539_ ), .ZN(_07201_ ) );
MUX2_X1 _15267_ ( .A(\myifu.myicache.data[0][31] ), .B(\myifu.myicache.data[1][31] ), .S(fanout_net_37 ), .Z(_07202_ ) );
MUX2_X1 _15268_ ( .A(\myifu.myicache.data[2][31] ), .B(\myifu.myicache.data[3][31] ), .S(fanout_net_37 ), .Z(_07203_ ) );
MUX2_X1 _15269_ ( .A(_07202_ ), .B(_07203_ ), .S(fanout_net_40 ), .Z(_07204_ ) );
NAND2_X1 _15270_ ( .A1(_07204_ ), .A2(_07198_ ), .ZN(_07205_ ) );
NAND2_X1 _15271_ ( .A1(_07201_ ), .A2(_07205_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
BUF_X4 _15272_ ( .A(_07176_ ), .Z(_07206_ ) );
BUF_X4 _15273_ ( .A(_07206_ ), .Z(_07207_ ) );
BUF_X4 _15274_ ( .A(_07186_ ), .Z(_07208_ ) );
BUF_X4 _15275_ ( .A(_07208_ ), .Z(_07209_ ) );
OAI21_X1 _15276_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07210_ ) );
CLKBUF_X2 _15277_ ( .A(_03226_ ), .Z(_07211_ ) );
CLKBUF_X2 _15278_ ( .A(_07174_ ), .Z(_07212_ ) );
OR4_X1 _15279_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [30] ), .ZN(_07213_ ) );
NAND3_X1 _15280_ ( .A1(_07210_ ), .A2(_07213_ ), .A3(fanout_net_41 ), .ZN(_07214_ ) );
MUX2_X1 _15281_ ( .A(\myifu.myicache.data[0][30] ), .B(\myifu.myicache.data[1][30] ), .S(fanout_net_37 ), .Z(_07215_ ) );
MUX2_X1 _15282_ ( .A(\myifu.myicache.data[2][30] ), .B(\myifu.myicache.data[3][30] ), .S(fanout_net_37 ), .Z(_07216_ ) );
MUX2_X1 _15283_ ( .A(_07215_ ), .B(_07216_ ), .S(fanout_net_40 ), .Z(_07217_ ) );
NAND2_X1 _15284_ ( .A1(_07217_ ), .A2(_07198_ ), .ZN(_07218_ ) );
NAND2_X1 _15285_ ( .A1(_07214_ ), .A2(_07218_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
OAI21_X1 _15286_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07219_ ) );
OR4_X1 _15287_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [21] ), .ZN(_07220_ ) );
NAND3_X1 _15288_ ( .A1(_07219_ ), .A2(_07220_ ), .A3(fanout_net_41 ), .ZN(_07221_ ) );
MUX2_X1 _15289_ ( .A(\myifu.myicache.data[0][21] ), .B(\myifu.myicache.data[1][21] ), .S(fanout_net_37 ), .Z(_07222_ ) );
MUX2_X1 _15290_ ( .A(\myifu.myicache.data[2][21] ), .B(\myifu.myicache.data[3][21] ), .S(fanout_net_37 ), .Z(_07223_ ) );
MUX2_X1 _15291_ ( .A(_07222_ ), .B(_07223_ ), .S(fanout_net_40 ), .Z(_07224_ ) );
NAND2_X1 _15292_ ( .A1(_07224_ ), .A2(_07198_ ), .ZN(_07225_ ) );
NAND2_X1 _15293_ ( .A1(_07221_ ), .A2(_07225_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
OAI21_X1 _15294_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07226_ ) );
OAI211_X1 _15295_ ( .A(fanout_net_41 ), .B(_07226_ ), .C1(_07192_ ), .C2(\myifu.data_in [20] ), .ZN(_07227_ ) );
MUX2_X1 _15296_ ( .A(\myifu.myicache.data[0][20] ), .B(\myifu.myicache.data[1][20] ), .S(fanout_net_37 ), .Z(_07228_ ) );
MUX2_X1 _15297_ ( .A(\myifu.myicache.data[2][20] ), .B(\myifu.myicache.data[3][20] ), .S(fanout_net_37 ), .Z(_07229_ ) );
MUX2_X1 _15298_ ( .A(_07228_ ), .B(_07229_ ), .S(fanout_net_40 ), .Z(_07230_ ) );
NAND2_X1 _15299_ ( .A1(_07230_ ), .A2(_07198_ ), .ZN(_07231_ ) );
NAND2_X1 _15300_ ( .A1(_07227_ ), .A2(_07231_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
OAI21_X1 _15301_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07232_ ) );
OR4_X1 _15302_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [19] ), .ZN(_07233_ ) );
NAND3_X1 _15303_ ( .A1(_07232_ ), .A2(_07233_ ), .A3(fanout_net_41 ), .ZN(_07234_ ) );
MUX2_X1 _15304_ ( .A(\myifu.myicache.data[0][19] ), .B(\myifu.myicache.data[1][19] ), .S(fanout_net_37 ), .Z(_07235_ ) );
MUX2_X1 _15305_ ( .A(\myifu.myicache.data[2][19] ), .B(\myifu.myicache.data[3][19] ), .S(fanout_net_37 ), .Z(_07236_ ) );
MUX2_X1 _15306_ ( .A(_07235_ ), .B(_07236_ ), .S(fanout_net_40 ), .Z(_07237_ ) );
NAND2_X1 _15307_ ( .A1(_07237_ ), .A2(_07198_ ), .ZN(_07238_ ) );
NAND2_X1 _15308_ ( .A1(_07234_ ), .A2(_07238_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
OAI21_X1 _15309_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07239_ ) );
OAI211_X1 _15310_ ( .A(fanout_net_41 ), .B(_07239_ ), .C1(_07192_ ), .C2(\myifu.data_in [18] ), .ZN(_07240_ ) );
MUX2_X1 _15311_ ( .A(\myifu.myicache.data[0][18] ), .B(\myifu.myicache.data[1][18] ), .S(fanout_net_37 ), .Z(_07241_ ) );
MUX2_X1 _15312_ ( .A(\myifu.myicache.data[2][18] ), .B(\myifu.myicache.data[3][18] ), .S(fanout_net_37 ), .Z(_07242_ ) );
MUX2_X1 _15313_ ( .A(_07241_ ), .B(_07242_ ), .S(fanout_net_40 ), .Z(_07243_ ) );
NAND2_X1 _15314_ ( .A1(_07243_ ), .A2(_07198_ ), .ZN(_07244_ ) );
NAND2_X1 _15315_ ( .A1(_07240_ ), .A2(_07244_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
OAI21_X1 _15316_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07245_ ) );
OAI211_X1 _15317_ ( .A(fanout_net_41 ), .B(_07245_ ), .C1(_07192_ ), .C2(\myifu.data_in [17] ), .ZN(_07246_ ) );
MUX2_X1 _15318_ ( .A(\myifu.myicache.data[0][17] ), .B(\myifu.myicache.data[1][17] ), .S(fanout_net_37 ), .Z(_07247_ ) );
MUX2_X1 _15319_ ( .A(\myifu.myicache.data[2][17] ), .B(\myifu.myicache.data[3][17] ), .S(fanout_net_37 ), .Z(_07248_ ) );
MUX2_X1 _15320_ ( .A(_07247_ ), .B(_07248_ ), .S(fanout_net_40 ), .Z(_07249_ ) );
NAND2_X1 _15321_ ( .A1(_07249_ ), .A2(_07198_ ), .ZN(_07250_ ) );
NAND2_X1 _15322_ ( .A1(_07246_ ), .A2(_07250_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
OAI21_X1 _15323_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07251_ ) );
OAI211_X1 _15324_ ( .A(fanout_net_41 ), .B(_07251_ ), .C1(_07192_ ), .C2(\myifu.data_in [16] ), .ZN(_07252_ ) );
MUX2_X1 _15325_ ( .A(\myifu.myicache.data[0][16] ), .B(\myifu.myicache.data[1][16] ), .S(fanout_net_37 ), .Z(_07253_ ) );
MUX2_X1 _15326_ ( .A(\myifu.myicache.data[2][16] ), .B(\myifu.myicache.data[3][16] ), .S(fanout_net_37 ), .Z(_07254_ ) );
MUX2_X1 _15327_ ( .A(_07253_ ), .B(_07254_ ), .S(fanout_net_40 ), .Z(_07255_ ) );
NAND2_X1 _15328_ ( .A1(_07255_ ), .A2(_07198_ ), .ZN(_07256_ ) );
NAND2_X1 _15329_ ( .A1(_07252_ ), .A2(_07256_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
OAI21_X1 _15330_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07257_ ) );
OAI211_X1 _15331_ ( .A(fanout_net_41 ), .B(_07257_ ), .C1(_07192_ ), .C2(\myifu.data_in [15] ), .ZN(_07258_ ) );
MUX2_X1 _15332_ ( .A(\myifu.myicache.data[0][15] ), .B(\myifu.myicache.data[1][15] ), .S(fanout_net_37 ), .Z(_07259_ ) );
MUX2_X1 _15333_ ( .A(\myifu.myicache.data[2][15] ), .B(\myifu.myicache.data[3][15] ), .S(fanout_net_37 ), .Z(_07260_ ) );
MUX2_X1 _15334_ ( .A(_07259_ ), .B(_07260_ ), .S(fanout_net_40 ), .Z(_07261_ ) );
NAND2_X1 _15335_ ( .A1(_07261_ ), .A2(_07198_ ), .ZN(_07262_ ) );
NAND2_X1 _15336_ ( .A1(_07258_ ), .A2(_07262_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
OAI21_X1 _15337_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07263_ ) );
OR4_X1 _15338_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [14] ), .ZN(_07264_ ) );
NAND3_X1 _15339_ ( .A1(_07263_ ), .A2(_07264_ ), .A3(fanout_net_41 ), .ZN(_07265_ ) );
MUX2_X1 _15340_ ( .A(\myifu.myicache.data[0][14] ), .B(\myifu.myicache.data[1][14] ), .S(fanout_net_37 ), .Z(_07266_ ) );
MUX2_X1 _15341_ ( .A(\myifu.myicache.data[2][14] ), .B(\myifu.myicache.data[3][14] ), .S(fanout_net_37 ), .Z(_07267_ ) );
MUX2_X1 _15342_ ( .A(_07266_ ), .B(_07267_ ), .S(fanout_net_40 ), .Z(_07268_ ) );
BUF_X4 _15343_ ( .A(_07197_ ), .Z(_07269_ ) );
NAND2_X1 _15344_ ( .A1(_07268_ ), .A2(_07269_ ), .ZN(_07270_ ) );
NAND2_X1 _15345_ ( .A1(_07265_ ), .A2(_07270_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
OAI21_X1 _15346_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07271_ ) );
OAI211_X1 _15347_ ( .A(fanout_net_41 ), .B(_07271_ ), .C1(_07192_ ), .C2(\myifu.data_in [13] ), .ZN(_07272_ ) );
MUX2_X1 _15348_ ( .A(\myifu.myicache.data[0][13] ), .B(\myifu.myicache.data[1][13] ), .S(fanout_net_37 ), .Z(_07273_ ) );
MUX2_X1 _15349_ ( .A(\myifu.myicache.data[2][13] ), .B(\myifu.myicache.data[3][13] ), .S(fanout_net_37 ), .Z(_07274_ ) );
MUX2_X1 _15350_ ( .A(_07273_ ), .B(_07274_ ), .S(fanout_net_40 ), .Z(_07275_ ) );
NAND2_X1 _15351_ ( .A1(_07275_ ), .A2(_07269_ ), .ZN(_07276_ ) );
NAND2_X1 _15352_ ( .A1(_07272_ ), .A2(_07276_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
OAI21_X1 _15353_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07277_ ) );
OR4_X1 _15354_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [12] ), .ZN(_07278_ ) );
NAND3_X1 _15355_ ( .A1(_07277_ ), .A2(_07278_ ), .A3(fanout_net_41 ), .ZN(_07279_ ) );
MUX2_X1 _15356_ ( .A(\myifu.myicache.data[0][12] ), .B(\myifu.myicache.data[1][12] ), .S(fanout_net_37 ), .Z(_07280_ ) );
MUX2_X1 _15357_ ( .A(\myifu.myicache.data[2][12] ), .B(\myifu.myicache.data[3][12] ), .S(fanout_net_37 ), .Z(_07281_ ) );
MUX2_X1 _15358_ ( .A(_07280_ ), .B(_07281_ ), .S(fanout_net_40 ), .Z(_07282_ ) );
NAND2_X1 _15359_ ( .A1(_07282_ ), .A2(_07269_ ), .ZN(_07283_ ) );
NAND2_X1 _15360_ ( .A1(_07279_ ), .A2(_07283_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
OAI21_X1 _15361_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07284_ ) );
OR4_X1 _15362_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [29] ), .ZN(_07285_ ) );
NAND3_X1 _15363_ ( .A1(_07284_ ), .A2(_07285_ ), .A3(fanout_net_41 ), .ZN(_07286_ ) );
MUX2_X1 _15364_ ( .A(\myifu.myicache.data[0][29] ), .B(\myifu.myicache.data[1][29] ), .S(fanout_net_37 ), .Z(_07287_ ) );
MUX2_X1 _15365_ ( .A(\myifu.myicache.data[2][29] ), .B(\myifu.myicache.data[3][29] ), .S(fanout_net_37 ), .Z(_07288_ ) );
MUX2_X1 _15366_ ( .A(_07287_ ), .B(_07288_ ), .S(fanout_net_40 ), .Z(_07289_ ) );
NAND2_X1 _15367_ ( .A1(_07289_ ), .A2(_07269_ ), .ZN(_07290_ ) );
NAND2_X1 _15368_ ( .A1(_07286_ ), .A2(_07290_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
OR4_X1 _15369_ ( .A1(_03226_ ), .A2(_07174_ ), .A3(_07186_ ), .A4(\myifu.data_in [11] ), .ZN(_07291_ ) );
OAI211_X1 _15370_ ( .A(_07291_ ), .B(fanout_net_41 ), .C1(_07190_ ), .C2(_02776_ ), .ZN(_07292_ ) );
MUX2_X1 _15371_ ( .A(\myifu.myicache.data[0][11] ), .B(\myifu.myicache.data[1][11] ), .S(fanout_net_37 ), .Z(_07293_ ) );
MUX2_X1 _15372_ ( .A(\myifu.myicache.data[2][11] ), .B(\myifu.myicache.data[3][11] ), .S(fanout_net_37 ), .Z(_07294_ ) );
MUX2_X1 _15373_ ( .A(_07293_ ), .B(_07294_ ), .S(fanout_net_40 ), .Z(_07295_ ) );
NAND2_X1 _15374_ ( .A1(_07295_ ), .A2(_07269_ ), .ZN(_07296_ ) );
NAND2_X1 _15375_ ( .A1(_07292_ ), .A2(_07296_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
OR4_X1 _15376_ ( .A1(_03226_ ), .A2(_07174_ ), .A3(_07186_ ), .A4(\myifu.data_in [10] ), .ZN(_07297_ ) );
OAI211_X1 _15377_ ( .A(_07297_ ), .B(fanout_net_41 ), .C1(_07190_ ), .C2(_02769_ ), .ZN(_07298_ ) );
MUX2_X1 _15378_ ( .A(\myifu.myicache.data[0][10] ), .B(\myifu.myicache.data[1][10] ), .S(fanout_net_37 ), .Z(_07299_ ) );
MUX2_X1 _15379_ ( .A(\myifu.myicache.data[2][10] ), .B(\myifu.myicache.data[3][10] ), .S(fanout_net_38 ), .Z(_07300_ ) );
MUX2_X1 _15380_ ( .A(_07299_ ), .B(_07300_ ), .S(fanout_net_40 ), .Z(_07301_ ) );
NAND2_X1 _15381_ ( .A1(_07301_ ), .A2(_07269_ ), .ZN(_07302_ ) );
NAND2_X1 _15382_ ( .A1(_07298_ ), .A2(_07302_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
OAI21_X1 _15383_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_07303_ ) );
OAI211_X1 _15384_ ( .A(fanout_net_41 ), .B(_07303_ ), .C1(_07192_ ), .C2(\myifu.data_in [9] ), .ZN(_07304_ ) );
MUX2_X1 _15385_ ( .A(\myifu.myicache.data[0][9] ), .B(\myifu.myicache.data[1][9] ), .S(fanout_net_38 ), .Z(_07305_ ) );
MUX2_X1 _15386_ ( .A(\myifu.myicache.data[2][9] ), .B(\myifu.myicache.data[3][9] ), .S(fanout_net_38 ), .Z(_07306_ ) );
MUX2_X1 _15387_ ( .A(_07305_ ), .B(_07306_ ), .S(fanout_net_40 ), .Z(_07307_ ) );
NAND2_X1 _15388_ ( .A1(_07307_ ), .A2(_07269_ ), .ZN(_07308_ ) );
NAND2_X1 _15389_ ( .A1(_07304_ ), .A2(_07308_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
OAI21_X1 _15390_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07309_ ) );
OR4_X1 _15391_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [7] ), .ZN(_07310_ ) );
NAND3_X1 _15392_ ( .A1(_07309_ ), .A2(_07310_ ), .A3(fanout_net_41 ), .ZN(_07311_ ) );
MUX2_X1 _15393_ ( .A(\myifu.myicache.data[0][7] ), .B(\myifu.myicache.data[1][7] ), .S(fanout_net_38 ), .Z(_07312_ ) );
MUX2_X1 _15394_ ( .A(\myifu.myicache.data[2][7] ), .B(\myifu.myicache.data[3][7] ), .S(fanout_net_38 ), .Z(_07313_ ) );
MUX2_X1 _15395_ ( .A(_07312_ ), .B(_07313_ ), .S(fanout_net_40 ), .Z(_07314_ ) );
NAND2_X1 _15396_ ( .A1(_07314_ ), .A2(_07269_ ), .ZN(_07315_ ) );
NAND2_X1 _15397_ ( .A1(_07311_ ), .A2(_07315_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
OAI21_X1 _15398_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_07316_ ) );
OR4_X1 _15399_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [6] ), .ZN(_07317_ ) );
NAND3_X1 _15400_ ( .A1(_07316_ ), .A2(_07317_ ), .A3(fanout_net_41 ), .ZN(_07318_ ) );
MUX2_X1 _15401_ ( .A(\myifu.myicache.data[0][6] ), .B(\myifu.myicache.data[1][6] ), .S(fanout_net_38 ), .Z(_07319_ ) );
MUX2_X1 _15402_ ( .A(\myifu.myicache.data[2][6] ), .B(\myifu.myicache.data[3][6] ), .S(fanout_net_38 ), .Z(_07320_ ) );
MUX2_X1 _15403_ ( .A(_07319_ ), .B(_07320_ ), .S(fanout_net_40 ), .Z(_07321_ ) );
NAND2_X1 _15404_ ( .A1(_07321_ ), .A2(_07269_ ), .ZN(_07322_ ) );
NAND2_X1 _15405_ ( .A1(_07318_ ), .A2(_07322_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
OAI21_X1 _15406_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_07323_ ) );
OAI211_X1 _15407_ ( .A(fanout_net_41 ), .B(_07323_ ), .C1(_07192_ ), .C2(\myifu.data_in [5] ), .ZN(_07324_ ) );
MUX2_X1 _15408_ ( .A(\myifu.myicache.data[0][5] ), .B(\myifu.myicache.data[1][5] ), .S(fanout_net_38 ), .Z(_07325_ ) );
MUX2_X1 _15409_ ( .A(\myifu.myicache.data[2][5] ), .B(\myifu.myicache.data[3][5] ), .S(fanout_net_38 ), .Z(_07326_ ) );
MUX2_X1 _15410_ ( .A(_07325_ ), .B(_07326_ ), .S(fanout_net_40 ), .Z(_07327_ ) );
NAND2_X1 _15411_ ( .A1(_07327_ ), .A2(_07269_ ), .ZN(_07328_ ) );
NAND2_X1 _15412_ ( .A1(_07324_ ), .A2(_07328_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
OAI21_X1 _15413_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_00271_ ) );
OR4_X1 _15414_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07187_ ), .A4(\myifu.data_in [4] ), .ZN(_00272_ ) );
NAND3_X1 _15415_ ( .A1(_00271_ ), .A2(_00272_ ), .A3(fanout_net_41 ), .ZN(_00273_ ) );
MUX2_X1 _15416_ ( .A(\myifu.myicache.data[0][4] ), .B(\myifu.myicache.data[1][4] ), .S(fanout_net_38 ), .Z(_00274_ ) );
MUX2_X1 _15417_ ( .A(\myifu.myicache.data[2][4] ), .B(\myifu.myicache.data[3][4] ), .S(fanout_net_38 ), .Z(_00275_ ) );
MUX2_X1 _15418_ ( .A(_00274_ ), .B(_00275_ ), .S(fanout_net_40 ), .Z(_00276_ ) );
BUF_X4 _15419_ ( .A(_07197_ ), .Z(_00277_ ) );
NAND2_X1 _15420_ ( .A1(_00276_ ), .A2(_00277_ ), .ZN(_00278_ ) );
NAND2_X1 _15421_ ( .A1(_00273_ ), .A2(_00278_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
OAI21_X1 _15422_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00279_ ) );
OAI211_X1 _15423_ ( .A(fanout_net_41 ), .B(_00279_ ), .C1(_07192_ ), .C2(\myifu.data_in [3] ), .ZN(_00280_ ) );
MUX2_X1 _15424_ ( .A(\myifu.myicache.data[0][3] ), .B(\myifu.myicache.data[1][3] ), .S(fanout_net_38 ), .Z(_00281_ ) );
MUX2_X1 _15425_ ( .A(\myifu.myicache.data[2][3] ), .B(\myifu.myicache.data[3][3] ), .S(fanout_net_38 ), .Z(_00282_ ) );
MUX2_X1 _15426_ ( .A(_00281_ ), .B(_00282_ ), .S(fanout_net_40 ), .Z(_00283_ ) );
NAND2_X1 _15427_ ( .A1(_00283_ ), .A2(_00277_ ), .ZN(_00284_ ) );
NAND2_X1 _15428_ ( .A1(_00280_ ), .A2(_00284_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
OAI21_X1 _15429_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00285_ ) );
OAI211_X1 _15430_ ( .A(fanout_net_41 ), .B(_00285_ ), .C1(_07191_ ), .C2(\myifu.data_in [2] ), .ZN(_00286_ ) );
MUX2_X1 _15431_ ( .A(\myifu.myicache.data[0][2] ), .B(\myifu.myicache.data[1][2] ), .S(fanout_net_38 ), .Z(_00287_ ) );
MUX2_X1 _15432_ ( .A(\myifu.myicache.data[2][2] ), .B(\myifu.myicache.data[3][2] ), .S(fanout_net_38 ), .Z(_00288_ ) );
MUX2_X1 _15433_ ( .A(_00287_ ), .B(_00288_ ), .S(fanout_net_40 ), .Z(_00289_ ) );
NAND2_X1 _15434_ ( .A1(_00289_ ), .A2(_00277_ ), .ZN(_00290_ ) );
NAND2_X1 _15435_ ( .A1(_00286_ ), .A2(_00290_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
OAI21_X1 _15436_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07207_ ), .B2(_07209_ ), .ZN(_00291_ ) );
OR4_X1 _15437_ ( .A1(_07211_ ), .A2(_07212_ ), .A3(_07186_ ), .A4(\myifu.data_in [1] ), .ZN(_00292_ ) );
NAND3_X1 _15438_ ( .A1(_00291_ ), .A2(_00292_ ), .A3(fanout_net_41 ), .ZN(_00293_ ) );
MUX2_X1 _15439_ ( .A(\myifu.myicache.data[0][1] ), .B(\myifu.myicache.data[1][1] ), .S(fanout_net_38 ), .Z(_00294_ ) );
MUX2_X1 _15440_ ( .A(\myifu.myicache.data[2][1] ), .B(\myifu.myicache.data[3][1] ), .S(fanout_net_38 ), .Z(_00295_ ) );
MUX2_X1 _15441_ ( .A(_00294_ ), .B(_00295_ ), .S(fanout_net_40 ), .Z(_00296_ ) );
NAND2_X1 _15442_ ( .A1(_00296_ ), .A2(_00277_ ), .ZN(_00297_ ) );
NAND2_X1 _15443_ ( .A1(_00293_ ), .A2(_00297_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
OAI21_X1 _15444_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_00298_ ) );
OR4_X1 _15445_ ( .A1(_03226_ ), .A2(_07174_ ), .A3(_07186_ ), .A4(\myifu.data_in [28] ), .ZN(_00299_ ) );
NAND3_X1 _15446_ ( .A1(_00298_ ), .A2(_00299_ ), .A3(fanout_net_41 ), .ZN(_00300_ ) );
MUX2_X1 _15447_ ( .A(\myifu.myicache.data[0][28] ), .B(\myifu.myicache.data[1][28] ), .S(fanout_net_38 ), .Z(_00301_ ) );
MUX2_X1 _15448_ ( .A(\myifu.myicache.data[2][28] ), .B(\myifu.myicache.data[3][28] ), .S(fanout_net_38 ), .Z(_00302_ ) );
MUX2_X1 _15449_ ( .A(_00301_ ), .B(_00302_ ), .S(fanout_net_40 ), .Z(_00303_ ) );
NAND2_X1 _15450_ ( .A1(_00303_ ), .A2(_00277_ ), .ZN(_00304_ ) );
NAND2_X1 _15451_ ( .A1(_00300_ ), .A2(_00304_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
OAI21_X1 _15452_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00305_ ) );
OAI211_X1 _15453_ ( .A(fanout_net_41 ), .B(_00305_ ), .C1(_07191_ ), .C2(\myifu.data_in [0] ), .ZN(_00306_ ) );
MUX2_X1 _15454_ ( .A(\myifu.myicache.data[0][0] ), .B(\myifu.myicache.data[1][0] ), .S(fanout_net_38 ), .Z(_00307_ ) );
MUX2_X1 _15455_ ( .A(\myifu.myicache.data[2][0] ), .B(\myifu.myicache.data[3][0] ), .S(fanout_net_38 ), .Z(_00308_ ) );
MUX2_X1 _15456_ ( .A(_00307_ ), .B(_00308_ ), .S(fanout_net_40 ), .Z(_00309_ ) );
NAND2_X1 _15457_ ( .A1(_00309_ ), .A2(_00277_ ), .ZN(_00310_ ) );
NAND2_X1 _15458_ ( .A1(_00306_ ), .A2(_00310_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
OAI21_X1 _15459_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00311_ ) );
OAI211_X1 _15460_ ( .A(fanout_net_41 ), .B(_00311_ ), .C1(_07191_ ), .C2(\myifu.data_in [27] ), .ZN(_00312_ ) );
MUX2_X1 _15461_ ( .A(\myifu.myicache.data[0][27] ), .B(\myifu.myicache.data[1][27] ), .S(fanout_net_38 ), .Z(_00313_ ) );
MUX2_X1 _15462_ ( .A(\myifu.myicache.data[2][27] ), .B(\myifu.myicache.data[3][27] ), .S(fanout_net_38 ), .Z(_00314_ ) );
MUX2_X1 _15463_ ( .A(_00313_ ), .B(_00314_ ), .S(fanout_net_40 ), .Z(_00315_ ) );
NAND2_X1 _15464_ ( .A1(_00315_ ), .A2(_00277_ ), .ZN(_00316_ ) );
NAND2_X1 _15465_ ( .A1(_00312_ ), .A2(_00316_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
OAI21_X1 _15466_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B1(_07177_ ), .B2(_07188_ ), .ZN(_00317_ ) );
OR4_X1 _15467_ ( .A1(_03226_ ), .A2(_07174_ ), .A3(_07186_ ), .A4(\myifu.data_in [26] ), .ZN(_00318_ ) );
NAND3_X1 _15468_ ( .A1(_00317_ ), .A2(_00318_ ), .A3(fanout_net_41 ), .ZN(_00319_ ) );
MUX2_X1 _15469_ ( .A(\myifu.myicache.data[0][26] ), .B(\myifu.myicache.data[1][26] ), .S(fanout_net_38 ), .Z(_00320_ ) );
MUX2_X1 _15470_ ( .A(\myifu.myicache.data[2][26] ), .B(\myifu.myicache.data[3][26] ), .S(fanout_net_38 ), .Z(_00321_ ) );
MUX2_X1 _15471_ ( .A(_00320_ ), .B(_00321_ ), .S(fanout_net_40 ), .Z(_00322_ ) );
NAND2_X1 _15472_ ( .A1(_00322_ ), .A2(_00277_ ), .ZN(_00323_ ) );
NAND2_X1 _15473_ ( .A1(_00319_ ), .A2(_00323_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
OAI21_X1 _15474_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00324_ ) );
OAI211_X1 _15475_ ( .A(\myifu.state [2] ), .B(_00324_ ), .C1(_07191_ ), .C2(\myifu.data_in [25] ), .ZN(_00325_ ) );
MUX2_X1 _15476_ ( .A(\myifu.myicache.data[0][25] ), .B(\myifu.myicache.data[1][25] ), .S(fanout_net_38 ), .Z(_00326_ ) );
MUX2_X1 _15477_ ( .A(\myifu.myicache.data[2][25] ), .B(\myifu.myicache.data[3][25] ), .S(fanout_net_38 ), .Z(_00327_ ) );
MUX2_X1 _15478_ ( .A(_00326_ ), .B(_00327_ ), .S(fanout_net_40 ), .Z(_00328_ ) );
NAND2_X1 _15479_ ( .A1(_00328_ ), .A2(_00277_ ), .ZN(_00329_ ) );
NAND2_X1 _15480_ ( .A1(_00325_ ), .A2(_00329_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
OAI21_X1 _15481_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00330_ ) );
OAI211_X1 _15482_ ( .A(\myifu.state [2] ), .B(_00330_ ), .C1(_07191_ ), .C2(\myifu.data_in [24] ), .ZN(_00331_ ) );
MUX2_X1 _15483_ ( .A(\myifu.myicache.data[0][24] ), .B(\myifu.myicache.data[1][24] ), .S(fanout_net_38 ), .Z(_00332_ ) );
MUX2_X1 _15484_ ( .A(\myifu.myicache.data[2][24] ), .B(\myifu.myicache.data[3][24] ), .S(fanout_net_38 ), .Z(_00333_ ) );
MUX2_X1 _15485_ ( .A(_00332_ ), .B(_00333_ ), .S(fanout_net_40 ), .Z(_00334_ ) );
NAND2_X1 _15486_ ( .A1(_00334_ ), .A2(_00277_ ), .ZN(_00335_ ) );
NAND2_X1 _15487_ ( .A1(_00331_ ), .A2(_00335_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
OAI21_X1 _15488_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00336_ ) );
OAI211_X1 _15489_ ( .A(\myifu.state [2] ), .B(_00336_ ), .C1(_07191_ ), .C2(\myifu.data_in [23] ), .ZN(_00337_ ) );
MUX2_X1 _15490_ ( .A(\myifu.myicache.data[0][23] ), .B(\myifu.myicache.data[1][23] ), .S(fanout_net_38 ), .Z(_00338_ ) );
MUX2_X1 _15491_ ( .A(\myifu.myicache.data[2][23] ), .B(\myifu.myicache.data[3][23] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_00339_ ) );
MUX2_X1 _15492_ ( .A(_00338_ ), .B(_00339_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_00340_ ) );
NAND2_X1 _15493_ ( .A1(_00340_ ), .A2(_07197_ ), .ZN(_00341_ ) );
NAND2_X1 _15494_ ( .A1(_00337_ ), .A2(_00341_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
OAI21_X1 _15495_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .B1(_07206_ ), .B2(_07208_ ), .ZN(_00342_ ) );
OAI211_X1 _15496_ ( .A(\myifu.state [2] ), .B(_00342_ ), .C1(_07191_ ), .C2(\myifu.data_in [22] ), .ZN(_00343_ ) );
MUX2_X1 _15497_ ( .A(\myifu.myicache.data[0][22] ), .B(\myifu.myicache.data[1][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_00344_ ) );
MUX2_X1 _15498_ ( .A(\myifu.myicache.data[2][22] ), .B(\myifu.myicache.data[3][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_00345_ ) );
MUX2_X1 _15499_ ( .A(_00344_ ), .B(_00345_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_00346_ ) );
NAND2_X1 _15500_ ( .A1(_00346_ ), .A2(_07197_ ), .ZN(_00347_ ) );
NAND2_X1 _15501_ ( .A1(_00343_ ), .A2(_00347_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
NOR3_X1 _15502_ ( .A1(_02741_ ), .A2(_07006_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_30_E_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_E ) );
AND3_X1 _15503_ ( .A1(_07175_ ), .A2(\myifu.state [2] ), .A3(_07183_ ), .ZN(_00348_ ) );
OAI21_X1 _15504_ ( .A(_00841_ ), .B1(_00348_ ), .B2(_07026_ ), .ZN(_00349_ ) );
NAND4_X1 _15505_ ( .A1(_01122_ ), .A2(_01199_ ), .A3(\myifu.state [0] ), .A4(_03151_ ), .ZN(_00350_ ) );
NAND2_X1 _15506_ ( .A1(_00349_ ), .A2(_00350_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
AOI21_X1 _15507_ ( .A(fanout_net_4 ), .B1(IDU_ready_IFU ), .B2(\myifu.state [1] ), .ZN(_00351_ ) );
AND2_X1 _15508_ ( .A1(_02362_ ), .A2(_01314_ ), .ZN(_00352_ ) );
OAI211_X1 _15509_ ( .A(_00351_ ), .B(_07029_ ), .C1(_00352_ ), .C2(_01316_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
AND2_X1 _15510_ ( .A1(_07175_ ), .A2(_07183_ ), .ZN(_00353_ ) );
INV_X1 _15511_ ( .A(_00353_ ), .ZN(_00354_ ) );
AOI22_X1 _15512_ ( .A1(_00354_ ), .A2(\myifu.state [2] ), .B1(_01315_ ), .B2(_00352_ ), .ZN(_00355_ ) );
NOR2_X1 _15513_ ( .A1(_00355_ ), .A2(fanout_net_4 ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND4_X1 _15514_ ( .A1(_02502_ ), .A2(_03151_ ), .A3(\IF_ID_pc [2] ), .A4(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND4_X1 _15515_ ( .A1(\IF_ID_pc [3] ), .A2(_03151_ ), .A3(_02503_ ), .A4(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
NOR3_X1 _15516_ ( .A1(_07135_ ), .A2(fanout_net_4 ), .A3(\myidu.stall_quest_fencei ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AOI21_X1 _15517_ ( .A(_01201_ ), .B1(_02362_ ), .B2(_01314_ ), .ZN(_00356_ ) );
AND2_X1 _15518_ ( .A1(_01200_ ), .A2(\myifu.state [0] ), .ZN(_00357_ ) );
OR4_X1 _15519_ ( .A1(_07026_ ), .A2(_00356_ ), .A3(_07030_ ), .A4(_00357_ ), .ZN(_00358_ ) );
AOI21_X1 _15520_ ( .A(_00358_ ), .B1(_00354_ ), .B2(\myifu.state [2] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _15521_ ( .A1(_02916_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_02524_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
INV_X1 _15522_ ( .A(fanout_net_43 ), .ZN(_00359_ ) );
MUX2_X1 _15523_ ( .A(_00359_ ), .B(_03153_ ), .S(\mylsu.state [0] ), .Z(_00360_ ) );
AOI21_X1 _15524_ ( .A(_00360_ ), .B1(_03233_ ), .B2(fanout_net_43 ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ) );
AOI211_X1 _15525_ ( .A(_03141_ ), .B(_00360_ ), .C1(_03233_ ), .C2(fanout_net_43 ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
INV_X1 _15526_ ( .A(_03088_ ), .ZN(_00361_ ) );
NAND2_X1 _15527_ ( .A1(_00361_ ), .A2(_03079_ ), .ZN(_00362_ ) );
NOR2_X1 _15528_ ( .A1(_01339_ ), .A2(_00362_ ), .ZN(_00363_ ) );
AND2_X1 _15529_ ( .A1(_01290_ ), .A2(_03128_ ), .ZN(_00364_ ) );
NAND4_X1 _15530_ ( .A1(_02365_ ), .A2(\mylsu.state [0] ), .A3(_00363_ ), .A4(_00364_ ), .ZN(_00365_ ) );
OAI21_X1 _15531_ ( .A(_00365_ ), .B1(_03232_ ), .B2(_03147_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND2_X1 _15532_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_00366_ ) );
AOI21_X1 _15533_ ( .A(_00366_ ), .B1(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .B2(_03087_ ), .ZN(_00367_ ) );
AND4_X1 _15534_ ( .A1(io_master_awready ), .A2(_03129_ ), .A3(_01303_ ), .A4(_00367_ ), .ZN(_00368_ ) );
NAND3_X1 _15535_ ( .A1(_03119_ ), .A2(\mylsu.state [0] ), .A3(_00368_ ), .ZN(_00369_ ) );
NAND3_X1 _15536_ ( .A1(_03140_ ), .A2(\mylsu.state [2] ), .A3(_03281_ ), .ZN(_00370_ ) );
NAND2_X1 _15537_ ( .A1(_00369_ ), .A2(_00370_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
BUF_X2 _15538_ ( .A(_00361_ ), .Z(_00371_ ) );
AND4_X1 _15539_ ( .A1(EXU_valid_LSU ), .A2(_00371_ ), .A3(_01303_ ), .A4(_00366_ ), .ZN(_00372_ ) );
NAND4_X1 _15540_ ( .A1(_03119_ ), .A2(\mylsu.state [0] ), .A3(_03140_ ), .A4(_00372_ ), .ZN(_00373_ ) );
NAND3_X1 _15541_ ( .A1(_03140_ ), .A2(\mylsu.state [4] ), .A3(io_master_awready ), .ZN(_00374_ ) );
NAND3_X1 _15542_ ( .A1(_03140_ ), .A2(\mylsu.state [2] ), .A3(io_master_wready ), .ZN(_00375_ ) );
OAI211_X1 _15543_ ( .A(_03140_ ), .B(\mylsu.state [1] ), .C1(_03216_ ), .C2(_03218_ ), .ZN(_00376_ ) );
NAND4_X1 _15544_ ( .A1(_00373_ ), .A2(_00374_ ), .A3(_00375_ ), .A4(_00376_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
AND4_X1 _15545_ ( .A1(_03281_ ), .A2(_01302_ ), .A3(_02369_ ), .A4(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_00377_ ) );
AND4_X1 _15546_ ( .A1(_03128_ ), .A2(_00377_ ), .A3(_03079_ ), .A4(_00367_ ), .ZN(_00378_ ) );
AND3_X1 _15547_ ( .A1(_01310_ ), .A2(\mylsu.state [0] ), .A3(_00378_ ), .ZN(_00379_ ) );
NAND3_X1 _15548_ ( .A1(_02367_ ), .A2(\mylsu.state [0] ), .A3(_00363_ ), .ZN(_00380_ ) );
NAND4_X1 _15549_ ( .A1(_03129_ ), .A2(\mylsu.state [0] ), .A3(_03081_ ), .A4(_03099_ ), .ZN(_00381_ ) );
NAND4_X1 _15550_ ( .A1(_01295_ ), .A2(_03079_ ), .A3(_01290_ ), .A4(_01296_ ), .ZN(_00382_ ) );
AOI21_X1 _15551_ ( .A(_00382_ ), .B1(_01288_ ), .B2(_01292_ ), .ZN(_00383_ ) );
NAND3_X1 _15552_ ( .A1(_00383_ ), .A2(\mylsu.state [0] ), .A3(_00364_ ), .ZN(_00384_ ) );
NAND3_X1 _15553_ ( .A1(_00380_ ), .A2(_00381_ ), .A3(_00384_ ), .ZN(_00385_ ) );
AND4_X1 _15554_ ( .A1(\io_master_arid [1] ), .A2(_03223_ ), .A3(_00250_ ), .A4(_03231_ ), .ZN(_00386_ ) );
NOR2_X1 _15555_ ( .A1(_00362_ ), .A2(_03280_ ), .ZN(_00387_ ) );
OAI21_X1 _15556_ ( .A(_00387_ ), .B1(_03146_ ), .B2(_01309_ ), .ZN(_00388_ ) );
NAND3_X1 _15557_ ( .A1(_01288_ ), .A2(_01292_ ), .A3(_00364_ ), .ZN(_00389_ ) );
AND4_X1 _15558_ ( .A1(EXU_valid_LSU ), .A2(_00388_ ), .A3(_00361_ ), .A4(_00389_ ), .ZN(_00390_ ) );
INV_X1 _15559_ ( .A(\mylsu.state [0] ), .ZN(_00391_ ) );
OAI221_X1 _15560_ ( .A(_03140_ ), .B1(_03213_ ), .B2(_03219_ ), .C1(_00390_ ), .C2(_00391_ ), .ZN(_00392_ ) );
OR4_X1 _15561_ ( .A1(_00379_ ), .A2(_00385_ ), .A3(_00386_ ), .A4(_00392_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND4_X1 _15562_ ( .A1(_03119_ ), .A2(io_master_wready ), .A3(_03205_ ), .A4(_00367_ ), .ZN(_00393_ ) );
AOI211_X1 _15563_ ( .A(io_master_awready ), .B(_03141_ ), .C1(_00393_ ), .C2(_03211_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
MUX2_X1 _15564_ ( .A(\LS_WB_wdata_csreg [21] ), .B(\EX_LS_result_csreg_mem [21] ), .S(_03097_ ), .Z(_00394_ ) );
MUX2_X1 _15565_ ( .A(_00394_ ), .B(\EX_LS_pc [21] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
BUF_X4 _15566_ ( .A(_03098_ ), .Z(_00395_ ) );
AOI21_X1 _15567_ ( .A(\EX_LS_pc [20] ), .B1(_00395_ ), .B2(_00371_ ), .ZN(_00396_ ) );
MUX2_X1 _15568_ ( .A(\LS_WB_wdata_csreg [20] ), .B(\EX_LS_result_csreg_mem [20] ), .S(_04077_ ), .Z(_00397_ ) );
BUF_X4 _15569_ ( .A(_03085_ ), .Z(_00398_ ) );
OAI22_X1 _15570_ ( .A1(_00397_ ), .A2(_03090_ ), .B1(\EX_LS_pc [20] ), .B2(_00398_ ), .ZN(_00399_ ) );
AOI21_X1 _15571_ ( .A(_00396_ ), .B1(_03142_ ), .B2(_00399_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
AOI21_X1 _15572_ ( .A(\EX_LS_pc [19] ), .B1(_00395_ ), .B2(_03089_ ), .ZN(_00400_ ) );
BUF_X4 _15573_ ( .A(_03538_ ), .Z(_00401_ ) );
AOI221_X4 _15574_ ( .A(_03086_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [19] ), .C1(\LS_WB_wdata_csreg [19] ), .C2(_00401_ ), .ZN(_00402_ ) );
AOI21_X1 _15575_ ( .A(_00400_ ), .B1(_03132_ ), .B2(_00402_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _15576_ ( .A(\LS_WB_wdata_csreg [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_03097_ ), .Z(_00403_ ) );
MUX2_X1 _15577_ ( .A(_00403_ ), .B(\EX_LS_pc [18] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _15578_ ( .A(\LS_WB_wdata_csreg [17] ), .B(\EX_LS_result_csreg_mem [17] ), .S(_03097_ ), .Z(_00404_ ) );
MUX2_X1 _15579_ ( .A(_00404_ ), .B(\EX_LS_pc [17] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _15580_ ( .A(\LS_WB_wdata_csreg [16] ), .B(\EX_LS_result_csreg_mem [16] ), .S(_03097_ ), .Z(_00405_ ) );
MUX2_X1 _15581_ ( .A(_00405_ ), .B(\EX_LS_pc [16] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
OAI21_X1 _15582_ ( .A(_00398_ ), .B1(_03097_ ), .B2(_01336_ ), .ZN(_00406_ ) );
AOI211_X1 _15583_ ( .A(_00406_ ), .B(_03137_ ), .C1(\EX_LS_result_csreg_mem [15] ), .C2(_03097_ ), .ZN(_00407_ ) );
AOI21_X1 _15584_ ( .A(\EX_LS_pc [15] ), .B1(_03142_ ), .B2(_03089_ ), .ZN(_00408_ ) );
NOR2_X1 _15585_ ( .A1(_00407_ ), .A2(_00408_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _15586_ ( .A(\EX_LS_pc [14] ), .B1(_00395_ ), .B2(_00371_ ), .ZN(_00409_ ) );
MUX2_X1 _15587_ ( .A(\LS_WB_wdata_csreg [14] ), .B(\EX_LS_result_csreg_mem [14] ), .S(_04077_ ), .Z(_00410_ ) );
OAI22_X1 _15588_ ( .A1(_00410_ ), .A2(_03090_ ), .B1(\EX_LS_pc [14] ), .B2(_00398_ ), .ZN(_00411_ ) );
AOI21_X1 _15589_ ( .A(_00409_ ), .B1(_03142_ ), .B2(_00411_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
AOI21_X1 _15590_ ( .A(\EX_LS_pc [13] ), .B1(_00395_ ), .B2(_03089_ ), .ZN(_00412_ ) );
AOI221_X4 _15591_ ( .A(_03086_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [13] ), .C1(\LS_WB_wdata_csreg [13] ), .C2(_00401_ ), .ZN(_00413_ ) );
AOI21_X1 _15592_ ( .A(_00412_ ), .B1(_03132_ ), .B2(_00413_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
AOI21_X1 _15593_ ( .A(\EX_LS_pc [12] ), .B1(_00395_ ), .B2(_03089_ ), .ZN(_00414_ ) );
AOI221_X4 _15594_ ( .A(_03086_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [12] ), .C1(\LS_WB_wdata_csreg [12] ), .C2(_00401_ ), .ZN(_00415_ ) );
AOI21_X1 _15595_ ( .A(_00414_ ), .B1(_03132_ ), .B2(_00415_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _15596_ ( .A(\EX_LS_pc [30] ), .B1(_00395_ ), .B2(_03089_ ), .ZN(_00416_ ) );
AOI221_X4 _15597_ ( .A(_03086_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [30] ), .C1(\LS_WB_wdata_csreg [30] ), .C2(_00401_ ), .ZN(_00417_ ) );
AOI21_X1 _15598_ ( .A(_00416_ ), .B1(_03132_ ), .B2(_00417_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _15599_ ( .A(\LS_WB_wdata_csreg [11] ), .B(\EX_LS_result_csreg_mem [11] ), .S(_03097_ ), .Z(_00418_ ) );
MUX2_X1 _15600_ ( .A(_00418_ ), .B(\EX_LS_pc [11] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
BUF_X4 _15601_ ( .A(_03096_ ), .Z(_00419_ ) );
MUX2_X1 _15602_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_00419_ ), .Z(_00420_ ) );
MUX2_X1 _15603_ ( .A(_00420_ ), .B(\EX_LS_pc [10] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
AOI21_X1 _15604_ ( .A(\EX_LS_pc [9] ), .B1(_00395_ ), .B2(_00371_ ), .ZN(_00421_ ) );
MUX2_X1 _15605_ ( .A(\LS_WB_wdata_csreg [9] ), .B(\EX_LS_result_csreg_mem [9] ), .S(_04077_ ), .Z(_00422_ ) );
OAI22_X1 _15606_ ( .A1(_00422_ ), .A2(_03090_ ), .B1(\EX_LS_pc [9] ), .B2(_00398_ ), .ZN(_00423_ ) );
AOI21_X1 _15607_ ( .A(_00421_ ), .B1(_03142_ ), .B2(_00423_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _15608_ ( .A(\LS_WB_wdata_csreg [8] ), .B(\EX_LS_result_csreg_mem [8] ), .S(_00419_ ), .Z(_00424_ ) );
MUX2_X1 _15609_ ( .A(_00424_ ), .B(\EX_LS_pc [8] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
AOI21_X1 _15610_ ( .A(\EX_LS_pc [7] ), .B1(_03142_ ), .B2(_03089_ ), .ZN(_00425_ ) );
OAI211_X1 _15611_ ( .A(_00371_ ), .B(_00398_ ), .C1(_00401_ ), .C2(_03250_ ), .ZN(_00426_ ) );
AOI221_X4 _15612_ ( .A(_00426_ ), .B1(\LS_WB_wdata_csreg [7] ), .B2(_00401_ ), .C1(_01341_ ), .C2(_01303_ ), .ZN(_00427_ ) );
NOR2_X1 _15613_ ( .A1(_00425_ ), .A2(_00427_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
AOI21_X1 _15614_ ( .A(\EX_LS_pc [6] ), .B1(_03142_ ), .B2(_03089_ ), .ZN(_00428_ ) );
OAI211_X1 _15615_ ( .A(_00371_ ), .B(_00398_ ), .C1(_00401_ ), .C2(_03251_ ), .ZN(_00429_ ) );
AOI221_X4 _15616_ ( .A(_00429_ ), .B1(\LS_WB_wdata_csreg [6] ), .B2(_00401_ ), .C1(_01341_ ), .C2(_01303_ ), .ZN(_00430_ ) );
NOR2_X1 _15617_ ( .A1(_00428_ ), .A2(_00430_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _15618_ ( .A(\LS_WB_wdata_csreg [5] ), .B(\EX_LS_result_csreg_mem [5] ), .S(_00419_ ), .Z(_00431_ ) );
MUX2_X1 _15619_ ( .A(_00431_ ), .B(\EX_LS_pc [5] ), .S(_03093_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _15620_ ( .A(\LS_WB_wdata_csreg [4] ), .B(\EX_LS_result_csreg_mem [4] ), .S(_00419_ ), .Z(_00432_ ) );
MUX2_X1 _15621_ ( .A(_00432_ ), .B(\EX_LS_pc [4] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _15622_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\EX_LS_result_csreg_mem [3] ), .S(_00419_ ), .Z(_00433_ ) );
MUX2_X1 _15623_ ( .A(_00433_ ), .B(\EX_LS_pc [3] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
OAI211_X1 _15624_ ( .A(_00371_ ), .B(_00398_ ), .C1(_03538_ ), .C2(_03241_ ), .ZN(_00434_ ) );
AOI221_X4 _15625_ ( .A(_00434_ ), .B1(\LS_WB_wdata_csreg [2] ), .B2(_00401_ ), .C1(_01341_ ), .C2(_01303_ ), .ZN(_00435_ ) );
AOI21_X1 _15626_ ( .A(_00435_ ), .B1(_03078_ ), .B2(_03093_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _15627_ ( .A(\LS_WB_wdata_csreg [29] ), .B(\EX_LS_result_csreg_mem [29] ), .S(_00419_ ), .Z(_00436_ ) );
MUX2_X1 _15628_ ( .A(_00436_ ), .B(\EX_LS_pc [29] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _15629_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\EX_LS_result_csreg_mem [1] ), .S(_00419_ ), .Z(_00437_ ) );
MUX2_X1 _15630_ ( .A(_00437_ ), .B(\EX_LS_pc [1] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _15631_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\EX_LS_result_csreg_mem [0] ), .S(_00419_ ), .Z(_00438_ ) );
MUX2_X1 _15632_ ( .A(_00438_ ), .B(\EX_LS_pc [0] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _15633_ ( .A(\LS_WB_wdata_csreg [28] ), .B(\EX_LS_result_csreg_mem [28] ), .S(_00419_ ), .Z(_00439_ ) );
MUX2_X1 _15634_ ( .A(_00439_ ), .B(\EX_LS_pc [28] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _15635_ ( .A(\EX_LS_pc [27] ), .B1(_00395_ ), .B2(_00371_ ), .ZN(_00440_ ) );
MUX2_X1 _15636_ ( .A(\LS_WB_wdata_csreg [27] ), .B(\EX_LS_result_csreg_mem [27] ), .S(_04077_ ), .Z(_00441_ ) );
OAI22_X1 _15637_ ( .A1(_00441_ ), .A2(_03090_ ), .B1(\EX_LS_pc [27] ), .B2(_00398_ ), .ZN(_00442_ ) );
AOI21_X1 _15638_ ( .A(_00440_ ), .B1(_03142_ ), .B2(_00442_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI21_X1 _15639_ ( .A(\EX_LS_pc [26] ), .B1(_00395_ ), .B2(_00371_ ), .ZN(_00443_ ) );
MUX2_X1 _15640_ ( .A(\LS_WB_wdata_csreg [26] ), .B(\EX_LS_result_csreg_mem [26] ), .S(_04077_ ), .Z(_00444_ ) );
OAI22_X1 _15641_ ( .A1(_00444_ ), .A2(_03090_ ), .B1(\EX_LS_pc [26] ), .B2(_00398_ ), .ZN(_00445_ ) );
AOI21_X1 _15642_ ( .A(_00443_ ), .B1(_03142_ ), .B2(_00445_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI21_X1 _15643_ ( .A(\EX_LS_pc [25] ), .B1(_00395_ ), .B2(_03089_ ), .ZN(_00446_ ) );
AOI221_X4 _15644_ ( .A(_03086_ ), .B1(\EX_LS_flag [2] ), .B2(\EX_LS_result_csreg_mem [25] ), .C1(\LS_WB_wdata_csreg [25] ), .C2(_00401_ ), .ZN(_00447_ ) );
AOI21_X1 _15645_ ( .A(_00446_ ), .B1(_03132_ ), .B2(_00447_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _15646_ ( .A(\EX_LS_pc [24] ), .B1(_03098_ ), .B2(_00371_ ), .ZN(_00448_ ) );
MUX2_X1 _15647_ ( .A(\LS_WB_wdata_csreg [24] ), .B(\EX_LS_result_csreg_mem [24] ), .S(_04077_ ), .Z(_00449_ ) );
OAI22_X1 _15648_ ( .A1(_00449_ ), .A2(_03090_ ), .B1(\EX_LS_pc [24] ), .B2(_00398_ ), .ZN(_00450_ ) );
AOI21_X1 _15649_ ( .A(_00448_ ), .B1(_03142_ ), .B2(_00450_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _15650_ ( .A(\EX_LS_pc [23] ), .B1(_03098_ ), .B2(_03089_ ), .ZN(_00451_ ) );
AOI221_X4 _15651_ ( .A(_03086_ ), .B1(\LS_WB_wdata_csreg [23] ), .B2(_03083_ ), .C1(\EX_LS_result_csreg_mem [23] ), .C2(_03097_ ), .ZN(_00452_ ) );
AOI21_X1 _15652_ ( .A(_00451_ ), .B1(_03132_ ), .B2(_00452_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _15653_ ( .A(\LS_WB_wdata_csreg [22] ), .B(\EX_LS_result_csreg_mem [22] ), .S(_00419_ ), .Z(_00453_ ) );
MUX2_X1 _15654_ ( .A(_00453_ ), .B(\EX_LS_pc [22] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _15655_ ( .A(\LS_WB_wdata_csreg [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_04077_ ), .Z(_00454_ ) );
MUX2_X1 _15656_ ( .A(_00454_ ), .B(\EX_LS_pc [31] ), .S(_03092_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _15657_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_00455_ ) );
INV_X1 _15658_ ( .A(_00455_ ), .ZN(_00456_ ) );
BUF_X2 _15659_ ( .A(_00456_ ), .Z(_00457_ ) );
NAND3_X1 _15660_ ( .A1(_07033_ ), .A2(_02364_ ), .A3(_00457_ ), .ZN(_00458_ ) );
OR3_X1 _15661_ ( .A1(_07064_ ), .A2(_03155_ ), .A3(_00456_ ), .ZN(_00459_ ) );
NAND2_X1 _15662_ ( .A1(_00458_ ), .A2(_00459_ ), .ZN(_00460_ ) );
AND2_X1 _15663_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_00461_ ) );
INV_X1 _15664_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_00462_ ) );
AND2_X2 _15665_ ( .A1(_00461_ ), .A2(_00462_ ), .ZN(_00463_ ) );
INV_X1 _15666_ ( .A(_00463_ ), .ZN(_00464_ ) );
NOR2_X2 _15667_ ( .A1(_00460_ ), .A2(_00464_ ), .ZN(_00465_ ) );
INV_X1 _15668_ ( .A(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_00466_ ) );
NOR2_X1 _15669_ ( .A1(_00466_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_00467_ ) );
INV_X1 _15670_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_00468_ ) );
AND2_X1 _15671_ ( .A1(_00467_ ), .A2(_00468_ ), .ZN(_00469_ ) );
NAND2_X1 _15672_ ( .A1(_00468_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_00470_ ) );
NOR2_X2 _15673_ ( .A1(_00470_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_00471_ ) );
OR2_X1 _15674_ ( .A1(_00469_ ), .A2(_00471_ ), .ZN(_00472_ ) );
NOR2_X2 _15675_ ( .A1(_00465_ ), .A2(_00472_ ), .ZN(_00473_ ) );
BUF_X4 _15676_ ( .A(_00473_ ), .Z(_00474_ ) );
BUF_X4 _15677_ ( .A(_00463_ ), .Z(_00475_ ) );
BUF_X4 _15678_ ( .A(_00475_ ), .Z(_00476_ ) );
NAND2_X1 _15679_ ( .A1(_07043_ ), .A2(_07045_ ), .ZN(_00477_ ) );
AND2_X2 _15680_ ( .A1(_00461_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_00478_ ) );
BUF_X4 _15681_ ( .A(_00478_ ), .Z(_00479_ ) );
NOR3_X1 _15682_ ( .A1(_00477_ ), .A2(_03158_ ), .A3(_00479_ ), .ZN(_00480_ ) );
OAI21_X1 _15683_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00480_ ), .ZN(_00481_ ) );
BUF_X2 _15684_ ( .A(_03155_ ), .Z(_00482_ ) );
NOR2_X1 _15685_ ( .A1(_03163_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_00483_ ) );
INV_X1 _15686_ ( .A(_00483_ ), .ZN(_00484_ ) );
NOR3_X1 _15687_ ( .A1(_07064_ ), .A2(_00482_ ), .A3(_00484_ ), .ZN(_00485_ ) );
NOR2_X1 _15688_ ( .A1(_03159_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_00486_ ) );
NOR2_X1 _15689_ ( .A1(_07130_ ), .A2(_03156_ ), .ZN(_00487_ ) );
AOI21_X1 _15690_ ( .A(_00485_ ), .B1(_00486_ ), .B2(_00487_ ), .ZN(_00488_ ) );
NAND4_X1 _15691_ ( .A1(_07033_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_02364_ ), .ZN(_00489_ ) );
OR3_X1 _15692_ ( .A1(_07091_ ), .A2(_00482_ ), .A3(_00457_ ), .ZN(_00490_ ) );
AND3_X2 _15693_ ( .A1(_00488_ ), .A2(_00489_ ), .A3(_00490_ ), .ZN(_00491_ ) );
BUF_X4 _15694_ ( .A(_00491_ ), .Z(_00492_ ) );
INV_X2 _15695_ ( .A(_00469_ ), .ZN(_00493_ ) );
BUF_X4 _15696_ ( .A(_00493_ ), .Z(_00494_ ) );
NOR2_X1 _15697_ ( .A1(_00492_ ), .A2(_00494_ ), .ZN(_00495_ ) );
NOR2_X1 _15698_ ( .A1(_00495_ ), .A2(_00359_ ), .ZN(_00496_ ) );
AOI22_X1 _15699_ ( .A1(_00481_ ), .A2(_00496_ ), .B1(_00359_ ), .B2(_03522_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
NAND3_X1 _15700_ ( .A1(_07046_ ), .A2(_07049_ ), .A3(_02363_ ), .ZN(_00497_ ) );
NOR2_X1 _15701_ ( .A1(_00497_ ), .A2(_00479_ ), .ZN(_00498_ ) );
OAI21_X1 _15702_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00498_ ), .ZN(_00499_ ) );
BUF_X4 _15703_ ( .A(_00493_ ), .Z(_00500_ ) );
BUF_X4 _15704_ ( .A(_00491_ ), .Z(_00501_ ) );
OAI21_X1 _15705_ ( .A(_00499_ ), .B1(_00500_ ), .B2(_00501_ ), .ZN(_00502_ ) );
MUX2_X1 _15706_ ( .A(\EX_LS_result_reg [20] ), .B(_00502_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _15707_ ( .A1(_07050_ ), .A2(\io_master_arid [1] ), .A3(_07052_ ), .ZN(_00503_ ) );
NOR2_X1 _15708_ ( .A1(_00503_ ), .A2(_00479_ ), .ZN(_00504_ ) );
OAI21_X1 _15709_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00504_ ), .ZN(_00505_ ) );
OAI21_X1 _15710_ ( .A(_00505_ ), .B1(_00500_ ), .B2(_00501_ ), .ZN(_00506_ ) );
MUX2_X1 _15711_ ( .A(\EX_LS_result_reg [19] ), .B(_00506_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _15712_ ( .A1(_07053_ ), .A2(_07055_ ), .A3(_02363_ ), .ZN(_00507_ ) );
NOR2_X1 _15713_ ( .A1(_00507_ ), .A2(_00479_ ), .ZN(_00508_ ) );
OAI21_X1 _15714_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00508_ ), .ZN(_00509_ ) );
OAI21_X1 _15715_ ( .A(_00509_ ), .B1(_00500_ ), .B2(_00501_ ), .ZN(_00510_ ) );
MUX2_X1 _15716_ ( .A(\EX_LS_result_reg [18] ), .B(_00510_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NOR4_X1 _15717_ ( .A1(_07056_ ), .A2(_03156_ ), .A3(_07058_ ), .A4(_00479_ ), .ZN(_00511_ ) );
OAI21_X1 _15718_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00511_ ), .ZN(_00512_ ) );
OAI21_X1 _15719_ ( .A(_00512_ ), .B1(_00500_ ), .B2(_00501_ ), .ZN(_00513_ ) );
MUX2_X1 _15720_ ( .A(\EX_LS_result_reg [17] ), .B(_00513_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _15721_ ( .A1(_07059_ ), .A2(_07061_ ), .A3(_02363_ ), .ZN(_00514_ ) );
NOR2_X1 _15722_ ( .A1(_00514_ ), .A2(_00479_ ), .ZN(_00515_ ) );
OAI21_X1 _15723_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00515_ ), .ZN(_00516_ ) );
OAI21_X1 _15724_ ( .A(_00516_ ), .B1(_00500_ ), .B2(_00501_ ), .ZN(_00517_ ) );
MUX2_X1 _15725_ ( .A(\EX_LS_result_reg [16] ), .B(_00517_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
BUF_X2 _15726_ ( .A(_00469_ ), .Z(_00518_ ) );
BUF_X2 _15727_ ( .A(_00461_ ), .Z(_00519_ ) );
OR3_X1 _15728_ ( .A1(_00518_ ), .A2(_00519_ ), .A3(_00471_ ), .ZN(_00520_ ) );
OR3_X1 _15729_ ( .A1(_07064_ ), .A2(_03157_ ), .A3(_00520_ ), .ZN(_00521_ ) );
NAND2_X1 _15730_ ( .A1(_00460_ ), .A2(_00519_ ), .ZN(_00522_ ) );
OAI211_X1 _15731_ ( .A(_00521_ ), .B(_00522_ ), .C1(_00501_ ), .C2(_00494_ ), .ZN(_00523_ ) );
MUX2_X1 _15732_ ( .A(\EX_LS_result_reg [15] ), .B(_00523_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
INV_X1 _15733_ ( .A(_00471_ ), .ZN(_00524_ ) );
NAND2_X1 _15734_ ( .A1(_00457_ ), .A2(_00461_ ), .ZN(_00525_ ) );
NAND3_X1 _15735_ ( .A1(_00493_ ), .A2(_00524_ ), .A3(_00525_ ), .ZN(_00526_ ) );
NOR2_X1 _15736_ ( .A1(_03156_ ), .A2(_00526_ ), .ZN(_00527_ ) );
OAI211_X1 _15737_ ( .A(_07067_ ), .B(_00527_ ), .C1(_03202_ ), .C2(\io_master_rdata [14] ), .ZN(_00528_ ) );
NAND2_X1 _15738_ ( .A1(_07034_ ), .A2(_07042_ ), .ZN(_00529_ ) );
OR3_X1 _15739_ ( .A1(_00529_ ), .A2(_03156_ ), .A3(_00525_ ), .ZN(_00530_ ) );
OAI211_X1 _15740_ ( .A(_00528_ ), .B(_00530_ ), .C1(_00501_ ), .C2(_00494_ ), .ZN(_00531_ ) );
MUX2_X1 _15741_ ( .A(\EX_LS_result_reg [14] ), .B(_00531_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
OR3_X1 _15742_ ( .A1(_07076_ ), .A2(_03157_ ), .A3(_00525_ ), .ZN(_00532_ ) );
OAI211_X1 _15743_ ( .A(_07070_ ), .B(_00527_ ), .C1(_03202_ ), .C2(\io_master_rdata [13] ), .ZN(_00533_ ) );
OAI211_X1 _15744_ ( .A(_00532_ ), .B(_00533_ ), .C1(_00501_ ), .C2(_00494_ ), .ZN(_00534_ ) );
MUX2_X1 _15745_ ( .A(\EX_LS_result_reg [13] ), .B(_00534_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _15746_ ( .A1(_07071_ ), .A2(_07073_ ), .A3(_00527_ ), .ZN(_00535_ ) );
NAND2_X1 _15747_ ( .A1(_07107_ ), .A2(_07109_ ), .ZN(_00536_ ) );
OR2_X2 _15748_ ( .A1(_00536_ ), .A2(_03155_ ), .ZN(_00537_ ) );
OAI221_X1 _15749_ ( .A(_00535_ ), .B1(_00525_ ), .B2(_00537_ ), .C1(_00492_ ), .C2(_00494_ ), .ZN(_00538_ ) );
MUX2_X1 _15750_ ( .A(\EX_LS_result_reg [12] ), .B(_00538_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
NOR3_X1 _15751_ ( .A1(_00529_ ), .A2(_03157_ ), .A3(_00519_ ), .ZN(_00539_ ) );
OAI21_X1 _15752_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00539_ ), .ZN(_00540_ ) );
OAI21_X1 _15753_ ( .A(_00540_ ), .B1(_00500_ ), .B2(_00492_ ), .ZN(_00541_ ) );
MUX2_X1 _15754_ ( .A(\EX_LS_result_reg [30] ), .B(_00541_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
OAI211_X1 _15755_ ( .A(_07079_ ), .B(_00527_ ), .C1(_03202_ ), .C2(\io_master_rdata [11] ), .ZN(_00542_ ) );
NAND2_X2 _15756_ ( .A1(_07116_ ), .A2(_07118_ ), .ZN(_00543_ ) );
OR2_X1 _15757_ ( .A1(_00543_ ), .A2(_03155_ ), .ZN(_00544_ ) );
OAI221_X1 _15758_ ( .A(_00542_ ), .B1(_00525_ ), .B2(_00544_ ), .C1(_00491_ ), .C2(_00493_ ), .ZN(_00545_ ) );
MUX2_X1 _15759_ ( .A(\EX_LS_result_reg [11] ), .B(_00545_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
OAI211_X1 _15760_ ( .A(_07082_ ), .B(_00527_ ), .C1(_03202_ ), .C2(\io_master_rdata [10] ), .ZN(_00546_ ) );
NAND2_X1 _15761_ ( .A1(_07119_ ), .A2(_07121_ ), .ZN(_00547_ ) );
OR2_X2 _15762_ ( .A1(_00547_ ), .A2(_03155_ ), .ZN(_00548_ ) );
OAI221_X1 _15763_ ( .A(_00546_ ), .B1(_00525_ ), .B2(_00548_ ), .C1(_00491_ ), .C2(_00493_ ), .ZN(_00549_ ) );
MUX2_X1 _15764_ ( .A(\EX_LS_result_reg [10] ), .B(_00549_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
OAI211_X1 _15765_ ( .A(_07085_ ), .B(_00527_ ), .C1(_03202_ ), .C2(\io_master_rdata [9] ), .ZN(_00550_ ) );
NAND2_X1 _15766_ ( .A1(_07122_ ), .A2(_07124_ ), .ZN(_00551_ ) );
OR3_X1 _15767_ ( .A1(_00551_ ), .A2(_03156_ ), .A3(_00525_ ), .ZN(_00552_ ) );
OAI211_X1 _15768_ ( .A(_00550_ ), .B(_00552_ ), .C1(_00501_ ), .C2(_00494_ ), .ZN(_00553_ ) );
MUX2_X1 _15769_ ( .A(\EX_LS_result_reg [9] ), .B(_00553_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _15770_ ( .A1(_07086_ ), .A2(_07088_ ), .A3(_00527_ ), .ZN(_00554_ ) );
NAND2_X1 _15771_ ( .A1(_07125_ ), .A2(_07127_ ), .ZN(_00555_ ) );
OR2_X2 _15772_ ( .A1(_00555_ ), .A2(_03155_ ), .ZN(_00556_ ) );
OAI221_X1 _15773_ ( .A(_00554_ ), .B1(_00525_ ), .B2(_00556_ ), .C1(_00491_ ), .C2(_00493_ ), .ZN(_00557_ ) );
MUX2_X1 _15774_ ( .A(\EX_LS_result_reg [8] ), .B(_00557_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
NOR2_X1 _15775_ ( .A1(_07091_ ), .A2(_03157_ ), .ZN(_00558_ ) );
OAI221_X1 _15776_ ( .A(fanout_net_43 ), .B1(_00558_ ), .B2(_00526_ ), .C1(_00487_ ), .C2(_00525_ ), .ZN(_00559_ ) );
AOI21_X1 _15777_ ( .A(_00559_ ), .B1(_00501_ ), .B2(_00472_ ), .ZN(_00560_ ) );
AND2_X1 _15778_ ( .A1(_00359_ ), .A2(\EX_LS_result_reg [7] ), .ZN(_00561_ ) );
OR2_X1 _15779_ ( .A1(_00560_ ), .A2(_00561_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
INV_X1 _15780_ ( .A(_00486_ ), .ZN(_00562_ ) );
AND4_X1 _15781_ ( .A1(_02364_ ), .A2(_07034_ ), .A3(_07042_ ), .A4(_00562_ ), .ZN(_00563_ ) );
AND4_X1 _15782_ ( .A1(_02364_ ), .A2(_07131_ ), .A3(_07133_ ), .A4(_00486_ ), .ZN(_00564_ ) );
OAI21_X1 _15783_ ( .A(_00484_ ), .B1(_00563_ ), .B2(_00564_ ), .ZN(_00565_ ) );
BUF_X2 _15784_ ( .A(_00483_ ), .Z(_00566_ ) );
NAND4_X1 _15785_ ( .A1(_07065_ ), .A2(\io_master_arid [1] ), .A3(_07067_ ), .A4(_00566_ ), .ZN(_00567_ ) );
AOI21_X1 _15786_ ( .A(_00455_ ), .B1(_00565_ ), .B2(_00567_ ), .ZN(_00568_ ) );
NOR3_X1 _15787_ ( .A1(_07094_ ), .A2(_00482_ ), .A3(_00457_ ), .ZN(_00569_ ) );
OAI21_X1 _15788_ ( .A(_00518_ ), .B1(_00568_ ), .B2(_00569_ ), .ZN(_00570_ ) );
AND4_X1 _15789_ ( .A1(_02363_ ), .A2(_07131_ ), .A3(_07133_ ), .A4(_00456_ ), .ZN(_00571_ ) );
OR2_X1 _15790_ ( .A1(_00569_ ), .A2(_00571_ ), .ZN(_00572_ ) );
AND2_X1 _15791_ ( .A1(_00572_ ), .A2(_00463_ ), .ZN(_00573_ ) );
OAI21_X1 _15792_ ( .A(_00479_ ), .B1(_00569_ ), .B2(_00571_ ), .ZN(_00574_ ) );
OR3_X1 _15793_ ( .A1(_07094_ ), .A2(_03156_ ), .A3(_00478_ ), .ZN(_00575_ ) );
AOI21_X1 _15794_ ( .A(_00475_ ), .B1(_00574_ ), .B2(_00575_ ), .ZN(_00576_ ) );
OAI21_X1 _15795_ ( .A(_00524_ ), .B1(_00573_ ), .B2(_00576_ ), .ZN(_00577_ ) );
OAI21_X1 _15796_ ( .A(_00471_ ), .B1(_00568_ ), .B2(_00569_ ), .ZN(_00578_ ) );
AND2_X1 _15797_ ( .A1(_00577_ ), .A2(_00578_ ), .ZN(_00579_ ) );
OAI21_X1 _15798_ ( .A(_00570_ ), .B1(_00579_ ), .B2(_00518_ ), .ZN(_00580_ ) );
MUX2_X1 _15799_ ( .A(\EX_LS_result_reg [6] ), .B(_00580_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _15800_ ( .A1(_00520_ ), .A2(_00457_ ), .ZN(_00581_ ) );
AOI21_X1 _15801_ ( .A(_03158_ ), .B1(_07097_ ), .B2(_00581_ ), .ZN(_00582_ ) );
NAND2_X1 _15802_ ( .A1(_07068_ ), .A2(_07070_ ), .ZN(_00583_ ) );
NAND2_X1 _15803_ ( .A1(_00583_ ), .A2(_00566_ ), .ZN(_00584_ ) );
NAND3_X1 _15804_ ( .A1(_07076_ ), .A2(_00484_ ), .A3(_00562_ ), .ZN(_00585_ ) );
AOI22_X1 _15805_ ( .A1(_00584_ ), .A2(_00585_ ), .B1(_00493_ ), .B2(_00524_ ), .ZN(_00586_ ) );
OAI21_X1 _15806_ ( .A(_00562_ ), .B1(_00518_ ), .B2(_00471_ ), .ZN(_00587_ ) );
AOI21_X1 _15807_ ( .A(_00586_ ), .B1(_00477_ ), .B2(_00587_ ), .ZN(_00588_ ) );
OAI211_X1 _15808_ ( .A(fanout_net_43 ), .B(_00582_ ), .C1(_00588_ ), .C2(_00581_ ), .ZN(_00589_ ) );
NAND2_X1 _15809_ ( .A1(_00359_ ), .A2(\EX_LS_result_reg [5] ), .ZN(_00590_ ) );
NAND2_X1 _15810_ ( .A1(_00589_ ), .A2(_00590_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
MUX2_X2 _15811_ ( .A(_00497_ ), .B(_00537_ ), .S(_00562_ ), .Z(_00591_ ) );
OR2_X2 _15812_ ( .A1(_00591_ ), .A2(_00566_ ), .ZN(_00592_ ) );
NAND4_X1 _15813_ ( .A1(_07071_ ), .A2(_07073_ ), .A3(\io_master_arid [1] ), .A4(_00566_ ), .ZN(_00593_ ) );
AOI21_X2 _15814_ ( .A(_00455_ ), .B1(_00592_ ), .B2(_00593_ ), .ZN(_00594_ ) );
NOR3_X1 _15815_ ( .A1(_07100_ ), .A2(_00482_ ), .A3(_00456_ ), .ZN(_00595_ ) );
OAI21_X1 _15816_ ( .A(_00518_ ), .B1(_00594_ ), .B2(_00595_ ), .ZN(_00596_ ) );
OAI21_X1 _15817_ ( .A(_00471_ ), .B1(_00594_ ), .B2(_00595_ ), .ZN(_00597_ ) );
AND4_X1 _15818_ ( .A1(_02363_ ), .A2(_07046_ ), .A3(_07049_ ), .A4(_00456_ ), .ZN(_00598_ ) );
OR2_X1 _15819_ ( .A1(_00595_ ), .A2(_00598_ ), .ZN(_00599_ ) );
AND2_X1 _15820_ ( .A1(_00599_ ), .A2(_00463_ ), .ZN(_00600_ ) );
OAI21_X1 _15821_ ( .A(_00479_ ), .B1(_00595_ ), .B2(_00598_ ), .ZN(_00601_ ) );
OR3_X1 _15822_ ( .A1(_07100_ ), .A2(_03156_ ), .A3(_00478_ ), .ZN(_00602_ ) );
AOI21_X1 _15823_ ( .A(_00475_ ), .B1(_00601_ ), .B2(_00602_ ), .ZN(_00603_ ) );
OAI21_X1 _15824_ ( .A(_00524_ ), .B1(_00600_ ), .B2(_00603_ ), .ZN(_00604_ ) );
AND2_X1 _15825_ ( .A1(_00597_ ), .A2(_00604_ ), .ZN(_00605_ ) );
OAI21_X1 _15826_ ( .A(_00596_ ), .B1(_00605_ ), .B2(_00518_ ), .ZN(_00606_ ) );
MUX2_X1 _15827_ ( .A(\EX_LS_result_reg [4] ), .B(_00606_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
NOR3_X1 _15828_ ( .A1(_07103_ ), .A2(_03155_ ), .A3(_00456_ ), .ZN(_00607_ ) );
INV_X1 _15829_ ( .A(_00607_ ), .ZN(_00608_ ) );
AND4_X1 _15830_ ( .A1(_02363_ ), .A2(_07077_ ), .A3(_07079_ ), .A4(_00483_ ), .ZN(_00609_ ) );
NAND4_X1 _15831_ ( .A1(_07050_ ), .A2(_02364_ ), .A3(_07052_ ), .A4(_00486_ ), .ZN(_00610_ ) );
OAI21_X1 _15832_ ( .A(_00610_ ), .B1(_00544_ ), .B2(_00486_ ), .ZN(_00611_ ) );
AOI21_X1 _15833_ ( .A(_00609_ ), .B1(_00611_ ), .B2(_00484_ ), .ZN(_00612_ ) );
OAI21_X1 _15834_ ( .A(_00608_ ), .B1(_00612_ ), .B2(_00455_ ), .ZN(_00613_ ) );
AND4_X1 _15835_ ( .A1(_02363_ ), .A2(_07050_ ), .A3(_07052_ ), .A4(_00456_ ), .ZN(_00614_ ) );
OAI21_X1 _15836_ ( .A(_00463_ ), .B1(_00614_ ), .B2(_00607_ ), .ZN(_00615_ ) );
OAI21_X1 _15837_ ( .A(_00478_ ), .B1(_00614_ ), .B2(_00607_ ), .ZN(_00616_ ) );
OR3_X1 _15838_ ( .A1(_07103_ ), .A2(_03155_ ), .A3(_00478_ ), .ZN(_00617_ ) );
AND2_X1 _15839_ ( .A1(_00616_ ), .A2(_00617_ ), .ZN(_00618_ ) );
OAI21_X1 _15840_ ( .A(_00615_ ), .B1(_00618_ ), .B2(_00463_ ), .ZN(_00619_ ) );
MUX2_X1 _15841_ ( .A(_00619_ ), .B(_00613_ ), .S(_00471_ ), .Z(_00620_ ) );
MUX2_X1 _15842_ ( .A(_00613_ ), .B(_00620_ ), .S(_00493_ ), .Z(_00621_ ) );
MUX2_X1 _15843_ ( .A(\EX_LS_result_reg [3] ), .B(_00621_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
MUX2_X1 _15844_ ( .A(_00507_ ), .B(_00548_ ), .S(_00562_ ), .Z(_00622_ ) );
OR2_X2 _15845_ ( .A1(_00622_ ), .A2(_00566_ ), .ZN(_00623_ ) );
NAND4_X1 _15846_ ( .A1(_07080_ ), .A2(\io_master_arid [1] ), .A3(_07082_ ), .A4(_00566_ ), .ZN(_00624_ ) );
AOI21_X2 _15847_ ( .A(_00455_ ), .B1(_00623_ ), .B2(_00624_ ), .ZN(_00625_ ) );
NOR3_X1 _15848_ ( .A1(_07106_ ), .A2(_03155_ ), .A3(_00456_ ), .ZN(_00626_ ) );
OAI21_X1 _15849_ ( .A(_00518_ ), .B1(_00625_ ), .B2(_00626_ ), .ZN(_00627_ ) );
OAI21_X1 _15850_ ( .A(_00471_ ), .B1(_00625_ ), .B2(_00626_ ), .ZN(_00628_ ) );
AND4_X1 _15851_ ( .A1(_02363_ ), .A2(_07053_ ), .A3(_07055_ ), .A4(_00456_ ), .ZN(_00629_ ) );
OR2_X1 _15852_ ( .A1(_00626_ ), .A2(_00629_ ), .ZN(_00630_ ) );
AND2_X1 _15853_ ( .A1(_00630_ ), .A2(_00463_ ), .ZN(_00631_ ) );
OAI21_X1 _15854_ ( .A(_00478_ ), .B1(_00626_ ), .B2(_00629_ ), .ZN(_00632_ ) );
OR3_X1 _15855_ ( .A1(_07106_ ), .A2(_00482_ ), .A3(_00478_ ), .ZN(_00633_ ) );
AOI21_X1 _15856_ ( .A(_00463_ ), .B1(_00632_ ), .B2(_00633_ ), .ZN(_00634_ ) );
OAI21_X1 _15857_ ( .A(_00524_ ), .B1(_00631_ ), .B2(_00634_ ), .ZN(_00635_ ) );
AND2_X1 _15858_ ( .A1(_00628_ ), .A2(_00635_ ), .ZN(_00636_ ) );
OAI21_X1 _15859_ ( .A(_00627_ ), .B1(_00636_ ), .B2(_00518_ ), .ZN(_00637_ ) );
MUX2_X1 _15860_ ( .A(\EX_LS_result_reg [2] ), .B(_00637_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
NOR3_X1 _15861_ ( .A1(_07076_ ), .A2(_03157_ ), .A3(_00519_ ), .ZN(_00638_ ) );
OAI21_X1 _15862_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00638_ ), .ZN(_00639_ ) );
OAI21_X1 _15863_ ( .A(_00639_ ), .B1(_00500_ ), .B2(_00492_ ), .ZN(_00640_ ) );
MUX2_X1 _15864_ ( .A(\EX_LS_result_reg [29] ), .B(_00640_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
NAND4_X1 _15865_ ( .A1(_07122_ ), .A2(_02364_ ), .A3(_07124_ ), .A4(_00562_ ), .ZN(_00641_ ) );
OR4_X2 _15866_ ( .A1(_00482_ ), .A2(_07056_ ), .A3(_07058_ ), .A4(_00562_ ), .ZN(_00642_ ) );
AOI21_X1 _15867_ ( .A(_00566_ ), .B1(_00641_ ), .B2(_00642_ ), .ZN(_00643_ ) );
AND4_X1 _15868_ ( .A1(_02364_ ), .A2(_07083_ ), .A3(_07085_ ), .A4(_00566_ ), .ZN(_00644_ ) );
OAI21_X1 _15869_ ( .A(_00457_ ), .B1(_00643_ ), .B2(_00644_ ), .ZN(_00645_ ) );
OR3_X1 _15870_ ( .A1(_07112_ ), .A2(_03156_ ), .A3(_00457_ ), .ZN(_00646_ ) );
AOI21_X1 _15871_ ( .A(_00524_ ), .B1(_00645_ ), .B2(_00646_ ), .ZN(_00647_ ) );
NOR4_X1 _15872_ ( .A1(_07056_ ), .A2(_00482_ ), .A3(_07058_ ), .A4(_00455_ ), .ZN(_00648_ ) );
NOR3_X1 _15873_ ( .A1(_07112_ ), .A2(_00482_ ), .A3(_00457_ ), .ZN(_00649_ ) );
OAI21_X1 _15874_ ( .A(_00478_ ), .B1(_00648_ ), .B2(_00649_ ), .ZN(_00650_ ) );
OR3_X1 _15875_ ( .A1(_07112_ ), .A2(_00482_ ), .A3(_00478_ ), .ZN(_00651_ ) );
NAND2_X1 _15876_ ( .A1(_00650_ ), .A2(_00651_ ), .ZN(_00652_ ) );
NAND2_X1 _15877_ ( .A1(_00652_ ), .A2(_00464_ ), .ZN(_00653_ ) );
OAI21_X1 _15878_ ( .A(_00475_ ), .B1(_00648_ ), .B2(_00649_ ), .ZN(_00654_ ) );
AOI21_X1 _15879_ ( .A(_00471_ ), .B1(_00653_ ), .B2(_00654_ ), .ZN(_00655_ ) );
OAI21_X1 _15880_ ( .A(_00493_ ), .B1(_00647_ ), .B2(_00655_ ), .ZN(_00656_ ) );
AND2_X1 _15881_ ( .A1(_00645_ ), .A2(_00646_ ), .ZN(_00657_ ) );
OAI21_X1 _15882_ ( .A(_00656_ ), .B1(_00500_ ), .B2(_00657_ ), .ZN(_00658_ ) );
MUX2_X1 _15883_ ( .A(\EX_LS_result_reg [1] ), .B(_00658_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _15884_ ( .A(_00514_ ), .B(_00556_ ), .S(_00562_ ), .Z(_00659_ ) );
OR2_X2 _15885_ ( .A1(_00659_ ), .A2(_00566_ ), .ZN(_00660_ ) );
NAND4_X1 _15886_ ( .A1(_07086_ ), .A2(_07088_ ), .A3(_02364_ ), .A4(_00566_ ), .ZN(_00661_ ) );
AOI21_X2 _15887_ ( .A(_00455_ ), .B1(_00660_ ), .B2(_00661_ ), .ZN(_00662_ ) );
NOR3_X1 _15888_ ( .A1(_07115_ ), .A2(_00482_ ), .A3(_00457_ ), .ZN(_00663_ ) );
OAI21_X1 _15889_ ( .A(_00518_ ), .B1(_00662_ ), .B2(_00663_ ), .ZN(_00664_ ) );
OAI21_X1 _15890_ ( .A(_00471_ ), .B1(_00662_ ), .B2(_00663_ ), .ZN(_00665_ ) );
AND4_X1 _15891_ ( .A1(_02364_ ), .A2(_07059_ ), .A3(_07061_ ), .A4(_00457_ ), .ZN(_00666_ ) );
OAI21_X1 _15892_ ( .A(_00479_ ), .B1(_00666_ ), .B2(_00663_ ), .ZN(_00667_ ) );
OR3_X1 _15893_ ( .A1(_07115_ ), .A2(_03156_ ), .A3(_00478_ ), .ZN(_00668_ ) );
AOI21_X1 _15894_ ( .A(_00475_ ), .B1(_00667_ ), .B2(_00668_ ), .ZN(_00669_ ) );
INV_X1 _15895_ ( .A(_00666_ ), .ZN(_00670_ ) );
INV_X1 _15896_ ( .A(_00663_ ), .ZN(_00671_ ) );
AOI21_X1 _15897_ ( .A(_00464_ ), .B1(_00670_ ), .B2(_00671_ ), .ZN(_00672_ ) );
OAI21_X1 _15898_ ( .A(_00524_ ), .B1(_00669_ ), .B2(_00672_ ), .ZN(_00673_ ) );
AND2_X1 _15899_ ( .A1(_00665_ ), .A2(_00673_ ), .ZN(_00674_ ) );
OAI21_X1 _15900_ ( .A(_00664_ ), .B1(_00674_ ), .B2(_00518_ ), .ZN(_00675_ ) );
MUX2_X1 _15901_ ( .A(\EX_LS_result_reg [0] ), .B(_00675_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
NOR3_X1 _15902_ ( .A1(_00536_ ), .A2(_03157_ ), .A3(_00519_ ), .ZN(_00676_ ) );
OAI21_X1 _15903_ ( .A(_00473_ ), .B1(_00475_ ), .B2(_00676_ ), .ZN(_00677_ ) );
OAI21_X1 _15904_ ( .A(_00677_ ), .B1(_00500_ ), .B2(_00492_ ), .ZN(_00678_ ) );
MUX2_X1 _15905_ ( .A(\EX_LS_result_reg [28] ), .B(_00678_ ), .S(fanout_net_43 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
NOR3_X1 _15906_ ( .A1(_00543_ ), .A2(_03158_ ), .A3(_00519_ ), .ZN(_00679_ ) );
OAI21_X1 _15907_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00679_ ), .ZN(_00680_ ) );
AOI22_X1 _15908_ ( .A1(_00680_ ), .A2(_00496_ ), .B1(_00359_ ), .B2(_04503_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
NOR3_X1 _15909_ ( .A1(_00547_ ), .A2(_03157_ ), .A3(_00519_ ), .ZN(_00681_ ) );
OAI21_X1 _15910_ ( .A(_00473_ ), .B1(_00475_ ), .B2(_00681_ ), .ZN(_00682_ ) );
OAI21_X1 _15911_ ( .A(_00682_ ), .B1(_00500_ ), .B2(_00492_ ), .ZN(_00683_ ) );
MUX2_X1 _15912_ ( .A(\EX_LS_result_reg [26] ), .B(_00683_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
NOR3_X1 _15913_ ( .A1(_00551_ ), .A2(_03158_ ), .A3(_00519_ ), .ZN(_00684_ ) );
OAI21_X1 _15914_ ( .A(_00474_ ), .B1(_00476_ ), .B2(_00684_ ), .ZN(_00685_ ) );
AOI22_X1 _15915_ ( .A1(_00685_ ), .A2(_00496_ ), .B1(_00359_ ), .B2(_04572_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
NOR3_X1 _15916_ ( .A1(_00555_ ), .A2(_03157_ ), .A3(_00519_ ), .ZN(_00686_ ) );
OAI21_X1 _15917_ ( .A(_00473_ ), .B1(_00475_ ), .B2(_00686_ ), .ZN(_00687_ ) );
OAI21_X1 _15918_ ( .A(_00687_ ), .B1(_00494_ ), .B2(_00492_ ), .ZN(_00688_ ) );
MUX2_X1 _15919_ ( .A(\EX_LS_result_reg [24] ), .B(_00688_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _15920_ ( .A1(_07130_ ), .A2(_03157_ ), .A3(_00519_ ), .ZN(_00689_ ) );
OAI21_X1 _15921_ ( .A(_00473_ ), .B1(_00475_ ), .B2(_00689_ ), .ZN(_00690_ ) );
OAI21_X1 _15922_ ( .A(_00690_ ), .B1(_00494_ ), .B2(_00492_ ), .ZN(_00691_ ) );
MUX2_X1 _15923_ ( .A(\EX_LS_result_reg [23] ), .B(_00691_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _15924_ ( .A1(_07131_ ), .A2(\io_master_arid [1] ), .A3(_07133_ ), .ZN(_00692_ ) );
NOR2_X1 _15925_ ( .A1(_00692_ ), .A2(_00479_ ), .ZN(_00693_ ) );
OAI21_X1 _15926_ ( .A(_00473_ ), .B1(_00475_ ), .B2(_00693_ ), .ZN(_00694_ ) );
OAI21_X1 _15927_ ( .A(_00694_ ), .B1(_00494_ ), .B2(_00492_ ), .ZN(_00695_ ) );
MUX2_X1 _15928_ ( .A(\EX_LS_result_reg [22] ), .B(_00695_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
OAI211_X1 _15929_ ( .A(_07033_ ), .B(\io_master_arid [1] ), .C1(_00466_ ), .C2(_00468_ ), .ZN(_00696_ ) );
AOI21_X1 _15930_ ( .A(_00465_ ), .B1(_00464_ ), .B2(_00696_ ), .ZN(_00697_ ) );
NAND3_X1 _15931_ ( .A1(_00697_ ), .A2(_00493_ ), .A3(_00524_ ), .ZN(_00698_ ) );
OAI21_X1 _15932_ ( .A(_00698_ ), .B1(_00494_ ), .B2(_00492_ ), .ZN(_00699_ ) );
MUX2_X1 _15933_ ( .A(\EX_LS_result_reg [31] ), .B(_00699_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR4_X1 _15934_ ( .A1(_01346_ ), .A2(_03077_ ), .A3(_00391_ ), .A4(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
CLKBUF_X1 _15935_ ( .A(fanout_net_4 ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
INV_X1 _15936_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_00700_ ) );
NOR2_X1 _15937_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(\LS_WB_waddr_reg [0] ), .ZN(_00701_ ) );
INV_X1 _15938_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_00702_ ) );
INV_X1 _15939_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_00703_ ) );
NAND3_X1 _15940_ ( .A1(_00701_ ), .A2(_00702_ ), .A3(_00703_ ), .ZN(_00704_ ) );
AND2_X1 _15941_ ( .A1(_00731_ ), .A2(LS_WB_wen_reg ), .ZN(_00705_ ) );
NAND2_X1 _15942_ ( .A1(_00704_ ), .A2(_00705_ ), .ZN(_00706_ ) );
BUF_X4 _15943_ ( .A(_00706_ ), .Z(_00707_ ) );
NOR2_X1 _15944_ ( .A1(_00707_ ), .A2(_00702_ ), .ZN(_00708_ ) );
INV_X1 _15945_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_00709_ ) );
NOR2_X1 _15946_ ( .A1(_00706_ ), .A2(_00709_ ), .ZN(_00710_ ) );
AND4_X1 _15947_ ( .A1(_00700_ ), .A2(_00708_ ), .A3(_00710_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
AOI21_X1 _15948_ ( .A(_00707_ ), .B1(_00700_ ), .B2(_00702_ ), .ZN(_00711_ ) );
NOR4_X1 _15949_ ( .A1(_00711_ ), .A2(_00710_ ), .A3(_00703_ ), .A4(_00707_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR2_X1 _15950_ ( .A1(_00707_ ), .A2(_00703_ ), .ZN(_00712_ ) );
NOR4_X1 _15951_ ( .A1(_00711_ ), .A2(_00712_ ), .A3(_00709_ ), .A4(_00707_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
NOR4_X1 _15952_ ( .A1(_00711_ ), .A2(_00703_ ), .A3(_00709_ ), .A4(_00707_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
AOI21_X1 _15953_ ( .A(_00707_ ), .B1(_00703_ ), .B2(_00709_ ), .ZN(_00713_ ) );
NOR2_X1 _15954_ ( .A1(_00706_ ), .A2(_00700_ ), .ZN(_00714_ ) );
NOR4_X1 _15955_ ( .A1(_00713_ ), .A2(_00714_ ), .A3(_00702_ ), .A4(_00707_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
AND4_X1 _15956_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_00714_ ), .A3(_00712_ ), .A4(_00709_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _15957_ ( .A1(_00700_ ), .A2(_00708_ ), .A3(_00712_ ), .A4(_00709_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
NOR4_X1 _15958_ ( .A1(_00713_ ), .A2(_00708_ ), .A3(_00700_ ), .A4(_00707_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
AND4_X1 _15959_ ( .A1(_00702_ ), .A2(_00714_ ), .A3(_00710_ ), .A4(_00703_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _15960_ ( .A1(_00700_ ), .A2(_00708_ ), .A3(_00710_ ), .A4(_00703_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _15961_ ( .A1(_00702_ ), .A2(_00714_ ), .A3(_00712_ ), .A4(_00709_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _15962_ ( .A1(_00702_ ), .A2(_00714_ ), .A3(_00710_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
NOR4_X1 _15963_ ( .A1(_00713_ ), .A2(_00700_ ), .A3(_00702_ ), .A4(_00707_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _15964_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_00714_ ), .A3(_00710_ ), .A4(_00703_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
AND4_X1 _15965_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_00714_ ), .A3(_00712_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _15966_ ( .A1(_01204_ ), .A2(_00841_ ), .A3(_01213_ ), .ZN(_00715_ ) );
NAND2_X1 _15967_ ( .A1(_00715_ ), .A2(_00841_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _15968_ ( .A(fanout_net_4 ), .B(_01204_ ), .C1(_01205_ ), .C2(_01239_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _15969_ ( .A(_00704_ ), .Z(_00716_ ) );
CLKBUF_X2 _15970_ ( .A(_00705_ ), .Z(_00717_ ) );
AND3_X1 _15971_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _15972_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _15973_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _15974_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _15975_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _15976_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _15977_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _15978_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _15979_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _15980_ ( .A1(_00716_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_00717_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _15981_ ( .A(_00704_ ), .Z(_00718_ ) );
CLKBUF_X2 _15982_ ( .A(_00705_ ), .Z(_00719_ ) );
AND3_X1 _15983_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _15984_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _15985_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _15986_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _15987_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _15988_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _15989_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _15990_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _15991_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _15992_ ( .A1(_00718_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_00719_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _15993_ ( .A(_00704_ ), .Z(_00720_ ) );
CLKBUF_X2 _15994_ ( .A(_00705_ ), .Z(_00721_ ) );
AND3_X1 _15995_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _15996_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _15997_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _15998_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _15999_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _16000_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _16001_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _16002_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _16003_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _16004_ ( .A1(_00720_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_00721_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _16005_ ( .A1(_00704_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_00705_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _16006_ ( .A1(_00704_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_00705_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_D ) );
AND3_X1 _16007_ ( .A1(_00841_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _16008_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_00722_ ) );
AND2_X1 _16009_ ( .A1(_00722_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_00723_ ) );
INV_X1 _16010_ ( .A(_00723_ ), .ZN(_00724_ ) );
NOR2_X1 _16011_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_00725_ ) );
OAI211_X1 _16012_ ( .A(_00731_ ), .B(\mysc.state [0] ), .C1(_00724_ ), .C2(_00725_ ), .ZN(_00726_ ) );
INV_X1 _16013_ ( .A(_00726_ ), .ZN(_00727_ ) );
OR3_X1 _16014_ ( .A1(_00727_ ), .A2(fanout_net_4 ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _16015_ ( .A1(_00724_ ), .A2(fanout_net_4 ), .A3(_00725_ ), .ZN(_00728_ ) );
NAND2_X1 _16016_ ( .A1(_00728_ ), .A2(\mysc.state [0] ), .ZN(_00729_ ) );
OR3_X1 _16017_ ( .A1(_03150_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_00730_ ) );
NAND2_X1 _16018_ ( .A1(_00729_ ), .A2(_00730_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _16019_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07329_ ) );
CLKGATE_X1 _16020_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07330_ ) );
CLKGATE_X1 _16021_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07331_ ) );
CLKGATE_X1 _16022_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07332_ ) );
CLKGATE_X1 _16023_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07333_ ) );
CLKGATE_X1 _16024_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07334_ ) );
CLKGATE_X1 _16025_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_07335_ ) );
CLKGATE_X1 _16026_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_07336_ ) );
CLKGATE_X1 _16027_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_07337_ ) );
CLKGATE_X1 _16028_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07338_ ) );
CLKGATE_X1 _16029_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_07339_ ) );
CLKGATE_X1 _16030_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_07340_ ) );
CLKGATE_X1 _16031_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_07341_ ) );
CLKGATE_X1 _16032_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_07342_ ) );
CLKGATE_X1 _16033_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07343_ ) );
CLKGATE_X1 _16034_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07344_ ) );
CLKGATE_X1 _16035_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_07345_ ) );
CLKGATE_X1 _16036_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_07346_ ) );
CLKGATE_X1 _16037_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_07347_ ) );
CLKGATE_X1 _16038_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ), .GCK(_07348_ ) );
CLKGATE_X1 _16039_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .GCK(_07349_ ) );
CLKGATE_X1 _16040_ ( .CK(clock ), .E(io_master_wready_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ), .GCK(_07350_ ) );
CLKGATE_X1 _16041_ ( .CK(clock ), .E(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_07351_ ) );
CLKGATE_X1 _16042_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_07352_ ) );
CLKGATE_X1 _16043_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_30_E ), .GCK(_07353_ ) );
CLKGATE_X1 _16044_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_07354_ ) );
CLKGATE_X1 _16045_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_07355_ ) );
CLKGATE_X1 _16046_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_07356_ ) );
CLKGATE_X1 _16047_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_07357_ ) );
CLKGATE_X1 _16048_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_07358_ ) );
CLKGATE_X1 _16049_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07359_ ) );
CLKGATE_X1 _16050_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07360_ ) );
CLKGATE_X1 _16051_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07361_ ) );
CLKGATE_X1 _16052_ ( .CK(clock ), .E(\myexu.check_quest_$_NAND__B_A_$_ORNOT__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_AND__A_Y ), .GCK(_07362_ ) );
CLKGATE_X1 _16053_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E_$_ANDNOT__Y_B_$_ANDNOT__B_Y_$_ANDNOT__A_Y ), .GCK(_07363_ ) );
CLKGATE_X1 _16054_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_07364_ ) );
CLKGATE_X1 _16055_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_07365_ ) );
CLKGATE_X1 _16056_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_07366_ ) );
CLKGATE_X1 _16057_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_07367_ ) );
CLKGATE_X1 _16058_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07368_ ) );
CLKGATE_X1 _16059_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07369_ ) );
CLKGATE_X1 _16060_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07370_ ) );
CLKGATE_X1 _16061_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_07371_ ) );
CLKGATE_X1 _16062_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07372_ ) );
CLKGATE_X1 _16063_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_07373_ ) );
CLKGATE_X1 _16064_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_07374_ ) );
CLKGATE_X1 _16065_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_B_$_OR__B_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07375_ ) );
CLKGATE_X1 _16066_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_07376_ ) );
CLKGATE_X1 _16067_ ( .CK(clock ), .E(\myexu.state_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_07377_ ) );
CLKGATE_X1 _16068_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_07378_ ) );
CLKGATE_X1 _16069_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07379_ ) );
CLKGATE_X1 _16070_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__B_Y_$_ORNOT__B_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07380_ ) );
CLKGATE_X1 _16071_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ), .GCK(_07381_ ) );
CLKGATE_X1 _16072_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ), .GCK(_07382_ ) );
CLKGATE_X1 _16073_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07383_ ) );
LOGIC1_X1 _16074_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _16075_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00000_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00064_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_07584_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_07585_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_07586_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_07587_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_07588_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_07589_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_07590_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_07591_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_07592_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_07593_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_07594_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_07595_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_07596_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_07597_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_07598_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_07599_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_07600_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_07601_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_07602_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_07603_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_07604_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_07605_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_07606_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_07607_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_07608_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_07609_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_07610_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_07611_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_07612_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_07613_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_07614_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07383_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_07615_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07382_ ), .Q(\mtvec [31] ), .QN(_07616_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07382_ ), .Q(\mtvec [30] ), .QN(_07617_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07382_ ), .Q(\mtvec [21] ), .QN(_07618_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07382_ ), .Q(\mtvec [20] ), .QN(_07619_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07382_ ), .Q(\mtvec [19] ), .QN(_07620_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07382_ ), .Q(\mtvec [18] ), .QN(_07621_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07382_ ), .Q(\mtvec [17] ), .QN(_07622_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07382_ ), .Q(\mtvec [16] ), .QN(_07623_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07382_ ), .Q(\mtvec [15] ), .QN(_07624_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07382_ ), .Q(\mtvec [14] ), .QN(_07625_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07382_ ), .Q(\mtvec [13] ), .QN(_07626_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07382_ ), .Q(\mtvec [12] ), .QN(_07627_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07382_ ), .Q(\mtvec [29] ), .QN(_07628_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07382_ ), .Q(\mtvec [11] ), .QN(_07629_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07382_ ), .Q(\mtvec [10] ), .QN(_07630_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07382_ ), .Q(\mtvec [9] ), .QN(_07631_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07382_ ), .Q(\mtvec [8] ), .QN(_07632_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07382_ ), .Q(\mtvec [7] ), .QN(_07633_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07382_ ), .Q(\mtvec [6] ), .QN(_07634_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07382_ ), .Q(\mtvec [5] ), .QN(_07635_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07382_ ), .Q(\mtvec [4] ), .QN(_07636_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07382_ ), .Q(\mtvec [3] ), .QN(_07637_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07382_ ), .Q(\mtvec [2] ), .QN(_07638_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07382_ ), .Q(\mtvec [28] ), .QN(_07639_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07382_ ), .Q(\mtvec [1] ), .QN(_07640_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07382_ ), .Q(\mtvec [0] ), .QN(_07641_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07382_ ), .Q(\mtvec [27] ), .QN(_07642_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07382_ ), .Q(\mtvec [26] ), .QN(_07643_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07382_ ), .Q(\mtvec [25] ), .QN(_07644_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07382_ ), .Q(\mtvec [24] ), .QN(_07645_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07382_ ), .Q(\mtvec [23] ), .QN(_07646_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07382_ ), .Q(\mtvec [22] ), .QN(_07647_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07381_ ), .Q(\mepc [31] ), .QN(_07648_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07381_ ), .Q(\mepc [30] ), .QN(_07649_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07381_ ), .Q(\mepc [21] ), .QN(_07650_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07381_ ), .Q(\mepc [20] ), .QN(_07651_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07381_ ), .Q(\mepc [19] ), .QN(_07652_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07381_ ), .Q(\mepc [18] ), .QN(_07653_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07381_ ), .Q(\mepc [17] ), .QN(_07654_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07381_ ), .Q(\mepc [16] ), .QN(_07655_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07381_ ), .Q(\mepc [15] ), .QN(_07656_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07381_ ), .Q(\mepc [14] ), .QN(_07657_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07381_ ), .Q(\mepc [13] ), .QN(_07658_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07381_ ), .Q(\mepc [12] ), .QN(_07659_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07381_ ), .Q(\mepc [29] ), .QN(_07660_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07381_ ), .Q(\mepc [11] ), .QN(_07661_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07381_ ), .Q(\mepc [10] ), .QN(_07662_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07381_ ), .Q(\mepc [9] ), .QN(_07663_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07381_ ), .Q(\mepc [8] ), .QN(_07664_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07381_ ), .Q(\mepc [7] ), .QN(_07665_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07381_ ), .Q(\mepc [6] ), .QN(_07666_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07381_ ), .Q(\mepc [5] ), .QN(_07667_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07381_ ), .Q(\mepc [4] ), .QN(_07668_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07381_ ), .Q(\mepc [3] ), .QN(_07669_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07381_ ), .Q(\mepc [2] ), .QN(_07670_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07381_ ), .Q(\mepc [28] ), .QN(_07671_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07381_ ), .Q(\mepc [1] ), .QN(_07672_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07381_ ), .Q(\mepc [0] ), .QN(_07673_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07381_ ), .Q(\mepc [27] ), .QN(_07674_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07381_ ), .Q(\mepc [26] ), .QN(_07675_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07381_ ), .Q(\mepc [25] ), .QN(_07676_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07381_ ), .Q(\mepc [24] ), .QN(_07677_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07381_ ), .Q(\mepc [23] ), .QN(_07678_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07381_ ), .Q(\mepc [22] ), .QN(_07679_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_07680_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_07681_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_07682_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_07583_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00065_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_07582_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00066_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_07581_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00067_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_07580_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00068_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_07579_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00069_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_07578_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00070_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_07577_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00071_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_07576_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00072_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_07575_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00073_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_07574_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00074_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_07573_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00075_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_07572_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00076_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_07571_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00077_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_07570_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00078_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_07569_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00079_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_07568_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00080_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_07567_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00081_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_07566_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00082_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_07565_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00083_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_07564_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00084_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_07563_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00085_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_07562_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00086_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_07561_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00087_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_07560_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00088_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_07559_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00089_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_07558_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00090_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_07557_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00091_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_07556_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00092_ ), .CK(_07380_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_07683_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PN0__Q ( .D(_00093_ ), .CK(clock ), .Q(excp_written ), .QN(_07684_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [31] ), .QN(_07555_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [30] ), .QN(_07685_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [21] ), .QN(_07686_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [20] ), .QN(_07687_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [19] ), .QN(_07688_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [18] ), .QN(_07689_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [17] ), .QN(_07690_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [16] ), .QN(_07691_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [15] ), .QN(_07692_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [14] ), .QN(_07693_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [13] ), .QN(_07694_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [12] ), .QN(_07695_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [29] ), .QN(_07696_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [11] ), .QN(_07697_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [10] ), .QN(_07698_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [9] ), .QN(_07699_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [8] ), .QN(_07700_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [7] ), .QN(_07701_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [6] ), .QN(_07702_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [5] ), .QN(_07703_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [4] ), .QN(_07704_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [3] ), .QN(_07705_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [2] ), .QN(_07706_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [28] ), .QN(_07707_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [1] ), .QN(_07708_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [0] ), .QN(_07709_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [27] ), .QN(_07710_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [26] ), .QN(_07711_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [25] ), .QN(_07712_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [24] ), .QN(_07713_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [23] ), .QN(_07714_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_07379_ ), .Q(\myec.mepc_tmp [22] ), .QN(_07554_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00094_ ), .CK(_07378_ ), .Q(\myec.state [1] ), .QN(_07553_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00095_ ), .CK(_07378_ ), .Q(\myec.state [0] ), .QN(_07715_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PP0__Q ( .D(_00096_ ), .CK(clock ), .Q(check_quest ), .QN(_07716_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_07552_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_07717_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_07718_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_07719_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_07720_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_07721_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_07722_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_07723_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_07724_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_07725_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_07726_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_07551_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00097_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_07550_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00098_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_07549_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00099_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_07548_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00100_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_07547_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00101_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_07546_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00102_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_07545_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00103_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_07544_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00104_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_07543_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00105_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_07542_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00106_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_07541_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00107_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_07540_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00108_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_07539_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00109_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_07538_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00110_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_07537_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00111_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_07536_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00112_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_07535_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00113_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_07534_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00114_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_07533_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00115_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_07532_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00116_ ), .CK(_07377_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_07531_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q ( .D(_00117_ ), .CK(_07376_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_07530_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_1 ( .D(_00118_ ), .CK(_07376_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_07529_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_2 ( .D(_00119_ ), .CK(_07376_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_07528_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_3 ( .D(_00120_ ), .CK(_07376_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_07527_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PP0P__Q_4 ( .D(_00121_ ), .CK(_07376_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_07526_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q ( .D(_00122_ ), .CK(_07376_ ), .Q(\EX_LS_pc [31] ), .QN(_07525_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_1 ( .D(_00123_ ), .CK(_07376_ ), .Q(\EX_LS_pc [30] ), .QN(_07524_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_10 ( .D(_00124_ ), .CK(_07376_ ), .Q(\EX_LS_pc [21] ), .QN(_07523_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_11 ( .D(_00125_ ), .CK(_07376_ ), .Q(\EX_LS_pc [20] ), .QN(_07522_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_12 ( .D(_00126_ ), .CK(_07376_ ), .Q(\EX_LS_pc [19] ), .QN(_07521_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_13 ( .D(_00127_ ), .CK(_07376_ ), .Q(\EX_LS_pc [18] ), .QN(_07520_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_14 ( .D(_00128_ ), .CK(_07376_ ), .Q(\EX_LS_pc [17] ), .QN(_07519_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_15 ( .D(_00129_ ), .CK(_07376_ ), .Q(\EX_LS_pc [16] ), .QN(_07518_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_16 ( .D(_00130_ ), .CK(_07376_ ), .Q(\EX_LS_pc [15] ), .QN(_07517_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_17 ( .D(_00131_ ), .CK(_07376_ ), .Q(\EX_LS_pc [14] ), .QN(_07516_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_18 ( .D(_00132_ ), .CK(_07376_ ), .Q(\EX_LS_pc [13] ), .QN(_07515_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_19 ( .D(_00133_ ), .CK(_07376_ ), .Q(\EX_LS_pc [12] ), .QN(_07514_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_2 ( .D(_00134_ ), .CK(_07376_ ), .Q(\EX_LS_pc [29] ), .QN(_07513_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_20 ( .D(_00135_ ), .CK(_07376_ ), .Q(\EX_LS_pc [11] ), .QN(_07512_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_21 ( .D(_00136_ ), .CK(_07376_ ), .Q(\EX_LS_pc [10] ), .QN(_07511_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_22 ( .D(_00137_ ), .CK(_07376_ ), .Q(\EX_LS_pc [9] ), .QN(_07510_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_23 ( .D(_00138_ ), .CK(_07376_ ), .Q(\EX_LS_pc [8] ), .QN(_07509_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_24 ( .D(_00139_ ), .CK(_07376_ ), .Q(\EX_LS_pc [7] ), .QN(_07508_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_25 ( .D(_00140_ ), .CK(_07376_ ), .Q(\EX_LS_pc [6] ), .QN(_07507_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_26 ( .D(_00141_ ), .CK(_07376_ ), .Q(\EX_LS_pc [5] ), .QN(_07506_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_27 ( .D(_00142_ ), .CK(_07376_ ), .Q(\EX_LS_pc [4] ), .QN(_07505_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_28 ( .D(_00143_ ), .CK(_07376_ ), .Q(\EX_LS_pc [3] ), .QN(_07504_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_29 ( .D(_00144_ ), .CK(_07376_ ), .Q(\EX_LS_pc [2] ), .QN(_07503_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_3 ( .D(_00145_ ), .CK(_07376_ ), .Q(\EX_LS_pc [28] ), .QN(_07502_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_30 ( .D(_00146_ ), .CK(_07376_ ), .Q(\EX_LS_pc [1] ), .QN(_07501_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_31 ( .D(_00147_ ), .CK(_07376_ ), .Q(\EX_LS_pc [0] ), .QN(_07500_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_4 ( .D(_00148_ ), .CK(_07376_ ), .Q(\EX_LS_pc [27] ), .QN(_07499_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_5 ( .D(_00149_ ), .CK(_07376_ ), .Q(\EX_LS_pc [26] ), .QN(_07498_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_6 ( .D(_00150_ ), .CK(_07376_ ), .Q(\EX_LS_pc [25] ), .QN(_07497_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_7 ( .D(_00151_ ), .CK(_07376_ ), .Q(\EX_LS_pc [24] ), .QN(_07496_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_8 ( .D(_00152_ ), .CK(_07376_ ), .Q(\EX_LS_pc [23] ), .QN(_07495_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PP0P__Q_9 ( .D(_00153_ ), .CK(_07376_ ), .Q(\EX_LS_pc [22] ), .QN(_07727_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_07728_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_07729_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_07730_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_07731_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_07732_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_07733_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_07734_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_07735_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_07736_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_07737_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_07738_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_07739_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_07740_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_07741_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_07742_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_07743_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_07744_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_07745_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_07746_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_07747_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_07748_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_07749_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_07750_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_07751_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_07752_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_07753_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_07754_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_07755_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_07756_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_07757_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_07758_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07377_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_07759_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_07377_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PP0__Q ( .D(_00155_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q ( .D(_00154_ ), .CK(_07376_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_1 ( .D(_00156_ ), .CK(_07376_ ), .Q(\EX_LS_flag [1] ), .QN(_07494_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_2 ( .D(_00157_ ), .CK(_07376_ ), .Q(\EX_LS_flag [0] ), .QN(_07493_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_3 ( .D(_00158_ ), .CK(_07376_ ), .Q(\EX_LS_typ [4] ), .QN(_07492_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_4 ( .D(_00159_ ), .CK(_07376_ ), .Q(\EX_LS_typ [3] ), .QN(_07491_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_5 ( .D(_00160_ ), .CK(_07376_ ), .Q(\EX_LS_typ [2] ), .QN(_07490_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_6 ( .D(_00161_ ), .CK(_07376_ ), .Q(\EX_LS_typ [1] ), .QN(_07489_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PP0P__Q_7 ( .D(_00162_ ), .CK(_07376_ ), .Q(\EX_LS_typ [0] ), .QN(_07488_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00163_ ), .CK(_07375_ ), .Q(\ID_EX_csr [11] ), .QN(_07487_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00164_ ), .CK(_07375_ ), .Q(\ID_EX_csr [10] ), .QN(_07486_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00165_ ), .CK(_07375_ ), .Q(\ID_EX_csr [1] ), .QN(_07485_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00166_ ), .CK(_07375_ ), .Q(\ID_EX_csr [0] ), .QN(_07484_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00167_ ), .CK(_07375_ ), .Q(\ID_EX_csr [9] ), .QN(_07483_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00168_ ), .CK(_07375_ ), .Q(\ID_EX_csr [8] ), .QN(_07482_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00169_ ), .CK(_07375_ ), .Q(\ID_EX_csr [7] ), .QN(_07481_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00170_ ), .CK(_07375_ ), .Q(\ID_EX_csr [6] ), .QN(_07480_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00171_ ), .CK(_07375_ ), .Q(\ID_EX_csr [5] ), .QN(_07479_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00172_ ), .CK(_07375_ ), .Q(\ID_EX_csr [4] ), .QN(_07478_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00173_ ), .CK(_07375_ ), .Q(\ID_EX_csr [3] ), .QN(_07477_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00174_ ), .CK(_07375_ ), .Q(\ID_EX_csr [2] ), .QN(_07476_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00175_ ), .CK(_07374_ ), .Q(exception_quest_IDU ), .QN(_07475_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00176_ ), .CK(_07373_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_07372_ ), .Q(\ID_EX_imm [31] ), .QN(_07760_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_07372_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_07372_ ), .Q(\ID_EX_imm [21] ), .QN(_07761_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_07372_ ), .Q(\ID_EX_imm [20] ), .QN(_07762_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_07372_ ), .Q(\ID_EX_imm [19] ), .QN(_07763_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_07372_ ), .Q(\ID_EX_imm [18] ), .QN(_07764_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_07372_ ), .Q(\ID_EX_imm [17] ), .QN(_07765_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_07372_ ), .Q(\ID_EX_imm [16] ), .QN(_07766_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_07372_ ), .Q(\ID_EX_imm [15] ), .QN(_07767_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_07372_ ), .Q(\ID_EX_imm [14] ), .QN(_07768_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_07372_ ), .Q(\ID_EX_imm [13] ), .QN(_07769_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_07372_ ), .Q(\ID_EX_imm [12] ), .QN(_07770_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_07372_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_07372_ ), .Q(\ID_EX_imm [11] ), .QN(_07771_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_07372_ ), .Q(\ID_EX_imm [10] ), .QN(_07772_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_07372_ ), .Q(\ID_EX_imm [9] ), .QN(_07773_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_07372_ ), .Q(\ID_EX_imm [8] ), .QN(_07774_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_07372_ ), .Q(\ID_EX_imm [7] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__B_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_07372_ ), .Q(\ID_EX_imm [6] ), .QN(_07775_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_07372_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_07372_ ), .Q(\ID_EX_imm [4] ), .QN(_07776_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_07372_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_07372_ ), .Q(\ID_EX_imm [2] ), .QN(_07777_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_07372_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_07372_ ), .Q(\ID_EX_imm [1] ), .QN(_07778_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_07372_ ), .Q(\ID_EX_imm [0] ), .QN(_07779_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_07372_ ), .Q(\ID_EX_imm [27] ), .QN(_07780_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_07372_ ), .Q(\ID_EX_imm [26] ), .QN(_07781_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_07372_ ), .Q(\ID_EX_imm [25] ), .QN(_07782_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_07372_ ), .Q(\ID_EX_imm [24] ), .QN(_07783_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_07372_ ), .Q(\ID_EX_imm [23] ), .QN(_07784_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_07372_ ), .Q(\ID_EX_imm [22] ), .QN(_07785_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07371_ ), .Q(\ID_EX_pc [31] ), .QN(_07786_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07371_ ), .Q(\ID_EX_pc [30] ), .QN(_07787_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07371_ ), .Q(\ID_EX_pc [21] ), .QN(_07788_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07371_ ), .Q(\ID_EX_pc [20] ), .QN(_07789_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07371_ ), .Q(\ID_EX_pc [19] ), .QN(_07790_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07371_ ), .Q(\ID_EX_pc [18] ), .QN(_07791_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07371_ ), .Q(\ID_EX_pc [17] ), .QN(_07792_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07371_ ), .Q(\ID_EX_pc [16] ), .QN(_07793_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07371_ ), .Q(\ID_EX_pc [15] ), .QN(_07794_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07371_ ), .Q(\ID_EX_pc [14] ), .QN(_07795_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07371_ ), .Q(\ID_EX_pc [13] ), .QN(_07796_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07371_ ), .Q(\ID_EX_pc [12] ), .QN(_07797_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07371_ ), .Q(\ID_EX_pc [29] ), .QN(_07798_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07371_ ), .Q(\ID_EX_pc [11] ), .QN(_07799_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07371_ ), .Q(\ID_EX_pc [10] ), .QN(_07800_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07371_ ), .Q(\ID_EX_pc [9] ), .QN(_07801_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07371_ ), .Q(\ID_EX_pc [8] ), .QN(_07802_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07371_ ), .Q(\ID_EX_pc [7] ), .QN(_07803_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07371_ ), .Q(\ID_EX_pc [6] ), .QN(_07804_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07371_ ), .Q(\ID_EX_pc [5] ), .QN(_07805_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07371_ ), .Q(\ID_EX_pc [4] ), .QN(_07806_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_07371_ ), .Q(\ID_EX_pc [3] ), .QN(_07807_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_07371_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07371_ ), .Q(\ID_EX_pc [28] ), .QN(_07808_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_07371_ ), .Q(\ID_EX_pc [1] ), .QN(_07809_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_07371_ ), .Q(\ID_EX_pc [0] ), .QN(_07810_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07371_ ), .Q(\ID_EX_pc [27] ), .QN(_07811_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07371_ ), .Q(\ID_EX_pc [26] ), .QN(_07812_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07371_ ), .Q(\ID_EX_pc [25] ), .QN(_07813_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07371_ ), .Q(\ID_EX_pc [24] ), .QN(_07814_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07371_ ), .Q(\ID_EX_pc [23] ), .QN(_07815_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07371_ ), .Q(\ID_EX_pc [22] ), .QN(_07474_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00177_ ), .CK(_07370_ ), .Q(\ID_EX_rd [4] ), .QN(_07473_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00178_ ), .CK(_07370_ ), .Q(\ID_EX_rd [3] ), .QN(_07472_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00179_ ), .CK(_07370_ ), .Q(\ID_EX_rd [2] ), .QN(_07471_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00180_ ), .CK(_07370_ ), .Q(\ID_EX_rd [1] ), .QN(_07470_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00181_ ), .CK(_07370_ ), .Q(\ID_EX_rd [0] ), .QN(_07469_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00182_ ), .CK(_07369_ ), .Q(\ID_EX_rs1 [4] ), .QN(_07468_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00183_ ), .CK(_07369_ ), .Q(\ID_EX_rs1 [3] ), .QN(_07467_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00185_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_07465_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00184_ ), .CK(_07369_ ), .Q(\ID_EX_rs1 [2] ), .QN(_07466_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00187_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_07463_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00186_ ), .CK(_07369_ ), .Q(\ID_EX_rs1 [1] ), .QN(_07464_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00189_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_07461_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00188_ ), .CK(_07369_ ), .Q(\ID_EX_rs1 [0] ), .QN(_07462_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00191_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_07459_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00190_ ), .CK(_07368_ ), .Q(\ID_EX_rs2 [4] ), .QN(_07460_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00192_ ), .CK(_07368_ ), .Q(\ID_EX_rs2 [3] ), .QN(_07458_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00194_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_07456_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00193_ ), .CK(_07368_ ), .Q(\ID_EX_rs2 [2] ), .QN(_07457_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00196_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_07454_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00195_ ), .CK(_07368_ ), .Q(\ID_EX_rs2 [1] ), .QN(_07455_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00198_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_07452_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00197_ ), .CK(_07368_ ), .Q(\ID_EX_rs2 [0] ), .QN(_07453_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00200_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_07450_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00199_ ), .CK(_07367_ ), .Q(\myidu.stall_quest_fencei ), .QN(_07451_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00201_ ), .CK(_07366_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_07449_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_07817_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00202_ ), .CK(_07365_ ), .Q(\ID_EX_typ [7] ), .QN(_07816_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00203_ ), .CK(_07365_ ), .Q(\ID_EX_typ [6] ), .QN(_07448_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00204_ ), .CK(_07365_ ), .Q(\ID_EX_typ [5] ), .QN(_07447_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00205_ ), .CK(_07365_ ), .Q(\ID_EX_typ [4] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00206_ ), .CK(_07365_ ), .Q(\ID_EX_typ [3] ), .QN(_07446_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00207_ ), .CK(_07365_ ), .Q(\ID_EX_typ [2] ), .QN(\myifu.check_assert_$_ANDNOT__B_Y_$_MUX__A_B_$_OR__B_A_$_OR__Y_B_$_ANDNOT__B_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00208_ ), .CK(_07365_ ), .Q(\ID_EX_typ [1] ), .QN(_07445_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00209_ ), .CK(_07365_ ), .Q(\ID_EX_typ [0] ), .QN(_07818_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_07364_ ), .Q(check_assert ), .QN(_07819_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_07363_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_07363_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_07363_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_07363_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_07363_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_07363_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_07363_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_07363_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_07363_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_07363_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_07363_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_07363_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_07363_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_07363_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_26_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_07363_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_07363_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_07363_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_07363_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_07363_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_07363_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_07363_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_07363_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_07363_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_07363_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_22_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ORNOT__Y_B_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_07363_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_07363_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_07363_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_07363_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_07363_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_07363_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_07363_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_07363_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_07820_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_07821_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_07822_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_07823_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_07824_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_07825_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_07826_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_07827_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_07828_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_07829_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_07830_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_07831_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_07832_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_07833_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_07834_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_07835_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_07836_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_07837_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_07838_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_07839_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_07840_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_07841_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_07842_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_07843_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_07844_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_07845_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_07846_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_07847_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_07848_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_07849_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_07850_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07362_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_07851_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_07852_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_07853_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_07854_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_07855_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_07856_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_07857_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_07858_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_07859_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_07860_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_07861_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_07862_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_07863_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_07864_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_07865_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_07866_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_07867_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_07868_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_07869_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_07870_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_07871_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_07872_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_07873_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_07874_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_07875_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_07876_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_07877_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_07878_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_07879_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_07880_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_07881_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_07882_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07361_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_07883_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_07884_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_07885_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_07886_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_07887_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_07888_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_07889_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_07890_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_07891_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_07892_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_07893_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_07894_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_07895_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_07896_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_07897_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_07898_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_07899_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_07900_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_07901_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_07902_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_07903_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_07904_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_07905_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_07906_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_07907_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_07908_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_07909_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_07910_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_07911_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_07912_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_07913_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_07914_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07360_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_07915_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_07916_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_07917_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_07918_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_07919_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_07920_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_07921_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_07922_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_07923_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_07924_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_07925_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_07926_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_07927_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_07928_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_07929_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_07930_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_07931_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_07932_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_07933_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_07934_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_07935_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_07936_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_07937_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_07938_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_07939_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_07940_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_07941_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_07942_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_07943_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_07944_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_07945_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_07946_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07359_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_07947_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][27] ), .QN(_07948_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_07949_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_07950_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_07951_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_07952_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_07953_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_07954_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_07955_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_07956_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_07957_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_07958_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_07959_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_07960_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_07961_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_07962_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_07963_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_07964_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_07965_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_07966_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_07967_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_07968_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_07969_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_07970_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_07971_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_07972_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_07973_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_07974_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07362_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_07975_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][27] ), .QN(_07976_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_07977_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_07978_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_07979_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_07980_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_07981_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_07982_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_07983_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_07984_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_07985_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_07986_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_07987_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_07988_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_07989_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_07990_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_07991_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_07992_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_07993_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_07994_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_07995_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_07996_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_07997_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_07998_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_07999_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08000_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08001_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08002_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07361_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08003_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][27] ), .QN(_08004_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08005_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08006_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08007_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08008_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08009_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08010_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08011_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08012_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08013_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08014_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08015_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08016_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08017_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08018_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08019_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08020_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08021_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08022_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08023_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08024_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08025_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08026_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08027_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08028_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08029_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08030_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07360_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08031_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][27] ), .QN(_08032_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08033_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08034_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08035_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08036_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08037_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08038_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08039_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08040_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08041_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08042_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08043_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08044_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08045_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08046_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08047_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08048_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08049_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08050_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08051_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08052_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08053_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08054_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08055_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08056_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08057_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08058_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07359_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_07444_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00210_ ), .CK(_07358_ ), .Q(\myifu.myicache.valid [0] ), .QN(_07443_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00211_ ), .CK(_07357_ ), .Q(\myifu.myicache.valid [1] ), .QN(_07442_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00212_ ), .CK(_07356_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08059_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_07355_ ), .Q(\myifu.myicache.valid [3] ), .QN(_07441_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00213_ ), .CK(_07354_ ), .Q(\IF_ID_pc [30] ), .QN(_07440_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00214_ ), .CK(_07354_ ), .Q(\IF_ID_pc [29] ), .QN(_07439_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00215_ ), .CK(_07354_ ), .Q(\IF_ID_pc [20] ), .QN(_07438_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00216_ ), .CK(_07354_ ), .Q(\IF_ID_pc [19] ), .QN(_07437_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00217_ ), .CK(_07354_ ), .Q(\IF_ID_pc [18] ), .QN(_07436_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00218_ ), .CK(_07354_ ), .Q(\IF_ID_pc [17] ), .QN(_07435_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00219_ ), .CK(_07354_ ), .Q(\IF_ID_pc [16] ), .QN(_07434_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00220_ ), .CK(_07354_ ), .Q(\IF_ID_pc [15] ), .QN(_07433_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00221_ ), .CK(_07354_ ), .Q(\IF_ID_pc [14] ), .QN(_07432_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00222_ ), .CK(_07354_ ), .Q(\IF_ID_pc [13] ), .QN(_07431_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00223_ ), .CK(_07354_ ), .Q(\IF_ID_pc [12] ), .QN(_07430_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00224_ ), .CK(_07354_ ), .Q(\IF_ID_pc [11] ), .QN(_07429_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00225_ ), .CK(_07354_ ), .Q(\IF_ID_pc [28] ), .QN(_07428_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00226_ ), .CK(_07354_ ), .Q(\IF_ID_pc [10] ), .QN(_07427_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00227_ ), .CK(_07354_ ), .Q(\IF_ID_pc [9] ), .QN(_07426_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00228_ ), .CK(_07354_ ), .Q(\IF_ID_pc [8] ), .QN(_07425_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00229_ ), .CK(_07354_ ), .Q(\IF_ID_pc [7] ), .QN(_07424_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00230_ ), .CK(_07354_ ), .Q(\IF_ID_pc [6] ), .QN(_07423_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00231_ ), .CK(_07354_ ), .Q(\IF_ID_pc [5] ), .QN(_07422_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00232_ ), .CK(_07354_ ), .Q(\IF_ID_pc [4] ), .QN(_07421_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00233_ ), .CK(_07354_ ), .Q(\IF_ID_pc [3] ), .QN(_07420_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00235_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_07418_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00234_ ), .CK(_07354_ ), .Q(\IF_ID_pc [2] ), .QN(_07419_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00237_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_07416_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00236_ ), .CK(_07354_ ), .Q(\IF_ID_pc [1] ), .QN(_07417_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00238_ ), .CK(_07354_ ), .Q(\IF_ID_pc [27] ), .QN(_07415_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00239_ ), .CK(_07353_ ), .Q(\IF_ID_pc [0] ), .QN(_07414_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00240_ ), .CK(_07354_ ), .Q(\IF_ID_pc [26] ), .QN(_07413_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00241_ ), .CK(_07354_ ), .Q(\IF_ID_pc [25] ), .QN(_07412_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00242_ ), .CK(_07354_ ), .Q(\IF_ID_pc [24] ), .QN(_07411_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00243_ ), .CK(_07354_ ), .Q(\IF_ID_pc [23] ), .QN(_07410_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00244_ ), .CK(_07354_ ), .Q(\IF_ID_pc [22] ), .QN(_07409_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00245_ ), .CK(_07354_ ), .Q(\IF_ID_pc [21] ), .QN(_07408_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00246_ ), .CK(_07354_ ), .Q(\IF_ID_pc [31] ), .QN(_07407_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_E_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_07406_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00248_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00247_ ), .CK(_07352_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08060_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08061_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08062_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08063_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08064_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08065_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08066_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08067_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08068_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08069_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08070_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08071_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08072_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08073_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08074_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08075_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08076_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08077_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08078_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08079_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08080_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08081_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08082_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08083_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08084_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08085_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08086_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08087_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08088_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08089_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08090_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08091_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07351_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08092_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08093_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08094_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08095_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08096_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08097_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08098_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08099_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08100_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08101_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08102_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08103_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08104_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08105_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08106_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08107_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08108_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08109_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08110_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08111_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08112_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08113_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08114_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08115_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08116_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08117_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08118_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08119_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08120_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08121_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08122_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08123_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07350_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_07405_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PP0P__Q ( .D(_00249_ ), .CK(_07349_ ), .Q(LS_WB_pc ), .QN(_07404_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PP0P__Q ( .D(_00250_ ), .CK(_07348_ ), .Q(\mylsu.previous_load_done ), .QN(_08124_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08125_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08126_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08127_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(io_master_wready_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_07351_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_07351_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08128_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_07351_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_07403_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00251_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_07402_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00252_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_07401_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00253_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_07400_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00254_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_07399_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00255_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_07398_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00256_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_07397_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00257_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_07396_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00258_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_07395_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00259_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_07394_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00260_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_07393_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00261_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_07392_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00262_ ), .CK(_07351_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08129_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_07351_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08130_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_07351_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08131_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_07351_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08132_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_07351_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08133_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08134_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08135_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08136_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08137_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08138_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08139_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08140_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08141_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08142_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08143_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08144_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08145_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08146_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08147_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08148_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08149_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08150_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08151_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08152_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08153_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08154_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08155_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08156_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08157_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08158_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08159_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08160_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08161_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08162_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08163_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08164_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_07351_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08165_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08166_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_08167_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_08168_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_08169_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_08170_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_08171_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_08172_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_08173_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_08174_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_08175_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_08176_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_08177_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_08178_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_08179_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_08180_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_08181_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_08182_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_08183_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_08184_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_08185_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_08186_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_08187_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_08188_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_08189_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_08190_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_08191_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_08192_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_08193_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_08194_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_08195_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_08196_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_07347_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_07391_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q ( .D(_00263_ ), .CK(_07346_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_07390_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_1 ( .D(_00264_ ), .CK(_07346_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_07389_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_2 ( .D(_00265_ ), .CK(_07346_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_07388_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_3 ( .D(_00266_ ), .CK(_07346_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_07387_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_4 ( .D(_00267_ ), .CK(_07346_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_07386_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_5 ( .D(_00268_ ), .CK(_07346_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_07385_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PP0P__Q ( .D(_00269_ ), .CK(_07346_ ), .Q(LS_WB_wen_reg ), .QN(_08197_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_08198_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_08199_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07345_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07344_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07343_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07342_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07341_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07340_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07339_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07338_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07337_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07336_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07335_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07334_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07333_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07332_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07331_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_OR__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07330_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00270_ ), .CK(_07329_ ), .Q(loaduse_clear ), .QN(_08200_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_08201_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_08202_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_07384_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\ID_EX_typ [2] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(excp_written ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myifu.state [2] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myifu.to_reset ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\mylsu.state [3] ), .Z(fanout_net_43 ) );

endmodule
