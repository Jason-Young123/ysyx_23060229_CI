//Generate the verilog at 2025-09-29T16:24:46 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire _08944_ ;
wire _08945_ ;
wire _08946_ ;
wire _08947_ ;
wire _08948_ ;
wire _08949_ ;
wire _08950_ ;
wire _08951_ ;
wire _08952_ ;
wire _08953_ ;
wire _08954_ ;
wire _08955_ ;
wire _08956_ ;
wire _08957_ ;
wire _08958_ ;
wire _08959_ ;
wire _08960_ ;
wire _08961_ ;
wire _08962_ ;
wire _08963_ ;
wire _08964_ ;
wire _08965_ ;
wire _08966_ ;
wire _08967_ ;
wire _08968_ ;
wire _08969_ ;
wire _08970_ ;
wire _08971_ ;
wire _08972_ ;
wire _08973_ ;
wire _08974_ ;
wire _08975_ ;
wire _08976_ ;
wire _08977_ ;
wire _08978_ ;
wire _08979_ ;
wire _08980_ ;
wire _08981_ ;
wire _08982_ ;
wire _08983_ ;
wire _08984_ ;
wire _08985_ ;
wire _08986_ ;
wire _08987_ ;
wire _08988_ ;
wire _08989_ ;
wire _08990_ ;
wire _08991_ ;
wire _08992_ ;
wire _08993_ ;
wire _08994_ ;
wire _08995_ ;
wire _08996_ ;
wire _08997_ ;
wire _08998_ ;
wire _08999_ ;
wire _09000_ ;
wire _09001_ ;
wire _09002_ ;
wire _09003_ ;
wire _09004_ ;
wire _09005_ ;
wire _09006_ ;
wire _09007_ ;
wire _09008_ ;
wire _09009_ ;
wire _09010_ ;
wire _09011_ ;
wire _09012_ ;
wire _09013_ ;
wire _09014_ ;
wire _09015_ ;
wire _09016_ ;
wire _09017_ ;
wire _09018_ ;
wire _09019_ ;
wire _09020_ ;
wire _09021_ ;
wire _09022_ ;
wire _09023_ ;
wire _09024_ ;
wire _09025_ ;
wire _09026_ ;
wire _09027_ ;
wire _09028_ ;
wire _09029_ ;
wire _09030_ ;
wire _09031_ ;
wire _09032_ ;
wire _09033_ ;
wire _09034_ ;
wire _09035_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.rst_logic_$_OR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__B_Y ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_ANDNOT__B_Y ;
wire \myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ;
wire \myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[4]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[5]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[6]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data[7]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[0]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[1]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[2]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.tag[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ;
wire \mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[1]_$_DFFE_PP__Q_D ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire fanout_net_45 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

INV_X1 _09036_ ( .A(\LS_WB_wdata_csreg [31] ), .ZN(_01584_ ) );
NOR2_X1 _09037_ ( .A1(_01584_ ), .A2(fanout_net_1 ), .ZN(_00000_ ) );
INV_X1 _09038_ ( .A(fanout_net_1 ), .ZN(_01585_ ) );
BUF_X4 _09039_ ( .A(_01585_ ), .Z(_01586_ ) );
BUF_X4 _09040_ ( .A(_01586_ ), .Z(_01587_ ) );
AND3_X4 _09041_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [0] ), .A3(\myclint.mtime [1] ), .ZN(_01588_ ) );
AND3_X4 _09042_ ( .A1(_01588_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01589_ ) );
AND3_X4 _09043_ ( .A1(_01589_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01590_ ) );
AND3_X4 _09044_ ( .A1(_01590_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01591_ ) );
AND3_X4 _09045_ ( .A1(_01591_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01592_ ) );
AND3_X4 _09046_ ( .A1(_01592_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01593_ ) );
AND3_X4 _09047_ ( .A1(_01593_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01594_ ) );
AND3_X4 _09048_ ( .A1(_01594_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01595_ ) );
AND3_X4 _09049_ ( .A1(_01595_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01596_ ) );
AND3_X4 _09050_ ( .A1(_01596_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01597_ ) );
AND3_X4 _09051_ ( .A1(_01597_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01598_ ) );
AND3_X4 _09052_ ( .A1(_01598_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01599_ ) );
AND3_X4 _09053_ ( .A1(_01599_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01600_ ) );
AND2_X4 _09054_ ( .A1(_01600_ ), .A2(\myclint.mtime [27] ), .ZN(_01601_ ) );
AND2_X1 _09055_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01602_ ) );
AND2_X2 _09056_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01603_ ) );
AND4_X4 _09057_ ( .A1(\myclint.mtime [33] ), .A2(_01601_ ), .A3(_01602_ ), .A4(_01603_ ), .ZN(_01604_ ) );
AND3_X4 _09058_ ( .A1(_01604_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01605_ ) );
AND2_X4 _09059_ ( .A1(_01605_ ), .A2(\myclint.mtime [35] ), .ZN(_01606_ ) );
AND2_X1 _09060_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [39] ), .ZN(_01607_ ) );
AND2_X1 _09061_ ( .A1(\myclint.mtime [36] ), .A2(\myclint.mtime [37] ), .ZN(_01608_ ) );
AND3_X4 _09062_ ( .A1(_01606_ ), .A2(_01607_ ), .A3(_01608_ ), .ZN(_01609_ ) );
NAND2_X1 _09063_ ( .A1(_01609_ ), .A2(\myclint.mtime [40] ), .ZN(_01610_ ) );
INV_X1 _09064_ ( .A(\myclint.mtime [41] ), .ZN(_01611_ ) );
NOR2_X2 _09065_ ( .A1(_01610_ ), .A2(_01611_ ), .ZN(_01612_ ) );
AND2_X2 _09066_ ( .A1(\myclint.mtime [42] ), .A2(\myclint.mtime [43] ), .ZN(_01613_ ) );
AND2_X2 _09067_ ( .A1(_01612_ ), .A2(_01613_ ), .ZN(_01614_ ) );
AND2_X1 _09068_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01615_ ) );
AND3_X1 _09069_ ( .A1(_01615_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01616_ ) );
AND2_X4 _09070_ ( .A1(_01614_ ), .A2(_01616_ ), .ZN(_01617_ ) );
AND2_X1 _09071_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01618_ ) );
AND2_X2 _09072_ ( .A1(_01617_ ), .A2(_01618_ ), .ZN(_01619_ ) );
AND2_X1 _09073_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01620_ ) );
AND2_X1 _09074_ ( .A1(_01619_ ), .A2(_01620_ ), .ZN(_01621_ ) );
AND2_X1 _09075_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01622_ ) );
AND2_X2 _09076_ ( .A1(_01621_ ), .A2(_01622_ ), .ZN(_01623_ ) );
AND2_X1 _09077_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01624_ ) );
AND2_X2 _09078_ ( .A1(_01623_ ), .A2(_01624_ ), .ZN(_01625_ ) );
AND2_X1 _09079_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01626_ ) );
AND2_X4 _09080_ ( .A1(_01625_ ), .A2(_01626_ ), .ZN(_01627_ ) );
AND2_X1 _09081_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01628_ ) );
AND2_X2 _09082_ ( .A1(_01627_ ), .A2(_01628_ ), .ZN(_01629_ ) );
NAND3_X1 _09083_ ( .A1(_01629_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01630_ ) );
NOR2_X2 _09084_ ( .A1(_01630_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01631_ ) );
OAI21_X1 _09085_ ( .A(_01587_ ), .B1(_01631_ ), .B2(\myclint.mtime [63] ), .ZN(_01632_ ) );
AND2_X1 _09086_ ( .A1(_01601_ ), .A2(_01603_ ), .ZN(_01633_ ) );
AND2_X1 _09087_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01634_ ) );
AND3_X1 _09088_ ( .A1(_01633_ ), .A2(_01634_ ), .A3(_01602_ ), .ZN(_01635_ ) );
AND2_X1 _09089_ ( .A1(_01635_ ), .A2(\myclint.mtime [34] ), .ZN(_01636_ ) );
AND2_X1 _09090_ ( .A1(_01636_ ), .A2(\myclint.mtime [35] ), .ZN(_01637_ ) );
AND3_X1 _09091_ ( .A1(_01637_ ), .A2(_01607_ ), .A3(_01608_ ), .ZN(_01638_ ) );
AND2_X1 _09092_ ( .A1(_01638_ ), .A2(\myclint.mtime [40] ), .ZN(_01639_ ) );
AND2_X2 _09093_ ( .A1(_01639_ ), .A2(\myclint.mtime [41] ), .ZN(_01640_ ) );
AND2_X2 _09094_ ( .A1(_01640_ ), .A2(_01613_ ), .ZN(_01641_ ) );
AND2_X1 _09095_ ( .A1(_01641_ ), .A2(_01616_ ), .ZN(_01642_ ) );
AND2_X2 _09096_ ( .A1(_01642_ ), .A2(_01618_ ), .ZN(_01643_ ) );
AND2_X1 _09097_ ( .A1(_01643_ ), .A2(_01620_ ), .ZN(_01644_ ) );
AND2_X1 _09098_ ( .A1(_01644_ ), .A2(_01622_ ), .ZN(_01645_ ) );
AND2_X1 _09099_ ( .A1(_01645_ ), .A2(_01624_ ), .ZN(_01646_ ) );
AND2_X2 _09100_ ( .A1(_01646_ ), .A2(_01626_ ), .ZN(_01647_ ) );
AND2_X1 _09101_ ( .A1(_01647_ ), .A2(_01628_ ), .ZN(_01648_ ) );
NAND3_X1 _09102_ ( .A1(_01648_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01649_ ) );
NOR2_X1 _09103_ ( .A1(_01649_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01650_ ) );
AOI21_X1 _09104_ ( .A(_01632_ ), .B1(_01650_ ), .B2(\myclint.mtime [63] ), .ZN(_00001_ ) );
AND2_X1 _09105_ ( .A1(_01588_ ), .A2(\myclint.mtime [3] ), .ZN(_01651_ ) );
AND4_X1 _09106_ ( .A1(\myclint.mtime [6] ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [5] ), .A4(\myclint.mtime [7] ), .ZN(_01652_ ) );
AND2_X1 _09107_ ( .A1(_01651_ ), .A2(_01652_ ), .ZN(_01653_ ) );
AND4_X1 _09108_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01654_ ) );
AND2_X1 _09109_ ( .A1(\myclint.mtime [8] ), .A2(\myclint.mtime [9] ), .ZN(_01655_ ) );
AND4_X1 _09110_ ( .A1(\myclint.mtime [10] ), .A2(_01654_ ), .A3(\myclint.mtime [11] ), .A4(_01655_ ), .ZN(_01656_ ) );
NAND2_X1 _09111_ ( .A1(_01653_ ), .A2(_01656_ ), .ZN(_01657_ ) );
AND2_X1 _09112_ ( .A1(\myclint.mtime [16] ), .A2(\myclint.mtime [17] ), .ZN(_01658_ ) );
NAND3_X1 _09113_ ( .A1(_01658_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [19] ), .ZN(_01659_ ) );
NAND4_X1 _09114_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01660_ ) );
NOR2_X1 _09115_ ( .A1(_01659_ ), .A2(_01660_ ), .ZN(_01661_ ) );
AND2_X1 _09116_ ( .A1(\myclint.mtime [24] ), .A2(\myclint.mtime [25] ), .ZN(_01662_ ) );
AND3_X1 _09117_ ( .A1(_01662_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [27] ), .ZN(_01663_ ) );
NAND4_X1 _09118_ ( .A1(_01661_ ), .A2(_01602_ ), .A3(_01603_ ), .A4(_01663_ ), .ZN(_01664_ ) );
NOR2_X1 _09119_ ( .A1(_01657_ ), .A2(_01664_ ), .ZN(_01665_ ) );
AND3_X1 _09120_ ( .A1(_01634_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01666_ ) );
AND3_X1 _09121_ ( .A1(_01666_ ), .A2(_01607_ ), .A3(_01608_ ), .ZN(_01667_ ) );
AND3_X1 _09122_ ( .A1(_01613_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01668_ ) );
AND3_X1 _09123_ ( .A1(_01667_ ), .A2(_01616_ ), .A3(_01668_ ), .ZN(_01669_ ) );
AND2_X1 _09124_ ( .A1(_01665_ ), .A2(_01669_ ), .ZN(_01670_ ) );
AND4_X1 _09125_ ( .A1(_01624_ ), .A2(_01622_ ), .A3(_01620_ ), .A4(_01618_ ), .ZN(_01671_ ) );
AND2_X1 _09126_ ( .A1(_01670_ ), .A2(_01671_ ), .ZN(_01672_ ) );
AND4_X1 _09127_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01673_ ) );
AND2_X1 _09128_ ( .A1(_01672_ ), .A2(_01673_ ), .ZN(_01674_ ) );
AND3_X1 _09129_ ( .A1(_01674_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01675_ ) );
XNOR2_X1 _09130_ ( .A(_01675_ ), .B(\myclint.mtime [62] ), .ZN(_01676_ ) );
NOR2_X1 _09131_ ( .A1(_01676_ ), .A2(fanout_net_1 ), .ZN(_00002_ ) );
INV_X1 _09132_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01677_ ) );
AND4_X1 _09133_ ( .A1(_01677_ ), .A2(_01643_ ), .A3(\myclint.mtime [53] ), .A4(_01620_ ), .ZN(_01678_ ) );
BUF_X4 _09134_ ( .A(_01586_ ), .Z(_01679_ ) );
AND3_X1 _09135_ ( .A1(_01619_ ), .A2(_01677_ ), .A3(_01620_ ), .ZN(_01680_ ) );
OAI21_X1 _09136_ ( .A(_01679_ ), .B1(_01680_ ), .B2(\myclint.mtime [53] ), .ZN(_01681_ ) );
NOR2_X1 _09137_ ( .A1(_01678_ ), .A2(_01681_ ), .ZN(_00003_ ) );
AND2_X1 _09138_ ( .A1(_01620_ ), .A2(_01618_ ), .ZN(_01682_ ) );
AND2_X1 _09139_ ( .A1(_01670_ ), .A2(_01682_ ), .ZN(_01683_ ) );
XNOR2_X1 _09140_ ( .A(_01683_ ), .B(\myclint.mtime [52] ), .ZN(_01684_ ) );
NOR2_X1 _09141_ ( .A1(_01684_ ), .A2(fanout_net_1 ), .ZN(_00004_ ) );
NAND2_X1 _09142_ ( .A1(_01617_ ), .A2(_01618_ ), .ZN(_01685_ ) );
NOR2_X1 _09143_ ( .A1(_01685_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01686_ ) );
OAI21_X1 _09144_ ( .A(_01587_ ), .B1(_01686_ ), .B2(\myclint.mtime [51] ), .ZN(_01687_ ) );
INV_X1 _09145_ ( .A(_01643_ ), .ZN(_01688_ ) );
NOR2_X1 _09146_ ( .A1(_01688_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01689_ ) );
AOI21_X1 _09147_ ( .A(_01687_ ), .B1(_01689_ ), .B2(\myclint.mtime [51] ), .ZN(_00005_ ) );
AND3_X1 _09148_ ( .A1(_01665_ ), .A2(_01618_ ), .A3(_01669_ ), .ZN(_01690_ ) );
XNOR2_X1 _09149_ ( .A(_01690_ ), .B(\myclint.mtime [50] ), .ZN(_01691_ ) );
NOR2_X1 _09150_ ( .A1(_01691_ ), .A2(fanout_net_1 ), .ZN(_00006_ ) );
NAND2_X1 _09151_ ( .A1(_01614_ ), .A2(_01616_ ), .ZN(_01692_ ) );
NOR2_X1 _09152_ ( .A1(_01692_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01693_ ) );
OAI21_X1 _09153_ ( .A(_01587_ ), .B1(_01693_ ), .B2(\myclint.mtime [49] ), .ZN(_01694_ ) );
INV_X1 _09154_ ( .A(_01641_ ), .ZN(_01695_ ) );
INV_X1 _09155_ ( .A(_01616_ ), .ZN(_01696_ ) );
NOR3_X1 _09156_ ( .A1(_01695_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01696_ ), .ZN(_01697_ ) );
AOI21_X1 _09157_ ( .A(_01694_ ), .B1(_01697_ ), .B2(\myclint.mtime [49] ), .ZN(_00007_ ) );
INV_X1 _09158_ ( .A(_01665_ ), .ZN(_01698_ ) );
INV_X1 _09159_ ( .A(_01669_ ), .ZN(_01699_ ) );
OR3_X1 _09160_ ( .A1(_01698_ ), .A2(_01699_ ), .A3(\myclint.mtime [48] ), .ZN(_01700_ ) );
OAI21_X1 _09161_ ( .A(\myclint.mtime [48] ), .B1(_01698_ ), .B2(_01699_ ), .ZN(_01701_ ) );
AOI21_X1 _09162_ ( .A(fanout_net_1 ), .B1(_01700_ ), .B2(_01701_ ), .ZN(_00008_ ) );
NAND3_X1 _09163_ ( .A1(_01612_ ), .A2(_01615_ ), .A3(_01613_ ), .ZN(_01702_ ) );
NOR2_X1 _09164_ ( .A1(_01702_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01703_ ) );
OAI21_X1 _09165_ ( .A(_01587_ ), .B1(_01703_ ), .B2(\myclint.mtime [47] ), .ZN(_01704_ ) );
NAND3_X1 _09166_ ( .A1(_01640_ ), .A2(\myclint.mtime [44] ), .A3(_01613_ ), .ZN(_01705_ ) );
INV_X1 _09167_ ( .A(\myclint.mtime [45] ), .ZN(_01706_ ) );
NOR3_X1 _09168_ ( .A1(_01705_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01706_ ), .ZN(_01707_ ) );
AOI21_X1 _09169_ ( .A(_01704_ ), .B1(_01707_ ), .B2(\myclint.mtime [47] ), .ZN(_00009_ ) );
AND2_X1 _09170_ ( .A1(_01665_ ), .A2(_01667_ ), .ZN(_01708_ ) );
AND3_X1 _09171_ ( .A1(_01708_ ), .A2(_01615_ ), .A3(_01668_ ), .ZN(_01709_ ) );
XNOR2_X1 _09172_ ( .A(_01709_ ), .B(\myclint.mtime [46] ), .ZN(_01710_ ) );
NOR2_X1 _09173_ ( .A1(_01710_ ), .A2(fanout_net_1 ), .ZN(_00010_ ) );
INV_X1 _09174_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01711_ ) );
NAND4_X1 _09175_ ( .A1(_01640_ ), .A2(\myclint.mtime [45] ), .A3(_01711_ ), .A4(_01613_ ), .ZN(_01712_ ) );
NAND3_X1 _09176_ ( .A1(_01612_ ), .A2(_01711_ ), .A3(_01613_ ), .ZN(_01713_ ) );
AOI21_X1 _09177_ ( .A(fanout_net_1 ), .B1(_01713_ ), .B2(_01706_ ), .ZN(_01714_ ) );
AND2_X1 _09178_ ( .A1(_01712_ ), .A2(_01714_ ), .ZN(_00011_ ) );
AND2_X1 _09179_ ( .A1(_01708_ ), .A2(_01668_ ), .ZN(_01715_ ) );
XNOR2_X1 _09180_ ( .A(_01715_ ), .B(\myclint.mtime [44] ), .ZN(_01716_ ) );
NOR2_X1 _09181_ ( .A1(_01716_ ), .A2(fanout_net_1 ), .ZN(_00012_ ) );
INV_X1 _09182_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01717_ ) );
AND4_X1 _09183_ ( .A1(\myclint.mtime [61] ), .A2(_01647_ ), .A3(_01717_ ), .A4(_01628_ ), .ZN(_01718_ ) );
AND3_X1 _09184_ ( .A1(_01627_ ), .A2(_01717_ ), .A3(_01628_ ), .ZN(_01719_ ) );
OAI21_X1 _09185_ ( .A(_01679_ ), .B1(_01719_ ), .B2(\myclint.mtime [61] ), .ZN(_01720_ ) );
NOR2_X1 _09186_ ( .A1(_01718_ ), .A2(_01720_ ), .ZN(_00013_ ) );
AND3_X1 _09187_ ( .A1(_01708_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01721_ ) );
INV_X1 _09188_ ( .A(_01721_ ), .ZN(_01722_ ) );
OR3_X1 _09189_ ( .A1(_01722_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [43] ), .ZN(_01723_ ) );
OAI21_X1 _09190_ ( .A(\myclint.mtime [43] ), .B1(_01722_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01724_ ) );
AOI21_X1 _09191_ ( .A(fanout_net_1 ), .B1(_01723_ ), .B2(_01724_ ), .ZN(_00014_ ) );
XNOR2_X1 _09192_ ( .A(_01721_ ), .B(\myclint.mtime [42] ), .ZN(_01725_ ) );
NOR2_X1 _09193_ ( .A1(_01725_ ), .A2(fanout_net_1 ), .ZN(_00015_ ) );
INV_X1 _09194_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01726_ ) );
AND3_X1 _09195_ ( .A1(_01638_ ), .A2(\myclint.mtime [41] ), .A3(_01726_ ), .ZN(_01727_ ) );
NAND3_X1 _09196_ ( .A1(_01606_ ), .A2(_01607_ ), .A3(_01608_ ), .ZN(_01728_ ) );
NOR2_X1 _09197_ ( .A1(_01728_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01729_ ) );
OAI21_X1 _09198_ ( .A(_01679_ ), .B1(_01729_ ), .B2(\myclint.mtime [41] ), .ZN(_01730_ ) );
NOR2_X1 _09199_ ( .A1(_01727_ ), .A2(_01730_ ), .ZN(_00016_ ) );
XNOR2_X1 _09200_ ( .A(_01708_ ), .B(\myclint.mtime [40] ), .ZN(_01731_ ) );
NOR2_X1 _09201_ ( .A1(_01731_ ), .A2(fanout_net_1 ), .ZN(_00017_ ) );
NAND3_X1 _09202_ ( .A1(_01665_ ), .A2(_01608_ ), .A3(_01666_ ), .ZN(_01732_ ) );
OR3_X1 _09203_ ( .A1(_01732_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [39] ), .ZN(_01733_ ) );
OAI21_X1 _09204_ ( .A(\myclint.mtime [39] ), .B1(_01732_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01734_ ) );
AOI21_X1 _09205_ ( .A(fanout_net_1 ), .B1(_01733_ ), .B2(_01734_ ), .ZN(_00018_ ) );
OR2_X1 _09206_ ( .A1(_01732_ ), .A2(\myclint.mtime [38] ), .ZN(_01735_ ) );
NAND2_X1 _09207_ ( .A1(_01732_ ), .A2(\myclint.mtime [38] ), .ZN(_01736_ ) );
AOI21_X1 _09208_ ( .A(fanout_net_1 ), .B1(_01735_ ), .B2(_01736_ ), .ZN(_00019_ ) );
INV_X1 _09209_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01737_ ) );
AND4_X1 _09210_ ( .A1(\myclint.mtime [37] ), .A2(_01636_ ), .A3(_01737_ ), .A4(\myclint.mtime [35] ), .ZN(_01738_ ) );
AND3_X1 _09211_ ( .A1(_01605_ ), .A2(_01737_ ), .A3(\myclint.mtime [35] ), .ZN(_01739_ ) );
OAI21_X1 _09212_ ( .A(_01679_ ), .B1(_01739_ ), .B2(\myclint.mtime [37] ), .ZN(_01740_ ) );
NOR2_X1 _09213_ ( .A1(_01738_ ), .A2(_01740_ ), .ZN(_00020_ ) );
AND2_X1 _09214_ ( .A1(_01665_ ), .A2(_01666_ ), .ZN(_01741_ ) );
XNOR2_X1 _09215_ ( .A(_01741_ ), .B(\myclint.mtime [36] ), .ZN(_01742_ ) );
NOR2_X1 _09216_ ( .A1(_01742_ ), .A2(fanout_net_1 ), .ZN(_00021_ ) );
AND2_X1 _09217_ ( .A1(_01653_ ), .A2(_01656_ ), .ZN(_01743_ ) );
AND4_X1 _09218_ ( .A1(_01602_ ), .A2(_01661_ ), .A3(_01603_ ), .A4(_01663_ ), .ZN(_01744_ ) );
NAND3_X1 _09219_ ( .A1(_01743_ ), .A2(_01634_ ), .A3(_01744_ ), .ZN(_01745_ ) );
OR3_X1 _09220_ ( .A1(_01745_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [35] ), .ZN(_01746_ ) );
OAI21_X1 _09221_ ( .A(\myclint.mtime [35] ), .B1(_01745_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01747_ ) );
AOI21_X1 _09222_ ( .A(fanout_net_1 ), .B1(_01746_ ), .B2(_01747_ ), .ZN(_00022_ ) );
CLKBUF_X2 _09223_ ( .A(_01586_ ), .Z(_01748_ ) );
NAND4_X1 _09224_ ( .A1(_01601_ ), .A2(\myclint.mtime [33] ), .A3(_01602_ ), .A4(_01603_ ), .ZN(_01749_ ) );
INV_X1 _09225_ ( .A(\myclint.mtime [32] ), .ZN(_01750_ ) );
NOR2_X1 _09226_ ( .A1(_01749_ ), .A2(_01750_ ), .ZN(_01751_ ) );
OAI21_X1 _09227_ ( .A(_01748_ ), .B1(_01751_ ), .B2(\myclint.mtime [34] ), .ZN(_01752_ ) );
NOR2_X1 _09228_ ( .A1(_01752_ ), .A2(_01605_ ), .ZN(_00023_ ) );
XNOR2_X1 _09229_ ( .A(_01674_ ), .B(\myclint.mtime [60] ), .ZN(_01753_ ) );
NOR2_X1 _09230_ ( .A1(_01753_ ), .A2(fanout_net_1 ), .ZN(_00024_ ) );
INV_X1 _09231_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .ZN(_01754_ ) );
AND3_X1 _09232_ ( .A1(_01633_ ), .A2(_01754_ ), .A3(_01602_ ), .ZN(_01755_ ) );
AND2_X1 _09233_ ( .A1(_01755_ ), .A2(\myclint.mtime [33] ), .ZN(_01756_ ) );
OAI21_X1 _09234_ ( .A(_01679_ ), .B1(_01755_ ), .B2(\myclint.mtime [33] ), .ZN(_01757_ ) );
NOR2_X1 _09235_ ( .A1(_01756_ ), .A2(_01757_ ), .ZN(_00025_ ) );
NAND4_X1 _09236_ ( .A1(_01744_ ), .A2(_01750_ ), .A3(_01653_ ), .A4(_01656_ ), .ZN(_01758_ ) );
OAI21_X1 _09237_ ( .A(\myclint.mtime [32] ), .B1(_01657_ ), .B2(_01664_ ), .ZN(_01759_ ) );
AOI21_X1 _09238_ ( .A(fanout_net_1 ), .B1(_01758_ ), .B2(_01759_ ), .ZN(_00026_ ) );
INV_X1 _09239_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01760_ ) );
AND3_X1 _09240_ ( .A1(_01601_ ), .A2(_01760_ ), .A3(_01603_ ), .ZN(_01761_ ) );
AND2_X1 _09241_ ( .A1(_01761_ ), .A2(\myclint.mtime [31] ), .ZN(_01762_ ) );
OAI21_X1 _09242_ ( .A(_01679_ ), .B1(_01761_ ), .B2(\myclint.mtime [31] ), .ZN(_01763_ ) );
NOR2_X1 _09243_ ( .A1(_01762_ ), .A2(_01763_ ), .ZN(_00027_ ) );
AND2_X1 _09244_ ( .A1(_01743_ ), .A2(_01661_ ), .ZN(_01764_ ) );
NAND3_X1 _09245_ ( .A1(_01764_ ), .A2(_01603_ ), .A3(_01663_ ), .ZN(_01765_ ) );
OR2_X1 _09246_ ( .A1(_01765_ ), .A2(\myclint.mtime [30] ), .ZN(_01766_ ) );
NAND2_X1 _09247_ ( .A1(_01765_ ), .A2(\myclint.mtime [30] ), .ZN(_01767_ ) );
AOI21_X1 _09248_ ( .A(fanout_net_1 ), .B1(_01766_ ), .B2(_01767_ ), .ZN(_00028_ ) );
INV_X1 _09249_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01768_ ) );
AND3_X1 _09250_ ( .A1(_01600_ ), .A2(_01768_ ), .A3(\myclint.mtime [27] ), .ZN(_01769_ ) );
AND2_X1 _09251_ ( .A1(_01769_ ), .A2(\myclint.mtime [29] ), .ZN(_01770_ ) );
OAI21_X1 _09252_ ( .A(_01679_ ), .B1(_01769_ ), .B2(\myclint.mtime [29] ), .ZN(_01771_ ) );
NOR2_X1 _09253_ ( .A1(_01770_ ), .A2(_01771_ ), .ZN(_00029_ ) );
NAND2_X1 _09254_ ( .A1(_01764_ ), .A2(_01663_ ), .ZN(_01772_ ) );
OR2_X1 _09255_ ( .A1(_01772_ ), .A2(\myclint.mtime [28] ), .ZN(_01773_ ) );
NAND2_X1 _09256_ ( .A1(_01772_ ), .A2(\myclint.mtime [28] ), .ZN(_01774_ ) );
AOI21_X1 _09257_ ( .A(fanout_net_1 ), .B1(_01773_ ), .B2(_01774_ ), .ZN(_00030_ ) );
NAND3_X1 _09258_ ( .A1(_01743_ ), .A2(_01662_ ), .A3(_01661_ ), .ZN(_01775_ ) );
OR3_X1 _09259_ ( .A1(_01775_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [27] ), .ZN(_01776_ ) );
OAI21_X1 _09260_ ( .A(\myclint.mtime [27] ), .B1(_01775_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01777_ ) );
AOI21_X1 _09261_ ( .A(fanout_net_1 ), .B1(_01776_ ), .B2(_01777_ ), .ZN(_00031_ ) );
BUF_X4 _09262_ ( .A(_01586_ ), .Z(_01778_ ) );
AND2_X1 _09263_ ( .A1(_01599_ ), .A2(\myclint.mtime [25] ), .ZN(_01779_ ) );
OAI21_X1 _09264_ ( .A(_01778_ ), .B1(_01779_ ), .B2(\myclint.mtime [26] ), .ZN(_01780_ ) );
NOR2_X1 _09265_ ( .A1(_01780_ ), .A2(_01600_ ), .ZN(_00032_ ) );
INV_X1 _09266_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01781_ ) );
AND3_X1 _09267_ ( .A1(_01598_ ), .A2(_01781_ ), .A3(\myclint.mtime [23] ), .ZN(_01782_ ) );
AND2_X1 _09268_ ( .A1(_01782_ ), .A2(\myclint.mtime [25] ), .ZN(_01783_ ) );
OAI21_X1 _09269_ ( .A(_01679_ ), .B1(_01782_ ), .B2(\myclint.mtime [25] ), .ZN(_01784_ ) );
NOR2_X1 _09270_ ( .A1(_01783_ ), .A2(_01784_ ), .ZN(_00033_ ) );
AND2_X1 _09271_ ( .A1(_01598_ ), .A2(\myclint.mtime [23] ), .ZN(_01785_ ) );
OAI21_X1 _09272_ ( .A(_01778_ ), .B1(_01785_ ), .B2(\myclint.mtime [24] ), .ZN(_01786_ ) );
NOR2_X1 _09273_ ( .A1(_01786_ ), .A2(_01599_ ), .ZN(_00034_ ) );
NAND2_X1 _09274_ ( .A1(_01625_ ), .A2(_01626_ ), .ZN(_01787_ ) );
NOR2_X1 _09275_ ( .A1(_01787_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01788_ ) );
OAI21_X1 _09276_ ( .A(_01587_ ), .B1(_01788_ ), .B2(\myclint.mtime [59] ), .ZN(_01789_ ) );
INV_X1 _09277_ ( .A(_01647_ ), .ZN(_01790_ ) );
NOR2_X1 _09278_ ( .A1(_01790_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01791_ ) );
AOI21_X1 _09279_ ( .A(_01789_ ), .B1(_01791_ ), .B2(\myclint.mtime [59] ), .ZN(_00035_ ) );
NOR2_X1 _09280_ ( .A1(_01657_ ), .A2(_01659_ ), .ZN(_01792_ ) );
NAND3_X1 _09281_ ( .A1(_01792_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01793_ ) );
OR3_X1 _09282_ ( .A1(_01793_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01794_ ) );
OAI21_X1 _09283_ ( .A(\myclint.mtime [23] ), .B1(_01793_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01795_ ) );
AOI21_X1 _09284_ ( .A(fanout_net_1 ), .B1(_01794_ ), .B2(_01795_ ), .ZN(_00036_ ) );
AND2_X1 _09285_ ( .A1(_01597_ ), .A2(\myclint.mtime [21] ), .ZN(_01796_ ) );
OAI21_X1 _09286_ ( .A(_01778_ ), .B1(_01796_ ), .B2(\myclint.mtime [22] ), .ZN(_01797_ ) );
NOR2_X1 _09287_ ( .A1(_01797_ ), .A2(_01598_ ), .ZN(_00037_ ) );
OR3_X1 _09288_ ( .A1(_01657_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01659_ ), .ZN(_01798_ ) );
NAND2_X1 _09289_ ( .A1(_01798_ ), .A2(\myclint.mtime [21] ), .ZN(_01799_ ) );
OR4_X1 _09290_ ( .A1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .A2(_01657_ ), .A3(\myclint.mtime [21] ), .A4(_01659_ ), .ZN(_01800_ ) );
AOI21_X1 _09291_ ( .A(fanout_net_1 ), .B1(_01799_ ), .B2(_01800_ ), .ZN(_00038_ ) );
AND2_X1 _09292_ ( .A1(_01596_ ), .A2(\myclint.mtime [19] ), .ZN(_01801_ ) );
OAI21_X1 _09293_ ( .A(_01778_ ), .B1(_01801_ ), .B2(\myclint.mtime [20] ), .ZN(_01802_ ) );
NOR2_X1 _09294_ ( .A1(_01802_ ), .A2(_01597_ ), .ZN(_00039_ ) );
NAND3_X1 _09295_ ( .A1(_01653_ ), .A2(_01656_ ), .A3(_01658_ ), .ZN(_01803_ ) );
OR3_X1 _09296_ ( .A1(_01803_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01804_ ) );
OAI21_X1 _09297_ ( .A(\myclint.mtime [19] ), .B1(_01803_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01805_ ) );
AOI21_X1 _09298_ ( .A(fanout_net_1 ), .B1(_01804_ ), .B2(_01805_ ), .ZN(_00040_ ) );
AND2_X1 _09299_ ( .A1(_01595_ ), .A2(\myclint.mtime [17] ), .ZN(_01806_ ) );
OAI21_X1 _09300_ ( .A(_01778_ ), .B1(_01806_ ), .B2(\myclint.mtime [18] ), .ZN(_01807_ ) );
NOR2_X1 _09301_ ( .A1(_01807_ ), .A2(_01596_ ), .ZN(_00041_ ) );
INV_X1 _09302_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01808_ ) );
AND3_X1 _09303_ ( .A1(_01594_ ), .A2(_01808_ ), .A3(\myclint.mtime [15] ), .ZN(_01809_ ) );
AND2_X1 _09304_ ( .A1(_01809_ ), .A2(\myclint.mtime [17] ), .ZN(_01810_ ) );
OAI21_X1 _09305_ ( .A(_01587_ ), .B1(_01809_ ), .B2(\myclint.mtime [17] ), .ZN(_01811_ ) );
NOR2_X1 _09306_ ( .A1(_01810_ ), .A2(_01811_ ), .ZN(_00042_ ) );
AND2_X1 _09307_ ( .A1(_01594_ ), .A2(\myclint.mtime [15] ), .ZN(_01812_ ) );
OAI21_X1 _09308_ ( .A(_01778_ ), .B1(_01812_ ), .B2(\myclint.mtime [16] ), .ZN(_01813_ ) );
NOR2_X1 _09309_ ( .A1(_01813_ ), .A2(_01595_ ), .ZN(_00043_ ) );
AND3_X1 _09310_ ( .A1(_01655_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [11] ), .ZN(_01814_ ) );
AND2_X1 _09311_ ( .A1(_01653_ ), .A2(_01814_ ), .ZN(_01815_ ) );
NAND3_X1 _09312_ ( .A1(_01815_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01816_ ) );
OR3_X1 _09313_ ( .A1(_01816_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01817_ ) );
OAI21_X1 _09314_ ( .A(\myclint.mtime [15] ), .B1(_01816_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01818_ ) );
AOI21_X1 _09315_ ( .A(fanout_net_1 ), .B1(_01817_ ), .B2(_01818_ ), .ZN(_00044_ ) );
AND2_X1 _09316_ ( .A1(_01593_ ), .A2(\myclint.mtime [13] ), .ZN(_01819_ ) );
OAI21_X1 _09317_ ( .A(_01778_ ), .B1(_01819_ ), .B2(\myclint.mtime [14] ), .ZN(_01820_ ) );
NOR2_X1 _09318_ ( .A1(_01820_ ), .A2(_01594_ ), .ZN(_00045_ ) );
NAND3_X1 _09319_ ( .A1(_01670_ ), .A2(_01626_ ), .A3(_01671_ ), .ZN(_01821_ ) );
OR2_X1 _09320_ ( .A1(_01821_ ), .A2(\myclint.mtime [58] ), .ZN(_01822_ ) );
NAND2_X1 _09321_ ( .A1(_01821_ ), .A2(\myclint.mtime [58] ), .ZN(_01823_ ) );
AOI21_X1 _09322_ ( .A(fanout_net_1 ), .B1(_01822_ ), .B2(_01823_ ), .ZN(_00046_ ) );
INV_X1 _09323_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01824_ ) );
AND3_X1 _09324_ ( .A1(_01592_ ), .A2(_01824_ ), .A3(\myclint.mtime [11] ), .ZN(_01825_ ) );
AND2_X1 _09325_ ( .A1(_01825_ ), .A2(\myclint.mtime [13] ), .ZN(_01826_ ) );
OAI21_X1 _09326_ ( .A(_01587_ ), .B1(_01825_ ), .B2(\myclint.mtime [13] ), .ZN(_01827_ ) );
NOR2_X1 _09327_ ( .A1(_01826_ ), .A2(_01827_ ), .ZN(_00047_ ) );
AND2_X1 _09328_ ( .A1(_01592_ ), .A2(\myclint.mtime [11] ), .ZN(_01828_ ) );
OAI21_X1 _09329_ ( .A(_01778_ ), .B1(_01828_ ), .B2(\myclint.mtime [12] ), .ZN(_01829_ ) );
NOR2_X1 _09330_ ( .A1(_01829_ ), .A2(_01593_ ), .ZN(_00048_ ) );
INV_X1 _09331_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01830_ ) );
AND3_X1 _09332_ ( .A1(_01591_ ), .A2(_01830_ ), .A3(\myclint.mtime [9] ), .ZN(_01831_ ) );
OAI21_X1 _09333_ ( .A(_01586_ ), .B1(_01831_ ), .B2(\myclint.mtime [11] ), .ZN(_01832_ ) );
AOI21_X1 _09334_ ( .A(_01832_ ), .B1(\myclint.mtime [11] ), .B2(_01831_ ), .ZN(_00049_ ) );
AOI21_X1 _09335_ ( .A(\myclint.mtime [10] ), .B1(_01591_ ), .B2(\myclint.mtime [9] ), .ZN(_01833_ ) );
NOR3_X1 _09336_ ( .A1(_01592_ ), .A2(_01833_ ), .A3(fanout_net_1 ), .ZN(_00050_ ) );
INV_X1 _09337_ ( .A(_01651_ ), .ZN(_01834_ ) );
NAND4_X1 _09338_ ( .A1(\myclint.mtime [6] ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [5] ), .A4(\myclint.mtime [7] ), .ZN(_01835_ ) );
OR3_X1 _09339_ ( .A1(_01834_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(_01835_ ), .ZN(_01836_ ) );
NAND2_X1 _09340_ ( .A1(_01836_ ), .A2(\myclint.mtime [9] ), .ZN(_01837_ ) );
OR4_X1 _09341_ ( .A1(\myclint.mtime [9] ), .A2(_01834_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .A4(_01835_ ), .ZN(_01838_ ) );
AOI21_X1 _09342_ ( .A(fanout_net_1 ), .B1(_01837_ ), .B2(_01838_ ), .ZN(_00051_ ) );
AND2_X1 _09343_ ( .A1(_01590_ ), .A2(\myclint.mtime [7] ), .ZN(_01839_ ) );
OAI21_X1 _09344_ ( .A(_01778_ ), .B1(_01839_ ), .B2(\myclint.mtime [8] ), .ZN(_01840_ ) );
NOR2_X1 _09345_ ( .A1(_01840_ ), .A2(_01591_ ), .ZN(_00052_ ) );
AND2_X1 _09346_ ( .A1(_01589_ ), .A2(\myclint.mtime [5] ), .ZN(_01841_ ) );
INV_X1 _09347_ ( .A(_01841_ ), .ZN(_01842_ ) );
OR3_X1 _09348_ ( .A1(_01842_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [7] ), .ZN(_01843_ ) );
OAI21_X1 _09349_ ( .A(\myclint.mtime [7] ), .B1(_01842_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01844_ ) );
AOI21_X1 _09350_ ( .A(fanout_net_1 ), .B1(_01843_ ), .B2(_01844_ ), .ZN(_00053_ ) );
OAI21_X1 _09351_ ( .A(_01778_ ), .B1(_01841_ ), .B2(\myclint.mtime [6] ), .ZN(_01845_ ) );
NOR2_X1 _09352_ ( .A1(_01845_ ), .A2(_01590_ ), .ZN(_00054_ ) );
OR3_X1 _09353_ ( .A1(_01834_ ), .A2(\myclint.mtime [5] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01846_ ) );
OAI21_X1 _09354_ ( .A(\myclint.mtime [5] ), .B1(_01834_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01847_ ) );
AOI21_X1 _09355_ ( .A(fanout_net_1 ), .B1(_01846_ ), .B2(_01847_ ), .ZN(_00055_ ) );
OAI21_X1 _09356_ ( .A(_01679_ ), .B1(_01651_ ), .B2(\myclint.mtime [4] ), .ZN(_01848_ ) );
NOR2_X1 _09357_ ( .A1(_01848_ ), .A2(_01589_ ), .ZN(_00056_ ) );
INV_X1 _09358_ ( .A(_01672_ ), .ZN(_01849_ ) );
OR3_X1 _09359_ ( .A1(_01849_ ), .A2(\myclint.mtime [57] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01850_ ) );
OAI21_X1 _09360_ ( .A(\myclint.mtime [57] ), .B1(_01849_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01851_ ) );
AOI21_X1 _09361_ ( .A(fanout_net_2 ), .B1(_01850_ ), .B2(_01851_ ), .ZN(_00057_ ) );
AND2_X1 _09362_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01852_ ) );
INV_X1 _09363_ ( .A(_01852_ ), .ZN(_01853_ ) );
OR3_X1 _09364_ ( .A1(_01853_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01854_ ) );
OAI21_X1 _09365_ ( .A(\myclint.mtime [3] ), .B1(_01853_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01855_ ) );
AOI21_X1 _09366_ ( .A(fanout_net_2 ), .B1(_01854_ ), .B2(_01855_ ), .ZN(_00058_ ) );
AOI21_X1 _09367_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [0] ), .B2(\myclint.mtime [1] ), .ZN(_01856_ ) );
NOR3_X1 _09368_ ( .A1(_01588_ ), .A2(_01856_ ), .A3(fanout_net_2 ), .ZN(_00059_ ) );
NOR2_X1 _09369_ ( .A1(\myclint.mtime [0] ), .A2(\myclint.mtime [1] ), .ZN(_01857_ ) );
NOR3_X1 _09370_ ( .A1(_01852_ ), .A2(_01857_ ), .A3(fanout_net_2 ), .ZN(_00060_ ) );
INV_X1 _09371_ ( .A(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_01858_ ) );
NOR2_X1 _09372_ ( .A1(_01858_ ), .A2(fanout_net_2 ), .ZN(_00061_ ) );
XNOR2_X1 _09373_ ( .A(_01672_ ), .B(\myclint.mtime [56] ), .ZN(_01859_ ) );
NOR2_X1 _09374_ ( .A1(_01859_ ), .A2(fanout_net_2 ), .ZN(_00062_ ) );
NAND3_X1 _09375_ ( .A1(_01670_ ), .A2(_01622_ ), .A3(_01682_ ), .ZN(_01860_ ) );
OR3_X1 _09376_ ( .A1(_01860_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01861_ ) );
OAI21_X1 _09377_ ( .A(\myclint.mtime [55] ), .B1(_01860_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01862_ ) );
AOI21_X1 _09378_ ( .A(fanout_net_2 ), .B1(_01861_ ), .B2(_01862_ ), .ZN(_00063_ ) );
OR2_X1 _09379_ ( .A1(_01860_ ), .A2(\myclint.mtime [54] ), .ZN(_01863_ ) );
NAND2_X1 _09380_ ( .A1(_01860_ ), .A2(\myclint.mtime [54] ), .ZN(_01864_ ) );
AOI21_X1 _09381_ ( .A(fanout_net_2 ), .B1(_01863_ ), .B2(_01864_ ), .ZN(_00064_ ) );
INV_X32 _09382_ ( .A(fanout_net_44 ), .ZN(_01865_ ) );
OR2_X1 _09383_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[3][1] ), .ZN(_01866_ ) );
OAI211_X1 _09384_ ( .A(_01866_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[2][1] ), .ZN(_01867_ ) );
OR2_X1 _09385_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_01868_ ) );
INV_X32 _09386_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01869_ ) );
BUF_X8 _09387_ ( .A(_01869_ ), .Z(_01870_ ) );
BUF_X16 _09388_ ( .A(_01865_ ), .Z(_01871_ ) );
BUF_X4 _09389_ ( .A(_01871_ ), .Z(_01872_ ) );
OAI211_X1 _09390_ ( .A(_01868_ ), .B(_01870_ ), .C1(_01872_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_01873_ ) );
NAND2_X1 _09391_ ( .A1(_01867_ ), .A2(_01873_ ), .ZN(_01874_ ) );
INV_X1 _09392_ ( .A(\IF_ID_pc [6] ), .ZN(_01875_ ) );
XNOR2_X1 _09393_ ( .A(_01874_ ), .B(_01875_ ), .ZN(_01876_ ) );
OR2_X4 _09394_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[1][17] ), .ZN(_01877_ ) );
OAI211_X1 _09395_ ( .A(_01877_ ), .B(_01870_ ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[0][17] ), .ZN(_01878_ ) );
OR2_X4 _09396_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][17] ), .ZN(_01879_ ) );
OAI211_X1 _09397_ ( .A(_01879_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01871_ ), .C2(\myifu.myicache.tag[3][17] ), .ZN(_01880_ ) );
INV_X1 _09398_ ( .A(\IF_ID_pc [22] ), .ZN(_01881_ ) );
AND3_X2 _09399_ ( .A1(_01878_ ), .A2(_01880_ ), .A3(_01881_ ), .ZN(_01882_ ) );
AOI21_X1 _09400_ ( .A(_01881_ ), .B1(_01878_ ), .B2(_01880_ ), .ZN(_01883_ ) );
OR2_X2 _09401_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[3][8] ), .ZN(_01884_ ) );
OAI211_X2 _09402_ ( .A(_01884_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[2][8] ), .ZN(_01885_ ) );
INV_X1 _09403_ ( .A(\IF_ID_pc [13] ), .ZN(_01886_ ) );
OR2_X4 _09404_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][8] ), .ZN(_01887_ ) );
OAI211_X1 _09405_ ( .A(_01887_ ), .B(_01869_ ), .C1(_01871_ ), .C2(\myifu.myicache.tag[1][8] ), .ZN(_01888_ ) );
AND3_X2 _09406_ ( .A1(_01885_ ), .A2(_01886_ ), .A3(_01888_ ), .ZN(_01889_ ) );
AOI21_X1 _09407_ ( .A(_01886_ ), .B1(_01885_ ), .B2(_01888_ ), .ZN(_01890_ ) );
OAI22_X1 _09408_ ( .A1(_01882_ ), .A2(_01883_ ), .B1(_01889_ ), .B2(_01890_ ), .ZN(_01891_ ) );
OR2_X4 _09409_ ( .A1(_01871_ ), .A2(\myifu.myicache.tag[1][4] ), .ZN(_01892_ ) );
OAI211_X1 _09410_ ( .A(_01892_ ), .B(_01870_ ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[0][4] ), .ZN(_01893_ ) );
OR2_X1 _09411_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[3][4] ), .ZN(_01894_ ) );
OAI211_X1 _09412_ ( .A(_01894_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[2][4] ), .ZN(_01895_ ) );
AND3_X1 _09413_ ( .A1(_01893_ ), .A2(_01895_ ), .A3(\IF_ID_pc [9] ), .ZN(_01896_ ) );
AOI21_X1 _09414_ ( .A(\IF_ID_pc [9] ), .B1(_01893_ ), .B2(_01895_ ), .ZN(_01897_ ) );
OR4_X2 _09415_ ( .A1(_01876_ ), .A2(_01891_ ), .A3(_01896_ ), .A4(_01897_ ), .ZN(_01898_ ) );
OR2_X2 _09416_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[1][21] ), .ZN(_01899_ ) );
OAI211_X1 _09417_ ( .A(_01899_ ), .B(_01870_ ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[0][21] ), .ZN(_01900_ ) );
OR2_X4 _09418_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[3][21] ), .ZN(_01901_ ) );
OAI211_X1 _09419_ ( .A(_01901_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[2][21] ), .ZN(_01902_ ) );
INV_X1 _09420_ ( .A(\IF_ID_pc [26] ), .ZN(_01903_ ) );
AND3_X1 _09421_ ( .A1(_01900_ ), .A2(_01902_ ), .A3(_01903_ ), .ZN(_01904_ ) );
AOI21_X1 _09422_ ( .A(_01903_ ), .B1(_01900_ ), .B2(_01902_ ), .ZN(_01905_ ) );
OR2_X2 _09423_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[1][0] ), .ZN(_01906_ ) );
OAI211_X1 _09424_ ( .A(_01906_ ), .B(_01869_ ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[0][0] ), .ZN(_01907_ ) );
OR2_X2 _09425_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[3][0] ), .ZN(_01908_ ) );
OAI211_X1 _09426_ ( .A(_01908_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[2][0] ), .ZN(_01909_ ) );
AND3_X2 _09427_ ( .A1(_01907_ ), .A2(_01909_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01910_ ) );
AOI21_X1 _09428_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_01907_ ), .B2(_01909_ ), .ZN(_01911_ ) );
OAI22_X1 _09429_ ( .A1(_01904_ ), .A2(_01905_ ), .B1(_01910_ ), .B2(_01911_ ), .ZN(_01912_ ) );
OR2_X1 _09430_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[0][26] ), .ZN(_01913_ ) );
OAI211_X1 _09431_ ( .A(_01913_ ), .B(_01869_ ), .C1(_01871_ ), .C2(\myifu.myicache.tag[1][26] ), .ZN(_01914_ ) );
OR2_X1 _09432_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][26] ), .ZN(_01915_ ) );
OAI211_X1 _09433_ ( .A(_01915_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01871_ ), .C2(\myifu.myicache.tag[3][26] ), .ZN(_01916_ ) );
NAND2_X1 _09434_ ( .A1(_01914_ ), .A2(_01916_ ), .ZN(_01917_ ) );
INV_X1 _09435_ ( .A(\IF_ID_pc [31] ), .ZN(_01918_ ) );
XNOR2_X1 _09436_ ( .A(_01917_ ), .B(_01918_ ), .ZN(_01919_ ) );
OR2_X1 _09437_ ( .A1(_01865_ ), .A2(\myifu.myicache.tag[1][10] ), .ZN(_01920_ ) );
OAI211_X1 _09438_ ( .A(_01920_ ), .B(_01870_ ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[0][10] ), .ZN(_01921_ ) );
OR2_X1 _09439_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][10] ), .ZN(_01922_ ) );
OAI211_X1 _09440_ ( .A(_01922_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01871_ ), .C2(\myifu.myicache.tag[3][10] ), .ZN(_01923_ ) );
AND3_X1 _09441_ ( .A1(_01921_ ), .A2(_01923_ ), .A3(\IF_ID_pc [15] ), .ZN(_01924_ ) );
AOI21_X1 _09442_ ( .A(\IF_ID_pc [15] ), .B1(_01921_ ), .B2(_01923_ ), .ZN(_01925_ ) );
OR4_X2 _09443_ ( .A1(_01912_ ), .A2(_01919_ ), .A3(_01924_ ), .A4(_01925_ ), .ZN(_01926_ ) );
MUX2_X1 _09444_ ( .A(\myifu.myicache.tag[2][3] ), .B(\myifu.myicache.tag[3][3] ), .S(fanout_net_44 ), .Z(_01927_ ) );
AND2_X1 _09445_ ( .A1(_01927_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01928_ ) );
BUF_X2 _09446_ ( .A(_01869_ ), .Z(_01929_ ) );
MUX2_X1 _09447_ ( .A(\myifu.myicache.tag[0][3] ), .B(\myifu.myicache.tag[1][3] ), .S(fanout_net_44 ), .Z(_01930_ ) );
AOI21_X1 _09448_ ( .A(_01928_ ), .B1(_01929_ ), .B2(_01930_ ), .ZN(_01931_ ) );
INV_X1 _09449_ ( .A(\IF_ID_pc [18] ), .ZN(_01932_ ) );
MUX2_X1 _09450_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(fanout_net_44 ), .Z(_01933_ ) );
MUX2_X1 _09451_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(fanout_net_44 ), .Z(_01934_ ) );
MUX2_X2 _09452_ ( .A(_01933_ ), .B(_01934_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01935_ ) );
AOI22_X1 _09453_ ( .A1(_01931_ ), .A2(\IF_ID_pc [8] ), .B1(_01932_ ), .B2(_01935_ ), .ZN(_01936_ ) );
MUX2_X1 _09454_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(fanout_net_44 ), .Z(_01937_ ) );
AND2_X1 _09455_ ( .A1(_01937_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01938_ ) );
MUX2_X1 _09456_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(fanout_net_44 ), .Z(_01939_ ) );
AOI21_X1 _09457_ ( .A(_01938_ ), .B1(_01929_ ), .B2(_01939_ ), .ZN(_01940_ ) );
NAND2_X1 _09458_ ( .A1(_01940_ ), .A2(\IF_ID_pc [16] ), .ZN(_01941_ ) );
MUX2_X1 _09459_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(fanout_net_44 ), .Z(_01942_ ) );
OR2_X1 _09460_ ( .A1(_01942_ ), .A2(_01870_ ), .ZN(_01943_ ) );
MUX2_X1 _09461_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(fanout_net_44 ), .Z(_01944_ ) );
OAI21_X1 _09462_ ( .A(_01943_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01944_ ), .ZN(_01945_ ) );
OAI211_X1 _09463_ ( .A(_01936_ ), .B(_01941_ ), .C1(\IF_ID_pc [27] ), .C2(_01945_ ), .ZN(_01946_ ) );
MUX2_X1 _09464_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(fanout_net_44 ), .Z(_01947_ ) );
MUX2_X1 _09465_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(fanout_net_44 ), .Z(_01948_ ) );
MUX2_X1 _09466_ ( .A(_01947_ ), .B(_01948_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01949_ ) );
OR2_X1 _09467_ ( .A1(_01871_ ), .A2(\myifu.myicache.tag[1][12] ), .ZN(_01950_ ) );
OAI211_X1 _09468_ ( .A(_01950_ ), .B(_01929_ ), .C1(fanout_net_44 ), .C2(\myifu.myicache.tag[0][12] ), .ZN(_01951_ ) );
INV_X1 _09469_ ( .A(\IF_ID_pc [17] ), .ZN(_01952_ ) );
OR2_X1 _09470_ ( .A1(fanout_net_44 ), .A2(\myifu.myicache.tag[2][12] ), .ZN(_01953_ ) );
OAI211_X1 _09471_ ( .A(_01953_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01872_ ), .C2(\myifu.myicache.tag[3][12] ), .ZN(_01954_ ) );
AND3_X1 _09472_ ( .A1(_01951_ ), .A2(_01952_ ), .A3(_01954_ ), .ZN(_01955_ ) );
AOI21_X1 _09473_ ( .A(_01952_ ), .B1(_01951_ ), .B2(_01954_ ), .ZN(_01956_ ) );
MUX2_X1 _09474_ ( .A(\myifu.myicache.tag[2][20] ), .B(\myifu.myicache.tag[3][20] ), .S(fanout_net_44 ), .Z(_01957_ ) );
OR2_X2 _09475_ ( .A1(_01957_ ), .A2(_01870_ ), .ZN(_01958_ ) );
MUX2_X1 _09476_ ( .A(\myifu.myicache.tag[0][20] ), .B(\myifu.myicache.tag[1][20] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01959_ ) );
OAI21_X2 _09477_ ( .A(_01958_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01959_ ), .ZN(_01960_ ) );
INV_X1 _09478_ ( .A(_01960_ ), .ZN(_01961_ ) );
INV_X1 _09479_ ( .A(\IF_ID_pc [25] ), .ZN(_01962_ ) );
OAI221_X1 _09480_ ( .A(_01949_ ), .B1(_01955_ ), .B2(_01956_ ), .C1(_01961_ ), .C2(_01962_ ), .ZN(_01963_ ) );
NOR4_X4 _09481_ ( .A1(_01898_ ), .A2(_01926_ ), .A3(_01946_ ), .A4(_01963_ ), .ZN(_01964_ ) );
AND2_X1 _09482_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[3][6] ), .ZN(_01965_ ) );
AOI211_X1 _09483_ ( .A(_01929_ ), .B(_01965_ ), .C1(_01872_ ), .C2(\myifu.myicache.tag[2][6] ), .ZN(_01966_ ) );
AND2_X1 _09484_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[1][6] ), .ZN(_01967_ ) );
AOI211_X1 _09485_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B(_01967_ ), .C1(_01872_ ), .C2(\myifu.myicache.tag[0][6] ), .ZN(_01968_ ) );
NOR2_X1 _09486_ ( .A1(_01966_ ), .A2(_01968_ ), .ZN(_01969_ ) );
XNOR2_X1 _09487_ ( .A(_01969_ ), .B(\IF_ID_pc [11] ), .ZN(_01970_ ) );
INV_X1 _09488_ ( .A(\IF_ID_pc [28] ), .ZN(_01971_ ) );
OR2_X1 _09489_ ( .A1(_01871_ ), .A2(\myifu.myicache.tag[3][23] ), .ZN(_01972_ ) );
OAI211_X1 _09490_ ( .A(_01972_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[2][23] ), .ZN(_01973_ ) );
OR2_X1 _09491_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][23] ), .ZN(_01974_ ) );
OAI211_X1 _09492_ ( .A(_01974_ ), .B(_01929_ ), .C1(_01872_ ), .C2(\myifu.myicache.tag[1][23] ), .ZN(_01975_ ) );
NAND2_X1 _09493_ ( .A1(_01973_ ), .A2(_01975_ ), .ZN(_01976_ ) );
MUX2_X1 _09494_ ( .A(\myifu.myicache.tag[2][5] ), .B(\myifu.myicache.tag[3][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01977_ ) );
OR2_X1 _09495_ ( .A1(_01977_ ), .A2(_01870_ ), .ZN(_01978_ ) );
MUX2_X1 _09496_ ( .A(\myifu.myicache.tag[0][5] ), .B(\myifu.myicache.tag[1][5] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01979_ ) );
OAI21_X1 _09497_ ( .A(_01978_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01979_ ), .ZN(_01980_ ) );
OAI221_X1 _09498_ ( .A(_01970_ ), .B1(_01971_ ), .B2(_01976_ ), .C1(\IF_ID_pc [10] ), .C2(_01980_ ), .ZN(_01981_ ) );
MUX2_X1 _09499_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01982_ ) );
AND2_X1 _09500_ ( .A1(_01982_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01983_ ) );
MUX2_X1 _09501_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01984_ ) );
AOI21_X1 _09502_ ( .A(_01983_ ), .B1(_01929_ ), .B2(_01984_ ), .ZN(_01985_ ) );
OR2_X1 _09503_ ( .A1(_01985_ ), .A2(\IF_ID_pc [23] ), .ZN(_01986_ ) );
OAI221_X1 _09504_ ( .A(_01986_ ), .B1(\IF_ID_pc [16] ), .B2(_01940_ ), .C1(\IF_ID_pc [8] ), .C2(_01931_ ), .ZN(_01987_ ) );
INV_X1 _09505_ ( .A(\IF_ID_pc [30] ), .ZN(_01988_ ) );
OR2_X4 _09506_ ( .A1(_01871_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_01989_ ) );
OAI211_X2 _09507_ ( .A(_01989_ ), .B(_01929_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_01990_ ) );
OR2_X1 _09508_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][25] ), .ZN(_01991_ ) );
OAI211_X1 _09509_ ( .A(_01991_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01872_ ), .C2(\myifu.myicache.tag[3][25] ), .ZN(_01992_ ) );
NAND2_X1 _09510_ ( .A1(_01990_ ), .A2(_01992_ ), .ZN(_01993_ ) );
AOI22_X1 _09511_ ( .A1(_01980_ ), .A2(\IF_ID_pc [10] ), .B1(_01988_ ), .B2(_01993_ ), .ZN(_01994_ ) );
NAND2_X1 _09512_ ( .A1(_01976_ ), .A2(_01971_ ), .ZN(_01995_ ) );
OAI211_X1 _09513_ ( .A(_01994_ ), .B(_01995_ ), .C1(_01988_ ), .C2(_01993_ ), .ZN(_01996_ ) );
MUX2_X1 _09514_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01997_ ) );
OR2_X1 _09515_ ( .A1(_01997_ ), .A2(_01870_ ), .ZN(_01998_ ) );
MUX2_X1 _09516_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01999_ ) );
OAI21_X1 _09517_ ( .A(_01998_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_01999_ ), .ZN(_02000_ ) );
MUX2_X1 _09518_ ( .A(\myifu.myicache.tag[0][7] ), .B(\myifu.myicache.tag[1][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02001_ ) );
MUX2_X1 _09519_ ( .A(\myifu.myicache.tag[2][7] ), .B(\myifu.myicache.tag[3][7] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02002_ ) );
MUX2_X2 _09520_ ( .A(_02001_ ), .B(_02002_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02003_ ) );
INV_X1 _09521_ ( .A(\IF_ID_pc [12] ), .ZN(_02004_ ) );
AOI22_X2 _09522_ ( .A1(_02000_ ), .A2(\IF_ID_pc [20] ), .B1(_02003_ ), .B2(_02004_ ), .ZN(_02005_ ) );
MUX2_X1 _09523_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02006_ ) );
OR2_X1 _09524_ ( .A1(_02006_ ), .A2(_01929_ ), .ZN(_02007_ ) );
MUX2_X1 _09525_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02008_ ) );
OAI21_X1 _09526_ ( .A(_02007_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B2(_02008_ ), .ZN(_02009_ ) );
NAND2_X1 _09527_ ( .A1(_02009_ ), .A2(\IF_ID_pc [14] ), .ZN(_02010_ ) );
OAI211_X1 _09528_ ( .A(_02005_ ), .B(_02010_ ), .C1(_01932_ ), .C2(_01935_ ), .ZN(_02011_ ) );
NOR4_X2 _09529_ ( .A1(_01981_ ), .A2(_01987_ ), .A3(_01996_ ), .A4(_02011_ ), .ZN(_02012_ ) );
NOR2_X1 _09530_ ( .A1(_02003_ ), .A2(_02004_ ), .ZN(_02013_ ) );
AOI21_X1 _09531_ ( .A(_02013_ ), .B1(\IF_ID_pc [23] ), .B2(_01985_ ), .ZN(_02014_ ) );
OAI221_X1 _09532_ ( .A(_02014_ ), .B1(\IF_ID_pc [14] ), .B2(_02009_ ), .C1(\IF_ID_pc [20] ), .C2(_02000_ ), .ZN(_02015_ ) );
MUX2_X1 _09533_ ( .A(\myifu.myicache.tag[0][2] ), .B(\myifu.myicache.tag[1][2] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02016_ ) );
NAND2_X1 _09534_ ( .A1(_02016_ ), .A2(_01929_ ), .ZN(_02017_ ) );
MUX2_X1 _09535_ ( .A(\myifu.myicache.tag[2][2] ), .B(\myifu.myicache.tag[3][2] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02018_ ) );
NAND2_X1 _09536_ ( .A1(_02018_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_02019_ ) );
NAND2_X1 _09537_ ( .A1(_02017_ ), .A2(_02019_ ), .ZN(_02020_ ) );
INV_X1 _09538_ ( .A(\IF_ID_pc [7] ), .ZN(_02021_ ) );
AOI22_X1 _09539_ ( .A1(_01961_ ), .A2(_01962_ ), .B1(_02020_ ), .B2(_02021_ ), .ZN(_02022_ ) );
OR2_X1 _09540_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][19] ), .ZN(_02023_ ) );
OAI211_X1 _09541_ ( .A(_02023_ ), .B(_01929_ ), .C1(_01872_ ), .C2(\myifu.myicache.tag[1][19] ), .ZN(_02024_ ) );
OR2_X1 _09542_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][19] ), .ZN(_02025_ ) );
OAI211_X1 _09543_ ( .A(_02025_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01872_ ), .C2(\myifu.myicache.tag[3][19] ), .ZN(_02026_ ) );
NAND2_X1 _09544_ ( .A1(_02024_ ), .A2(_02026_ ), .ZN(_02027_ ) );
INV_X1 _09545_ ( .A(\IF_ID_pc [24] ), .ZN(_02028_ ) );
NAND2_X1 _09546_ ( .A1(_02027_ ), .A2(_02028_ ), .ZN(_02029_ ) );
OAI211_X1 _09547_ ( .A(_02022_ ), .B(_02029_ ), .C1(_02021_ ), .C2(_02020_ ), .ZN(_02030_ ) );
INV_X1 _09548_ ( .A(\IF_ID_pc [21] ), .ZN(_02031_ ) );
MUX2_X1 _09549_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02032_ ) );
MUX2_X1 _09550_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02033_ ) );
MUX2_X2 _09551_ ( .A(_02032_ ), .B(_02033_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02034_ ) );
AOI22_X1 _09552_ ( .A1(_01945_ ), .A2(\IF_ID_pc [27] ), .B1(_02031_ ), .B2(_02034_ ), .ZN(_02035_ ) );
MUX2_X1 _09553_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02036_ ) );
MUX2_X1 _09554_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02037_ ) );
MUX2_X1 _09555_ ( .A(_02036_ ), .B(_02037_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02038_ ) );
INV_X1 _09556_ ( .A(\IF_ID_pc [29] ), .ZN(_02039_ ) );
NAND2_X1 _09557_ ( .A1(_02038_ ), .A2(_02039_ ), .ZN(_02040_ ) );
OAI211_X1 _09558_ ( .A(_02035_ ), .B(_02040_ ), .C1(_02028_ ), .C2(_02027_ ), .ZN(_02041_ ) );
OR2_X1 _09559_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][14] ), .ZN(_02042_ ) );
OAI211_X1 _09560_ ( .A(_02042_ ), .B(_01870_ ), .C1(_01872_ ), .C2(\myifu.myicache.tag[1][14] ), .ZN(_02043_ ) );
OR2_X1 _09561_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][14] ), .ZN(_02044_ ) );
OAI211_X1 _09562_ ( .A(_02044_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01872_ ), .C2(\myifu.myicache.tag[3][14] ), .ZN(_02045_ ) );
NAND2_X1 _09563_ ( .A1(_02043_ ), .A2(_02045_ ), .ZN(_02046_ ) );
XNOR2_X1 _09564_ ( .A(_02046_ ), .B(\IF_ID_pc [19] ), .ZN(_02047_ ) );
OAI221_X1 _09565_ ( .A(_02047_ ), .B1(_02039_ ), .B2(_02038_ ), .C1(_02031_ ), .C2(_02034_ ), .ZN(_02048_ ) );
NOR4_X2 _09566_ ( .A1(_02015_ ), .A2(_02030_ ), .A3(_02041_ ), .A4(_02048_ ), .ZN(_02049_ ) );
NAND3_X2 _09567_ ( .A1(_01964_ ), .A2(_02012_ ), .A3(_02049_ ), .ZN(_02050_ ) );
AND2_X4 _09568_ ( .A1(_02050_ ), .A2(\myifu.state [0] ), .ZN(_02051_ ) );
INV_X1 _09569_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_02052_ ) );
NOR2_X4 _09570_ ( .A1(_02051_ ), .A2(_02052_ ), .ZN(_02053_ ) );
NOR2_X1 _09571_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_02054_ ) );
NOR2_X4 _09572_ ( .A1(_02053_ ), .A2(_02054_ ), .ZN(_02055_ ) );
INV_X1 _09573_ ( .A(\EX_LS_flag [2] ), .ZN(_02056_ ) );
NAND4_X1 _09574_ ( .A1(_02056_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(EXU_valid_LSU ), .ZN(_02057_ ) );
NOR2_X1 _09575_ ( .A1(_02057_ ), .A2(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02058_ ) );
INV_X1 _09576_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_02059_ ) );
NOR2_X1 _09577_ ( .A1(_02058_ ), .A2(_02059_ ), .ZN(_02060_ ) );
NOR2_X4 _09578_ ( .A1(_02055_ ), .A2(_02060_ ), .ZN(_02061_ ) );
BUF_X8 _09579_ ( .A(_02061_ ), .Z(_02062_ ) );
OR3_X1 _09580_ ( .A1(_02057_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02063_ ) );
BUF_X4 _09581_ ( .A(_02058_ ), .Z(_02064_ ) );
OAI211_X1 _09582_ ( .A(_02062_ ), .B(_02063_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_02064_ ), .ZN(_02065_ ) );
INV_X4 _09583_ ( .A(_02055_ ), .ZN(_02066_ ) );
OAI21_X1 _09584_ ( .A(_02065_ ), .B1(_01952_ ), .B2(_02066_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09585_ ( .A1(_02057_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02067_ ) );
OAI211_X1 _09586_ ( .A(_02062_ ), .B(_02067_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_02064_ ), .ZN(_02068_ ) );
OAI21_X1 _09587_ ( .A(_02068_ ), .B1(_01932_ ), .B2(_02066_ ), .ZN(\io_master_araddr [18] ) );
OR3_X1 _09588_ ( .A1(_02057_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02069_ ) );
OAI211_X1 _09589_ ( .A(_02062_ ), .B(_02069_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_02064_ ), .ZN(_02070_ ) );
INV_X1 _09590_ ( .A(\IF_ID_pc [20] ), .ZN(_02071_ ) );
OAI21_X1 _09591_ ( .A(_02070_ ), .B1(_02071_ ), .B2(_02066_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09592_ ( .A1(_02057_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02072_ ) );
OAI211_X1 _09593_ ( .A(_02061_ ), .B(_02072_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_02064_ ), .ZN(_02073_ ) );
INV_X1 _09594_ ( .A(\IF_ID_pc [23] ), .ZN(_02074_ ) );
OAI21_X2 _09595_ ( .A(_02073_ ), .B1(_02074_ ), .B2(_02066_ ), .ZN(\io_master_araddr [23] ) );
OR4_X2 _09596_ ( .A1(\io_master_araddr [17] ), .A2(\io_master_araddr [18] ), .A3(\io_master_araddr [20] ), .A4(\io_master_araddr [23] ), .ZN(_02075_ ) );
BUF_X4 _09597_ ( .A(_02062_ ), .Z(_02076_ ) );
CLKBUF_X2 _09598_ ( .A(_02057_ ), .Z(_02077_ ) );
OR3_X1 _09599_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02078_ ) );
BUF_X4 _09600_ ( .A(_02064_ ), .Z(_02079_ ) );
OAI211_X1 _09601_ ( .A(_02076_ ), .B(_02078_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_02079_ ), .ZN(_02080_ ) );
OAI21_X1 _09602_ ( .A(_02080_ ), .B1(_01881_ ), .B2(_02066_ ), .ZN(\io_master_araddr [22] ) );
OR3_X1 _09603_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02081_ ) );
OAI211_X1 _09604_ ( .A(_02062_ ), .B(_02081_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_02064_ ), .ZN(_02082_ ) );
OAI21_X1 _09605_ ( .A(_02082_ ), .B1(_02031_ ), .B2(_02066_ ), .ZN(\io_master_araddr [21] ) );
OR3_X2 _09606_ ( .A1(_02075_ ), .A2(\io_master_araddr [22] ), .A3(\io_master_araddr [21] ), .ZN(_02083_ ) );
OR3_X1 _09607_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02084_ ) );
OAI211_X1 _09608_ ( .A(_02076_ ), .B(_02084_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_02079_ ), .ZN(_02085_ ) );
INV_X1 _09609_ ( .A(\IF_ID_pc [16] ), .ZN(_02086_ ) );
BUF_X4 _09610_ ( .A(_02066_ ), .Z(_02087_ ) );
OAI21_X1 _09611_ ( .A(_02085_ ), .B1(_02086_ ), .B2(_02087_ ), .ZN(\io_master_araddr [16] ) );
OR3_X1 _09612_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02088_ ) );
OAI211_X1 _09613_ ( .A(_02076_ ), .B(_02088_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_02079_ ), .ZN(_02089_ ) );
INV_X1 _09614_ ( .A(\IF_ID_pc [19] ), .ZN(_02090_ ) );
OAI21_X1 _09615_ ( .A(_02089_ ), .B1(_02090_ ), .B2(_02087_ ), .ZN(\io_master_araddr [19] ) );
OR3_X4 _09616_ ( .A1(_02083_ ), .A2(\io_master_araddr [16] ), .A3(\io_master_araddr [19] ), .ZN(_02091_ ) );
NOR3_X1 _09617_ ( .A1(_02053_ ), .A2(_01962_ ), .A3(_02054_ ), .ZN(_02092_ ) );
MUX2_X1 _09618_ ( .A(\mylsu.araddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_02058_ ), .Z(_02093_ ) );
AOI21_X2 _09619_ ( .A(_02092_ ), .B1(_02062_ ), .B2(_02093_ ), .ZN(_02094_ ) );
INV_X2 _09620_ ( .A(_02094_ ), .ZN(\io_master_araddr [25] ) );
OR3_X1 _09621_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02095_ ) );
OAI211_X1 _09622_ ( .A(_02062_ ), .B(_02095_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_02064_ ), .ZN(_02096_ ) );
OAI221_X1 _09623_ ( .A(\IF_ID_pc [27] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02051_ ), .C2(_02052_ ), .ZN(_02097_ ) );
NAND3_X2 _09624_ ( .A1(\io_master_araddr [25] ), .A2(_02096_ ), .A3(_02097_ ), .ZN(_02098_ ) );
OR3_X1 _09625_ ( .A1(_02057_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02099_ ) );
OAI211_X1 _09626_ ( .A(_02062_ ), .B(_02099_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_02064_ ), .ZN(_02100_ ) );
OAI21_X1 _09627_ ( .A(_02100_ ), .B1(_01903_ ), .B2(_02066_ ), .ZN(\io_master_araddr [26] ) );
OR3_X1 _09628_ ( .A1(_02057_ ), .A2(\EX_LS_dest_csreg_mem [24] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02101_ ) );
OAI211_X1 _09629_ ( .A(_02062_ ), .B(_02101_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_02064_ ), .ZN(_02102_ ) );
OAI21_X1 _09630_ ( .A(_02102_ ), .B1(_02028_ ), .B2(_02066_ ), .ZN(\io_master_araddr [24] ) );
OR3_X4 _09631_ ( .A1(_02098_ ), .A2(\io_master_araddr [26] ), .A3(\io_master_araddr [24] ), .ZN(_02103_ ) );
OR3_X1 _09632_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02104_ ) );
OAI211_X1 _09633_ ( .A(_02076_ ), .B(_02104_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_02079_ ), .ZN(_02105_ ) );
OAI21_X1 _09634_ ( .A(_02105_ ), .B1(_01918_ ), .B2(_02066_ ), .ZN(\io_master_araddr [31] ) );
OR3_X1 _09635_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02106_ ) );
OAI211_X1 _09636_ ( .A(_02062_ ), .B(_02106_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_02064_ ), .ZN(_02107_ ) );
OAI221_X1 _09637_ ( .A(\IF_ID_pc [28] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02051_ ), .C2(_02052_ ), .ZN(_02108_ ) );
AND2_X1 _09638_ ( .A1(_02107_ ), .A2(_02108_ ), .ZN(_02109_ ) );
INV_X1 _09639_ ( .A(_02109_ ), .ZN(\io_master_araddr [28] ) );
OR3_X4 _09640_ ( .A1(_02103_ ), .A2(\io_master_araddr [31] ), .A3(\io_master_araddr [28] ), .ZN(_02110_ ) );
OR3_X1 _09641_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02111_ ) );
OAI211_X1 _09642_ ( .A(_02076_ ), .B(_02111_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_02079_ ), .ZN(_02112_ ) );
OAI21_X1 _09643_ ( .A(_02112_ ), .B1(_01988_ ), .B2(_02087_ ), .ZN(\io_master_araddr [30] ) );
OR3_X1 _09644_ ( .A1(_02077_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_02113_ ) );
OAI211_X1 _09645_ ( .A(_02076_ ), .B(_02113_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_02079_ ), .ZN(_02114_ ) );
OAI221_X1 _09646_ ( .A(\IF_ID_pc [29] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_02051_ ), .C2(_02052_ ), .ZN(_02115_ ) );
AND2_X1 _09647_ ( .A1(_02114_ ), .A2(_02115_ ), .ZN(_02116_ ) );
INV_X1 _09648_ ( .A(_02116_ ), .ZN(\io_master_araddr [29] ) );
OR3_X4 _09649_ ( .A1(_02110_ ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [29] ), .ZN(_02117_ ) );
NOR2_X4 _09650_ ( .A1(_02091_ ), .A2(_02117_ ), .ZN(_02118_ ) );
BUF_X8 _09651_ ( .A(_02118_ ), .Z(_02119_ ) );
BUF_X2 _09652_ ( .A(_02119_ ), .Z(_02120_ ) );
BUF_X2 _09653_ ( .A(_02120_ ), .Z(_02121_ ) );
BUF_X2 _09654_ ( .A(_02121_ ), .Z(_02122_ ) );
CLKBUF_X2 _09655_ ( .A(_02055_ ), .Z(_02123_ ) );
CLKBUF_X2 _09656_ ( .A(_02123_ ), .Z(_02124_ ) );
CLKBUF_X2 _09657_ ( .A(_02124_ ), .Z(_02125_ ) );
OR2_X1 _09658_ ( .A1(\EX_LS_dest_csreg_mem [26] ), .A2(\EX_LS_dest_csreg_mem [24] ), .ZN(_02126_ ) );
OR3_X1 _09659_ ( .A1(_02126_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\EX_LS_dest_csreg_mem [25] ), .ZN(_02127_ ) );
OR4_X1 _09660_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(_02127_ ), .A3(\EX_LS_dest_csreg_mem [30] ), .A4(\EX_LS_dest_csreg_mem [29] ), .ZN(_02128_ ) );
OR2_X1 _09661_ ( .A1(_02128_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .ZN(_02129_ ) );
AND2_X4 _09662_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02130_ ) );
AND2_X4 _09663_ ( .A1(_02130_ ), .A2(_02056_ ), .ZN(_02131_ ) );
INV_X1 _09664_ ( .A(_02131_ ), .ZN(_02132_ ) );
NOR2_X1 _09665_ ( .A1(_02129_ ), .A2(_02132_ ), .ZN(_02133_ ) );
BUF_X4 _09666_ ( .A(_02131_ ), .Z(_02134_ ) );
NOR2_X1 _09667_ ( .A1(fanout_net_5 ), .A2(fanout_net_6 ), .ZN(_02135_ ) );
INV_X1 _09668_ ( .A(_02135_ ), .ZN(_02136_ ) );
INV_X1 _09669_ ( .A(\EX_LS_typ [1] ), .ZN(_02137_ ) );
INV_X1 _09670_ ( .A(\EX_LS_typ [3] ), .ZN(_02138_ ) );
NAND4_X1 _09671_ ( .A1(_02136_ ), .A2(_02137_ ), .A3(_02138_ ), .A4(\EX_LS_typ [2] ), .ZN(_02139_ ) );
AND2_X1 _09672_ ( .A1(fanout_net_5 ), .A2(\EX_LS_typ [1] ), .ZN(_02140_ ) );
NOR2_X1 _09673_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02141_ ) );
NAND2_X1 _09674_ ( .A1(_02140_ ), .A2(_02141_ ), .ZN(_02142_ ) );
AOI21_X1 _09675_ ( .A(\EX_LS_typ [0] ), .B1(_02139_ ), .B2(_02142_ ), .ZN(_02143_ ) );
AND3_X1 _09676_ ( .A1(_02140_ ), .A2(\EX_LS_typ [0] ), .A3(_02141_ ), .ZN(_02144_ ) );
OAI21_X1 _09677_ ( .A(_02134_ ), .B1(_02143_ ), .B2(_02144_ ), .ZN(_02145_ ) );
NOR2_X1 _09678_ ( .A1(_02145_ ), .A2(\EX_LS_typ [4] ), .ZN(_02146_ ) );
NOR2_X1 _09679_ ( .A1(_02133_ ), .A2(_02146_ ), .ZN(_02147_ ) );
INV_X32 _09680_ ( .A(\EX_LS_flag [1] ), .ZN(_02148_ ) );
NOR2_X4 _09681_ ( .A1(_02148_ ), .A2(\EX_LS_flag [0] ), .ZN(_02149_ ) );
AND2_X1 _09682_ ( .A1(_02149_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02150_ ) );
INV_X1 _09683_ ( .A(_02150_ ), .ZN(_02151_ ) );
NOR2_X1 _09684_ ( .A1(_02129_ ), .A2(_02151_ ), .ZN(_02152_ ) );
NAND3_X1 _09685_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02153_ ) );
OAI21_X1 _09686_ ( .A(_02142_ ), .B1(_02135_ ), .B2(_02153_ ), .ZN(_02154_ ) );
INV_X1 _09687_ ( .A(\EX_LS_typ [4] ), .ZN(_02155_ ) );
NAND3_X1 _09688_ ( .A1(_02056_ ), .A2(_02155_ ), .A3(\EX_LS_typ [0] ), .ZN(_02156_ ) );
NOR3_X1 _09689_ ( .A1(_02156_ ), .A2(_02148_ ), .A3(\EX_LS_flag [0] ), .ZN(_02157_ ) );
AND2_X1 _09690_ ( .A1(_02154_ ), .A2(_02157_ ), .ZN(_02158_ ) );
NOR2_X1 _09691_ ( .A1(_02152_ ), .A2(_02158_ ), .ZN(_02159_ ) );
AND2_X1 _09692_ ( .A1(_02147_ ), .A2(_02159_ ), .ZN(_02160_ ) );
AOI211_X1 _09693_ ( .A(_02059_ ), .B(_02125_ ), .C1(_02079_ ), .C2(_02160_ ), .ZN(_02161_ ) );
NOR2_X1 _09694_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02162_ ) );
AND3_X1 _09695_ ( .A1(_02050_ ), .A2(\myifu.state [0] ), .A3(_02162_ ), .ZN(_02163_ ) );
NOR4_X1 _09696_ ( .A1(_02053_ ), .A2(_02052_ ), .A3(_02054_ ), .A4(_02163_ ), .ZN(_02164_ ) );
NOR2_X1 _09697_ ( .A1(_02161_ ), .A2(_02164_ ), .ZN(_02165_ ) );
AND3_X1 _09698_ ( .A1(_02122_ ), .A2(\myclint.rvalid ), .A3(_02165_ ), .ZN(_02166_ ) );
AND2_X1 _09699_ ( .A1(_02096_ ), .A2(_02097_ ), .ZN(_02167_ ) );
INV_X1 _09700_ ( .A(_02167_ ), .ZN(\io_master_araddr [27] ) );
NOR4_X1 _09701_ ( .A1(\io_master_araddr [27] ), .A2(\io_master_araddr [28] ), .A3(\io_master_araddr [21] ), .A4(\io_master_araddr [18] ), .ZN(_02168_ ) );
NOR4_X1 _09702_ ( .A1(\io_master_araddr [24] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [23] ), .A4(\io_master_araddr [19] ), .ZN(_02169_ ) );
AND2_X1 _09703_ ( .A1(_02168_ ), .A2(_02169_ ), .ZN(_02170_ ) );
OR4_X1 _09704_ ( .A1(\io_master_araddr [29] ), .A2(\io_master_araddr [17] ), .A3(\io_master_araddr [22] ), .A4(\io_master_araddr [16] ), .ZN(_02171_ ) );
OR4_X1 _09705_ ( .A1(\io_master_araddr [31] ), .A2(\io_master_araddr [30] ), .A3(\io_master_araddr [26] ), .A4(_02094_ ), .ZN(_02172_ ) );
NOR2_X1 _09706_ ( .A1(_02171_ ), .A2(_02172_ ), .ZN(_02173_ ) );
AND2_X2 _09707_ ( .A1(_02170_ ), .A2(_02173_ ), .ZN(_02174_ ) );
INV_X1 _09708_ ( .A(_02174_ ), .ZN(_02175_ ) );
CLKBUF_X2 _09709_ ( .A(_02125_ ), .Z(_02176_ ) );
CLKBUF_X2 _09710_ ( .A(_02079_ ), .Z(_02177_ ) );
AOI21_X1 _09711_ ( .A(_02176_ ), .B1(_02177_ ), .B2(_02160_ ), .ZN(_02178_ ) );
AOI211_X1 _09712_ ( .A(_02054_ ), .B(_02053_ ), .C1(\myifu.state [0] ), .C2(_02162_ ), .ZN(_02179_ ) );
NOR3_X1 _09713_ ( .A1(_02175_ ), .A2(_02178_ ), .A3(_02179_ ), .ZN(_02180_ ) );
OAI21_X1 _09714_ ( .A(_01587_ ), .B1(_02180_ ), .B2(\myclint.rvalid ), .ZN(_02181_ ) );
NOR2_X1 _09715_ ( .A1(_02166_ ), .A2(_02181_ ), .ZN(_00065_ ) );
INV_X1 _09716_ ( .A(\LS_WB_wdata_csreg [30] ), .ZN(_02182_ ) );
NOR2_X1 _09717_ ( .A1(_02182_ ), .A2(fanout_net_2 ), .ZN(_00066_ ) );
INV_X1 _09718_ ( .A(\LS_WB_wdata_csreg [21] ), .ZN(_02183_ ) );
NOR2_X1 _09719_ ( .A1(_02183_ ), .A2(fanout_net_2 ), .ZN(_00067_ ) );
INV_X1 _09720_ ( .A(\LS_WB_wdata_csreg [20] ), .ZN(_02184_ ) );
NOR2_X1 _09721_ ( .A1(_02184_ ), .A2(fanout_net_2 ), .ZN(_00068_ ) );
INV_X1 _09722_ ( .A(\LS_WB_wdata_csreg [19] ), .ZN(_02185_ ) );
NOR2_X1 _09723_ ( .A1(_02185_ ), .A2(fanout_net_2 ), .ZN(_00069_ ) );
INV_X1 _09724_ ( .A(\LS_WB_wdata_csreg [18] ), .ZN(_02186_ ) );
NOR2_X1 _09725_ ( .A1(_02186_ ), .A2(fanout_net_2 ), .ZN(_00070_ ) );
INV_X1 _09726_ ( .A(\LS_WB_wdata_csreg [17] ), .ZN(_02187_ ) );
NOR2_X1 _09727_ ( .A1(_02187_ ), .A2(fanout_net_2 ), .ZN(_00071_ ) );
INV_X1 _09728_ ( .A(\LS_WB_wdata_csreg [16] ), .ZN(_02188_ ) );
NOR2_X1 _09729_ ( .A1(_02188_ ), .A2(fanout_net_2 ), .ZN(_00072_ ) );
INV_X1 _09730_ ( .A(\LS_WB_wdata_csreg [15] ), .ZN(_02189_ ) );
NOR2_X1 _09731_ ( .A1(_02189_ ), .A2(fanout_net_2 ), .ZN(_00073_ ) );
INV_X1 _09732_ ( .A(\LS_WB_wdata_csreg [14] ), .ZN(_02190_ ) );
NOR2_X1 _09733_ ( .A1(_02190_ ), .A2(fanout_net_2 ), .ZN(_00074_ ) );
INV_X1 _09734_ ( .A(\LS_WB_wdata_csreg [13] ), .ZN(_02191_ ) );
NOR2_X1 _09735_ ( .A1(_02191_ ), .A2(fanout_net_2 ), .ZN(_00075_ ) );
INV_X1 _09736_ ( .A(\LS_WB_wdata_csreg [12] ), .ZN(_02192_ ) );
NOR2_X1 _09737_ ( .A1(_02192_ ), .A2(fanout_net_2 ), .ZN(_00076_ ) );
INV_X1 _09738_ ( .A(\LS_WB_wdata_csreg [29] ), .ZN(_02193_ ) );
NOR2_X1 _09739_ ( .A1(_02193_ ), .A2(fanout_net_2 ), .ZN(_00077_ ) );
INV_X1 _09740_ ( .A(\LS_WB_wdata_csreg [11] ), .ZN(_02194_ ) );
NOR2_X1 _09741_ ( .A1(_02194_ ), .A2(fanout_net_2 ), .ZN(_00078_ ) );
INV_X1 _09742_ ( .A(\LS_WB_wdata_csreg [10] ), .ZN(_02195_ ) );
NOR2_X1 _09743_ ( .A1(_02195_ ), .A2(fanout_net_2 ), .ZN(_00079_ ) );
INV_X1 _09744_ ( .A(\LS_WB_wdata_csreg [9] ), .ZN(_02196_ ) );
NOR2_X1 _09745_ ( .A1(_02196_ ), .A2(fanout_net_2 ), .ZN(_00080_ ) );
INV_X1 _09746_ ( .A(\LS_WB_wdata_csreg [8] ), .ZN(_02197_ ) );
NOR2_X1 _09747_ ( .A1(_02197_ ), .A2(fanout_net_2 ), .ZN(_00081_ ) );
INV_X1 _09748_ ( .A(\LS_WB_wdata_csreg [7] ), .ZN(_02198_ ) );
NOR2_X1 _09749_ ( .A1(_02198_ ), .A2(fanout_net_2 ), .ZN(_00082_ ) );
INV_X1 _09750_ ( .A(\LS_WB_wdata_csreg [6] ), .ZN(_02199_ ) );
NOR2_X1 _09751_ ( .A1(_02199_ ), .A2(fanout_net_2 ), .ZN(_00083_ ) );
INV_X1 _09752_ ( .A(\LS_WB_wdata_csreg [5] ), .ZN(_02200_ ) );
NOR2_X1 _09753_ ( .A1(_02200_ ), .A2(fanout_net_2 ), .ZN(_00084_ ) );
INV_X1 _09754_ ( .A(\LS_WB_wdata_csreg [4] ), .ZN(_02201_ ) );
NOR2_X1 _09755_ ( .A1(_02201_ ), .A2(fanout_net_2 ), .ZN(_00085_ ) );
INV_X1 _09756_ ( .A(\LS_WB_wdata_csreg [3] ), .ZN(_02202_ ) );
NOR2_X1 _09757_ ( .A1(_02202_ ), .A2(fanout_net_2 ), .ZN(_00086_ ) );
INV_X1 _09758_ ( .A(\LS_WB_wdata_csreg [2] ), .ZN(_02203_ ) );
NOR2_X1 _09759_ ( .A1(_02203_ ), .A2(fanout_net_3 ), .ZN(_00087_ ) );
INV_X1 _09760_ ( .A(\LS_WB_wdata_csreg [28] ), .ZN(_02204_ ) );
NOR2_X1 _09761_ ( .A1(_02204_ ), .A2(fanout_net_3 ), .ZN(_00088_ ) );
INV_X1 _09762_ ( .A(\LS_WB_wdata_csreg [1] ), .ZN(_02205_ ) );
NOR2_X1 _09763_ ( .A1(_02205_ ), .A2(fanout_net_3 ), .ZN(_00089_ ) );
INV_X1 _09764_ ( .A(\LS_WB_wdata_csreg [0] ), .ZN(_02206_ ) );
NOR2_X1 _09765_ ( .A1(_02206_ ), .A2(fanout_net_3 ), .ZN(_00090_ ) );
INV_X1 _09766_ ( .A(\LS_WB_wdata_csreg [27] ), .ZN(_02207_ ) );
NOR2_X1 _09767_ ( .A1(_02207_ ), .A2(fanout_net_3 ), .ZN(_00091_ ) );
INV_X1 _09768_ ( .A(\LS_WB_wdata_csreg [26] ), .ZN(_02208_ ) );
NOR2_X1 _09769_ ( .A1(_02208_ ), .A2(fanout_net_3 ), .ZN(_00092_ ) );
INV_X1 _09770_ ( .A(\LS_WB_wdata_csreg [25] ), .ZN(_02209_ ) );
NOR2_X1 _09771_ ( .A1(_02209_ ), .A2(fanout_net_3 ), .ZN(_00093_ ) );
INV_X1 _09772_ ( .A(\LS_WB_wdata_csreg [24] ), .ZN(_02210_ ) );
NOR2_X1 _09773_ ( .A1(_02210_ ), .A2(fanout_net_3 ), .ZN(_00094_ ) );
INV_X1 _09774_ ( .A(\LS_WB_wdata_csreg [23] ), .ZN(_02211_ ) );
NOR2_X1 _09775_ ( .A1(_02211_ ), .A2(fanout_net_3 ), .ZN(_00095_ ) );
INV_X1 _09776_ ( .A(\LS_WB_wdata_csreg [22] ), .ZN(_02212_ ) );
NOR2_X1 _09777_ ( .A1(_02212_ ), .A2(fanout_net_3 ), .ZN(_00096_ ) );
NOR3_X1 _09778_ ( .A1(_01584_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00097_ ) );
NOR3_X1 _09779_ ( .A1(_02182_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00098_ ) );
NOR3_X1 _09780_ ( .A1(_02183_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00099_ ) );
NOR3_X1 _09781_ ( .A1(_02184_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00100_ ) );
NOR3_X1 _09782_ ( .A1(_02185_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00101_ ) );
NOR3_X1 _09783_ ( .A1(_02186_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00102_ ) );
NOR3_X1 _09784_ ( .A1(_02187_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00103_ ) );
NOR3_X1 _09785_ ( .A1(_02188_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00104_ ) );
NOR3_X1 _09786_ ( .A1(_02189_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00105_ ) );
NOR3_X1 _09787_ ( .A1(_02190_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00106_ ) );
NOR3_X1 _09788_ ( .A1(_02191_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00107_ ) );
NOR3_X1 _09789_ ( .A1(_02192_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00108_ ) );
NOR3_X1 _09790_ ( .A1(_02193_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00109_ ) );
NOR3_X1 _09791_ ( .A1(_02194_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00110_ ) );
NOR3_X1 _09792_ ( .A1(_02195_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00111_ ) );
NOR3_X1 _09793_ ( .A1(_02196_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00112_ ) );
NOR3_X1 _09794_ ( .A1(_02197_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00113_ ) );
NOR3_X1 _09795_ ( .A1(_02198_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00114_ ) );
NOR3_X1 _09796_ ( .A1(_02199_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00115_ ) );
NOR3_X1 _09797_ ( .A1(_02200_ ), .A2(fanout_net_3 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00116_ ) );
NOR3_X1 _09798_ ( .A1(_02201_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00117_ ) );
INV_X1 _09799_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02213_ ) );
NOR2_X1 _09800_ ( .A1(_02213_ ), .A2(\LS_WB_wen_csreg [3] ), .ZN(_02214_ ) );
AOI211_X1 _09801_ ( .A(fanout_net_4 ), .B(_02214_ ), .C1(_02202_ ), .C2(_02213_ ), .ZN(_00118_ ) );
NOR2_X1 _09802_ ( .A1(_02213_ ), .A2(\LS_WB_wen_csreg [2] ), .ZN(_02215_ ) );
AOI211_X1 _09803_ ( .A(fanout_net_4 ), .B(_02215_ ), .C1(_02203_ ), .C2(_02213_ ), .ZN(_00119_ ) );
NOR3_X1 _09804_ ( .A1(_02204_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00120_ ) );
NOR2_X1 _09805_ ( .A1(_02213_ ), .A2(\LS_WB_wen_csreg [1] ), .ZN(_02216_ ) );
AOI211_X1 _09806_ ( .A(fanout_net_4 ), .B(_02216_ ), .C1(_02205_ ), .C2(_02213_ ), .ZN(_00121_ ) );
NOR2_X1 _09807_ ( .A1(_02213_ ), .A2(\LS_WB_wen_csreg [0] ), .ZN(_02217_ ) );
AOI211_X1 _09808_ ( .A(fanout_net_4 ), .B(_02217_ ), .C1(_02206_ ), .C2(_02213_ ), .ZN(_00122_ ) );
NOR3_X1 _09809_ ( .A1(_02207_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00123_ ) );
NOR3_X1 _09810_ ( .A1(_02208_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00124_ ) );
NOR3_X1 _09811_ ( .A1(_02209_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00125_ ) );
NOR3_X1 _09812_ ( .A1(_02210_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00126_ ) );
NOR3_X1 _09813_ ( .A1(_02211_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00127_ ) );
NOR3_X1 _09814_ ( .A1(_02212_ ), .A2(fanout_net_4 ), .A3(\LS_WB_wen_csreg [6] ), .ZN(_00128_ ) );
AND3_X1 _09815_ ( .A1(_01748_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00129_ ) );
INV_X1 _09816_ ( .A(_02147_ ), .ZN(_02218_ ) );
INV_X1 _09817_ ( .A(_02159_ ), .ZN(_02219_ ) );
BUF_X2 _09818_ ( .A(_02219_ ), .Z(_02220_ ) );
NOR2_X1 _09819_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02221_ ) );
NAND2_X1 _09820_ ( .A1(_02221_ ), .A2(_01586_ ), .ZN(_02222_ ) );
OR2_X1 _09821_ ( .A1(\myexu.pc_jump [26] ), .A2(\myexu.pc_jump [25] ), .ZN(_02223_ ) );
OR3_X1 _09822_ ( .A1(_02223_ ), .A2(\myexu.pc_jump [27] ), .A3(\myexu.pc_jump [24] ), .ZN(_02224_ ) );
OR4_X1 _09823_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02225_ ) );
NOR2_X1 _09824_ ( .A1(_02224_ ), .A2(_02225_ ), .ZN(_02226_ ) );
NOR2_X1 _09825_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02227_ ) );
INV_X1 _09826_ ( .A(_02227_ ), .ZN(_02228_ ) );
NOR3_X1 _09827_ ( .A1(_02226_ ), .A2(exception_quest_IDU ), .A3(_02228_ ), .ZN(_02229_ ) );
NOR4_X1 _09828_ ( .A1(_02218_ ), .A2(_02220_ ), .A3(_02222_ ), .A4(_02229_ ), .ZN(_00130_ ) );
AOI21_X1 _09829_ ( .A(_02222_ ), .B1(_02160_ ), .B2(exception_quest_IDU ), .ZN(_00131_ ) );
AND2_X4 _09830_ ( .A1(_02148_ ), .A2(\EX_LS_flag [0] ), .ZN(_02230_ ) );
AND2_X1 _09831_ ( .A1(_02230_ ), .A2(\EX_LS_flag [2] ), .ZN(_02231_ ) );
AOI211_X2 _09832_ ( .A(_02131_ ), .B(_02231_ ), .C1(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .C2(_02230_ ), .ZN(_02232_ ) );
AND2_X2 _09833_ ( .A1(_02149_ ), .A2(\EX_LS_flag [2] ), .ZN(_02233_ ) );
INV_X4 _09834_ ( .A(_02233_ ), .ZN(_02234_ ) );
NAND2_X4 _09835_ ( .A1(_02232_ ), .A2(_02234_ ), .ZN(_02235_ ) );
XNOR2_X1 _09836_ ( .A(\ID_EX_rs1 [2] ), .B(\EX_LS_dest_reg [2] ), .ZN(_02236_ ) );
INV_X1 _09837_ ( .A(\EX_LS_dest_reg [3] ), .ZN(_02237_ ) );
NAND2_X1 _09838_ ( .A1(_02237_ ), .A2(\ID_EX_rs1 [3] ), .ZN(_02238_ ) );
INV_X16 _09839_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02239_ ) );
OR2_X1 _09840_ ( .A1(_02239_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02240_ ) );
NAND3_X1 _09841_ ( .A1(_02236_ ), .A2(_02238_ ), .A3(_02240_ ), .ZN(_02241_ ) );
XOR2_X2 _09842_ ( .A(\ID_EX_rs1 [4] ), .B(\EX_LS_dest_reg [4] ), .Z(_02242_ ) );
INV_X1 _09843_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .ZN(_02243_ ) );
NOR2_X1 _09844_ ( .A1(_02237_ ), .A2(\ID_EX_rs1 [3] ), .ZN(_02244_ ) );
NOR4_X2 _09845_ ( .A1(_02241_ ), .A2(_02242_ ), .A3(_02243_ ), .A4(_02244_ ), .ZN(_02245_ ) );
NAND2_X2 _09846_ ( .A1(_02235_ ), .A2(_02245_ ), .ZN(_02246_ ) );
CLKBUF_X3 _09847_ ( .A(_02246_ ), .Z(_02247_ ) );
XNOR2_X1 _09848_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .ZN(_02248_ ) );
NAND2_X1 _09849_ ( .A1(_02239_ ), .A2(\ID_EX_rs1 [1] ), .ZN(_02249_ ) );
OR3_X1 _09850_ ( .A1(\EX_LS_dest_reg [2] ), .A2(\EX_LS_dest_reg [1] ), .A3(\EX_LS_dest_reg [0] ), .ZN(_02250_ ) );
OR2_X1 _09851_ ( .A1(\EX_LS_dest_reg [4] ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02251_ ) );
OAI211_X1 _09852_ ( .A(_02248_ ), .B(_02249_ ), .C1(_02250_ ), .C2(_02251_ ), .ZN(_02252_ ) );
BUF_X2 _09853_ ( .A(_02252_ ), .Z(_02253_ ) );
NOR2_X1 _09854_ ( .A1(_02247_ ), .A2(_02253_ ), .ZN(_02254_ ) );
MUX2_X1 _09855_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02255_ ) );
MUX2_X1 _09856_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02256_ ) );
MUX2_X1 _09857_ ( .A(_02255_ ), .B(_02256_ ), .S(fanout_net_25 ), .Z(_02257_ ) );
INV_X1 _09858_ ( .A(fanout_net_28 ), .ZN(_02258_ ) );
BUF_X4 _09859_ ( .A(_02258_ ), .Z(_02259_ ) );
BUF_X4 _09860_ ( .A(_02259_ ), .Z(_02260_ ) );
BUF_X4 _09861_ ( .A(_02260_ ), .Z(_02261_ ) );
BUF_X4 _09862_ ( .A(_02261_ ), .Z(_02262_ ) );
NOR2_X1 _09863_ ( .A1(_02257_ ), .A2(_02262_ ), .ZN(_02263_ ) );
BUF_X4 _09864_ ( .A(_02262_ ), .Z(_02264_ ) );
OAI21_X1 _09865_ ( .A(fanout_net_25 ), .B1(fanout_net_17 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02265_ ) );
INV_X1 _09866_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02266_ ) );
AOI21_X1 _09867_ ( .A(_02265_ ), .B1(fanout_net_17 ), .B2(_02266_ ), .ZN(_02267_ ) );
INV_X1 _09868_ ( .A(fanout_net_25 ), .ZN(_02268_ ) );
BUF_X4 _09869_ ( .A(_02268_ ), .Z(_02269_ ) );
BUF_X4 _09870_ ( .A(_02269_ ), .Z(_02270_ ) );
BUF_X4 _09871_ ( .A(_02270_ ), .Z(_02271_ ) );
BUF_X4 _09872_ ( .A(_02271_ ), .Z(_02272_ ) );
BUF_X4 _09873_ ( .A(_02272_ ), .Z(_02273_ ) );
MUX2_X1 _09874_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02274_ ) );
AOI21_X1 _09875_ ( .A(_02267_ ), .B1(_02273_ ), .B2(_02274_ ), .ZN(_02275_ ) );
AOI211_X1 _09876_ ( .A(fanout_net_30 ), .B(_02263_ ), .C1(_02264_ ), .C2(_02275_ ), .ZN(_02276_ ) );
AND2_X1 _09877_ ( .A1(fanout_net_28 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02277_ ) );
BUF_X4 _09878_ ( .A(_02259_ ), .Z(_02278_ ) );
BUF_X4 _09879_ ( .A(_02278_ ), .Z(_02279_ ) );
AOI211_X1 _09880_ ( .A(fanout_net_17 ), .B(_02277_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02280_ ) );
INV_X1 _09881_ ( .A(fanout_net_17 ), .ZN(_02281_ ) );
BUF_X2 _09882_ ( .A(_02281_ ), .Z(_02282_ ) );
BUF_X4 _09883_ ( .A(_02282_ ), .Z(_02283_ ) );
BUF_X2 _09884_ ( .A(_02283_ ), .Z(_02284_ ) );
BUF_X2 _09885_ ( .A(_02284_ ), .Z(_02285_ ) );
AND2_X1 _09886_ ( .A1(fanout_net_28 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02286_ ) );
AOI211_X1 _09887_ ( .A(_02285_ ), .B(_02286_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02287_ ) );
OAI21_X1 _09888_ ( .A(fanout_net_25 ), .B1(_02280_ ), .B2(_02287_ ), .ZN(_02288_ ) );
AND2_X1 _09889_ ( .A1(fanout_net_28 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02289_ ) );
AOI211_X1 _09890_ ( .A(fanout_net_17 ), .B(_02289_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02290_ ) );
AND2_X1 _09891_ ( .A1(fanout_net_28 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02291_ ) );
AOI211_X1 _09892_ ( .A(_02285_ ), .B(_02291_ ), .C1(_02279_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02292_ ) );
OAI21_X1 _09893_ ( .A(_02273_ ), .B1(_02290_ ), .B2(_02292_ ), .ZN(_02293_ ) );
AND3_X1 _09894_ ( .A1(_02288_ ), .A2(_02293_ ), .A3(fanout_net_30 ), .ZN(_02294_ ) );
OR3_X1 _09895_ ( .A1(_02254_ ), .A2(_02276_ ), .A3(_02294_ ), .ZN(_02295_ ) );
OR3_X1 _09896_ ( .A1(_02247_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02253_ ), .ZN(_02296_ ) );
AND2_X2 _09897_ ( .A1(_02295_ ), .A2(_02296_ ), .ZN(_02297_ ) );
XOR2_X1 _09898_ ( .A(_02297_ ), .B(\ID_EX_imm [30] ), .Z(_02298_ ) );
OR2_X1 _09899_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02299_ ) );
BUF_X4 _09900_ ( .A(_02269_ ), .Z(_02300_ ) );
BUF_X4 _09901_ ( .A(_02300_ ), .Z(_02301_ ) );
BUF_X4 _09902_ ( .A(_02301_ ), .Z(_02302_ ) );
CLKBUF_X2 _09903_ ( .A(_02281_ ), .Z(_02303_ ) );
BUF_X2 _09904_ ( .A(_02303_ ), .Z(_02304_ ) );
BUF_X2 _09905_ ( .A(_02304_ ), .Z(_02305_ ) );
BUF_X4 _09906_ ( .A(_02305_ ), .Z(_02306_ ) );
OAI211_X1 _09907_ ( .A(_02299_ ), .B(_02302_ ), .C1(_02306_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02307_ ) );
INV_X1 _09908_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02308_ ) );
NAND2_X1 _09909_ ( .A1(_02308_ ), .A2(fanout_net_17 ), .ZN(_02309_ ) );
OAI211_X1 _09910_ ( .A(_02309_ ), .B(fanout_net_25 ), .C1(fanout_net_17 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02310_ ) );
NAND3_X1 _09911_ ( .A1(_02307_ ), .A2(_02310_ ), .A3(_02262_ ), .ZN(_02311_ ) );
MUX2_X1 _09912_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02312_ ) );
MUX2_X1 _09913_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02313_ ) );
MUX2_X1 _09914_ ( .A(_02312_ ), .B(_02313_ ), .S(_02272_ ), .Z(_02314_ ) );
BUF_X4 _09915_ ( .A(_02279_ ), .Z(_02315_ ) );
OAI211_X1 _09916_ ( .A(fanout_net_30 ), .B(_02311_ ), .C1(_02314_ ), .C2(_02315_ ), .ZN(_02316_ ) );
INV_X1 _09917_ ( .A(fanout_net_30 ), .ZN(_02317_ ) );
BUF_X4 _09918_ ( .A(_02317_ ), .Z(_02318_ ) );
BUF_X4 _09919_ ( .A(_02318_ ), .Z(_02319_ ) );
BUF_X4 _09920_ ( .A(_02319_ ), .Z(_02320_ ) );
OR2_X1 _09921_ ( .A1(fanout_net_17 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02321_ ) );
OAI211_X1 _09922_ ( .A(_02321_ ), .B(_02272_ ), .C1(_02306_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02322_ ) );
INV_X1 _09923_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02323_ ) );
NAND2_X1 _09924_ ( .A1(_02323_ ), .A2(fanout_net_17 ), .ZN(_02324_ ) );
OAI211_X1 _09925_ ( .A(_02324_ ), .B(fanout_net_25 ), .C1(fanout_net_17 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02325_ ) );
NAND3_X1 _09926_ ( .A1(_02322_ ), .A2(_02325_ ), .A3(_02262_ ), .ZN(_02326_ ) );
MUX2_X1 _09927_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02327_ ) );
MUX2_X1 _09928_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02328_ ) );
MUX2_X1 _09929_ ( .A(_02327_ ), .B(_02328_ ), .S(_02272_ ), .Z(_02329_ ) );
OAI211_X1 _09930_ ( .A(_02320_ ), .B(_02326_ ), .C1(_02329_ ), .C2(_02315_ ), .ZN(_02330_ ) );
NAND2_X1 _09931_ ( .A1(_02316_ ), .A2(_02330_ ), .ZN(_02331_ ) );
OR2_X1 _09932_ ( .A1(_02237_ ), .A2(\ID_EX_rs1 [3] ), .ZN(_02332_ ) );
NAND3_X1 _09933_ ( .A1(_02236_ ), .A2(_02332_ ), .A3(_02238_ ), .ZN(_02333_ ) );
NAND3_X1 _09934_ ( .A1(_02248_ ), .A2(_02249_ ), .A3(_02240_ ), .ZN(_02334_ ) );
NOR2_X1 _09935_ ( .A1(_02250_ ), .A2(_02251_ ), .ZN(_02335_ ) );
NOR4_X4 _09936_ ( .A1(_02333_ ), .A2(_02334_ ), .A3(_02335_ ), .A4(_02242_ ), .ZN(_02336_ ) );
NAND2_X2 _09937_ ( .A1(_02235_ ), .A2(_02336_ ), .ZN(_02337_ ) );
BUF_X4 _09938_ ( .A(_02337_ ), .Z(_02338_ ) );
BUF_X4 _09939_ ( .A(_02338_ ), .Z(_02339_ ) );
BUF_X4 _09940_ ( .A(_02243_ ), .Z(_02340_ ) );
BUF_X4 _09941_ ( .A(_02340_ ), .Z(_02341_ ) );
OAI21_X1 _09942_ ( .A(_02331_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_02342_ ) );
BUF_X4 _09943_ ( .A(_02235_ ), .Z(_02343_ ) );
BUF_X4 _09944_ ( .A(_02343_ ), .Z(_02344_ ) );
BUF_X4 _09945_ ( .A(_02336_ ), .Z(_02345_ ) );
BUF_X4 _09946_ ( .A(_02345_ ), .Z(_02346_ ) );
NAND4_X1 _09947_ ( .A1(_02344_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_02347_ ) );
AND2_X2 _09948_ ( .A1(_02342_ ), .A2(_02347_ ), .ZN(_02348_ ) );
INV_X1 _09949_ ( .A(\ID_EX_imm [27] ), .ZN(_02349_ ) );
XNOR2_X1 _09950_ ( .A(_02348_ ), .B(_02349_ ), .ZN(_02350_ ) );
OR3_X1 _09951_ ( .A1(_02246_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02252_ ), .ZN(_02351_ ) );
BUF_X2 _09952_ ( .A(_02282_ ), .Z(_02352_ ) );
BUF_X2 _09953_ ( .A(_02352_ ), .Z(_02353_ ) );
OR2_X1 _09954_ ( .A1(_02353_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02354_ ) );
OAI211_X1 _09955_ ( .A(_02354_ ), .B(_02272_ ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02355_ ) );
OR2_X1 _09956_ ( .A1(_02353_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02356_ ) );
OAI211_X1 _09957_ ( .A(_02356_ ), .B(fanout_net_25 ), .C1(fanout_net_17 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02357_ ) );
NAND3_X1 _09958_ ( .A1(_02355_ ), .A2(_02357_ ), .A3(fanout_net_28 ), .ZN(_02358_ ) );
MUX2_X1 _09959_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02359_ ) );
MUX2_X1 _09960_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02360_ ) );
MUX2_X1 _09961_ ( .A(_02359_ ), .B(_02360_ ), .S(_02272_ ), .Z(_02361_ ) );
OAI211_X1 _09962_ ( .A(_02319_ ), .B(_02358_ ), .C1(_02361_ ), .C2(fanout_net_28 ), .ZN(_02362_ ) );
NOR2_X1 _09963_ ( .A1(_02285_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02363_ ) );
OAI21_X1 _09964_ ( .A(fanout_net_25 ), .B1(fanout_net_17 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02364_ ) );
NOR2_X1 _09965_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02365_ ) );
OAI21_X1 _09966_ ( .A(_02272_ ), .B1(_02285_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02366_ ) );
OAI221_X1 _09967_ ( .A(_02279_ ), .B1(_02363_ ), .B2(_02364_ ), .C1(_02365_ ), .C2(_02366_ ), .ZN(_02367_ ) );
MUX2_X1 _09968_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02368_ ) );
MUX2_X1 _09969_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02369_ ) );
MUX2_X1 _09970_ ( .A(_02368_ ), .B(_02369_ ), .S(fanout_net_25 ), .Z(_02370_ ) );
OAI211_X1 _09971_ ( .A(fanout_net_30 ), .B(_02367_ ), .C1(_02370_ ), .C2(_02262_ ), .ZN(_02371_ ) );
OAI211_X1 _09972_ ( .A(_02362_ ), .B(_02371_ ), .C1(_02246_ ), .C2(_02253_ ), .ZN(_02372_ ) );
NAND2_X1 _09973_ ( .A1(_02351_ ), .A2(_02372_ ), .ZN(_02373_ ) );
XOR2_X1 _09974_ ( .A(_02373_ ), .B(\ID_EX_imm [22] ), .Z(_02374_ ) );
NOR2_X1 _09975_ ( .A1(_02305_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02375_ ) );
OAI21_X1 _09976_ ( .A(fanout_net_25 ), .B1(fanout_net_17 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02376_ ) );
NOR2_X1 _09977_ ( .A1(fanout_net_17 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02377_ ) );
OAI21_X1 _09978_ ( .A(_02301_ ), .B1(_02305_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02378_ ) );
OAI221_X1 _09979_ ( .A(_02261_ ), .B1(_02375_ ), .B2(_02376_ ), .C1(_02377_ ), .C2(_02378_ ), .ZN(_02379_ ) );
MUX2_X1 _09980_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02380_ ) );
MUX2_X1 _09981_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_17 ), .Z(_02381_ ) );
MUX2_X1 _09982_ ( .A(_02380_ ), .B(_02381_ ), .S(fanout_net_25 ), .Z(_02382_ ) );
OAI211_X1 _09983_ ( .A(fanout_net_30 ), .B(_02379_ ), .C1(_02382_ ), .C2(_02262_ ), .ZN(_02383_ ) );
OR2_X1 _09984_ ( .A1(_02284_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02384_ ) );
OAI211_X1 _09985_ ( .A(_02384_ ), .B(_02301_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02385_ ) );
OR2_X1 _09986_ ( .A1(_02284_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02386_ ) );
OAI211_X1 _09987_ ( .A(_02386_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02387_ ) );
NAND3_X1 _09988_ ( .A1(_02385_ ), .A2(_02387_ ), .A3(fanout_net_28 ), .ZN(_02388_ ) );
MUX2_X1 _09989_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02389_ ) );
MUX2_X1 _09990_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02390_ ) );
MUX2_X1 _09991_ ( .A(_02389_ ), .B(_02390_ ), .S(_02301_ ), .Z(_02391_ ) );
OAI211_X1 _09992_ ( .A(_02319_ ), .B(_02388_ ), .C1(_02391_ ), .C2(fanout_net_28 ), .ZN(_02392_ ) );
NAND2_X1 _09993_ ( .A1(_02383_ ), .A2(_02392_ ), .ZN(_02393_ ) );
OAI21_X1 _09994_ ( .A(_02393_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_02394_ ) );
NAND4_X1 _09995_ ( .A1(_02344_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_02395_ ) );
AND2_X2 _09996_ ( .A1(_02394_ ), .A2(_02395_ ), .ZN(_02396_ ) );
INV_X1 _09997_ ( .A(\ID_EX_imm [23] ), .ZN(_02397_ ) );
XNOR2_X1 _09998_ ( .A(_02396_ ), .B(_02397_ ), .ZN(_02398_ ) );
AND2_X1 _09999_ ( .A1(_02374_ ), .A2(_02398_ ), .ZN(_02399_ ) );
OR2_X1 _10000_ ( .A1(_02285_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02400_ ) );
BUF_X4 _10001_ ( .A(_02272_ ), .Z(_02401_ ) );
OAI211_X1 _10002_ ( .A(_02400_ ), .B(_02401_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02402_ ) );
OR2_X1 _10003_ ( .A1(_02305_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02403_ ) );
OAI211_X1 _10004_ ( .A(_02403_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02404_ ) );
NAND3_X1 _10005_ ( .A1(_02402_ ), .A2(_02404_ ), .A3(_02315_ ), .ZN(_02405_ ) );
MUX2_X1 _10006_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02406_ ) );
MUX2_X1 _10007_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02407_ ) );
MUX2_X1 _10008_ ( .A(_02406_ ), .B(_02407_ ), .S(_02302_ ), .Z(_02408_ ) );
OAI211_X1 _10009_ ( .A(fanout_net_30 ), .B(_02405_ ), .C1(_02408_ ), .C2(_02264_ ), .ZN(_02409_ ) );
OR2_X1 _10010_ ( .A1(_02285_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02410_ ) );
OAI211_X1 _10011_ ( .A(_02410_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02411_ ) );
OR2_X1 _10012_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02412_ ) );
OAI211_X1 _10013_ ( .A(_02412_ ), .B(_02302_ ), .C1(_02306_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02413_ ) );
NAND3_X1 _10014_ ( .A1(_02411_ ), .A2(_02262_ ), .A3(_02413_ ), .ZN(_02414_ ) );
MUX2_X1 _10015_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02415_ ) );
MUX2_X1 _10016_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02416_ ) );
MUX2_X1 _10017_ ( .A(_02415_ ), .B(_02416_ ), .S(_02302_ ), .Z(_02417_ ) );
OAI211_X1 _10018_ ( .A(_02320_ ), .B(_02414_ ), .C1(_02417_ ), .C2(_02315_ ), .ZN(_02418_ ) );
NAND2_X1 _10019_ ( .A1(_02409_ ), .A2(_02418_ ), .ZN(_02419_ ) );
OAI21_X1 _10020_ ( .A(_02419_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_02420_ ) );
NAND4_X1 _10021_ ( .A1(_02344_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_02421_ ) );
AND2_X2 _10022_ ( .A1(_02420_ ), .A2(_02421_ ), .ZN(_02422_ ) );
XOR2_X1 _10023_ ( .A(_02422_ ), .B(\ID_EX_imm [20] ), .Z(_02423_ ) );
OR2_X1 _10024_ ( .A1(_02305_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02424_ ) );
OAI211_X1 _10025_ ( .A(_02424_ ), .B(_02302_ ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02425_ ) );
OR2_X1 _10026_ ( .A1(_02305_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02426_ ) );
OAI211_X1 _10027_ ( .A(_02426_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02427_ ) );
NAND3_X1 _10028_ ( .A1(_02425_ ), .A2(_02427_ ), .A3(_02262_ ), .ZN(_02428_ ) );
MUX2_X1 _10029_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02429_ ) );
MUX2_X1 _10030_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02430_ ) );
MUX2_X1 _10031_ ( .A(_02429_ ), .B(_02430_ ), .S(_02302_ ), .Z(_02431_ ) );
OAI211_X1 _10032_ ( .A(_02320_ ), .B(_02428_ ), .C1(_02431_ ), .C2(_02315_ ), .ZN(_02432_ ) );
OR2_X1 _10033_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02433_ ) );
OAI211_X1 _10034_ ( .A(_02433_ ), .B(fanout_net_25 ), .C1(_02306_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02434_ ) );
OR2_X1 _10035_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02435_ ) );
OAI211_X1 _10036_ ( .A(_02435_ ), .B(_02302_ ), .C1(_02306_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02436_ ) );
NAND3_X1 _10037_ ( .A1(_02434_ ), .A2(_02436_ ), .A3(fanout_net_28 ), .ZN(_02437_ ) );
MUX2_X1 _10038_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02438_ ) );
MUX2_X1 _10039_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02439_ ) );
MUX2_X1 _10040_ ( .A(_02438_ ), .B(_02439_ ), .S(fanout_net_25 ), .Z(_02440_ ) );
OAI211_X1 _10041_ ( .A(fanout_net_30 ), .B(_02437_ ), .C1(_02440_ ), .C2(fanout_net_28 ), .ZN(_02441_ ) );
NAND2_X1 _10042_ ( .A1(_02432_ ), .A2(_02441_ ), .ZN(_02442_ ) );
OAI21_X1 _10043_ ( .A(_02442_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_02443_ ) );
NAND4_X1 _10044_ ( .A1(_02344_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_02444_ ) );
AND3_X1 _10045_ ( .A1(_02443_ ), .A2(\ID_EX_imm [21] ), .A3(_02444_ ), .ZN(_02445_ ) );
AOI21_X1 _10046_ ( .A(\ID_EX_imm [21] ), .B1(_02443_ ), .B2(_02444_ ), .ZN(_02446_ ) );
NOR2_X1 _10047_ ( .A1(_02445_ ), .A2(_02446_ ), .ZN(_02447_ ) );
AND2_X1 _10048_ ( .A1(_02423_ ), .A2(_02447_ ), .ZN(_02448_ ) );
AND2_X1 _10049_ ( .A1(_02399_ ), .A2(_02448_ ), .ZN(_02449_ ) );
OR2_X1 _10050_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02450_ ) );
BUF_X2 _10051_ ( .A(_02353_ ), .Z(_02451_ ) );
OAI211_X1 _10052_ ( .A(_02450_ ), .B(_02272_ ), .C1(_02451_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02452_ ) );
OR2_X1 _10053_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02453_ ) );
OAI211_X1 _10054_ ( .A(_02453_ ), .B(fanout_net_25 ), .C1(_02285_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02454_ ) );
NAND3_X1 _10055_ ( .A1(_02452_ ), .A2(_02454_ ), .A3(_02279_ ), .ZN(_02455_ ) );
MUX2_X1 _10056_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02456_ ) );
MUX2_X1 _10057_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02457_ ) );
MUX2_X1 _10058_ ( .A(_02456_ ), .B(_02457_ ), .S(_02301_ ), .Z(_02458_ ) );
OAI211_X1 _10059_ ( .A(_02319_ ), .B(_02455_ ), .C1(_02458_ ), .C2(_02262_ ), .ZN(_02459_ ) );
OR2_X1 _10060_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02460_ ) );
OAI211_X1 _10061_ ( .A(_02460_ ), .B(fanout_net_25 ), .C1(_02285_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02461_ ) );
OR2_X1 _10062_ ( .A1(fanout_net_18 ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02462_ ) );
OAI211_X1 _10063_ ( .A(_02462_ ), .B(_02272_ ), .C1(_02285_ ), .C2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02463_ ) );
NAND3_X1 _10064_ ( .A1(_02461_ ), .A2(_02463_ ), .A3(fanout_net_28 ), .ZN(_02464_ ) );
MUX2_X1 _10065_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02465_ ) );
MUX2_X1 _10066_ ( .A(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_18 ), .Z(_02466_ ) );
MUX2_X1 _10067_ ( .A(_02465_ ), .B(_02466_ ), .S(fanout_net_25 ), .Z(_02467_ ) );
OAI211_X1 _10068_ ( .A(fanout_net_30 ), .B(_02464_ ), .C1(_02467_ ), .C2(fanout_net_28 ), .ZN(_02468_ ) );
NAND2_X1 _10069_ ( .A1(_02459_ ), .A2(_02468_ ), .ZN(_02469_ ) );
OAI21_X1 _10070_ ( .A(_02469_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_02470_ ) );
NAND4_X1 _10071_ ( .A1(_02344_ ), .A2(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_02471_ ) );
AND2_X2 _10072_ ( .A1(_02470_ ), .A2(_02471_ ), .ZN(_02472_ ) );
INV_X1 _10073_ ( .A(\ID_EX_imm [16] ), .ZN(_02473_ ) );
XNOR2_X1 _10074_ ( .A(_02472_ ), .B(_02473_ ), .ZN(_02474_ ) );
INV_X1 _10075_ ( .A(_02474_ ), .ZN(_02475_ ) );
OR2_X1 _10076_ ( .A1(_02282_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02476_ ) );
OAI211_X1 _10077_ ( .A(_02476_ ), .B(fanout_net_25 ), .C1(fanout_net_18 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02477_ ) );
OR2_X1 _10078_ ( .A1(fanout_net_18 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02478_ ) );
BUF_X4 _10079_ ( .A(_02268_ ), .Z(_02479_ ) );
OAI211_X1 _10080_ ( .A(_02478_ ), .B(_02479_ ), .C1(_02283_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02480_ ) );
NAND3_X1 _10081_ ( .A1(_02477_ ), .A2(_02259_ ), .A3(_02480_ ), .ZN(_02481_ ) );
MUX2_X1 _10082_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02482_ ) );
MUX2_X1 _10083_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02483_ ) );
MUX2_X1 _10084_ ( .A(_02482_ ), .B(_02483_ ), .S(_02269_ ), .Z(_02484_ ) );
OAI211_X1 _10085_ ( .A(_02318_ ), .B(_02481_ ), .C1(_02484_ ), .C2(_02260_ ), .ZN(_02485_ ) );
OR2_X1 _10086_ ( .A1(_02282_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02486_ ) );
OAI211_X1 _10087_ ( .A(_02486_ ), .B(fanout_net_25 ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02487_ ) );
OR2_X1 _10088_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02488_ ) );
OAI211_X1 _10089_ ( .A(_02488_ ), .B(_02479_ ), .C1(_02283_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02489_ ) );
NAND3_X1 _10090_ ( .A1(_02487_ ), .A2(fanout_net_28 ), .A3(_02489_ ), .ZN(_02490_ ) );
MUX2_X1 _10091_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02491_ ) );
MUX2_X1 _10092_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02492_ ) );
MUX2_X1 _10093_ ( .A(_02491_ ), .B(_02492_ ), .S(fanout_net_25 ), .Z(_02493_ ) );
OAI211_X1 _10094_ ( .A(fanout_net_30 ), .B(_02490_ ), .C1(_02493_ ), .C2(fanout_net_28 ), .ZN(_02494_ ) );
NAND2_X1 _10095_ ( .A1(_02485_ ), .A2(_02494_ ), .ZN(_02495_ ) );
OAI21_X1 _10096_ ( .A(_02495_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02496_ ) );
NAND4_X1 _10097_ ( .A1(_02343_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02497_ ) );
AND2_X2 _10098_ ( .A1(_02496_ ), .A2(_02497_ ), .ZN(_02498_ ) );
INV_X1 _10099_ ( .A(\ID_EX_imm [8] ), .ZN(_02499_ ) );
XNOR2_X1 _10100_ ( .A(_02498_ ), .B(_02499_ ), .ZN(_02500_ ) );
OR2_X1 _10101_ ( .A1(_02282_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02501_ ) );
OAI211_X1 _10102_ ( .A(_02501_ ), .B(fanout_net_25 ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02502_ ) );
OR2_X1 _10103_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02503_ ) );
OAI211_X1 _10104_ ( .A(_02503_ ), .B(_02270_ ), .C1(_02352_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02504_ ) );
NAND3_X1 _10105_ ( .A1(_02502_ ), .A2(_02260_ ), .A3(_02504_ ), .ZN(_02505_ ) );
MUX2_X1 _10106_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02506_ ) );
MUX2_X1 _10107_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02507_ ) );
MUX2_X1 _10108_ ( .A(_02506_ ), .B(_02507_ ), .S(_02479_ ), .Z(_02508_ ) );
OAI211_X1 _10109_ ( .A(fanout_net_30 ), .B(_02505_ ), .C1(_02508_ ), .C2(_02278_ ), .ZN(_02509_ ) );
OR2_X1 _10110_ ( .A1(_02282_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02510_ ) );
OAI211_X1 _10111_ ( .A(_02510_ ), .B(_02270_ ), .C1(fanout_net_19 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02511_ ) );
OR2_X1 _10112_ ( .A1(fanout_net_19 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02512_ ) );
OAI211_X1 _10113_ ( .A(_02512_ ), .B(fanout_net_25 ), .C1(_02352_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02513_ ) );
NAND3_X1 _10114_ ( .A1(_02511_ ), .A2(_02260_ ), .A3(_02513_ ), .ZN(_02514_ ) );
MUX2_X1 _10115_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02515_ ) );
MUX2_X1 _10116_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02516_ ) );
MUX2_X1 _10117_ ( .A(_02515_ ), .B(_02516_ ), .S(_02479_ ), .Z(_02517_ ) );
OAI211_X1 _10118_ ( .A(_02318_ ), .B(_02514_ ), .C1(_02517_ ), .C2(_02278_ ), .ZN(_02518_ ) );
NAND2_X1 _10119_ ( .A1(_02509_ ), .A2(_02518_ ), .ZN(_02519_ ) );
OAI21_X4 _10120_ ( .A(_02519_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02520_ ) );
NAND4_X4 _10121_ ( .A1(_02343_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02521_ ) );
AND3_X1 _10122_ ( .A1(_02520_ ), .A2(\ID_EX_imm [9] ), .A3(_02521_ ), .ZN(_02522_ ) );
AOI21_X1 _10123_ ( .A(\ID_EX_imm [9] ), .B1(_02520_ ), .B2(_02521_ ), .ZN(_02523_ ) );
NOR2_X2 _10124_ ( .A1(_02522_ ), .A2(_02523_ ), .ZN(_02524_ ) );
AND2_X1 _10125_ ( .A1(_02500_ ), .A2(_02524_ ), .ZN(_02525_ ) );
OR2_X1 _10126_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02526_ ) );
OAI211_X1 _10127_ ( .A(_02526_ ), .B(_02300_ ), .C1(_02304_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02527_ ) );
OR2_X1 _10128_ ( .A1(fanout_net_19 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02528_ ) );
OAI211_X1 _10129_ ( .A(_02528_ ), .B(fanout_net_25 ), .C1(_02304_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02529_ ) );
NAND3_X1 _10130_ ( .A1(_02527_ ), .A2(_02529_ ), .A3(_02260_ ), .ZN(_02530_ ) );
MUX2_X1 _10131_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02531_ ) );
MUX2_X1 _10132_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02532_ ) );
MUX2_X1 _10133_ ( .A(_02531_ ), .B(_02532_ ), .S(_02270_ ), .Z(_02533_ ) );
OAI211_X1 _10134_ ( .A(_02318_ ), .B(_02530_ ), .C1(_02533_ ), .C2(_02261_ ), .ZN(_02534_ ) );
OR2_X1 _10135_ ( .A1(_02303_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02535_ ) );
OAI211_X1 _10136_ ( .A(_02535_ ), .B(fanout_net_25 ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02536_ ) );
OR2_X1 _10137_ ( .A1(_02303_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02537_ ) );
OAI211_X1 _10138_ ( .A(_02537_ ), .B(_02300_ ), .C1(fanout_net_19 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02538_ ) );
NAND3_X1 _10139_ ( .A1(_02536_ ), .A2(_02538_ ), .A3(fanout_net_28 ), .ZN(_02539_ ) );
MUX2_X1 _10140_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02540_ ) );
MUX2_X1 _10141_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02541_ ) );
MUX2_X1 _10142_ ( .A(_02540_ ), .B(_02541_ ), .S(fanout_net_25 ), .Z(_02542_ ) );
OAI211_X1 _10143_ ( .A(fanout_net_30 ), .B(_02539_ ), .C1(_02542_ ), .C2(fanout_net_28 ), .ZN(_02543_ ) );
NAND2_X1 _10144_ ( .A1(_02534_ ), .A2(_02543_ ), .ZN(_02544_ ) );
OAI21_X1 _10145_ ( .A(_02544_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02545_ ) );
NAND4_X1 _10146_ ( .A1(_02343_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02546_ ) );
AND3_X1 _10147_ ( .A1(_02545_ ), .A2(\ID_EX_imm [11] ), .A3(_02546_ ), .ZN(_02547_ ) );
AOI21_X1 _10148_ ( .A(\ID_EX_imm [11] ), .B1(_02545_ ), .B2(_02546_ ), .ZN(_02548_ ) );
NOR2_X1 _10149_ ( .A1(_02547_ ), .A2(_02548_ ), .ZN(_02549_ ) );
OR2_X1 _10150_ ( .A1(_02303_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02550_ ) );
OAI211_X1 _10151_ ( .A(_02550_ ), .B(_02300_ ), .C1(fanout_net_19 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02551_ ) );
OR2_X1 _10152_ ( .A1(_02303_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02552_ ) );
OAI211_X1 _10153_ ( .A(_02552_ ), .B(fanout_net_25 ), .C1(fanout_net_19 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02553_ ) );
NAND3_X1 _10154_ ( .A1(_02551_ ), .A2(_02553_ ), .A3(_02260_ ), .ZN(_02554_ ) );
MUX2_X1 _10155_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02555_ ) );
MUX2_X1 _10156_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02556_ ) );
MUX2_X1 _10157_ ( .A(_02555_ ), .B(_02556_ ), .S(_02270_ ), .Z(_02557_ ) );
OAI211_X1 _10158_ ( .A(_02318_ ), .B(_02554_ ), .C1(_02557_ ), .C2(_02278_ ), .ZN(_02558_ ) );
OR2_X1 _10159_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02559_ ) );
OAI211_X1 _10160_ ( .A(_02559_ ), .B(fanout_net_25 ), .C1(_02304_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02560_ ) );
OR2_X1 _10161_ ( .A1(fanout_net_19 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02561_ ) );
OAI211_X1 _10162_ ( .A(_02561_ ), .B(_02270_ ), .C1(_02304_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02562_ ) );
NAND3_X1 _10163_ ( .A1(_02560_ ), .A2(_02562_ ), .A3(fanout_net_28 ), .ZN(_02563_ ) );
MUX2_X1 _10164_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02564_ ) );
MUX2_X1 _10165_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_19 ), .Z(_02565_ ) );
MUX2_X1 _10166_ ( .A(_02564_ ), .B(_02565_ ), .S(fanout_net_26 ), .Z(_02566_ ) );
OAI211_X1 _10167_ ( .A(fanout_net_30 ), .B(_02563_ ), .C1(_02566_ ), .C2(fanout_net_28 ), .ZN(_02567_ ) );
NAND2_X1 _10168_ ( .A1(_02558_ ), .A2(_02567_ ), .ZN(_02568_ ) );
OAI21_X1 _10169_ ( .A(_02568_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02569_ ) );
NAND4_X1 _10170_ ( .A1(_02343_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02570_ ) );
AND2_X2 _10171_ ( .A1(_02569_ ), .A2(_02570_ ), .ZN(_02571_ ) );
INV_X1 _10172_ ( .A(\ID_EX_imm [10] ), .ZN(_02572_ ) );
XNOR2_X1 _10173_ ( .A(_02571_ ), .B(_02572_ ), .ZN(_02573_ ) );
AND3_X1 _10174_ ( .A1(_02525_ ), .A2(_02549_ ), .A3(_02573_ ), .ZN(_02574_ ) );
INV_X1 _10175_ ( .A(_02574_ ), .ZN(_02575_ ) );
OR2_X1 _10176_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02576_ ) );
OAI211_X1 _10177_ ( .A(_02576_ ), .B(fanout_net_26 ), .C1(_02303_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02577_ ) );
INV_X1 _10178_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02578_ ) );
NAND2_X1 _10179_ ( .A1(_02578_ ), .A2(fanout_net_20 ), .ZN(_02579_ ) );
OAI211_X1 _10180_ ( .A(_02579_ ), .B(_02269_ ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02580_ ) );
NAND3_X1 _10181_ ( .A1(_02577_ ), .A2(_02580_ ), .A3(_02259_ ), .ZN(_02581_ ) );
MUX2_X1 _10182_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02582_ ) );
MUX2_X1 _10183_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02583_ ) );
MUX2_X1 _10184_ ( .A(_02582_ ), .B(_02583_ ), .S(_02268_ ), .Z(_02584_ ) );
OAI211_X1 _10185_ ( .A(_02317_ ), .B(_02581_ ), .C1(_02584_ ), .C2(_02259_ ), .ZN(_02585_ ) );
OR2_X1 _10186_ ( .A1(_02281_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02586_ ) );
OAI211_X1 _10187_ ( .A(_02586_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02587_ ) );
OR2_X1 _10188_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02588_ ) );
OAI211_X1 _10189_ ( .A(_02588_ ), .B(_02269_ ), .C1(_02282_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02589_ ) );
NAND3_X1 _10190_ ( .A1(_02587_ ), .A2(fanout_net_28 ), .A3(_02589_ ), .ZN(_02590_ ) );
MUX2_X1 _10191_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02591_ ) );
MUX2_X1 _10192_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02592_ ) );
MUX2_X1 _10193_ ( .A(_02591_ ), .B(_02592_ ), .S(fanout_net_26 ), .Z(_02593_ ) );
OAI211_X1 _10194_ ( .A(fanout_net_30 ), .B(_02590_ ), .C1(_02593_ ), .C2(fanout_net_28 ), .ZN(_02594_ ) );
NAND2_X1 _10195_ ( .A1(_02585_ ), .A2(_02594_ ), .ZN(_02595_ ) );
OAI21_X1 _10196_ ( .A(_02595_ ), .B1(_02337_ ), .B2(_02243_ ), .ZN(_02596_ ) );
NAND4_X1 _10197_ ( .A1(_02235_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02336_ ), .ZN(_02597_ ) );
AND2_X2 _10198_ ( .A1(_02596_ ), .A2(_02597_ ), .ZN(_02598_ ) );
XNOR2_X2 _10199_ ( .A(_02598_ ), .B(\ID_EX_imm [5] ), .ZN(_02599_ ) );
INV_X1 _10200_ ( .A(\ID_EX_imm [4] ), .ZN(_02600_ ) );
OR2_X1 _10201_ ( .A1(_02281_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02601_ ) );
OAI211_X1 _10202_ ( .A(_02601_ ), .B(_02269_ ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02602_ ) );
OR2_X1 _10203_ ( .A1(_02281_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02603_ ) );
OAI211_X1 _10204_ ( .A(_02603_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02604_ ) );
NAND3_X1 _10205_ ( .A1(_02602_ ), .A2(_02604_ ), .A3(_02259_ ), .ZN(_02605_ ) );
MUX2_X1 _10206_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02606_ ) );
MUX2_X1 _10207_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02607_ ) );
MUX2_X1 _10208_ ( .A(_02606_ ), .B(_02607_ ), .S(_02269_ ), .Z(_02608_ ) );
OAI211_X1 _10209_ ( .A(_02317_ ), .B(_02605_ ), .C1(_02608_ ), .C2(_02260_ ), .ZN(_02609_ ) );
OR2_X1 _10210_ ( .A1(_02281_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02610_ ) );
OAI211_X1 _10211_ ( .A(_02610_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02611_ ) );
OR2_X1 _10212_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02612_ ) );
OAI211_X1 _10213_ ( .A(_02612_ ), .B(_02269_ ), .C1(_02303_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02613_ ) );
NAND3_X1 _10214_ ( .A1(_02611_ ), .A2(fanout_net_28 ), .A3(_02613_ ), .ZN(_02614_ ) );
MUX2_X1 _10215_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02615_ ) );
MUX2_X1 _10216_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02616_ ) );
MUX2_X1 _10217_ ( .A(_02615_ ), .B(_02616_ ), .S(fanout_net_26 ), .Z(_02617_ ) );
OAI211_X1 _10218_ ( .A(fanout_net_30 ), .B(_02614_ ), .C1(_02617_ ), .C2(fanout_net_28 ), .ZN(_02618_ ) );
NAND2_X1 _10219_ ( .A1(_02609_ ), .A2(_02618_ ), .ZN(_02619_ ) );
OAI21_X1 _10220_ ( .A(_02619_ ), .B1(_02337_ ), .B2(_02243_ ), .ZN(_02620_ ) );
NAND4_X1 _10221_ ( .A1(_02235_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02336_ ), .ZN(_02621_ ) );
AND2_X2 _10222_ ( .A1(_02620_ ), .A2(_02621_ ), .ZN(_02622_ ) );
INV_X1 _10223_ ( .A(_02622_ ), .ZN(_02623_ ) );
NOR3_X1 _10224_ ( .A1(_02599_ ), .A2(_02600_ ), .A3(_02623_ ), .ZN(_02624_ ) );
INV_X1 _10225_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02625_ ) );
AOI21_X1 _10226_ ( .A(_02624_ ), .B1(_02625_ ), .B2(_02598_ ), .ZN(_02626_ ) );
NOR2_X1 _10227_ ( .A1(_02352_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02627_ ) );
OAI21_X1 _10228_ ( .A(fanout_net_26 ), .B1(fanout_net_20 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02628_ ) );
NOR2_X1 _10229_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02629_ ) );
OAI21_X1 _10230_ ( .A(_02270_ ), .B1(_02352_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02630_ ) );
OAI221_X1 _10231_ ( .A(_02260_ ), .B1(_02627_ ), .B2(_02628_ ), .C1(_02629_ ), .C2(_02630_ ), .ZN(_02631_ ) );
MUX2_X1 _10232_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02632_ ) );
MUX2_X1 _10233_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02633_ ) );
MUX2_X1 _10234_ ( .A(_02632_ ), .B(_02633_ ), .S(fanout_net_26 ), .Z(_02634_ ) );
OAI211_X1 _10235_ ( .A(fanout_net_30 ), .B(_02631_ ), .C1(_02634_ ), .C2(_02278_ ), .ZN(_02635_ ) );
OR2_X1 _10236_ ( .A1(_02303_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02636_ ) );
OAI211_X1 _10237_ ( .A(_02636_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02637_ ) );
OR2_X1 _10238_ ( .A1(fanout_net_20 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02638_ ) );
OAI211_X1 _10239_ ( .A(_02638_ ), .B(_02300_ ), .C1(_02304_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02639_ ) );
NAND3_X1 _10240_ ( .A1(_02637_ ), .A2(fanout_net_28 ), .A3(_02639_ ), .ZN(_02640_ ) );
MUX2_X1 _10241_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02641_ ) );
MUX2_X1 _10242_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02642_ ) );
MUX2_X1 _10243_ ( .A(_02641_ ), .B(_02642_ ), .S(_02270_ ), .Z(_02643_ ) );
OAI211_X1 _10244_ ( .A(_02318_ ), .B(_02640_ ), .C1(_02643_ ), .C2(fanout_net_28 ), .ZN(_02644_ ) );
NAND2_X1 _10245_ ( .A1(_02635_ ), .A2(_02644_ ), .ZN(_02645_ ) );
OAI21_X1 _10246_ ( .A(_02645_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02646_ ) );
NAND4_X1 _10247_ ( .A1(_02343_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02647_ ) );
AND3_X1 _10248_ ( .A1(_02646_ ), .A2(\ID_EX_imm [7] ), .A3(_02647_ ), .ZN(_02648_ ) );
AOI21_X1 _10249_ ( .A(\ID_EX_imm [7] ), .B1(_02646_ ), .B2(_02647_ ), .ZN(_02649_ ) );
OR3_X1 _10250_ ( .A1(_02246_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02252_ ), .ZN(_02650_ ) );
OR2_X1 _10251_ ( .A1(_02282_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02651_ ) );
OAI211_X1 _10252_ ( .A(_02651_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02652_ ) );
OR2_X1 _10253_ ( .A1(fanout_net_20 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02653_ ) );
OAI211_X1 _10254_ ( .A(_02653_ ), .B(_02479_ ), .C1(_02283_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02654_ ) );
NAND3_X1 _10255_ ( .A1(_02652_ ), .A2(_02259_ ), .A3(_02654_ ), .ZN(_02655_ ) );
MUX2_X1 _10256_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02656_ ) );
MUX2_X1 _10257_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_20 ), .Z(_02657_ ) );
MUX2_X1 _10258_ ( .A(_02656_ ), .B(_02657_ ), .S(_02479_ ), .Z(_02658_ ) );
OAI211_X1 _10259_ ( .A(_02318_ ), .B(_02655_ ), .C1(_02658_ ), .C2(_02278_ ), .ZN(_02659_ ) );
OR2_X1 _10260_ ( .A1(_02282_ ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02660_ ) );
OAI211_X1 _10261_ ( .A(_02660_ ), .B(fanout_net_26 ), .C1(fanout_net_20 ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02661_ ) );
OR2_X1 _10262_ ( .A1(fanout_net_21 ), .A2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02662_ ) );
OAI211_X1 _10263_ ( .A(_02662_ ), .B(_02479_ ), .C1(_02283_ ), .C2(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02663_ ) );
NAND3_X1 _10264_ ( .A1(_02661_ ), .A2(fanout_net_28 ), .A3(_02663_ ), .ZN(_02664_ ) );
MUX2_X1 _10265_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02665_ ) );
MUX2_X1 _10266_ ( .A(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02666_ ) );
MUX2_X1 _10267_ ( .A(_02665_ ), .B(_02666_ ), .S(fanout_net_26 ), .Z(_02667_ ) );
OAI211_X1 _10268_ ( .A(fanout_net_30 ), .B(_02664_ ), .C1(_02667_ ), .C2(fanout_net_28 ), .ZN(_02668_ ) );
OAI211_X1 _10269_ ( .A(_02659_ ), .B(_02668_ ), .C1(_02246_ ), .C2(_02252_ ), .ZN(_02669_ ) );
NAND2_X1 _10270_ ( .A1(_02650_ ), .A2(_02669_ ), .ZN(_02670_ ) );
INV_X1 _10271_ ( .A(\ID_EX_imm [6] ), .ZN(_02671_ ) );
XNOR2_X1 _10272_ ( .A(_02670_ ), .B(_02671_ ), .ZN(_02672_ ) );
INV_X1 _10273_ ( .A(_02672_ ), .ZN(_02673_ ) );
NOR4_X2 _10274_ ( .A1(_02626_ ), .A2(_02648_ ), .A3(_02649_ ), .A4(_02673_ ), .ZN(_02674_ ) );
NAND2_X1 _10275_ ( .A1(_02670_ ), .A2(\ID_EX_imm [6] ), .ZN(_02675_ ) );
NOR3_X1 _10276_ ( .A1(_02675_ ), .A2(_02648_ ), .A3(_02649_ ), .ZN(_02676_ ) );
NOR3_X1 _10277_ ( .A1(_02674_ ), .A2(_02648_ ), .A3(_02676_ ), .ZN(_02677_ ) );
XNOR2_X1 _10278_ ( .A(_02622_ ), .B(_02600_ ), .ZN(_02678_ ) );
INV_X1 _10279_ ( .A(_02678_ ), .ZN(_02679_ ) );
NOR2_X1 _10280_ ( .A1(_02679_ ), .A2(_02599_ ), .ZN(_02680_ ) );
NOR2_X1 _10281_ ( .A1(_02648_ ), .A2(_02649_ ), .ZN(_02681_ ) );
AND3_X1 _10282_ ( .A1(_02680_ ), .A2(_02681_ ), .A3(_02672_ ), .ZN(_02682_ ) );
OR2_X1 _10283_ ( .A1(_02281_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02683_ ) );
OAI211_X1 _10284_ ( .A(_02683_ ), .B(_02268_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02684_ ) );
OR2_X1 _10285_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02685_ ) );
OAI211_X1 _10286_ ( .A(_02685_ ), .B(fanout_net_26 ), .C1(_02281_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02686_ ) );
NAND3_X1 _10287_ ( .A1(_02684_ ), .A2(_02258_ ), .A3(_02686_ ), .ZN(_02687_ ) );
MUX2_X1 _10288_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02688_ ) );
MUX2_X1 _10289_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02689_ ) );
MUX2_X1 _10290_ ( .A(_02688_ ), .B(_02689_ ), .S(_02268_ ), .Z(_02690_ ) );
OAI211_X1 _10291_ ( .A(_02317_ ), .B(_02687_ ), .C1(_02690_ ), .C2(_02259_ ), .ZN(_02691_ ) );
OR2_X1 _10292_ ( .A1(_02281_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02692_ ) );
OAI211_X1 _10293_ ( .A(_02692_ ), .B(fanout_net_26 ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02693_ ) );
OR2_X1 _10294_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02694_ ) );
OAI211_X1 _10295_ ( .A(_02694_ ), .B(_02268_ ), .C1(_02281_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02695_ ) );
NAND3_X1 _10296_ ( .A1(_02693_ ), .A2(fanout_net_28 ), .A3(_02695_ ), .ZN(_02696_ ) );
MUX2_X1 _10297_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02697_ ) );
MUX2_X1 _10298_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02698_ ) );
MUX2_X1 _10299_ ( .A(_02697_ ), .B(_02698_ ), .S(fanout_net_26 ), .Z(_02699_ ) );
OAI211_X1 _10300_ ( .A(fanout_net_30 ), .B(_02696_ ), .C1(_02699_ ), .C2(fanout_net_28 ), .ZN(_02700_ ) );
NAND2_X1 _10301_ ( .A1(_02691_ ), .A2(_02700_ ), .ZN(_02701_ ) );
OAI21_X1 _10302_ ( .A(_02701_ ), .B1(_02337_ ), .B2(_02243_ ), .ZN(_02702_ ) );
NAND4_X1 _10303_ ( .A1(_02235_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02336_ ), .ZN(_02703_ ) );
AND2_X2 _10304_ ( .A1(_02702_ ), .A2(_02703_ ), .ZN(_02704_ ) );
INV_X1 _10305_ ( .A(\ID_EX_imm [1] ), .ZN(_02705_ ) );
XNOR2_X2 _10306_ ( .A(_02704_ ), .B(_02705_ ), .ZN(_02706_ ) );
OR2_X1 _10307_ ( .A1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .A2(fanout_net_21 ), .ZN(_02707_ ) );
OAI211_X1 _10308_ ( .A(_02707_ ), .B(_02479_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .C2(_02303_ ), .ZN(_02708_ ) );
OR2_X1 _10309_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02709_ ) );
OAI211_X1 _10310_ ( .A(_02709_ ), .B(fanout_net_26 ), .C1(_02283_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02710_ ) );
NAND3_X1 _10311_ ( .A1(_02708_ ), .A2(_02710_ ), .A3(_02259_ ), .ZN(_02711_ ) );
MUX2_X1 _10312_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02712_ ) );
MUX2_X1 _10313_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02713_ ) );
MUX2_X1 _10314_ ( .A(_02712_ ), .B(_02713_ ), .S(_02269_ ), .Z(_02714_ ) );
OAI211_X1 _10315_ ( .A(_02318_ ), .B(_02711_ ), .C1(_02714_ ), .C2(_02260_ ), .ZN(_02715_ ) );
OR2_X1 _10316_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02716_ ) );
OAI211_X1 _10317_ ( .A(_02716_ ), .B(fanout_net_26 ), .C1(_02283_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02717_ ) );
OR2_X1 _10318_ ( .A1(fanout_net_21 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02718_ ) );
OAI211_X1 _10319_ ( .A(_02718_ ), .B(_02269_ ), .C1(_02283_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02719_ ) );
NAND3_X1 _10320_ ( .A1(_02717_ ), .A2(_02719_ ), .A3(fanout_net_28 ), .ZN(_02720_ ) );
MUX2_X1 _10321_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02721_ ) );
MUX2_X1 _10322_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02722_ ) );
MUX2_X1 _10323_ ( .A(_02721_ ), .B(_02722_ ), .S(fanout_net_26 ), .Z(_02723_ ) );
OAI211_X1 _10324_ ( .A(fanout_net_30 ), .B(_02720_ ), .C1(_02723_ ), .C2(fanout_net_29 ), .ZN(_02724_ ) );
NAND2_X1 _10325_ ( .A1(_02715_ ), .A2(_02724_ ), .ZN(_02725_ ) );
OAI21_X1 _10326_ ( .A(_02725_ ), .B1(_02337_ ), .B2(_02243_ ), .ZN(_02726_ ) );
NAND4_X1 _10327_ ( .A1(_02235_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02336_ ), .ZN(_02727_ ) );
AND3_X1 _10328_ ( .A1(_02726_ ), .A2(\ID_EX_imm [0] ), .A3(_02727_ ), .ZN(_02728_ ) );
AND2_X1 _10329_ ( .A1(_02706_ ), .A2(_02728_ ), .ZN(_02729_ ) );
AOI21_X2 _10330_ ( .A(_02729_ ), .B1(\ID_EX_imm [1] ), .B2(_02704_ ), .ZN(_02730_ ) );
OR3_X1 _10331_ ( .A1(_02246_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02252_ ), .ZN(_02731_ ) );
OR2_X1 _10332_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02732_ ) );
OAI211_X1 _10333_ ( .A(_02732_ ), .B(_02300_ ), .C1(_02304_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02733_ ) );
OR2_X1 _10334_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02734_ ) );
OAI211_X1 _10335_ ( .A(_02734_ ), .B(fanout_net_26 ), .C1(_02304_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02735_ ) );
NAND3_X1 _10336_ ( .A1(_02733_ ), .A2(_02735_ ), .A3(fanout_net_29 ), .ZN(_02736_ ) );
MUX2_X1 _10337_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02737_ ) );
MUX2_X1 _10338_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02738_ ) );
MUX2_X1 _10339_ ( .A(_02737_ ), .B(_02738_ ), .S(_02270_ ), .Z(_02739_ ) );
OAI211_X1 _10340_ ( .A(_02318_ ), .B(_02736_ ), .C1(_02739_ ), .C2(fanout_net_29 ), .ZN(_02740_ ) );
NOR2_X1 _10341_ ( .A1(_02352_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02741_ ) );
OAI21_X1 _10342_ ( .A(fanout_net_26 ), .B1(fanout_net_21 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02742_ ) );
INV_X1 _10343_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02743_ ) );
INV_X1 _10344_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02744_ ) );
MUX2_X1 _10345_ ( .A(_02743_ ), .B(_02744_ ), .S(fanout_net_21 ), .Z(_02745_ ) );
OAI221_X1 _10346_ ( .A(_02260_ ), .B1(_02741_ ), .B2(_02742_ ), .C1(_02745_ ), .C2(fanout_net_26 ), .ZN(_02746_ ) );
MUX2_X1 _10347_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02747_ ) );
MUX2_X1 _10348_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02748_ ) );
MUX2_X1 _10349_ ( .A(_02747_ ), .B(_02748_ ), .S(fanout_net_26 ), .Z(_02749_ ) );
OAI211_X1 _10350_ ( .A(fanout_net_30 ), .B(_02746_ ), .C1(_02749_ ), .C2(_02278_ ), .ZN(_02750_ ) );
OAI211_X1 _10351_ ( .A(_02740_ ), .B(_02750_ ), .C1(_02246_ ), .C2(_02252_ ), .ZN(_02751_ ) );
NAND2_X4 _10352_ ( .A1(_02731_ ), .A2(_02751_ ), .ZN(_02752_ ) );
XNOR2_X1 _10353_ ( .A(_02752_ ), .B(\ID_EX_imm [3] ), .ZN(_02753_ ) );
OR3_X1 _10354_ ( .A1(_02246_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02252_ ), .ZN(_02754_ ) );
OR2_X1 _10355_ ( .A1(_02303_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02755_ ) );
OAI211_X1 _10356_ ( .A(_02755_ ), .B(_02270_ ), .C1(fanout_net_21 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02756_ ) );
OR2_X1 _10357_ ( .A1(_02282_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02757_ ) );
OAI211_X1 _10358_ ( .A(_02757_ ), .B(fanout_net_26 ), .C1(fanout_net_21 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02758_ ) );
NAND3_X1 _10359_ ( .A1(_02756_ ), .A2(_02758_ ), .A3(fanout_net_29 ), .ZN(_02759_ ) );
MUX2_X1 _10360_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02760_ ) );
MUX2_X1 _10361_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02761_ ) );
MUX2_X1 _10362_ ( .A(_02760_ ), .B(_02761_ ), .S(_02479_ ), .Z(_02762_ ) );
OAI211_X1 _10363_ ( .A(_02318_ ), .B(_02759_ ), .C1(_02762_ ), .C2(fanout_net_29 ), .ZN(_02763_ ) );
NOR2_X1 _10364_ ( .A1(_02283_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02764_ ) );
OAI21_X1 _10365_ ( .A(fanout_net_26 ), .B1(fanout_net_22 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02765_ ) );
NOR2_X1 _10366_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02766_ ) );
OAI21_X1 _10367_ ( .A(_02479_ ), .B1(_02283_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02767_ ) );
OAI221_X1 _10368_ ( .A(_02259_ ), .B1(_02764_ ), .B2(_02765_ ), .C1(_02766_ ), .C2(_02767_ ), .ZN(_02768_ ) );
MUX2_X1 _10369_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02769_ ) );
MUX2_X1 _10370_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02770_ ) );
MUX2_X1 _10371_ ( .A(_02769_ ), .B(_02770_ ), .S(fanout_net_26 ), .Z(_02771_ ) );
OAI211_X1 _10372_ ( .A(fanout_net_30 ), .B(_02768_ ), .C1(_02771_ ), .C2(_02278_ ), .ZN(_02772_ ) );
OAI211_X1 _10373_ ( .A(_02763_ ), .B(_02772_ ), .C1(_02246_ ), .C2(_02252_ ), .ZN(_02773_ ) );
NAND2_X2 _10374_ ( .A1(_02754_ ), .A2(_02773_ ), .ZN(_02774_ ) );
INV_X1 _10375_ ( .A(\ID_EX_imm [2] ), .ZN(_02775_ ) );
XNOR2_X1 _10376_ ( .A(_02774_ ), .B(_02775_ ), .ZN(_02776_ ) );
INV_X1 _10377_ ( .A(_02776_ ), .ZN(_02777_ ) );
NOR3_X2 _10378_ ( .A1(_02730_ ), .A2(_02753_ ), .A3(_02777_ ), .ZN(_02778_ ) );
AND2_X1 _10379_ ( .A1(_02774_ ), .A2(\ID_EX_imm [2] ), .ZN(_02779_ ) );
INV_X1 _10380_ ( .A(_02779_ ), .ZN(_02780_ ) );
INV_X1 _10381_ ( .A(_02752_ ), .ZN(_02781_ ) );
OAI22_X1 _10382_ ( .A1(_02753_ ), .A2(_02780_ ), .B1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B2(_02781_ ), .ZN(_02782_ ) );
OAI21_X1 _10383_ ( .A(_02682_ ), .B1(_02778_ ), .B2(_02782_ ), .ZN(_02783_ ) );
AOI21_X2 _10384_ ( .A(_02575_ ), .B1(_02677_ ), .B2(_02783_ ), .ZN(_02784_ ) );
AND2_X1 _10385_ ( .A1(_02498_ ), .A2(\ID_EX_imm [8] ), .ZN(_02785_ ) );
AOI21_X1 _10386_ ( .A(_02522_ ), .B1(_02785_ ), .B2(_02524_ ), .ZN(_02786_ ) );
INV_X1 _10387_ ( .A(_02786_ ), .ZN(_02787_ ) );
NAND3_X1 _10388_ ( .A1(_02787_ ), .A2(_02549_ ), .A3(_02573_ ), .ZN(_02788_ ) );
AND2_X1 _10389_ ( .A1(_02571_ ), .A2(\ID_EX_imm [10] ), .ZN(_02789_ ) );
AOI21_X1 _10390_ ( .A(_02547_ ), .B1(_02789_ ), .B2(_02549_ ), .ZN(_02790_ ) );
AND2_X1 _10391_ ( .A1(_02788_ ), .A2(_02790_ ), .ZN(_02791_ ) );
INV_X1 _10392_ ( .A(_02791_ ), .ZN(_02792_ ) );
NOR2_X2 _10393_ ( .A1(_02784_ ), .A2(_02792_ ), .ZN(_02793_ ) );
NOR2_X1 _10394_ ( .A1(_02284_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02794_ ) );
OAI21_X1 _10395_ ( .A(fanout_net_26 ), .B1(fanout_net_22 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02795_ ) );
NOR2_X1 _10396_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02796_ ) );
OAI21_X1 _10397_ ( .A(_02300_ ), .B1(_02284_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02797_ ) );
OAI221_X1 _10398_ ( .A(_02278_ ), .B1(_02794_ ), .B2(_02795_ ), .C1(_02796_ ), .C2(_02797_ ), .ZN(_02798_ ) );
MUX2_X1 _10399_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02799_ ) );
MUX2_X1 _10400_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02800_ ) );
MUX2_X1 _10401_ ( .A(_02799_ ), .B(_02800_ ), .S(fanout_net_26 ), .Z(_02801_ ) );
OAI211_X1 _10402_ ( .A(fanout_net_30 ), .B(_02798_ ), .C1(_02801_ ), .C2(_02261_ ), .ZN(_02802_ ) );
OR2_X1 _10403_ ( .A1(_02352_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02803_ ) );
OAI211_X1 _10404_ ( .A(_02803_ ), .B(fanout_net_26 ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02804_ ) );
OR2_X1 _10405_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02805_ ) );
OAI211_X1 _10406_ ( .A(_02805_ ), .B(_02271_ ), .C1(_02284_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02806_ ) );
NAND3_X1 _10407_ ( .A1(_02804_ ), .A2(fanout_net_29 ), .A3(_02806_ ), .ZN(_02807_ ) );
MUX2_X1 _10408_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02808_ ) );
MUX2_X1 _10409_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02809_ ) );
MUX2_X1 _10410_ ( .A(_02808_ ), .B(_02809_ ), .S(_02300_ ), .Z(_02810_ ) );
OAI211_X1 _10411_ ( .A(_02319_ ), .B(_02807_ ), .C1(_02810_ ), .C2(fanout_net_29 ), .ZN(_02811_ ) );
NAND2_X1 _10412_ ( .A1(_02802_ ), .A2(_02811_ ), .ZN(_02812_ ) );
OAI21_X1 _10413_ ( .A(_02812_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02813_ ) );
NAND4_X1 _10414_ ( .A1(_02343_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02814_ ) );
AND2_X2 _10415_ ( .A1(_02813_ ), .A2(_02814_ ), .ZN(_02815_ ) );
XOR2_X1 _10416_ ( .A(_02815_ ), .B(\ID_EX_imm [15] ), .Z(_02816_ ) );
OR2_X1 _10417_ ( .A1(_02352_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02817_ ) );
OAI211_X1 _10418_ ( .A(_02817_ ), .B(_02271_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02818_ ) );
OR2_X1 _10419_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02819_ ) );
OAI211_X1 _10420_ ( .A(_02819_ ), .B(fanout_net_26 ), .C1(_02353_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02820_ ) );
NAND3_X1 _10421_ ( .A1(_02818_ ), .A2(_02261_ ), .A3(_02820_ ), .ZN(_02821_ ) );
MUX2_X1 _10422_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02822_ ) );
MUX2_X1 _10423_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02823_ ) );
MUX2_X1 _10424_ ( .A(_02822_ ), .B(_02823_ ), .S(_02271_ ), .Z(_02824_ ) );
OAI211_X1 _10425_ ( .A(_02319_ ), .B(_02821_ ), .C1(_02824_ ), .C2(_02279_ ), .ZN(_02825_ ) );
OR2_X1 _10426_ ( .A1(_02352_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02826_ ) );
OAI211_X1 _10427_ ( .A(_02826_ ), .B(_02271_ ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02827_ ) );
OR2_X1 _10428_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02828_ ) );
OAI211_X1 _10429_ ( .A(_02828_ ), .B(fanout_net_27 ), .C1(_02353_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02829_ ) );
NAND3_X1 _10430_ ( .A1(_02827_ ), .A2(fanout_net_29 ), .A3(_02829_ ), .ZN(_02830_ ) );
MUX2_X1 _10431_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02831_ ) );
MUX2_X1 _10432_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02832_ ) );
MUX2_X1 _10433_ ( .A(_02831_ ), .B(_02832_ ), .S(fanout_net_27 ), .Z(_02833_ ) );
OAI211_X1 _10434_ ( .A(fanout_net_30 ), .B(_02830_ ), .C1(_02833_ ), .C2(fanout_net_29 ), .ZN(_02834_ ) );
NAND2_X1 _10435_ ( .A1(_02825_ ), .A2(_02834_ ), .ZN(_02835_ ) );
OAI21_X1 _10436_ ( .A(_02835_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02836_ ) );
NAND4_X1 _10437_ ( .A1(_02343_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02837_ ) );
AND2_X2 _10438_ ( .A1(_02836_ ), .A2(_02837_ ), .ZN(_02838_ ) );
XOR2_X1 _10439_ ( .A(_02838_ ), .B(\ID_EX_imm [14] ), .Z(_02839_ ) );
AND2_X1 _10440_ ( .A1(_02816_ ), .A2(_02839_ ), .ZN(_02840_ ) );
NOR2_X1 _10441_ ( .A1(_02304_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02841_ ) );
OAI21_X1 _10442_ ( .A(fanout_net_27 ), .B1(fanout_net_22 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02842_ ) );
NOR2_X1 _10443_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02843_ ) );
OAI21_X1 _10444_ ( .A(_02300_ ), .B1(_02284_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02844_ ) );
OAI221_X1 _10445_ ( .A(_02278_ ), .B1(_02841_ ), .B2(_02842_ ), .C1(_02843_ ), .C2(_02844_ ), .ZN(_02845_ ) );
MUX2_X1 _10446_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02846_ ) );
MUX2_X1 _10447_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02847_ ) );
MUX2_X1 _10448_ ( .A(_02846_ ), .B(_02847_ ), .S(fanout_net_27 ), .Z(_02848_ ) );
OAI211_X1 _10449_ ( .A(fanout_net_30 ), .B(_02845_ ), .C1(_02848_ ), .C2(_02261_ ), .ZN(_02849_ ) );
OR2_X1 _10450_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02850_ ) );
OAI211_X1 _10451_ ( .A(_02850_ ), .B(_02271_ ), .C1(_02284_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02851_ ) );
OR2_X1 _10452_ ( .A1(fanout_net_22 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02852_ ) );
OAI211_X1 _10453_ ( .A(_02852_ ), .B(fanout_net_27 ), .C1(_02284_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02853_ ) );
NAND3_X1 _10454_ ( .A1(_02851_ ), .A2(_02853_ ), .A3(fanout_net_29 ), .ZN(_02854_ ) );
MUX2_X1 _10455_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02855_ ) );
MUX2_X1 _10456_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02856_ ) );
MUX2_X1 _10457_ ( .A(_02855_ ), .B(_02856_ ), .S(_02300_ ), .Z(_02857_ ) );
OAI211_X1 _10458_ ( .A(_02319_ ), .B(_02854_ ), .C1(_02857_ ), .C2(fanout_net_29 ), .ZN(_02858_ ) );
NAND2_X1 _10459_ ( .A1(_02849_ ), .A2(_02858_ ), .ZN(_02859_ ) );
OAI21_X1 _10460_ ( .A(_02859_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02860_ ) );
NAND4_X1 _10461_ ( .A1(_02343_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02861_ ) );
AND3_X1 _10462_ ( .A1(_02860_ ), .A2(\ID_EX_imm [13] ), .A3(_02861_ ), .ZN(_02862_ ) );
AOI21_X1 _10463_ ( .A(\ID_EX_imm [13] ), .B1(_02860_ ), .B2(_02861_ ), .ZN(_02863_ ) );
NOR2_X1 _10464_ ( .A1(_02862_ ), .A2(_02863_ ), .ZN(_02864_ ) );
OR2_X1 _10465_ ( .A1(_02352_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02865_ ) );
OAI211_X1 _10466_ ( .A(_02865_ ), .B(fanout_net_27 ), .C1(fanout_net_22 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02866_ ) );
OR2_X1 _10467_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02867_ ) );
OAI211_X1 _10468_ ( .A(_02867_ ), .B(_02271_ ), .C1(_02353_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02868_ ) );
NAND3_X1 _10469_ ( .A1(_02866_ ), .A2(_02261_ ), .A3(_02868_ ), .ZN(_02869_ ) );
MUX2_X1 _10470_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02870_ ) );
MUX2_X1 _10471_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02871_ ) );
MUX2_X1 _10472_ ( .A(_02870_ ), .B(_02871_ ), .S(_02271_ ), .Z(_02872_ ) );
OAI211_X1 _10473_ ( .A(_02319_ ), .B(_02869_ ), .C1(_02872_ ), .C2(_02261_ ), .ZN(_02873_ ) );
OR2_X1 _10474_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02874_ ) );
OAI211_X1 _10475_ ( .A(_02874_ ), .B(fanout_net_27 ), .C1(_02353_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02875_ ) );
OR2_X1 _10476_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02876_ ) );
OAI211_X1 _10477_ ( .A(_02876_ ), .B(_02271_ ), .C1(_02284_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02877_ ) );
NAND3_X1 _10478_ ( .A1(_02875_ ), .A2(_02877_ ), .A3(fanout_net_29 ), .ZN(_02878_ ) );
MUX2_X1 _10479_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02879_ ) );
MUX2_X1 _10480_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02880_ ) );
MUX2_X1 _10481_ ( .A(_02879_ ), .B(_02880_ ), .S(fanout_net_27 ), .Z(_02881_ ) );
OAI211_X1 _10482_ ( .A(fanout_net_30 ), .B(_02878_ ), .C1(_02881_ ), .C2(fanout_net_29 ), .ZN(_02882_ ) );
NAND2_X1 _10483_ ( .A1(_02873_ ), .A2(_02882_ ), .ZN(_02883_ ) );
OAI21_X1 _10484_ ( .A(_02883_ ), .B1(_02338_ ), .B2(_02340_ ), .ZN(_02884_ ) );
NAND4_X1 _10485_ ( .A1(_02343_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02345_ ), .ZN(_02885_ ) );
AND2_X2 _10486_ ( .A1(_02884_ ), .A2(_02885_ ), .ZN(_02886_ ) );
XOR2_X1 _10487_ ( .A(_02886_ ), .B(\ID_EX_imm [12] ), .Z(_02887_ ) );
NAND3_X1 _10488_ ( .A1(_02840_ ), .A2(_02864_ ), .A3(_02887_ ), .ZN(_02888_ ) );
OR2_X4 _10489_ ( .A1(_02793_ ), .A2(_02888_ ), .ZN(_02889_ ) );
NAND2_X1 _10490_ ( .A1(_02886_ ), .A2(\ID_EX_imm [12] ), .ZN(_02890_ ) );
NOR3_X1 _10491_ ( .A1(_02890_ ), .A2(_02863_ ), .A3(_02862_ ), .ZN(_02891_ ) );
OAI211_X1 _10492_ ( .A(_02816_ ), .B(_02839_ ), .C1(_02891_ ), .C2(_02862_ ), .ZN(_02892_ ) );
NAND2_X1 _10493_ ( .A1(_02815_ ), .A2(\ID_EX_imm [15] ), .ZN(_02893_ ) );
NAND4_X1 _10494_ ( .A1(_02816_ ), .A2(\ID_EX_imm [14] ), .A3(_02836_ ), .A4(_02837_ ), .ZN(_02894_ ) );
AND3_X1 _10495_ ( .A1(_02892_ ), .A2(_02893_ ), .A3(_02894_ ), .ZN(_02895_ ) );
AOI21_X4 _10496_ ( .A(_02475_ ), .B1(_02889_ ), .B2(_02895_ ), .ZN(_02896_ ) );
OR3_X1 _10497_ ( .A1(_02247_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02252_ ), .ZN(_02897_ ) );
OR2_X1 _10498_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02898_ ) );
OAI211_X1 _10499_ ( .A(_02898_ ), .B(_02302_ ), .C1(_02306_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02899_ ) );
OR2_X1 _10500_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02900_ ) );
OAI211_X1 _10501_ ( .A(_02900_ ), .B(fanout_net_27 ), .C1(_02306_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02901_ ) );
NAND3_X1 _10502_ ( .A1(_02899_ ), .A2(_02901_ ), .A3(fanout_net_29 ), .ZN(_02902_ ) );
MUX2_X1 _10503_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02903_ ) );
MUX2_X1 _10504_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02904_ ) );
MUX2_X1 _10505_ ( .A(_02903_ ), .B(_02904_ ), .S(_02302_ ), .Z(_02905_ ) );
OAI211_X1 _10506_ ( .A(_02320_ ), .B(_02902_ ), .C1(_02905_ ), .C2(fanout_net_29 ), .ZN(_02906_ ) );
NOR2_X1 _10507_ ( .A1(_02451_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02907_ ) );
OAI21_X1 _10508_ ( .A(fanout_net_27 ), .B1(fanout_net_23 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02908_ ) );
NOR2_X1 _10509_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02909_ ) );
OAI21_X1 _10510_ ( .A(_02302_ ), .B1(_02306_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02910_ ) );
OAI221_X1 _10511_ ( .A(_02262_ ), .B1(_02907_ ), .B2(_02908_ ), .C1(_02909_ ), .C2(_02910_ ), .ZN(_02911_ ) );
MUX2_X1 _10512_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02912_ ) );
MUX2_X1 _10513_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02913_ ) );
MUX2_X1 _10514_ ( .A(_02912_ ), .B(_02913_ ), .S(fanout_net_27 ), .Z(_02914_ ) );
OAI211_X1 _10515_ ( .A(fanout_net_30 ), .B(_02911_ ), .C1(_02914_ ), .C2(_02315_ ), .ZN(_02915_ ) );
OAI211_X1 _10516_ ( .A(_02906_ ), .B(_02915_ ), .C1(_02247_ ), .C2(_02253_ ), .ZN(_02916_ ) );
NAND2_X2 _10517_ ( .A1(_02897_ ), .A2(_02916_ ), .ZN(_02917_ ) );
XOR2_X1 _10518_ ( .A(_02917_ ), .B(\ID_EX_imm [18] ), .Z(_02918_ ) );
OR2_X1 _10519_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02919_ ) );
OAI211_X1 _10520_ ( .A(_02919_ ), .B(_02301_ ), .C1(_02305_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02920_ ) );
OR2_X1 _10521_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02921_ ) );
OAI211_X1 _10522_ ( .A(_02921_ ), .B(fanout_net_27 ), .C1(_02305_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02922_ ) );
NAND3_X1 _10523_ ( .A1(_02920_ ), .A2(_02922_ ), .A3(_02261_ ), .ZN(_02923_ ) );
MUX2_X1 _10524_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02924_ ) );
MUX2_X1 _10525_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02925_ ) );
MUX2_X1 _10526_ ( .A(_02924_ ), .B(_02925_ ), .S(_02301_ ), .Z(_02926_ ) );
OAI211_X1 _10527_ ( .A(_02319_ ), .B(_02923_ ), .C1(_02926_ ), .C2(_02279_ ), .ZN(_02927_ ) );
OR2_X1 _10528_ ( .A1(_02304_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02928_ ) );
OAI211_X1 _10529_ ( .A(_02928_ ), .B(_02301_ ), .C1(fanout_net_23 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02929_ ) );
OR2_X1 _10530_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02930_ ) );
OAI211_X1 _10531_ ( .A(_02930_ ), .B(fanout_net_27 ), .C1(_02353_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02931_ ) );
NAND3_X1 _10532_ ( .A1(_02929_ ), .A2(fanout_net_29 ), .A3(_02931_ ), .ZN(_02932_ ) );
MUX2_X1 _10533_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02933_ ) );
MUX2_X1 _10534_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02934_ ) );
MUX2_X1 _10535_ ( .A(_02933_ ), .B(_02934_ ), .S(fanout_net_27 ), .Z(_02935_ ) );
OAI211_X1 _10536_ ( .A(fanout_net_30 ), .B(_02932_ ), .C1(_02935_ ), .C2(fanout_net_29 ), .ZN(_02936_ ) );
NAND2_X1 _10537_ ( .A1(_02927_ ), .A2(_02936_ ), .ZN(_02937_ ) );
OAI21_X1 _10538_ ( .A(_02937_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_02938_ ) );
NAND4_X1 _10539_ ( .A1(_02344_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_02939_ ) );
AND2_X2 _10540_ ( .A1(_02938_ ), .A2(_02939_ ), .ZN(_02940_ ) );
INV_X1 _10541_ ( .A(\ID_EX_imm [19] ), .ZN(_02941_ ) );
XNOR2_X1 _10542_ ( .A(_02940_ ), .B(_02941_ ), .ZN(_02942_ ) );
AND2_X1 _10543_ ( .A1(_02918_ ), .A2(_02942_ ), .ZN(_02943_ ) );
NOR2_X1 _10544_ ( .A1(_02353_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02944_ ) );
OAI21_X1 _10545_ ( .A(fanout_net_27 ), .B1(fanout_net_23 ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02945_ ) );
NOR2_X1 _10546_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02946_ ) );
OAI21_X1 _10547_ ( .A(_02301_ ), .B1(_02353_ ), .B2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02947_ ) );
OAI221_X1 _10548_ ( .A(_02261_ ), .B1(_02944_ ), .B2(_02945_ ), .C1(_02946_ ), .C2(_02947_ ), .ZN(_02948_ ) );
MUX2_X1 _10549_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02949_ ) );
MUX2_X1 _10550_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02950_ ) );
MUX2_X1 _10551_ ( .A(_02949_ ), .B(_02950_ ), .S(fanout_net_27 ), .Z(_02951_ ) );
OAI211_X1 _10552_ ( .A(fanout_net_30 ), .B(_02948_ ), .C1(_02951_ ), .C2(_02279_ ), .ZN(_02952_ ) );
OR2_X1 _10553_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02953_ ) );
OAI211_X1 _10554_ ( .A(_02953_ ), .B(_02301_ ), .C1(_02305_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02954_ ) );
OR2_X1 _10555_ ( .A1(fanout_net_23 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02955_ ) );
OAI211_X1 _10556_ ( .A(_02955_ ), .B(fanout_net_27 ), .C1(_02305_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02956_ ) );
NAND3_X1 _10557_ ( .A1(_02954_ ), .A2(_02956_ ), .A3(fanout_net_29 ), .ZN(_02957_ ) );
MUX2_X1 _10558_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02958_ ) );
MUX2_X1 _10559_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02959_ ) );
MUX2_X1 _10560_ ( .A(_02958_ ), .B(_02959_ ), .S(_02271_ ), .Z(_02960_ ) );
OAI211_X1 _10561_ ( .A(_02319_ ), .B(_02957_ ), .C1(_02960_ ), .C2(fanout_net_29 ), .ZN(_02961_ ) );
NAND2_X1 _10562_ ( .A1(_02952_ ), .A2(_02961_ ), .ZN(_02962_ ) );
OAI21_X1 _10563_ ( .A(_02962_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_02963_ ) );
NAND4_X1 _10564_ ( .A1(_02344_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_02964_ ) );
AND2_X2 _10565_ ( .A1(_02963_ ), .A2(_02964_ ), .ZN(_02965_ ) );
INV_X1 _10566_ ( .A(\ID_EX_imm [17] ), .ZN(_02966_ ) );
XNOR2_X1 _10567_ ( .A(_02965_ ), .B(_02966_ ), .ZN(_02967_ ) );
AND4_X2 _10568_ ( .A1(_02449_ ), .A2(_02896_ ), .A3(_02943_ ), .A4(_02967_ ), .ZN(_02968_ ) );
INV_X1 _10569_ ( .A(_02968_ ), .ZN(_02969_ ) );
AND2_X1 _10570_ ( .A1(_02472_ ), .A2(\ID_EX_imm [16] ), .ZN(_02970_ ) );
AND2_X1 _10571_ ( .A1(_02967_ ), .A2(_02970_ ), .ZN(_02971_ ) );
AOI21_X1 _10572_ ( .A(_02971_ ), .B1(\ID_EX_imm [17] ), .B2(_02965_ ), .ZN(_02972_ ) );
INV_X1 _10573_ ( .A(_02972_ ), .ZN(_02973_ ) );
NAND2_X1 _10574_ ( .A1(_02973_ ), .A2(_02943_ ), .ZN(_02974_ ) );
AND2_X1 _10575_ ( .A1(_02917_ ), .A2(\ID_EX_imm [18] ), .ZN(_02975_ ) );
AND2_X1 _10576_ ( .A1(_02942_ ), .A2(_02975_ ), .ZN(_02976_ ) );
AOI21_X1 _10577_ ( .A(_02976_ ), .B1(\ID_EX_imm [19] ), .B2(_02940_ ), .ZN(_02977_ ) );
AND2_X1 _10578_ ( .A1(_02974_ ), .A2(_02977_ ), .ZN(_02978_ ) );
INV_X1 _10579_ ( .A(_02978_ ), .ZN(_02979_ ) );
AND3_X1 _10580_ ( .A1(_02979_ ), .A2(_02399_ ), .A3(_02448_ ), .ZN(_02980_ ) );
AND2_X1 _10581_ ( .A1(_02396_ ), .A2(\ID_EX_imm [23] ), .ZN(_02981_ ) );
NAND2_X1 _10582_ ( .A1(_02422_ ), .A2(\ID_EX_imm [20] ), .ZN(_02982_ ) );
NOR3_X1 _10583_ ( .A1(_02982_ ), .A2(_02445_ ), .A3(_02446_ ), .ZN(_02983_ ) );
OR2_X1 _10584_ ( .A1(_02983_ ), .A2(_02445_ ), .ZN(_02984_ ) );
AND3_X1 _10585_ ( .A1(_02984_ ), .A2(_02398_ ), .A3(_02374_ ), .ZN(_02985_ ) );
AND2_X1 _10586_ ( .A1(_02373_ ), .A2(\ID_EX_imm [22] ), .ZN(_02986_ ) );
AND2_X1 _10587_ ( .A1(_02398_ ), .A2(_02986_ ), .ZN(_02987_ ) );
NOR4_X1 _10588_ ( .A1(_02980_ ), .A2(_02981_ ), .A3(_02985_ ), .A4(_02987_ ), .ZN(_02988_ ) );
AND2_X2 _10589_ ( .A1(_02969_ ), .A2(_02988_ ), .ZN(_02989_ ) );
OR2_X1 _10590_ ( .A1(_02451_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02990_ ) );
OAI211_X1 _10591_ ( .A(_02990_ ), .B(_02273_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02991_ ) );
BUF_X4 _10592_ ( .A(_02451_ ), .Z(_02992_ ) );
NOR2_X1 _10593_ ( .A1(_02992_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02993_ ) );
OAI21_X1 _10594_ ( .A(fanout_net_27 ), .B1(fanout_net_24 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02994_ ) );
OAI211_X1 _10595_ ( .A(_02991_ ), .B(fanout_net_29 ), .C1(_02993_ ), .C2(_02994_ ), .ZN(_02995_ ) );
MUX2_X1 _10596_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02996_ ) );
MUX2_X1 _10597_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02997_ ) );
MUX2_X1 _10598_ ( .A(_02996_ ), .B(_02997_ ), .S(fanout_net_27 ), .Z(_02998_ ) );
OAI211_X1 _10599_ ( .A(_02995_ ), .B(fanout_net_30 ), .C1(_02998_ ), .C2(fanout_net_29 ), .ZN(_02999_ ) );
OR2_X1 _10600_ ( .A1(_02451_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03000_ ) );
OAI211_X1 _10601_ ( .A(_03000_ ), .B(fanout_net_27 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03001_ ) );
OR2_X1 _10602_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03002_ ) );
OAI211_X1 _10603_ ( .A(_03002_ ), .B(_02273_ ), .C1(_02992_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03003_ ) );
NAND3_X1 _10604_ ( .A1(_03001_ ), .A2(_02264_ ), .A3(_03003_ ), .ZN(_03004_ ) );
MUX2_X1 _10605_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03005_ ) );
MUX2_X1 _10606_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03006_ ) );
MUX2_X1 _10607_ ( .A(_03005_ ), .B(_03006_ ), .S(_02401_ ), .Z(_03007_ ) );
OAI211_X1 _10608_ ( .A(_02320_ ), .B(_03004_ ), .C1(_03007_ ), .C2(_02264_ ), .ZN(_03008_ ) );
NAND2_X1 _10609_ ( .A1(_02999_ ), .A2(_03008_ ), .ZN(_03009_ ) );
OAI21_X1 _10610_ ( .A(_03009_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_03010_ ) );
NAND4_X1 _10611_ ( .A1(_02344_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_03011_ ) );
AND3_X1 _10612_ ( .A1(_03010_ ), .A2(\ID_EX_imm [24] ), .A3(_03011_ ), .ZN(_03012_ ) );
AOI21_X1 _10613_ ( .A(\ID_EX_imm [24] ), .B1(_03010_ ), .B2(_03011_ ), .ZN(_03013_ ) );
NOR3_X2 _10614_ ( .A1(_02989_ ), .A2(_03012_ ), .A3(_03013_ ), .ZN(_03014_ ) );
NOR2_X1 _10615_ ( .A1(_03014_ ), .A2(_03012_ ), .ZN(_03015_ ) );
INV_X1 _10616_ ( .A(\ID_EX_imm [25] ), .ZN(_03016_ ) );
OR2_X1 _10617_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03017_ ) );
OAI211_X1 _10618_ ( .A(_03017_ ), .B(_02273_ ), .C1(_02992_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03018_ ) );
INV_X1 _10619_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03019_ ) );
NAND2_X1 _10620_ ( .A1(_03019_ ), .A2(fanout_net_24 ), .ZN(_03020_ ) );
OAI211_X1 _10621_ ( .A(_03020_ ), .B(fanout_net_27 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03021_ ) );
NAND3_X1 _10622_ ( .A1(_03018_ ), .A2(_03021_ ), .A3(_02315_ ), .ZN(_03022_ ) );
MUX2_X1 _10623_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03023_ ) );
MUX2_X1 _10624_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03024_ ) );
MUX2_X1 _10625_ ( .A(_03023_ ), .B(_03024_ ), .S(_02401_ ), .Z(_03025_ ) );
OAI211_X1 _10626_ ( .A(_02320_ ), .B(_03022_ ), .C1(_03025_ ), .C2(_02264_ ), .ZN(_03026_ ) );
OR2_X1 _10627_ ( .A1(_02451_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03027_ ) );
OAI211_X1 _10628_ ( .A(_03027_ ), .B(fanout_net_27 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03028_ ) );
OR2_X1 _10629_ ( .A1(fanout_net_24 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03029_ ) );
OAI211_X1 _10630_ ( .A(_03029_ ), .B(_02401_ ), .C1(_02992_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03030_ ) );
NAND3_X1 _10631_ ( .A1(_03028_ ), .A2(_03030_ ), .A3(fanout_net_29 ), .ZN(_03031_ ) );
MUX2_X1 _10632_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03032_ ) );
MUX2_X1 _10633_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03033_ ) );
MUX2_X1 _10634_ ( .A(_03032_ ), .B(_03033_ ), .S(fanout_net_27 ), .Z(_03034_ ) );
OAI211_X1 _10635_ ( .A(fanout_net_30 ), .B(_03031_ ), .C1(_03034_ ), .C2(fanout_net_29 ), .ZN(_03035_ ) );
NAND2_X1 _10636_ ( .A1(_03026_ ), .A2(_03035_ ), .ZN(_03036_ ) );
OAI21_X1 _10637_ ( .A(_03036_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_03037_ ) );
NAND4_X1 _10638_ ( .A1(_02344_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_03038_ ) );
AND2_X2 _10639_ ( .A1(_03037_ ), .A2(_03038_ ), .ZN(_03039_ ) );
INV_X1 _10640_ ( .A(_03039_ ), .ZN(_03040_ ) );
OAI21_X1 _10641_ ( .A(_03015_ ), .B1(_03016_ ), .B2(_03040_ ), .ZN(_03041_ ) );
OR3_X1 _10642_ ( .A1(_02247_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02253_ ), .ZN(_03042_ ) );
OR2_X1 _10643_ ( .A1(_02451_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03043_ ) );
OAI211_X1 _10644_ ( .A(_03043_ ), .B(_02401_ ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03044_ ) );
OR2_X1 _10645_ ( .A1(_02285_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03045_ ) );
OAI211_X1 _10646_ ( .A(_03045_ ), .B(fanout_net_27 ), .C1(fanout_net_24 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03046_ ) );
NAND3_X1 _10647_ ( .A1(_03044_ ), .A2(_03046_ ), .A3(fanout_net_29 ), .ZN(_03047_ ) );
MUX2_X1 _10648_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03048_ ) );
MUX2_X1 _10649_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03049_ ) );
MUX2_X1 _10650_ ( .A(_03048_ ), .B(_03049_ ), .S(_02401_ ), .Z(_03050_ ) );
OAI211_X1 _10651_ ( .A(_02320_ ), .B(_03047_ ), .C1(_03050_ ), .C2(fanout_net_29 ), .ZN(_03051_ ) );
NOR2_X1 _10652_ ( .A1(_02306_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03052_ ) );
OAI21_X1 _10653_ ( .A(fanout_net_27 ), .B1(fanout_net_24 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03053_ ) );
INV_X1 _10654_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03054_ ) );
INV_X1 _10655_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03055_ ) );
MUX2_X1 _10656_ ( .A(_03054_ ), .B(_03055_ ), .S(fanout_net_24 ), .Z(_03056_ ) );
OAI221_X1 _10657_ ( .A(_02315_ ), .B1(_03052_ ), .B2(_03053_ ), .C1(_03056_ ), .C2(fanout_net_27 ), .ZN(_03057_ ) );
MUX2_X1 _10658_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03058_ ) );
MUX2_X1 _10659_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_03059_ ) );
MUX2_X1 _10660_ ( .A(_03058_ ), .B(_03059_ ), .S(fanout_net_27 ), .Z(_03060_ ) );
OAI211_X1 _10661_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03057_ ), .C1(_03060_ ), .C2(_02264_ ), .ZN(_03061_ ) );
OAI211_X1 _10662_ ( .A(_03051_ ), .B(_03061_ ), .C1(_02247_ ), .C2(_02253_ ), .ZN(_03062_ ) );
NAND2_X2 _10663_ ( .A1(_03042_ ), .A2(_03062_ ), .ZN(_03063_ ) );
INV_X1 _10664_ ( .A(\ID_EX_imm [26] ), .ZN(_03064_ ) );
XNOR2_X1 _10665_ ( .A(_03063_ ), .B(_03064_ ), .ZN(_03065_ ) );
OR2_X1 _10666_ ( .A1(_03039_ ), .A2(\ID_EX_imm [25] ), .ZN(_03066_ ) );
AND4_X2 _10667_ ( .A1(_02350_ ), .A2(_03041_ ), .A3(_03065_ ), .A4(_03066_ ), .ZN(_03067_ ) );
AND2_X1 _10668_ ( .A1(_03063_ ), .A2(\ID_EX_imm [26] ), .ZN(_03068_ ) );
AND2_X1 _10669_ ( .A1(_02350_ ), .A2(_03068_ ), .ZN(_03069_ ) );
AOI21_X1 _10670_ ( .A(_03069_ ), .B1(\ID_EX_imm [27] ), .B2(_02348_ ), .ZN(_03070_ ) );
INV_X1 _10671_ ( .A(_03070_ ), .ZN(_03071_ ) );
NOR2_X2 _10672_ ( .A1(_03067_ ), .A2(_03071_ ), .ZN(_03072_ ) );
OR3_X1 _10673_ ( .A1(_02247_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02253_ ), .ZN(_03073_ ) );
INV_X1 _10674_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03074_ ) );
NAND2_X1 _10675_ ( .A1(_03074_ ), .A2(fanout_net_24 ), .ZN(_03075_ ) );
OAI211_X1 _10676_ ( .A(_03075_ ), .B(_02273_ ), .C1(fanout_net_24 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03076_ ) );
INV_X1 _10677_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03077_ ) );
NAND2_X1 _10678_ ( .A1(_03077_ ), .A2(fanout_net_24 ), .ZN(_03078_ ) );
OAI211_X1 _10679_ ( .A(_03078_ ), .B(fanout_net_27 ), .C1(fanout_net_24 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03079_ ) );
NAND3_X1 _10680_ ( .A1(_03076_ ), .A2(_03079_ ), .A3(_02315_ ), .ZN(_03080_ ) );
MUX2_X1 _10681_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03081_ ) );
MUX2_X1 _10682_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03082_ ) );
MUX2_X1 _10683_ ( .A(_03081_ ), .B(_03082_ ), .S(_02401_ ), .Z(_03083_ ) );
OAI211_X1 _10684_ ( .A(_02320_ ), .B(_03080_ ), .C1(_03083_ ), .C2(_02264_ ), .ZN(_03084_ ) );
OR2_X1 _10685_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03085_ ) );
OAI211_X1 _10686_ ( .A(_03085_ ), .B(fanout_net_27 ), .C1(_02992_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03086_ ) );
OR2_X1 _10687_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03087_ ) );
OAI211_X1 _10688_ ( .A(_03087_ ), .B(_02401_ ), .C1(_02306_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03088_ ) );
NAND3_X1 _10689_ ( .A1(_03086_ ), .A2(_03088_ ), .A3(fanout_net_29 ), .ZN(_03089_ ) );
MUX2_X1 _10690_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03090_ ) );
MUX2_X1 _10691_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03091_ ) );
MUX2_X1 _10692_ ( .A(_03090_ ), .B(_03091_ ), .S(fanout_net_27 ), .Z(_03092_ ) );
OAI211_X1 _10693_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_03089_ ), .C1(_03092_ ), .C2(fanout_net_29 ), .ZN(_03093_ ) );
OAI211_X1 _10694_ ( .A(_03084_ ), .B(_03093_ ), .C1(_02247_ ), .C2(_02253_ ), .ZN(_03094_ ) );
NAND2_X1 _10695_ ( .A1(_03073_ ), .A2(_03094_ ), .ZN(_03095_ ) );
XNOR2_X1 _10696_ ( .A(_03095_ ), .B(\ID_EX_imm [28] ), .ZN(_03096_ ) );
NOR2_X2 _10697_ ( .A1(_03072_ ), .A2(_03096_ ), .ZN(_03097_ ) );
OR3_X1 _10698_ ( .A1(_02247_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02253_ ), .ZN(_03098_ ) );
OR2_X1 _10699_ ( .A1(_02451_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03099_ ) );
OAI211_X1 _10700_ ( .A(_03099_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03100_ ) );
OR2_X1 _10701_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03101_ ) );
OAI211_X1 _10702_ ( .A(_03101_ ), .B(_02273_ ), .C1(_02992_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03102_ ) );
NAND3_X1 _10703_ ( .A1(_03100_ ), .A2(_02315_ ), .A3(_03102_ ), .ZN(_03103_ ) );
MUX2_X1 _10704_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03104_ ) );
MUX2_X1 _10705_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03105_ ) );
MUX2_X1 _10706_ ( .A(_03104_ ), .B(_03105_ ), .S(_02401_ ), .Z(_03106_ ) );
OAI211_X1 _10707_ ( .A(_02320_ ), .B(_03103_ ), .C1(_03106_ ), .C2(_02264_ ), .ZN(_03107_ ) );
OR2_X1 _10708_ ( .A1(_02451_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03108_ ) );
OAI211_X1 _10709_ ( .A(_03108_ ), .B(_02401_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03109_ ) );
NOR2_X1 _10710_ ( .A1(_02992_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03110_ ) );
OAI21_X1 _10711_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03111_ ) );
OAI211_X1 _10712_ ( .A(_03109_ ), .B(fanout_net_29 ), .C1(_03110_ ), .C2(_03111_ ), .ZN(_03112_ ) );
MUX2_X1 _10713_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03113_ ) );
MUX2_X1 _10714_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03114_ ) );
MUX2_X1 _10715_ ( .A(_03113_ ), .B(_03114_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03115_ ) );
OAI211_X1 _10716_ ( .A(_03112_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .C1(_03115_ ), .C2(fanout_net_29 ), .ZN(_03116_ ) );
OAI211_X1 _10717_ ( .A(_03107_ ), .B(_03116_ ), .C1(_02247_ ), .C2(_02253_ ), .ZN(_03117_ ) );
NAND2_X2 _10718_ ( .A1(_03098_ ), .A2(_03117_ ), .ZN(_03118_ ) );
INV_X1 _10719_ ( .A(\ID_EX_imm [29] ), .ZN(_03119_ ) );
XNOR2_X1 _10720_ ( .A(_03118_ ), .B(_03119_ ), .ZN(_03120_ ) );
NAND2_X1 _10721_ ( .A1(_03097_ ), .A2(_03120_ ), .ZN(_03121_ ) );
AOI21_X1 _10722_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_03073_ ), .B2(_03094_ ), .ZN(_03122_ ) );
INV_X1 _10723_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03123_ ) );
AOI22_X1 _10724_ ( .A1(_03120_ ), .A2(_03122_ ), .B1(_03123_ ), .B2(_03118_ ), .ZN(_03124_ ) );
AOI21_X1 _10725_ ( .A(_02298_ ), .B1(_03121_ ), .B2(_03124_ ), .ZN(_03125_ ) );
AOI21_X1 _10726_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_02295_ ), .B2(_02296_ ), .ZN(_03126_ ) );
NOR2_X1 _10727_ ( .A1(_03125_ ), .A2(_03126_ ), .ZN(_03127_ ) );
OR2_X1 _10728_ ( .A1(_02451_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03128_ ) );
OAI211_X1 _10729_ ( .A(_03128_ ), .B(_02273_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03129_ ) );
NOR2_X1 _10730_ ( .A1(_02992_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03130_ ) );
OAI21_X1 _10731_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03131_ ) );
OAI211_X1 _10732_ ( .A(_03129_ ), .B(fanout_net_29 ), .C1(_03130_ ), .C2(_03131_ ), .ZN(_03132_ ) );
MUX2_X1 _10733_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03133_ ) );
MUX2_X1 _10734_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03134_ ) );
MUX2_X1 _10735_ ( .A(_03133_ ), .B(_03134_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_03135_ ) );
OAI211_X1 _10736_ ( .A(_03132_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .C1(_03135_ ), .C2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_03136_ ) );
OR2_X1 _10737_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_03137_ ) );
OAI211_X1 _10738_ ( .A(_03137_ ), .B(_02273_ ), .C1(_02992_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_03138_ ) );
OR2_X1 _10739_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03139_ ) );
OAI211_X1 _10740_ ( .A(_03139_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_02992_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_03140_ ) );
NAND3_X1 _10741_ ( .A1(_03138_ ), .A2(_03140_ ), .A3(_02264_ ), .ZN(_03141_ ) );
MUX2_X1 _10742_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03142_ ) );
MUX2_X1 _10743_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_03143_ ) );
MUX2_X1 _10744_ ( .A(_03142_ ), .B(_03143_ ), .S(_02273_ ), .Z(_03144_ ) );
OAI211_X1 _10745_ ( .A(_02320_ ), .B(_03141_ ), .C1(_03144_ ), .C2(_02264_ ), .ZN(_03145_ ) );
NAND2_X1 _10746_ ( .A1(_03136_ ), .A2(_03145_ ), .ZN(_03146_ ) );
OAI21_X1 _10747_ ( .A(_03146_ ), .B1(_02339_ ), .B2(_02341_ ), .ZN(_03147_ ) );
NAND4_X1 _10748_ ( .A1(_02344_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(\myidu.fc_disenable_$_NOT__A_Y ), .A4(_02346_ ), .ZN(_03148_ ) );
AND2_X1 _10749_ ( .A1(_03147_ ), .A2(_03148_ ), .ZN(_03149_ ) );
BUF_X2 _10750_ ( .A(_03149_ ), .Z(_03150_ ) );
XNOR2_X1 _10751_ ( .A(_03150_ ), .B(\ID_EX_imm [31] ), .ZN(_03151_ ) );
XNOR2_X1 _10752_ ( .A(_03127_ ), .B(_03151_ ), .ZN(_03152_ ) );
AND2_X2 _10753_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_03153_ ) );
BUF_X4 _10754_ ( .A(_03153_ ), .Z(_03154_ ) );
NOR2_X1 _10755_ ( .A1(_03152_ ), .A2(_03154_ ), .ZN(_00133_ ) );
NAND2_X1 _10756_ ( .A1(_03121_ ), .A2(_03124_ ), .ZN(_03155_ ) );
XNOR2_X1 _10757_ ( .A(_03155_ ), .B(_02298_ ), .ZN(_03156_ ) );
INV_X1 _10758_ ( .A(_03153_ ), .ZN(_03157_ ) );
CLKBUF_X2 _10759_ ( .A(_03157_ ), .Z(_03158_ ) );
AND2_X1 _10760_ ( .A1(_03156_ ), .A2(_03158_ ), .ZN(_00134_ ) );
AND3_X1 _10761_ ( .A1(_02896_ ), .A2(_02943_ ), .A3(_02967_ ), .ZN(_03159_ ) );
OAI21_X1 _10762_ ( .A(_02423_ ), .B1(_03159_ ), .B2(_02979_ ), .ZN(_03160_ ) );
NAND2_X1 _10763_ ( .A1(_03160_ ), .A2(_02982_ ), .ZN(_03161_ ) );
XNOR2_X1 _10764_ ( .A(_03161_ ), .B(_02447_ ), .ZN(_03162_ ) );
NOR2_X1 _10765_ ( .A1(_03162_ ), .A2(_03154_ ), .ZN(_00135_ ) );
OR3_X1 _10766_ ( .A1(_03159_ ), .A2(_02423_ ), .A3(_02979_ ), .ZN(_03163_ ) );
AND3_X1 _10767_ ( .A1(_03163_ ), .A2(_03158_ ), .A3(_03160_ ), .ZN(_00136_ ) );
AND2_X1 _10768_ ( .A1(_02896_ ), .A2(_02967_ ), .ZN(_03164_ ) );
NOR2_X1 _10769_ ( .A1(_03164_ ), .A2(_02973_ ), .ZN(_03165_ ) );
NOR2_X1 _10770_ ( .A1(_02917_ ), .A2(\ID_EX_imm [18] ), .ZN(_03166_ ) );
NOR3_X1 _10771_ ( .A1(_03165_ ), .A2(_02975_ ), .A3(_03166_ ), .ZN(_03167_ ) );
OR2_X1 _10772_ ( .A1(_03167_ ), .A2(_02975_ ), .ZN(_03168_ ) );
XNOR2_X1 _10773_ ( .A(_03168_ ), .B(_02942_ ), .ZN(_03169_ ) );
NOR2_X1 _10774_ ( .A1(_03169_ ), .A2(_03154_ ), .ZN(_00137_ ) );
XNOR2_X1 _10775_ ( .A(_03165_ ), .B(_02918_ ), .ZN(_03170_ ) );
AND2_X1 _10776_ ( .A1(_03170_ ), .A2(_03158_ ), .ZN(_00138_ ) );
OR2_X1 _10777_ ( .A1(_02896_ ), .A2(_02970_ ), .ZN(_03171_ ) );
XNOR2_X1 _10778_ ( .A(_03171_ ), .B(_02967_ ), .ZN(_03172_ ) );
NOR2_X1 _10779_ ( .A1(_03172_ ), .A2(_03154_ ), .ZN(_00139_ ) );
AND3_X1 _10780_ ( .A1(_02889_ ), .A2(_02895_ ), .A3(_02475_ ), .ZN(_03173_ ) );
NOR3_X1 _10781_ ( .A1(_03173_ ), .A2(_02896_ ), .A3(_03153_ ), .ZN(_00140_ ) );
INV_X1 _10782_ ( .A(_02864_ ), .ZN(_03174_ ) );
INV_X1 _10783_ ( .A(_02887_ ), .ZN(_03175_ ) );
NOR3_X1 _10784_ ( .A1(_02793_ ), .A2(_03174_ ), .A3(_03175_ ), .ZN(_03176_ ) );
OR2_X1 _10785_ ( .A1(_02891_ ), .A2(_02862_ ), .ZN(_03177_ ) );
OAI21_X1 _10786_ ( .A(_02839_ ), .B1(_03176_ ), .B2(_03177_ ), .ZN(_03178_ ) );
NAND2_X1 _10787_ ( .A1(_02838_ ), .A2(\ID_EX_imm [14] ), .ZN(_03179_ ) );
NAND2_X1 _10788_ ( .A1(_03178_ ), .A2(_03179_ ), .ZN(_03180_ ) );
XNOR2_X1 _10789_ ( .A(_03180_ ), .B(_02816_ ), .ZN(_03181_ ) );
NOR2_X1 _10790_ ( .A1(_03181_ ), .A2(_03154_ ), .ZN(_00141_ ) );
OR3_X1 _10791_ ( .A1(_03176_ ), .A2(_02839_ ), .A3(_03177_ ), .ZN(_03182_ ) );
AND3_X1 _10792_ ( .A1(_03182_ ), .A2(_03158_ ), .A3(_03178_ ), .ZN(_00142_ ) );
OAI21_X1 _10793_ ( .A(_02887_ ), .B1(_02784_ ), .B2(_02792_ ), .ZN(_03183_ ) );
NAND2_X1 _10794_ ( .A1(_03183_ ), .A2(_02890_ ), .ZN(_03184_ ) );
XNOR2_X1 _10795_ ( .A(_03184_ ), .B(_03174_ ), .ZN(_03185_ ) );
AND2_X1 _10796_ ( .A1(_03185_ ), .A2(_03158_ ), .ZN(_00143_ ) );
XNOR2_X1 _10797_ ( .A(_02793_ ), .B(_02887_ ), .ZN(_03186_ ) );
AND2_X1 _10798_ ( .A1(_03186_ ), .A2(_03158_ ), .ZN(_00144_ ) );
OR2_X1 _10799_ ( .A1(_03097_ ), .A2(_03122_ ), .ZN(_03187_ ) );
XNOR2_X1 _10800_ ( .A(_03187_ ), .B(_03120_ ), .ZN(_03188_ ) );
NOR2_X1 _10801_ ( .A1(_03188_ ), .A2(_03154_ ), .ZN(_00145_ ) );
XNOR2_X1 _10802_ ( .A(_03072_ ), .B(_03096_ ), .ZN(_03189_ ) );
NOR2_X1 _10803_ ( .A1(_03189_ ), .A2(_03154_ ), .ZN(_00146_ ) );
AND3_X1 _10804_ ( .A1(_03041_ ), .A2(_03065_ ), .A3(_03066_ ), .ZN(_03190_ ) );
OR2_X1 _10805_ ( .A1(_03190_ ), .A2(_03068_ ), .ZN(_03191_ ) );
XNOR2_X1 _10806_ ( .A(_03191_ ), .B(_02350_ ), .ZN(_03192_ ) );
NOR2_X1 _10807_ ( .A1(_03192_ ), .A2(_03154_ ), .ZN(_00147_ ) );
AOI21_X1 _10808_ ( .A(_03065_ ), .B1(_03041_ ), .B2(_03066_ ), .ZN(_03193_ ) );
NOR3_X1 _10809_ ( .A1(_03190_ ), .A2(_03193_ ), .A3(_03153_ ), .ZN(_00148_ ) );
XNOR2_X1 _10810_ ( .A(_03039_ ), .B(\ID_EX_imm [25] ), .ZN(_03194_ ) );
XNOR2_X1 _10811_ ( .A(_03015_ ), .B(_03194_ ), .ZN(_03195_ ) );
NOR2_X1 _10812_ ( .A1(_03195_ ), .A2(_03154_ ), .ZN(_00149_ ) );
AND2_X2 _10813_ ( .A1(_03010_ ), .A2(_03011_ ), .ZN(_03196_ ) );
INV_X1 _10814_ ( .A(\ID_EX_imm [24] ), .ZN(_03197_ ) );
XNOR2_X1 _10815_ ( .A(_03196_ ), .B(_03197_ ), .ZN(_03198_ ) );
XNOR2_X1 _10816_ ( .A(_02989_ ), .B(_03198_ ), .ZN(_03199_ ) );
AND2_X1 _10817_ ( .A1(_03199_ ), .A2(_03158_ ), .ZN(_00150_ ) );
OAI21_X1 _10818_ ( .A(_02448_ ), .B1(_03159_ ), .B2(_02979_ ), .ZN(_03200_ ) );
INV_X1 _10819_ ( .A(_03200_ ), .ZN(_03201_ ) );
OR2_X1 _10820_ ( .A1(_03201_ ), .A2(_02984_ ), .ZN(_03202_ ) );
AND2_X1 _10821_ ( .A1(_03202_ ), .A2(_02374_ ), .ZN(_03203_ ) );
OR2_X1 _10822_ ( .A1(_03203_ ), .A2(_02986_ ), .ZN(_03204_ ) );
XNOR2_X1 _10823_ ( .A(_03204_ ), .B(_02398_ ), .ZN(_03205_ ) );
NOR2_X1 _10824_ ( .A1(_03205_ ), .A2(_03154_ ), .ZN(_00151_ ) );
XOR2_X1 _10825_ ( .A(_03202_ ), .B(_02374_ ), .Z(_03206_ ) );
AND2_X1 _10826_ ( .A1(_03206_ ), .A2(_03158_ ), .ZN(_00152_ ) );
AND2_X1 _10827_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_03207_ ) );
NOR2_X1 _10828_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_03208_ ) );
AND2_X1 _10829_ ( .A1(_03207_ ), .A2(_03208_ ), .ZN(_03209_ ) );
CLKBUF_X2 _10830_ ( .A(_03209_ ), .Z(_03210_ ) );
INV_X1 _10831_ ( .A(_03210_ ), .ZN(_03211_ ) );
AND2_X2 _10832_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03212_ ) );
INV_X1 _10833_ ( .A(\IF_ID_inst [12] ), .ZN(_03213_ ) );
NAND4_X1 _10834_ ( .A1(_03212_ ), .A2(\IF_ID_inst [13] ), .A3(_03213_ ), .A4(\IF_ID_inst [6] ), .ZN(_03214_ ) );
NOR2_X1 _10835_ ( .A1(_03211_ ), .A2(_03214_ ), .ZN(_03215_ ) );
AND4_X1 _10836_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03216_ ) );
AND2_X1 _10837_ ( .A1(_03210_ ), .A2(_03216_ ), .ZN(_03217_ ) );
NOR2_X2 _10838_ ( .A1(_03215_ ), .A2(_03217_ ), .ZN(_03218_ ) );
BUF_X4 _10839_ ( .A(_03218_ ), .Z(_03219_ ) );
INV_X1 _10840_ ( .A(\IF_ID_inst [31] ), .ZN(_03220_ ) );
NOR2_X1 _10841_ ( .A1(fanout_net_4 ), .A2(excp_written ), .ZN(_03221_ ) );
AND2_X2 _10842_ ( .A1(_02221_ ), .A2(_03221_ ), .ZN(_03222_ ) );
INV_X2 _10843_ ( .A(_03222_ ), .ZN(_03223_ ) );
BUF_X4 _10844_ ( .A(_03223_ ), .Z(_03224_ ) );
NOR3_X1 _10845_ ( .A1(_03219_ ), .A2(_03220_ ), .A3(_03224_ ), .ZN(_00231_ ) );
INV_X1 _10846_ ( .A(\IF_ID_inst [30] ), .ZN(_03225_ ) );
NOR3_X1 _10847_ ( .A1(_03219_ ), .A2(_03225_ ), .A3(_03224_ ), .ZN(_00232_ ) );
INV_X1 _10848_ ( .A(\IF_ID_inst [21] ), .ZN(_03226_ ) );
NOR3_X1 _10849_ ( .A1(_03219_ ), .A2(_03226_ ), .A3(_03224_ ), .ZN(_00233_ ) );
BUF_X4 _10850_ ( .A(_03223_ ), .Z(_03227_ ) );
INV_X1 _10851_ ( .A(_03218_ ), .ZN(_03228_ ) );
INV_X1 _10852_ ( .A(\IF_ID_inst [20] ), .ZN(_03229_ ) );
AOI21_X1 _10853_ ( .A(_03227_ ), .B1(_03228_ ), .B2(_03229_ ), .ZN(_00234_ ) );
INV_X1 _10854_ ( .A(\IF_ID_inst [29] ), .ZN(_03230_ ) );
AOI21_X1 _10855_ ( .A(_03227_ ), .B1(_03228_ ), .B2(_03230_ ), .ZN(_00235_ ) );
INV_X1 _10856_ ( .A(\IF_ID_inst [28] ), .ZN(_03231_ ) );
AOI21_X1 _10857_ ( .A(_03227_ ), .B1(_03228_ ), .B2(_03231_ ), .ZN(_00236_ ) );
INV_X1 _10858_ ( .A(\IF_ID_inst [27] ), .ZN(_03232_ ) );
BUF_X4 _10859_ ( .A(_03223_ ), .Z(_03233_ ) );
NOR3_X1 _10860_ ( .A1(_03219_ ), .A2(_03232_ ), .A3(_03233_ ), .ZN(_00237_ ) );
INV_X1 _10861_ ( .A(\IF_ID_inst [26] ), .ZN(_03234_ ) );
AOI21_X1 _10862_ ( .A(_03227_ ), .B1(_03228_ ), .B2(_03234_ ), .ZN(_00238_ ) );
INV_X1 _10863_ ( .A(\IF_ID_inst [25] ), .ZN(_03235_ ) );
NOR3_X1 _10864_ ( .A1(_03219_ ), .A2(_03235_ ), .A3(_03233_ ), .ZN(_00239_ ) );
INV_X1 _10865_ ( .A(\IF_ID_inst [24] ), .ZN(_03236_ ) );
NOR3_X1 _10866_ ( .A1(_03219_ ), .A2(_03236_ ), .A3(_03233_ ), .ZN(_00240_ ) );
INV_X1 _10867_ ( .A(\IF_ID_inst [23] ), .ZN(_03237_ ) );
NOR3_X1 _10868_ ( .A1(_03219_ ), .A2(_03237_ ), .A3(_03233_ ), .ZN(_00241_ ) );
INV_X1 _10869_ ( .A(\IF_ID_inst [22] ), .ZN(_03238_ ) );
NOR3_X1 _10870_ ( .A1(_03219_ ), .A2(_03238_ ), .A3(_03233_ ), .ZN(_00242_ ) );
CLKBUF_X2 _10871_ ( .A(_03221_ ), .Z(_03239_ ) );
AND3_X1 _10872_ ( .A1(_02221_ ), .A2(_03239_ ), .A3(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00243_ ) );
AND3_X1 _10873_ ( .A1(_02221_ ), .A2(_03239_ ), .A3(\myidu.state [2] ), .ZN(_00244_ ) );
INV_X1 _10874_ ( .A(\IF_ID_inst [7] ), .ZN(_03240_ ) );
AND4_X1 _10875_ ( .A1(\IF_ID_inst [6] ), .A2(_03210_ ), .A3(_03240_ ), .A4(_03212_ ), .ZN(_03241_ ) );
OR3_X1 _10876_ ( .A1(\IF_ID_inst [11] ), .A2(\IF_ID_inst [10] ), .A3(\IF_ID_inst [9] ), .ZN(_03242_ ) );
NOR2_X1 _10877_ ( .A1(_03242_ ), .A2(\IF_ID_inst [8] ), .ZN(_03243_ ) );
NOR4_X1 _10878_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_03244_ ) );
AND3_X1 _10879_ ( .A1(_03241_ ), .A2(_03243_ ), .A3(_03244_ ), .ZN(_03245_ ) );
NOR2_X1 _10880_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [18] ), .ZN(_03246_ ) );
NOR2_X1 _10881_ ( .A1(\IF_ID_inst [17] ), .A2(\IF_ID_inst [16] ), .ZN(_03247_ ) );
NOR2_X1 _10882_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_03248_ ) );
AND3_X1 _10883_ ( .A1(_03246_ ), .A2(_03247_ ), .A3(_03248_ ), .ZN(_03249_ ) );
NAND3_X1 _10884_ ( .A1(_03249_ ), .A2(_03226_ ), .A3(\IF_ID_inst [20] ), .ZN(_03250_ ) );
NOR2_X1 _10885_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_03251_ ) );
NOR2_X1 _10886_ ( .A1(\IF_ID_inst [27] ), .A2(\IF_ID_inst [24] ), .ZN(_03252_ ) );
AND2_X1 _10887_ ( .A1(_03251_ ), .A2(_03252_ ), .ZN(_03253_ ) );
INV_X1 _10888_ ( .A(_03253_ ), .ZN(_03254_ ) );
NAND4_X1 _10889_ ( .A1(_03225_ ), .A2(_03230_ ), .A3(_03231_ ), .A4(_03220_ ), .ZN(_03255_ ) );
NOR3_X1 _10890_ ( .A1(_03250_ ), .A2(_03254_ ), .A3(_03255_ ), .ZN(_03256_ ) );
NAND2_X1 _10891_ ( .A1(_03245_ ), .A2(_03256_ ), .ZN(_03257_ ) );
NOR2_X1 _10892_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03258_ ) );
BUF_X2 _10893_ ( .A(_03258_ ), .Z(_03259_ ) );
INV_X1 _10894_ ( .A(_03259_ ), .ZN(_03260_ ) );
AND3_X1 _10895_ ( .A1(_03207_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_03261_ ) );
NOR2_X1 _10896_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03262_ ) );
INV_X1 _10897_ ( .A(\IF_ID_inst [6] ), .ZN(_03263_ ) );
AND3_X1 _10898_ ( .A1(_03262_ ), .A2(\IF_ID_inst [12] ), .A3(_03263_ ), .ZN(_03264_ ) );
NAND2_X1 _10899_ ( .A1(_03261_ ), .A2(_03264_ ), .ZN(_03265_ ) );
OAI21_X1 _10900_ ( .A(_03257_ ), .B1(_03260_ ), .B2(_03265_ ), .ZN(_03266_ ) );
AND2_X1 _10901_ ( .A1(_03246_ ), .A2(_03247_ ), .ZN(_03267_ ) );
NAND2_X1 _10902_ ( .A1(_03220_ ), .A2(\IF_ID_inst [28] ), .ZN(_03268_ ) );
NOR3_X1 _10903_ ( .A1(_03268_ ), .A2(\IF_ID_inst [30] ), .A3(_03230_ ), .ZN(_03269_ ) );
AND3_X1 _10904_ ( .A1(_03248_ ), .A2(\IF_ID_inst [21] ), .A3(_03229_ ), .ZN(_03270_ ) );
AND4_X1 _10905_ ( .A1(_03267_ ), .A2(_03269_ ), .A3(_03270_ ), .A4(_03253_ ), .ZN(_03271_ ) );
AND2_X1 _10906_ ( .A1(_03245_ ), .A2(_03271_ ), .ZN(_03272_ ) );
INV_X1 _10907_ ( .A(\IF_ID_inst [4] ), .ZN(_03273_ ) );
NAND4_X1 _10908_ ( .A1(_03273_ ), .A2(\IF_ID_inst [5] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [6] ), .ZN(_03274_ ) );
NOR2_X1 _10909_ ( .A1(_03211_ ), .A2(_03274_ ), .ZN(_03275_ ) );
AND2_X1 _10910_ ( .A1(\IF_ID_inst [14] ), .A2(\IF_ID_inst [13] ), .ZN(_03276_ ) );
AND2_X1 _10911_ ( .A1(_03275_ ), .A2(_03276_ ), .ZN(_03277_ ) );
NOR3_X1 _10912_ ( .A1(_03266_ ), .A2(_03272_ ), .A3(_03277_ ), .ZN(_03278_ ) );
NOR2_X1 _10913_ ( .A1(_03263_ ), .A2(\IF_ID_inst [12] ), .ZN(_03279_ ) );
INV_X1 _10914_ ( .A(\IF_ID_inst [5] ), .ZN(_03280_ ) );
NOR2_X1 _10915_ ( .A1(_03280_ ), .A2(\IF_ID_inst [4] ), .ZN(_03281_ ) );
AND2_X1 _10916_ ( .A1(_03279_ ), .A2(_03281_ ), .ZN(_03282_ ) );
BUF_X2 _10917_ ( .A(_03210_ ), .Z(_03283_ ) );
AND2_X1 _10918_ ( .A1(_03282_ ), .A2(_03283_ ), .ZN(_03284_ ) );
NAND2_X1 _10919_ ( .A1(_03284_ ), .A2(_03259_ ), .ZN(_03285_ ) );
AND2_X1 _10920_ ( .A1(_03284_ ), .A2(\IF_ID_inst [14] ), .ZN(_03286_ ) );
NOR3_X1 _10921_ ( .A1(_03211_ ), .A2(\IF_ID_inst [13] ), .A3(_03274_ ), .ZN(_03287_ ) );
NOR2_X1 _10922_ ( .A1(_03286_ ), .A2(_03287_ ), .ZN(_03288_ ) );
NOR2_X1 _10923_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03289_ ) );
AND3_X1 _10924_ ( .A1(_03210_ ), .A2(_03281_ ), .A3(_03289_ ), .ZN(_03290_ ) );
INV_X1 _10925_ ( .A(\IF_ID_inst [13] ), .ZN(_03291_ ) );
NOR2_X1 _10926_ ( .A1(_03291_ ), .A2(\IF_ID_inst [14] ), .ZN(_03292_ ) );
AND2_X1 _10927_ ( .A1(_03290_ ), .A2(_03292_ ), .ZN(_03293_ ) );
INV_X1 _10928_ ( .A(_03293_ ), .ZN(_03294_ ) );
AND2_X1 _10929_ ( .A1(_03290_ ), .A2(_03259_ ), .ZN(_03295_ ) );
AND4_X1 _10930_ ( .A1(_03273_ ), .A2(_03263_ ), .A3(\IF_ID_inst [5] ), .A4(\IF_ID_inst [12] ), .ZN(_03296_ ) );
AND2_X1 _10931_ ( .A1(_03283_ ), .A2(_03296_ ), .ZN(_03297_ ) );
AND2_X1 _10932_ ( .A1(_03297_ ), .A2(_03259_ ), .ZN(_03298_ ) );
NOR2_X1 _10933_ ( .A1(_03295_ ), .A2(_03298_ ), .ZN(_03299_ ) );
AND4_X1 _10934_ ( .A1(_03285_ ), .A2(_03288_ ), .A3(_03294_ ), .A4(_03299_ ), .ZN(_03300_ ) );
AND4_X1 _10935_ ( .A1(\IF_ID_inst [11] ), .A2(_03278_ ), .A3(_03300_ ), .A4(_03222_ ), .ZN(_00245_ ) );
AND4_X1 _10936_ ( .A1(\IF_ID_inst [10] ), .A2(_03278_ ), .A3(_03300_ ), .A4(_03222_ ), .ZN(_00246_ ) );
AND4_X1 _10937_ ( .A1(\IF_ID_inst [9] ), .A2(_03278_ ), .A3(_03300_ ), .A4(_03222_ ), .ZN(_00247_ ) );
AND4_X1 _10938_ ( .A1(\IF_ID_inst [8] ), .A2(_03278_ ), .A3(_03300_ ), .A4(_03222_ ), .ZN(_00248_ ) );
AND4_X1 _10939_ ( .A1(\IF_ID_inst [7] ), .A2(_03278_ ), .A3(_03300_ ), .A4(_03222_ ), .ZN(_00249_ ) );
INV_X1 _10940_ ( .A(\IF_ID_inst [19] ), .ZN(_03301_ ) );
INV_X1 _10941_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03302_ ) );
AND2_X1 _10942_ ( .A1(_03281_ ), .A2(_03302_ ), .ZN(_03303_ ) );
AND2_X2 _10943_ ( .A1(_03303_ ), .A2(_03261_ ), .ZN(_03304_ ) );
CLKBUF_X2 _10944_ ( .A(_03304_ ), .Z(_03305_ ) );
CLKBUF_X2 _10945_ ( .A(_03305_ ), .Z(_03306_ ) );
NAND3_X1 _10946_ ( .A1(\IF_ID_inst [2] ), .A2(\IF_ID_inst [0] ), .A3(\IF_ID_inst [1] ), .ZN(_03307_ ) );
NOR2_X1 _10947_ ( .A1(_03307_ ), .A2(\IF_ID_inst [3] ), .ZN(_03308_ ) );
NOR2_X1 _10948_ ( .A1(_03273_ ), .A2(\IF_ID_inst [6] ), .ZN(_03309_ ) );
AND2_X1 _10949_ ( .A1(_03308_ ), .A2(_03309_ ), .ZN(_03310_ ) );
NOR2_X1 _10950_ ( .A1(_03306_ ), .A2(_03310_ ), .ZN(_03311_ ) );
INV_X1 _10951_ ( .A(\IF_ID_inst [15] ), .ZN(_03312_ ) );
AND4_X1 _10952_ ( .A1(_03213_ ), .A2(_03240_ ), .A3(_03312_ ), .A4(\IF_ID_inst [6] ), .ZN(_03313_ ) );
AND3_X1 _10953_ ( .A1(_03313_ ), .A2(_03212_ ), .A3(_03258_ ), .ZN(_03314_ ) );
NAND3_X1 _10954_ ( .A1(_03314_ ), .A2(_03283_ ), .A3(_03243_ ), .ZN(_03315_ ) );
NAND4_X1 _10955_ ( .A1(_03269_ ), .A2(_03270_ ), .A3(_03267_ ), .A4(_03253_ ), .ZN(_03316_ ) );
OAI21_X1 _10956_ ( .A(_03311_ ), .B1(_03315_ ), .B2(_03316_ ), .ZN(_03317_ ) );
NOR4_X1 _10957_ ( .A1(_03266_ ), .A2(_03301_ ), .A3(_03233_ ), .A4(_03317_ ), .ZN(_00250_ ) );
INV_X1 _10958_ ( .A(\IF_ID_inst [18] ), .ZN(_03318_ ) );
NOR4_X1 _10959_ ( .A1(_03266_ ), .A2(_03318_ ), .A3(_03233_ ), .A4(_03317_ ), .ZN(_00251_ ) );
INV_X1 _10960_ ( .A(\IF_ID_inst [17] ), .ZN(_03319_ ) );
NOR4_X1 _10961_ ( .A1(_03266_ ), .A2(_03319_ ), .A3(_03233_ ), .A4(_03317_ ), .ZN(_00252_ ) );
NOR2_X1 _10962_ ( .A1(_03266_ ), .A2(_03317_ ), .ZN(_03320_ ) );
NOR3_X1 _10963_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_03321_ ) );
AND2_X1 _10964_ ( .A1(_03321_ ), .A2(_03232_ ), .ZN(_03322_ ) );
INV_X1 _10965_ ( .A(\IF_ID_inst [14] ), .ZN(_03323_ ) );
AND3_X1 _10966_ ( .A1(_03251_ ), .A2(_03323_ ), .A3(\IF_ID_inst [13] ), .ZN(_03324_ ) );
AND3_X1 _10967_ ( .A1(_03322_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03324_ ), .ZN(_03325_ ) );
AND2_X2 _10968_ ( .A1(_03210_ ), .A2(_03289_ ), .ZN(_03326_ ) );
AND3_X1 _10969_ ( .A1(_03325_ ), .A2(_03212_ ), .A3(_03326_ ), .ZN(_03327_ ) );
AND2_X1 _10970_ ( .A1(_03258_ ), .A2(_03251_ ), .ZN(_03328_ ) );
NOR2_X1 _10971_ ( .A1(_03225_ ), .A2(\IF_ID_inst [29] ), .ZN(_03329_ ) );
NOR2_X1 _10972_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_03330_ ) );
AND3_X1 _10973_ ( .A1(_03329_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03330_ ), .ZN(_03331_ ) );
AND4_X1 _10974_ ( .A1(_03212_ ), .A2(_03326_ ), .A3(_03328_ ), .A4(_03331_ ), .ZN(_03332_ ) );
NOR2_X1 _10975_ ( .A1(_03327_ ), .A2(_03332_ ), .ZN(_03333_ ) );
INV_X1 _10976_ ( .A(_03333_ ), .ZN(_03334_ ) );
AND4_X1 _10977_ ( .A1(\IF_ID_inst [4] ), .A2(_03280_ ), .A3(_03263_ ), .A4(\IF_ID_inst [12] ), .ZN(_03335_ ) );
AND2_X1 _10978_ ( .A1(_03210_ ), .A2(_03335_ ), .ZN(_03336_ ) );
AND3_X1 _10979_ ( .A1(_03321_ ), .A2(_03232_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03337_ ) );
AND3_X1 _10980_ ( .A1(_03336_ ), .A2(_03328_ ), .A3(_03337_ ), .ZN(_03338_ ) );
NOR2_X1 _10981_ ( .A1(_03273_ ), .A2(\IF_ID_inst [5] ), .ZN(_03339_ ) );
AND2_X1 _10982_ ( .A1(_03326_ ), .A2(_03339_ ), .ZN(_03340_ ) );
INV_X1 _10983_ ( .A(_03292_ ), .ZN(_03341_ ) );
AND2_X1 _10984_ ( .A1(_03340_ ), .A2(_03341_ ), .ZN(_03342_ ) );
AND3_X1 _10985_ ( .A1(_03210_ ), .A2(_03335_ ), .A3(\IF_ID_inst [13] ), .ZN(_03343_ ) );
AND2_X1 _10986_ ( .A1(_03343_ ), .A2(\IF_ID_inst [14] ), .ZN(_03344_ ) );
NOR4_X1 _10987_ ( .A1(_03334_ ), .A2(_03338_ ), .A3(_03342_ ), .A4(_03344_ ), .ZN(_03345_ ) );
AND2_X1 _10988_ ( .A1(_03326_ ), .A2(_03262_ ), .ZN(_03346_ ) );
AND2_X1 _10989_ ( .A1(_03346_ ), .A2(_03292_ ), .ZN(_03347_ ) );
INV_X1 _10990_ ( .A(_03347_ ), .ZN(_03348_ ) );
AND3_X1 _10991_ ( .A1(_03279_ ), .A2(_03281_ ), .A3(_03258_ ), .ZN(_03349_ ) );
AND2_X1 _10992_ ( .A1(_03349_ ), .A2(_03308_ ), .ZN(_03350_ ) );
INV_X1 _10993_ ( .A(_03350_ ), .ZN(_03351_ ) );
AND4_X1 _10994_ ( .A1(_03218_ ), .A2(_03348_ ), .A3(_03285_ ), .A4(_03351_ ), .ZN(_03352_ ) );
AND2_X1 _10995_ ( .A1(_03340_ ), .A2(_03292_ ), .ZN(_03353_ ) );
INV_X1 _10996_ ( .A(_03353_ ), .ZN(_03354_ ) );
AND3_X1 _10997_ ( .A1(_03326_ ), .A2(_03291_ ), .A3(_03262_ ), .ZN(_03355_ ) );
AND2_X1 _10998_ ( .A1(_03264_ ), .A2(_03210_ ), .ZN(_03356_ ) );
AND2_X1 _10999_ ( .A1(_03356_ ), .A2(_03291_ ), .ZN(_03357_ ) );
NOR2_X1 _11000_ ( .A1(_03355_ ), .A2(_03357_ ), .ZN(_03358_ ) );
NAND2_X1 _11001_ ( .A1(_03343_ ), .A2(_03323_ ), .ZN(_03359_ ) );
AND3_X1 _11002_ ( .A1(_03354_ ), .A2(_03358_ ), .A3(_03359_ ), .ZN(_03360_ ) );
AND4_X1 _11003_ ( .A1(_03320_ ), .A2(_03345_ ), .A3(_03352_ ), .A4(_03360_ ), .ZN(_03361_ ) );
INV_X1 _11004_ ( .A(_03277_ ), .ZN(_03362_ ) );
AND2_X1 _11005_ ( .A1(_03337_ ), .A2(_03328_ ), .ZN(_03363_ ) );
NOR2_X1 _11006_ ( .A1(_03323_ ), .A2(\IF_ID_inst [13] ), .ZN(_03364_ ) );
AND2_X1 _11007_ ( .A1(_03364_ ), .A2(_03251_ ), .ZN(_03365_ ) );
AND2_X1 _11008_ ( .A1(_03337_ ), .A2(_03365_ ), .ZN(_03366_ ) );
OAI211_X1 _11009_ ( .A(_03212_ ), .B(_03326_ ), .C1(_03363_ ), .C2(_03366_ ), .ZN(_03367_ ) );
AND3_X1 _11010_ ( .A1(_03276_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03251_ ), .ZN(_03368_ ) );
AND3_X1 _11011_ ( .A1(_03368_ ), .A2(_03232_ ), .A3(_03321_ ), .ZN(_03369_ ) );
AND3_X1 _11012_ ( .A1(_03207_ ), .A2(\IF_ID_inst [12] ), .A3(_03208_ ), .ZN(_03370_ ) );
AND3_X1 _11013_ ( .A1(_03263_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_03371_ ) );
AND2_X1 _11014_ ( .A1(_03370_ ), .A2(_03371_ ), .ZN(_03372_ ) );
NAND2_X1 _11015_ ( .A1(_03369_ ), .A2(_03372_ ), .ZN(_03373_ ) );
NAND3_X1 _11016_ ( .A1(_03372_ ), .A2(_03331_ ), .A3(_03365_ ), .ZN(_03374_ ) );
NAND3_X1 _11017_ ( .A1(_03369_ ), .A2(_03212_ ), .A3(_03326_ ), .ZN(_03375_ ) );
NAND4_X1 _11018_ ( .A1(_03367_ ), .A2(_03373_ ), .A3(_03374_ ), .A4(_03375_ ), .ZN(_03376_ ) );
INV_X1 _11019_ ( .A(_03372_ ), .ZN(_03377_ ) );
NOR2_X1 _11020_ ( .A1(_03325_ ), .A2(_03366_ ), .ZN(_03378_ ) );
INV_X1 _11021_ ( .A(_03363_ ), .ZN(_03379_ ) );
AOI21_X1 _11022_ ( .A(_03377_ ), .B1(_03378_ ), .B2(_03379_ ), .ZN(_03380_ ) );
NOR2_X1 _11023_ ( .A1(_03376_ ), .A2(_03380_ ), .ZN(_03381_ ) );
OAI21_X1 _11024_ ( .A(_03259_ ), .B1(_03290_ ), .B2(_03297_ ), .ZN(_03382_ ) );
AND2_X1 _11025_ ( .A1(_03331_ ), .A2(_03365_ ), .ZN(_03383_ ) );
OAI21_X1 _11026_ ( .A(_03336_ ), .B1(_03366_ ), .B2(_03383_ ), .ZN(_03384_ ) );
AND3_X1 _11027_ ( .A1(_03294_ ), .A2(_03382_ ), .A3(_03384_ ), .ZN(_03385_ ) );
AND4_X1 _11028_ ( .A1(_03362_ ), .A2(_03381_ ), .A3(_03288_ ), .A4(_03385_ ), .ZN(_03386_ ) );
AND2_X1 _11029_ ( .A1(_03361_ ), .A2(_03386_ ), .ZN(_03387_ ) );
BUF_X4 _11030_ ( .A(_03387_ ), .Z(_03388_ ) );
INV_X1 _11031_ ( .A(_03388_ ), .ZN(_03389_ ) );
XNOR2_X1 _11032_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_03390_ ) );
XNOR2_X1 _11033_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_03391_ ) );
XNOR2_X1 _11034_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_03392_ ) );
XNOR2_X1 _11035_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_03393_ ) );
AND4_X1 _11036_ ( .A1(_03390_ ), .A2(_03391_ ), .A3(_03392_ ), .A4(_03393_ ), .ZN(_03394_ ) );
XNOR2_X1 _11037_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .ZN(_03395_ ) );
XNOR2_X1 _11038_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .ZN(_03396_ ) );
XNOR2_X1 _11039_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_03397_ ) );
XNOR2_X1 _11040_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_03398_ ) );
AND4_X1 _11041_ ( .A1(_03395_ ), .A2(_03396_ ), .A3(_03397_ ), .A4(_03398_ ), .ZN(_03399_ ) );
XNOR2_X1 _11042_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_03400_ ) );
XNOR2_X1 _11043_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_03401_ ) );
XNOR2_X1 _11044_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_03402_ ) );
XNOR2_X1 _11045_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_03403_ ) );
AND4_X1 _11046_ ( .A1(_03400_ ), .A2(_03401_ ), .A3(_03402_ ), .A4(_03403_ ), .ZN(_03404_ ) );
XNOR2_X1 _11047_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_03405_ ) );
XNOR2_X1 _11048_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_03406_ ) );
XNOR2_X1 _11049_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_03407_ ) );
XNOR2_X1 _11050_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .ZN(_03408_ ) );
AND4_X1 _11051_ ( .A1(_03405_ ), .A2(_03406_ ), .A3(_03407_ ), .A4(_03408_ ), .ZN(_03409_ ) );
AND4_X1 _11052_ ( .A1(_03394_ ), .A2(_03399_ ), .A3(_03404_ ), .A4(_03409_ ), .ZN(_03410_ ) );
XNOR2_X1 _11053_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_03411_ ) );
XNOR2_X1 _11054_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_03412_ ) );
XNOR2_X1 _11055_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .ZN(_03413_ ) );
XNOR2_X1 _11056_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .ZN(_03414_ ) );
AND4_X1 _11057_ ( .A1(_03411_ ), .A2(_03412_ ), .A3(_03413_ ), .A4(_03414_ ), .ZN(_03415_ ) );
XNOR2_X1 _11058_ ( .A(fanout_net_9 ), .B(\myexu.pc_jump [3] ), .ZN(_03416_ ) );
XNOR2_X1 _11059_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .ZN(_03417_ ) );
XNOR2_X1 _11060_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .ZN(_03418_ ) );
INV_X1 _11061_ ( .A(\IF_ID_pc [2] ), .ZN(_03419_ ) );
AOI22_X1 _11062_ ( .A1(_01962_ ), .A2(\myexu.pc_jump [25] ), .B1(_03419_ ), .B2(\myexu.pc_jump [2] ), .ZN(_03420_ ) );
AND4_X1 _11063_ ( .A1(_03416_ ), .A2(_03417_ ), .A3(_03418_ ), .A4(_03420_ ), .ZN(_03421_ ) );
XNOR2_X1 _11064_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .ZN(_03422_ ) );
INV_X1 _11065_ ( .A(\myexu.pc_jump [21] ), .ZN(_03423_ ) );
OAI221_X1 _11066_ ( .A(_03422_ ), .B1(\IF_ID_pc [21] ), .B2(_03423_ ), .C1(_01962_ ), .C2(\myexu.pc_jump [25] ), .ZN(_03424_ ) );
AOI22_X1 _11067_ ( .A1(_02039_ ), .A2(\myexu.pc_jump [29] ), .B1(_03423_ ), .B2(\IF_ID_pc [21] ), .ZN(_03425_ ) );
INV_X1 _11068_ ( .A(fanout_net_13 ), .ZN(_03426_ ) );
OAI221_X1 _11069_ ( .A(_03425_ ), .B1(_03426_ ), .B2(\myexu.pc_jump [4] ), .C1(_02039_ ), .C2(\myexu.pc_jump [29] ), .ZN(_03427_ ) );
XNOR2_X1 _11070_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_03428_ ) );
XNOR2_X1 _11071_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .ZN(_03429_ ) );
INV_X1 _11072_ ( .A(\IF_ID_pc [1] ), .ZN(_03430_ ) );
AOI22_X1 _11073_ ( .A1(_03426_ ), .A2(\myexu.pc_jump [4] ), .B1(_03430_ ), .B2(\myexu.pc_jump [1] ), .ZN(_03431_ ) );
INV_X1 _11074_ ( .A(\myexu.pc_jump [1] ), .ZN(_03432_ ) );
INV_X1 _11075_ ( .A(\myexu.pc_jump [2] ), .ZN(_03433_ ) );
AOI22_X1 _11076_ ( .A1(_03432_ ), .A2(\IF_ID_pc [1] ), .B1(_03433_ ), .B2(\IF_ID_pc [2] ), .ZN(_03434_ ) );
NAND4_X1 _11077_ ( .A1(_03428_ ), .A2(_03429_ ), .A3(_03431_ ), .A4(_03434_ ), .ZN(_03435_ ) );
NOR3_X1 _11078_ ( .A1(_03424_ ), .A2(_03427_ ), .A3(_03435_ ), .ZN(_03436_ ) );
AND4_X1 _11079_ ( .A1(_03410_ ), .A2(_03415_ ), .A3(_03421_ ), .A4(_03436_ ), .ZN(_03437_ ) );
INV_X1 _11080_ ( .A(check_quest ), .ZN(_03438_ ) );
NOR2_X2 _11081_ ( .A1(_03437_ ), .A2(_03438_ ), .ZN(_03439_ ) );
INV_X1 _11082_ ( .A(\myifu.state [1] ), .ZN(_03440_ ) );
NOR2_X1 _11083_ ( .A1(_03440_ ), .A2(\myifu.to_reset ), .ZN(_03441_ ) );
INV_X1 _11084_ ( .A(_03441_ ), .ZN(_03442_ ) );
NOR2_X1 _11085_ ( .A1(_03439_ ), .A2(_03442_ ), .ZN(_03443_ ) );
AND2_X2 _11086_ ( .A1(_03443_ ), .A2(IDU_ready_IFU ), .ZN(_03444_ ) );
NAND4_X1 _11087_ ( .A1(_03389_ ), .A2(\IF_ID_inst [18] ), .A3(_03320_ ), .A4(_03444_ ), .ZN(_03445_ ) );
INV_X1 _11088_ ( .A(_03444_ ), .ZN(_03446_ ) );
BUF_X4 _11089_ ( .A(_03446_ ), .Z(_03447_ ) );
OAI21_X1 _11090_ ( .A(\ID_EX_rs1 [3] ), .B1(_03388_ ), .B2(_03447_ ), .ZN(_03448_ ) );
AOI21_X1 _11091_ ( .A(_03227_ ), .B1(_03445_ ), .B2(_03448_ ), .ZN(_00253_ ) );
INV_X1 _11092_ ( .A(\IF_ID_inst [16] ), .ZN(_03449_ ) );
NOR4_X1 _11093_ ( .A1(_03266_ ), .A2(_03449_ ), .A3(_03233_ ), .A4(_03317_ ), .ZN(_00254_ ) );
NAND4_X1 _11094_ ( .A1(_03389_ ), .A2(\IF_ID_inst [17] ), .A3(_03320_ ), .A4(_03444_ ), .ZN(_03450_ ) );
OAI21_X1 _11095_ ( .A(\ID_EX_rs1 [2] ), .B1(_03388_ ), .B2(_03447_ ), .ZN(_03451_ ) );
AOI21_X1 _11096_ ( .A(_03227_ ), .B1(_03450_ ), .B2(_03451_ ), .ZN(_00255_ ) );
NOR4_X1 _11097_ ( .A1(_03266_ ), .A2(_03312_ ), .A3(_03223_ ), .A4(_03317_ ), .ZN(_00256_ ) );
BUF_X2 _11098_ ( .A(_03222_ ), .Z(_03452_ ) );
NOR2_X1 _11099_ ( .A1(_03388_ ), .A2(_03447_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OAI21_X1 _11100_ ( .A(_03452_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [1] ), .ZN(_03453_ ) );
AOI221_X4 _11101_ ( .A(_03447_ ), .B1(\IF_ID_inst [16] ), .B2(_03320_ ), .C1(_03361_ ), .C2(_03386_ ), .ZN(_03454_ ) );
NOR2_X1 _11102_ ( .A1(_03453_ ), .A2(_03454_ ), .ZN(_00257_ ) );
NOR2_X1 _11103_ ( .A1(_03342_ ), .A2(_03343_ ), .ZN(_03455_ ) );
OR2_X1 _11104_ ( .A1(_03350_ ), .A2(_03306_ ), .ZN(_03456_ ) );
AOI21_X1 _11105_ ( .A(_03456_ ), .B1(_03292_ ), .B2(_03346_ ), .ZN(_03457_ ) );
NAND3_X1 _11106_ ( .A1(_03455_ ), .A2(_03457_ ), .A3(_03358_ ), .ZN(_03458_ ) );
AND3_X1 _11107_ ( .A1(_03314_ ), .A2(_03210_ ), .A3(_03243_ ), .ZN(_03459_ ) );
AND4_X1 _11108_ ( .A1(_03267_ ), .A2(_03269_ ), .A3(_03270_ ), .A4(_03253_ ), .ZN(_03460_ ) );
AND2_X1 _11109_ ( .A1(_03459_ ), .A2(_03460_ ), .ZN(_03461_ ) );
INV_X1 _11110_ ( .A(_03261_ ), .ZN(_03462_ ) );
NAND4_X1 _11111_ ( .A1(_03259_ ), .A2(_03262_ ), .A3(\IF_ID_inst [12] ), .A4(_03263_ ), .ZN(_03463_ ) );
NOR2_X1 _11112_ ( .A1(_03462_ ), .A2(_03463_ ), .ZN(_03464_ ) );
OR2_X1 _11113_ ( .A1(_03461_ ), .A2(_03464_ ), .ZN(_03465_ ) );
NAND4_X1 _11114_ ( .A1(_03283_ ), .A2(_03313_ ), .A3(_03212_ ), .A4(_03259_ ), .ZN(_03466_ ) );
NOR4_X1 _11115_ ( .A1(_03466_ ), .A2(_03250_ ), .A3(\IF_ID_inst [8] ), .A4(_03242_ ), .ZN(_03467_ ) );
NOR2_X1 _11116_ ( .A1(_03254_ ), .A2(_03255_ ), .ZN(_03468_ ) );
AND2_X1 _11117_ ( .A1(_03467_ ), .A2(_03468_ ), .ZN(_03469_ ) );
NOR4_X1 _11118_ ( .A1(_03458_ ), .A2(_03465_ ), .A3(_03228_ ), .A4(_03469_ ), .ZN(_03470_ ) );
NOR2_X1 _11119_ ( .A1(_03353_ ), .A2(_03310_ ), .ZN(_03471_ ) );
OR2_X1 _11120_ ( .A1(_03366_ ), .A2(_03383_ ), .ZN(_03472_ ) );
AOI21_X1 _11121_ ( .A(_03338_ ), .B1(_03472_ ), .B2(_03336_ ), .ZN(_03473_ ) );
AND2_X1 _11122_ ( .A1(_03471_ ), .A2(_03473_ ), .ZN(_03474_ ) );
AND4_X1 _11123_ ( .A1(\IF_ID_inst [24] ), .A2(_03470_ ), .A3(_03452_ ), .A4(_03474_ ), .ZN(_00258_ ) );
NAND4_X1 _11124_ ( .A1(_03389_ ), .A2(\IF_ID_inst [15] ), .A3(_03320_ ), .A4(_03444_ ), .ZN(_03475_ ) );
OAI21_X1 _11125_ ( .A(\ID_EX_rs1 [0] ), .B1(_03388_ ), .B2(_03447_ ), .ZN(_03476_ ) );
AOI21_X1 _11126_ ( .A(_03227_ ), .B1(_03475_ ), .B2(_03476_ ), .ZN(_00259_ ) );
AND4_X1 _11127_ ( .A1(\IF_ID_inst [23] ), .A2(_03470_ ), .A3(_03452_ ), .A4(_03474_ ), .ZN(_00260_ ) );
AND4_X1 _11128_ ( .A1(\IF_ID_inst [22] ), .A2(_03470_ ), .A3(_03452_ ), .A4(_03474_ ), .ZN(_00261_ ) );
AND2_X1 _11129_ ( .A1(_03470_ ), .A2(_03474_ ), .ZN(_03477_ ) );
AOI221_X4 _11130_ ( .A(_03446_ ), .B1(_03361_ ), .B2(_03386_ ), .C1(\IF_ID_inst [23] ), .C2(_03477_ ), .ZN(_03478_ ) );
INV_X1 _11131_ ( .A(\ID_EX_rs2 [3] ), .ZN(_03479_ ) );
INV_X1 _11132_ ( .A(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .ZN(_03480_ ) );
AOI211_X1 _11133_ ( .A(_03223_ ), .B(_03478_ ), .C1(_03479_ ), .C2(_03480_ ), .ZN(_00262_ ) );
AND4_X1 _11134_ ( .A1(\IF_ID_inst [21] ), .A2(_03470_ ), .A3(_03222_ ), .A4(_03474_ ), .ZN(_00263_ ) );
NAND4_X1 _11135_ ( .A1(_03389_ ), .A2(\IF_ID_inst [22] ), .A3(_03444_ ), .A4(_03477_ ), .ZN(_03481_ ) );
OAI21_X1 _11136_ ( .A(\ID_EX_rs2 [2] ), .B1(_03388_ ), .B2(_03447_ ), .ZN(_03482_ ) );
AOI21_X1 _11137_ ( .A(_03227_ ), .B1(_03481_ ), .B2(_03482_ ), .ZN(_00264_ ) );
AND4_X1 _11138_ ( .A1(\IF_ID_inst [20] ), .A2(_03470_ ), .A3(_03222_ ), .A4(_03474_ ), .ZN(_00265_ ) );
OAI21_X1 _11139_ ( .A(_03452_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs2 [1] ), .ZN(_03483_ ) );
AOI221_X4 _11140_ ( .A(_03446_ ), .B1(_03361_ ), .B2(_03386_ ), .C1(\IF_ID_inst [21] ), .C2(_03477_ ), .ZN(_03484_ ) );
NOR2_X1 _11141_ ( .A1(_03483_ ), .A2(_03484_ ), .ZN(_00266_ ) );
NOR4_X1 _11142_ ( .A1(_03462_ ), .A2(_03233_ ), .A3(IDU_valid_EXU ), .A4(_03463_ ), .ZN(_00267_ ) );
NAND4_X1 _11143_ ( .A1(_03389_ ), .A2(\IF_ID_inst [20] ), .A3(_03444_ ), .A4(_03477_ ), .ZN(_03485_ ) );
OAI21_X1 _11144_ ( .A(\ID_EX_rs2 [0] ), .B1(_03388_ ), .B2(_03447_ ), .ZN(_03486_ ) );
AOI21_X1 _11145_ ( .A(_03227_ ), .B1(_03485_ ), .B2(_03486_ ), .ZN(_00268_ ) );
XNOR2_X1 _11146_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_03487_ ) );
XNOR2_X1 _11147_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_03488_ ) );
XNOR2_X1 _11148_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_03489_ ) );
XNOR2_X1 _11149_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_03490_ ) );
AND4_X1 _11150_ ( .A1(_03487_ ), .A2(_03488_ ), .A3(_03489_ ), .A4(_03490_ ), .ZN(_03491_ ) );
XNOR2_X1 _11151_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_03492_ ) );
AND2_X1 _11152_ ( .A1(_03491_ ), .A2(_03492_ ), .ZN(_03493_ ) );
AND2_X1 _11153_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03494_ ) );
INV_X1 _11154_ ( .A(\ID_EX_typ [7] ), .ZN(_03495_ ) );
AND2_X1 _11155_ ( .A1(_03494_ ), .A2(_03495_ ), .ZN(_03496_ ) );
AND2_X1 _11156_ ( .A1(_03493_ ), .A2(_03496_ ), .ZN(_03497_ ) );
INV_X1 _11157_ ( .A(_03497_ ), .ZN(_03498_ ) );
XNOR2_X1 _11158_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_03499_ ) );
XNOR2_X1 _11159_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_03500_ ) );
XNOR2_X1 _11160_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_03501_ ) );
XNOR2_X1 _11161_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_03502_ ) );
AND4_X1 _11162_ ( .A1(_03499_ ), .A2(_03500_ ), .A3(_03501_ ), .A4(_03502_ ), .ZN(_03503_ ) );
XNOR2_X1 _11163_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_03504_ ) );
NAND3_X1 _11164_ ( .A1(_03503_ ), .A2(_03496_ ), .A3(_03504_ ), .ZN(_03505_ ) );
AND2_X1 _11165_ ( .A1(_03498_ ), .A2(_03505_ ), .ZN(_03506_ ) );
NOR3_X1 _11166_ ( .A1(_03506_ ), .A2(_03266_ ), .A3(_03317_ ), .ZN(_03507_ ) );
OR2_X1 _11167_ ( .A1(_03342_ ), .A2(_03344_ ), .ZN(_03508_ ) );
OAI21_X1 _11168_ ( .A(_03346_ ), .B1(_03323_ ), .B2(_03291_ ), .ZN(_03509_ ) );
AOI22_X1 _11169_ ( .A1(_03356_ ), .A2(_03291_ ), .B1(_03349_ ), .B2(_03308_ ), .ZN(_03510_ ) );
NAND4_X1 _11170_ ( .A1(_03354_ ), .A2(_03359_ ), .A3(_03509_ ), .A4(_03510_ ), .ZN(_03511_ ) );
OR4_X1 _11171_ ( .A1(_03228_ ), .A2(_03507_ ), .A3(_03508_ ), .A4(_03511_ ), .ZN(_03512_ ) );
NAND3_X1 _11172_ ( .A1(_03512_ ), .A2(IDU_ready_IFU ), .A3(_03452_ ), .ZN(_03513_ ) );
NOR2_X2 _11173_ ( .A1(_03511_ ), .A2(_03508_ ), .ZN(_03514_ ) );
AOI21_X1 _11174_ ( .A(_03497_ ), .B1(_03514_ ), .B2(_03218_ ), .ZN(_03515_ ) );
NOR2_X1 _11175_ ( .A1(_03513_ ), .A2(_03515_ ), .ZN(_00269_ ) );
NAND4_X1 _11176_ ( .A1(_03314_ ), .A2(_03229_ ), .A3(_03283_ ), .A4(_03243_ ), .ZN(_03516_ ) );
NAND3_X1 _11177_ ( .A1(_03468_ ), .A2(_03226_ ), .A3(_03249_ ), .ZN(_03517_ ) );
NOR2_X1 _11178_ ( .A1(_03516_ ), .A2(_03517_ ), .ZN(_03518_ ) );
NOR4_X1 _11179_ ( .A1(_03465_ ), .A2(_03518_ ), .A3(_03228_ ), .A4(_03456_ ), .ZN(_03519_ ) );
NOR2_X1 _11180_ ( .A1(_03275_ ), .A2(_03284_ ), .ZN(_03520_ ) );
NOR2_X1 _11181_ ( .A1(_03520_ ), .A2(_03292_ ), .ZN(_03521_ ) );
INV_X1 _11182_ ( .A(_03521_ ), .ZN(_03522_ ) );
AOI21_X1 _11183_ ( .A(_03227_ ), .B1(_03519_ ), .B2(_03522_ ), .ZN(_00270_ ) );
AND2_X1 _11184_ ( .A1(_03294_ ), .A2(_03382_ ), .ZN(_03523_ ) );
AND2_X1 _11185_ ( .A1(_03356_ ), .A2(_03364_ ), .ZN(_03524_ ) );
INV_X1 _11186_ ( .A(_03524_ ), .ZN(_03525_ ) );
NAND2_X1 _11187_ ( .A1(_03356_ ), .A2(_03259_ ), .ZN(_03526_ ) );
AND4_X1 _11188_ ( .A1(_03523_ ), .A2(_03525_ ), .A3(_03526_ ), .A4(_03509_ ), .ZN(_03527_ ) );
NOR2_X1 _11189_ ( .A1(_03518_ ), .A2(_03228_ ), .ZN(_03528_ ) );
AOI21_X1 _11190_ ( .A(_03224_ ), .B1(_03527_ ), .B2(_03528_ ), .ZN(_00271_ ) );
NAND4_X1 _11191_ ( .A1(_03322_ ), .A2(_03365_ ), .A3(_03283_ ), .A4(_03335_ ), .ZN(_03529_ ) );
INV_X1 _11192_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03530_ ) );
NOR2_X1 _11193_ ( .A1(_03529_ ), .A2(_03530_ ), .ZN(_03531_ ) );
NAND4_X1 _11194_ ( .A1(_03322_ ), .A2(_03283_ ), .A3(_03335_ ), .A4(_03328_ ), .ZN(_03532_ ) );
NOR2_X1 _11195_ ( .A1(_03532_ ), .A2(_03530_ ), .ZN(_03533_ ) );
NOR2_X1 _11196_ ( .A1(_03531_ ), .A2(_03533_ ), .ZN(_03534_ ) );
AND4_X1 _11197_ ( .A1(_03336_ ), .A2(_03330_ ), .A3(_03329_ ), .A4(_03365_ ), .ZN(_03535_ ) );
NAND2_X1 _11198_ ( .A1(_03535_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03536_ ) );
INV_X1 _11199_ ( .A(_03340_ ), .ZN(_03537_ ) );
OAI211_X1 _11200_ ( .A(_03534_ ), .B(_03536_ ), .C1(_03341_ ), .C2(_03537_ ), .ZN(_03538_ ) );
AND3_X1 _11201_ ( .A1(_03249_ ), .A2(_03226_ ), .A3(_03229_ ), .ZN(_03539_ ) );
AND3_X1 _11202_ ( .A1(_03459_ ), .A2(_03468_ ), .A3(_03539_ ), .ZN(_03540_ ) );
NOR4_X1 _11203_ ( .A1(_03458_ ), .A2(_03310_ ), .A3(_03538_ ), .A4(_03540_ ), .ZN(_03541_ ) );
NOR3_X1 _11204_ ( .A1(_03334_ ), .A2(_03376_ ), .A3(_03380_ ), .ZN(_03542_ ) );
AOI21_X1 _11205_ ( .A(_03224_ ), .B1(_03541_ ), .B2(_03542_ ), .ZN(_00272_ ) );
AOI211_X1 _11206_ ( .A(_03464_ ), .B(_03343_ ), .C1(_03340_ ), .C2(_03341_ ), .ZN(_03543_ ) );
AOI21_X1 _11207_ ( .A(_03224_ ), .B1(_03474_ ), .B2(_03543_ ), .ZN(_00273_ ) );
NAND2_X1 _11208_ ( .A1(_03459_ ), .A2(_03460_ ), .ZN(_03544_ ) );
INV_X1 _11209_ ( .A(_03327_ ), .ZN(_03545_ ) );
NAND4_X1 _11210_ ( .A1(_03326_ ), .A2(_03212_ ), .A3(_03328_ ), .A4(_03331_ ), .ZN(_03546_ ) );
AND4_X1 _11211_ ( .A1(_03544_ ), .A2(_03545_ ), .A3(_03294_ ), .A4(_03546_ ), .ZN(_03547_ ) );
AOI21_X1 _11212_ ( .A(_03224_ ), .B1(_03547_ ), .B2(_03471_ ), .ZN(_00274_ ) );
NAND3_X1 _11213_ ( .A1(_03348_ ), .A2(_03374_ ), .A3(_03359_ ), .ZN(_03548_ ) );
AND2_X1 _11214_ ( .A1(_03275_ ), .A2(\IF_ID_inst [14] ), .ZN(_03549_ ) );
AND3_X1 _11215_ ( .A1(_03283_ ), .A2(\IF_ID_inst [13] ), .A3(_03216_ ), .ZN(_03550_ ) );
OR2_X1 _11216_ ( .A1(_03293_ ), .A2(_03310_ ), .ZN(_03551_ ) );
NOR4_X1 _11217_ ( .A1(_03548_ ), .A2(_03549_ ), .A3(_03550_ ), .A4(_03551_ ), .ZN(_03552_ ) );
AND2_X1 _11218_ ( .A1(_03472_ ), .A2(_03336_ ), .ZN(_03553_ ) );
NOR3_X1 _11219_ ( .A1(_03553_ ), .A2(_03380_ ), .A3(_03338_ ), .ZN(_03554_ ) );
AOI21_X1 _11220_ ( .A(_03224_ ), .B1(_03552_ ), .B2(_03554_ ), .ZN(_00275_ ) );
AND2_X1 _11221_ ( .A1(_03340_ ), .A2(\IF_ID_inst [14] ), .ZN(_03555_ ) );
INV_X1 _11222_ ( .A(_03555_ ), .ZN(_03556_ ) );
OAI22_X1 _11223_ ( .A1(_03366_ ), .A2(_03383_ ), .B1(_03336_ ), .B2(_03372_ ), .ZN(_03557_ ) );
AND4_X1 _11224_ ( .A1(_03525_ ), .A2(_03556_ ), .A3(_03375_ ), .A4(_03557_ ), .ZN(_03558_ ) );
NAND2_X1 _11225_ ( .A1(_03308_ ), .A2(_03371_ ), .ZN(_03559_ ) );
AOI221_X4 _11226_ ( .A(_03215_ ), .B1(_03290_ ), .B2(_03292_ ), .C1(\IF_ID_inst [14] ), .C2(_03284_ ), .ZN(_03560_ ) );
AND3_X1 _11227_ ( .A1(_03366_ ), .A2(_03212_ ), .A3(_03326_ ), .ZN(_03561_ ) );
INV_X1 _11228_ ( .A(_03561_ ), .ZN(_03562_ ) );
OAI211_X1 _11229_ ( .A(_03283_ ), .B(_03259_ ), .C1(_03264_ ), .C2(_03296_ ), .ZN(_03563_ ) );
AND4_X1 _11230_ ( .A1(_03559_ ), .A2(_03560_ ), .A3(_03562_ ), .A4(_03563_ ), .ZN(_03564_ ) );
AOI21_X1 _11231_ ( .A(_03224_ ), .B1(_03558_ ), .B2(_03564_ ), .ZN(_00276_ ) );
OR4_X1 _11232_ ( .A1(_03293_ ), .A2(_03327_ ), .A3(_03344_ ), .A4(_03350_ ), .ZN(_03565_ ) );
NAND2_X1 _11233_ ( .A1(_03275_ ), .A2(_03259_ ), .ZN(_03566_ ) );
INV_X1 _11234_ ( .A(_03338_ ), .ZN(_03567_ ) );
NAND3_X1 _11235_ ( .A1(_03562_ ), .A2(_03566_ ), .A3(_03567_ ), .ZN(_03568_ ) );
NAND2_X1 _11236_ ( .A1(_03459_ ), .A2(_03468_ ), .ZN(_03569_ ) );
OAI21_X1 _11237_ ( .A(_03382_ ), .B1(_03569_ ), .B2(_03250_ ), .ZN(_03570_ ) );
OAI21_X1 _11238_ ( .A(_03372_ ), .B1(_03363_ ), .B2(_03383_ ), .ZN(_03571_ ) );
NAND4_X1 _11239_ ( .A1(_03331_ ), .A2(_03365_ ), .A3(_03283_ ), .A4(_03335_ ), .ZN(_03572_ ) );
NAND4_X1 _11240_ ( .A1(_03525_ ), .A2(_03571_ ), .A3(_03373_ ), .A4(_03572_ ), .ZN(_03573_ ) );
NOR4_X1 _11241_ ( .A1(_03565_ ), .A2(_03568_ ), .A3(_03570_ ), .A4(_03573_ ), .ZN(_03574_ ) );
INV_X1 _11242_ ( .A(_03355_ ), .ZN(_03575_ ) );
OAI211_X1 _11243_ ( .A(_03575_ ), .B(_03218_ ), .C1(_03537_ ), .C2(\IF_ID_inst [13] ), .ZN(_03576_ ) );
NOR2_X1 _11244_ ( .A1(_03520_ ), .A2(_03291_ ), .ZN(_03577_ ) );
OAI21_X1 _11245_ ( .A(\IF_ID_inst [14] ), .B1(_03576_ ), .B2(_03577_ ), .ZN(_03578_ ) );
AOI21_X1 _11246_ ( .A(_03224_ ), .B1(_03574_ ), .B2(_03578_ ), .ZN(_00277_ ) );
INV_X1 _11247_ ( .A(_03437_ ), .ZN(_03579_ ) );
INV_X1 _11248_ ( .A(\myifu.to_reset ), .ZN(_03580_ ) );
BUF_X4 _11249_ ( .A(_03580_ ), .Z(_03581_ ) );
NAND4_X1 _11250_ ( .A1(_03579_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_03581_ ), .ZN(_03582_ ) );
NAND2_X1 _11251_ ( .A1(\mtvec [0] ), .A2(\myifu.to_reset ), .ZN(_03583_ ) );
AOI21_X1 _11252_ ( .A(fanout_net_4 ), .B1(_03582_ ), .B2(_03583_ ), .ZN(_00281_ ) );
AND4_X1 _11253_ ( .A1(\IF_ID_inst [31] ), .A2(_03273_ ), .A3(_03302_ ), .A4(\IF_ID_inst [5] ), .ZN(_03584_ ) );
AND2_X2 _11254_ ( .A1(_03209_ ), .A2(_03584_ ), .ZN(_03585_ ) );
AOI21_X1 _11255_ ( .A(_03585_ ), .B1(_03306_ ), .B2(\IF_ID_inst [31] ), .ZN(_03586_ ) );
NAND4_X1 _11256_ ( .A1(_03281_ ), .A2(_03302_ ), .A3(_03207_ ), .A4(_03208_ ), .ZN(_03587_ ) );
NOR2_X1 _11257_ ( .A1(_03587_ ), .A2(_03220_ ), .ZN(_03588_ ) );
AND2_X1 _11258_ ( .A1(_03588_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03589_ ) );
NOR3_X1 _11259_ ( .A1(_03586_ ), .A2(_03589_ ), .A3(_02039_ ), .ZN(_03590_ ) );
AND2_X1 _11260_ ( .A1(_03585_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03591_ ) );
NOR2_X1 _11261_ ( .A1(_03586_ ), .A2(_03591_ ), .ZN(_03592_ ) );
BUF_X4 _11262_ ( .A(_03592_ ), .Z(_03593_ ) );
BUF_X2 _11263_ ( .A(_03593_ ), .Z(_03594_ ) );
XNOR2_X1 _11264_ ( .A(_03594_ ), .B(_02039_ ), .ZN(_03595_ ) );
INV_X1 _11265_ ( .A(_03595_ ), .ZN(_03596_ ) );
XNOR2_X1 _11266_ ( .A(_03593_ ), .B(_01971_ ), .ZN(_03597_ ) );
XOR2_X1 _11267_ ( .A(_03593_ ), .B(\IF_ID_pc [27] ), .Z(_03598_ ) );
XNOR2_X1 _11268_ ( .A(_03593_ ), .B(_01903_ ), .ZN(_03599_ ) );
XNOR2_X1 _11269_ ( .A(_03593_ ), .B(_01962_ ), .ZN(_03600_ ) );
AND4_X1 _11270_ ( .A1(_03597_ ), .A2(_03598_ ), .A3(_03599_ ), .A4(_03600_ ), .ZN(_03601_ ) );
AND2_X1 _11271_ ( .A1(_03305_ ), .A2(\IF_ID_inst [27] ), .ZN(_03602_ ) );
INV_X1 _11272_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03603_ ) );
AOI21_X1 _11273_ ( .A(_03602_ ), .B1(_03603_ ), .B2(_03585_ ), .ZN(_03604_ ) );
XNOR2_X1 _11274_ ( .A(_03604_ ), .B(\IF_ID_pc [7] ), .ZN(_03605_ ) );
INV_X1 _11275_ ( .A(_03585_ ), .ZN(_03606_ ) );
NOR2_X1 _11276_ ( .A1(_03606_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03607_ ) );
AND2_X1 _11277_ ( .A1(_03305_ ), .A2(\IF_ID_inst [25] ), .ZN(_03608_ ) );
NOR2_X1 _11278_ ( .A1(_03607_ ), .A2(_03608_ ), .ZN(_03609_ ) );
INV_X1 _11279_ ( .A(\IF_ID_pc [5] ), .ZN(_03610_ ) );
XNOR2_X1 _11280_ ( .A(_03609_ ), .B(_03610_ ), .ZN(_03611_ ) );
AND2_X1 _11281_ ( .A1(_03304_ ), .A2(\IF_ID_inst [26] ), .ZN(_03612_ ) );
INV_X1 _11282_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03613_ ) );
AOI21_X1 _11283_ ( .A(_03612_ ), .B1(_03613_ ), .B2(_03585_ ), .ZN(_03614_ ) );
XNOR2_X1 _11284_ ( .A(_03614_ ), .B(\IF_ID_pc [6] ), .ZN(_03615_ ) );
INV_X1 _11285_ ( .A(_03615_ ), .ZN(_03616_ ) );
INV_X1 _11286_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03617_ ) );
NOR3_X1 _11287_ ( .A1(_03587_ ), .A2(_03220_ ), .A3(_03617_ ), .ZN(_03618_ ) );
AOI21_X1 _11288_ ( .A(_03618_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .B2(_03304_ ), .ZN(_03619_ ) );
XNOR2_X1 _11289_ ( .A(_03619_ ), .B(_03419_ ), .ZN(_03620_ ) );
INV_X1 _11290_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03621_ ) );
AND3_X1 _11291_ ( .A1(_03209_ ), .A2(_03584_ ), .A3(_03621_ ), .ZN(_03622_ ) );
AOI21_X1 _11292_ ( .A(_03622_ ), .B1(\IF_ID_inst [21] ), .B2(_03304_ ), .ZN(_03623_ ) );
NOR2_X1 _11293_ ( .A1(_03623_ ), .A2(_03430_ ), .ZN(_03624_ ) );
AND2_X1 _11294_ ( .A1(_03620_ ), .A2(_03624_ ), .ZN(_03625_ ) );
AND2_X1 _11295_ ( .A1(_03619_ ), .A2(\IF_ID_pc [2] ), .ZN(_03626_ ) );
NOR2_X1 _11296_ ( .A1(_03625_ ), .A2(_03626_ ), .ZN(_03627_ ) );
AOI21_X1 _11297_ ( .A(_03588_ ), .B1(_03304_ ), .B2(\IF_ID_inst [23] ), .ZN(_03628_ ) );
INV_X1 _11298_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03629_ ) );
NOR3_X1 _11299_ ( .A1(_03587_ ), .A2(_03220_ ), .A3(_03629_ ), .ZN(_03630_ ) );
NOR2_X1 _11300_ ( .A1(_03628_ ), .A2(_03630_ ), .ZN(_03631_ ) );
XNOR2_X1 _11301_ ( .A(_03631_ ), .B(fanout_net_9 ), .ZN(_03632_ ) );
INV_X1 _11302_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03633_ ) );
NAND3_X1 _11303_ ( .A1(_03209_ ), .A2(_03584_ ), .A3(_03633_ ), .ZN(_03634_ ) );
INV_X1 _11304_ ( .A(_03304_ ), .ZN(_03635_ ) );
OAI21_X1 _11305_ ( .A(_03634_ ), .B1(_03635_ ), .B2(_03236_ ), .ZN(_03636_ ) );
XNOR2_X1 _11306_ ( .A(_03636_ ), .B(fanout_net_13 ), .ZN(_03637_ ) );
OR3_X1 _11307_ ( .A1(_03627_ ), .A2(_03632_ ), .A3(_03637_ ), .ZN(_03638_ ) );
OR3_X1 _11308_ ( .A1(_03628_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .A3(_03630_ ), .ZN(_03639_ ) );
NOR2_X1 _11309_ ( .A1(_03637_ ), .A2(_03639_ ), .ZN(_03640_ ) );
AOI21_X1 _11310_ ( .A(_03640_ ), .B1(fanout_net_13 ), .B2(_03636_ ), .ZN(_03641_ ) );
AOI211_X1 _11311_ ( .A(_03611_ ), .B(_03616_ ), .C1(_03638_ ), .C2(_03641_ ), .ZN(_03642_ ) );
NOR2_X1 _11312_ ( .A1(_03609_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03643_ ) );
NAND2_X1 _11313_ ( .A1(_03615_ ), .A2(_03643_ ), .ZN(_03644_ ) );
OAI21_X1 _11314_ ( .A(_03644_ ), .B1(_01875_ ), .B2(_03614_ ), .ZN(_03645_ ) );
OAI21_X1 _11315_ ( .A(_03605_ ), .B1(_03642_ ), .B2(_03645_ ), .ZN(_03646_ ) );
INV_X1 _11316_ ( .A(_03646_ ), .ZN(_03647_ ) );
NOR2_X1 _11317_ ( .A1(_03604_ ), .A2(_02021_ ), .ZN(_03648_ ) );
AND2_X1 _11318_ ( .A1(_03306_ ), .A2(\IF_ID_inst [28] ), .ZN(_03649_ ) );
INV_X1 _11319_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03650_ ) );
AOI21_X1 _11320_ ( .A(_03649_ ), .B1(_03650_ ), .B2(_03585_ ), .ZN(_03651_ ) );
INV_X1 _11321_ ( .A(_03651_ ), .ZN(_03652_ ) );
OAI22_X1 _11322_ ( .A1(_03647_ ), .A2(_03648_ ), .B1(\IF_ID_pc [8] ), .B2(_03652_ ), .ZN(_03653_ ) );
INV_X1 _11323_ ( .A(\IF_ID_pc [8] ), .ZN(_03654_ ) );
NOR2_X1 _11324_ ( .A1(_03651_ ), .A2(_03654_ ), .ZN(_03655_ ) );
INV_X1 _11325_ ( .A(_03655_ ), .ZN(_03656_ ) );
NAND2_X1 _11326_ ( .A1(_03653_ ), .A2(_03656_ ), .ZN(_03657_ ) );
AND2_X1 _11327_ ( .A1(_03305_ ), .A2(\IF_ID_inst [15] ), .ZN(_03658_ ) );
MUX2_X1 _11328_ ( .A(_03530_ ), .B(_03658_ ), .S(_03606_ ), .Z(_03659_ ) );
INV_X1 _11329_ ( .A(\IF_ID_pc [15] ), .ZN(_03660_ ) );
XNOR2_X1 _11330_ ( .A(_03659_ ), .B(_03660_ ), .ZN(_03661_ ) );
AND2_X1 _11331_ ( .A1(_03305_ ), .A2(\IF_ID_inst [16] ), .ZN(_03662_ ) );
INV_X1 _11332_ ( .A(_03662_ ), .ZN(_03663_ ) );
INV_X1 _11333_ ( .A(_03588_ ), .ZN(_03664_ ) );
AOI21_X1 _11334_ ( .A(_03589_ ), .B1(_03663_ ), .B2(_03664_ ), .ZN(_03665_ ) );
XNOR2_X1 _11335_ ( .A(_03665_ ), .B(_02086_ ), .ZN(_03666_ ) );
AND2_X1 _11336_ ( .A1(_03661_ ), .A2(_03666_ ), .ZN(_03667_ ) );
AND2_X1 _11337_ ( .A1(_03305_ ), .A2(\IF_ID_inst [14] ), .ZN(_03668_ ) );
MUX2_X1 _11338_ ( .A(_03530_ ), .B(_03668_ ), .S(_03606_ ), .Z(_03669_ ) );
INV_X1 _11339_ ( .A(\IF_ID_pc [14] ), .ZN(_03670_ ) );
XNOR2_X1 _11340_ ( .A(_03669_ ), .B(_03670_ ), .ZN(_03671_ ) );
INV_X1 _11341_ ( .A(_03589_ ), .ZN(_03672_ ) );
AND2_X1 _11342_ ( .A1(_03305_ ), .A2(\IF_ID_inst [13] ), .ZN(_03673_ ) );
OAI21_X1 _11343_ ( .A(_03672_ ), .B1(_03673_ ), .B2(_03588_ ), .ZN(_03674_ ) );
XNOR2_X1 _11344_ ( .A(_03674_ ), .B(\IF_ID_pc [13] ), .ZN(_03675_ ) );
AND2_X1 _11345_ ( .A1(_03671_ ), .A2(_03675_ ), .ZN(_03676_ ) );
AND2_X1 _11346_ ( .A1(_03667_ ), .A2(_03676_ ), .ZN(_03677_ ) );
INV_X1 _11347_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03678_ ) );
AND3_X1 _11348_ ( .A1(_03209_ ), .A2(_03584_ ), .A3(_03678_ ), .ZN(_03679_ ) );
AOI21_X1 _11349_ ( .A(_03679_ ), .B1(\IF_ID_inst [20] ), .B2(_03305_ ), .ZN(_03680_ ) );
XNOR2_X1 _11350_ ( .A(_03680_ ), .B(\IF_ID_pc [11] ), .ZN(_03681_ ) );
AOI21_X1 _11351_ ( .A(_03585_ ), .B1(_03305_ ), .B2(\IF_ID_inst [12] ), .ZN(_03682_ ) );
NOR3_X1 _11352_ ( .A1(_03682_ ), .A2(_03589_ ), .A3(_02004_ ), .ZN(_03683_ ) );
INV_X1 _11353_ ( .A(_03683_ ), .ZN(_03684_ ) );
OAI21_X1 _11354_ ( .A(_02004_ ), .B1(_03682_ ), .B2(_03591_ ), .ZN(_03685_ ) );
AND3_X1 _11355_ ( .A1(_03681_ ), .A2(_03684_ ), .A3(_03685_ ), .ZN(_03686_ ) );
AND2_X1 _11356_ ( .A1(_03305_ ), .A2(\IF_ID_inst [30] ), .ZN(_03687_ ) );
INV_X1 _11357_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03688_ ) );
AOI21_X1 _11358_ ( .A(_03687_ ), .B1(_03688_ ), .B2(_03585_ ), .ZN(_03689_ ) );
XNOR2_X1 _11359_ ( .A(_03689_ ), .B(\IF_ID_pc [10] ), .ZN(_03690_ ) );
AND2_X1 _11360_ ( .A1(_03306_ ), .A2(\IF_ID_inst [29] ), .ZN(_03691_ ) );
INV_X1 _11361_ ( .A(_03691_ ), .ZN(_03692_ ) );
INV_X1 _11362_ ( .A(\IF_ID_pc [9] ), .ZN(_03693_ ) );
INV_X1 _11363_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03694_ ) );
NAND4_X1 _11364_ ( .A1(_03303_ ), .A2(\IF_ID_inst [31] ), .A3(_03209_ ), .A4(_03694_ ), .ZN(_03695_ ) );
AND3_X1 _11365_ ( .A1(_03692_ ), .A2(_03693_ ), .A3(_03695_ ), .ZN(_03696_ ) );
AOI21_X1 _11366_ ( .A(_03693_ ), .B1(_03692_ ), .B2(_03695_ ), .ZN(_03697_ ) );
NOR2_X1 _11367_ ( .A1(_03696_ ), .A2(_03697_ ), .ZN(_03698_ ) );
AND3_X1 _11368_ ( .A1(_03686_ ), .A2(_03690_ ), .A3(_03698_ ), .ZN(_03699_ ) );
AND3_X1 _11369_ ( .A1(_03657_ ), .A2(_03677_ ), .A3(_03699_ ), .ZN(_03700_ ) );
INV_X1 _11370_ ( .A(\IF_ID_pc [10] ), .ZN(_03701_ ) );
NOR2_X1 _11371_ ( .A1(_03689_ ), .A2(_03701_ ), .ZN(_03702_ ) );
AND2_X1 _11372_ ( .A1(_03689_ ), .A2(_03701_ ), .ZN(_03703_ ) );
INV_X1 _11373_ ( .A(_03703_ ), .ZN(_03704_ ) );
AOI21_X1 _11374_ ( .A(_03702_ ), .B1(_03704_ ), .B2(_03697_ ), .ZN(_03705_ ) );
INV_X1 _11375_ ( .A(_03686_ ), .ZN(_03706_ ) );
OR2_X1 _11376_ ( .A1(_03705_ ), .A2(_03706_ ), .ZN(_03707_ ) );
INV_X1 _11377_ ( .A(\IF_ID_pc [11] ), .ZN(_03708_ ) );
NOR2_X1 _11378_ ( .A1(_03680_ ), .A2(_03708_ ), .ZN(_03709_ ) );
NAND3_X1 _11379_ ( .A1(_03684_ ), .A2(_03685_ ), .A3(_03709_ ), .ZN(_03710_ ) );
NAND3_X1 _11380_ ( .A1(_03707_ ), .A2(_03684_ ), .A3(_03710_ ), .ZN(_03711_ ) );
NAND2_X1 _11381_ ( .A1(_03711_ ), .A2(_03677_ ), .ZN(_03712_ ) );
AND2_X1 _11382_ ( .A1(_03659_ ), .A2(\IF_ID_pc [15] ), .ZN(_03713_ ) );
AND2_X1 _11383_ ( .A1(_03666_ ), .A2(_03713_ ), .ZN(_03714_ ) );
AOI21_X1 _11384_ ( .A(_03714_ ), .B1(\IF_ID_pc [16] ), .B2(_03665_ ), .ZN(_03715_ ) );
INV_X1 _11385_ ( .A(_03667_ ), .ZN(_03716_ ) );
AND2_X1 _11386_ ( .A1(_03669_ ), .A2(\IF_ID_pc [14] ), .ZN(_03717_ ) );
NOR2_X1 _11387_ ( .A1(_03674_ ), .A2(_01886_ ), .ZN(_03718_ ) );
AOI21_X1 _11388_ ( .A(_03717_ ), .B1(_03671_ ), .B2(_03718_ ), .ZN(_03719_ ) );
OAI211_X1 _11389_ ( .A(_03712_ ), .B(_03715_ ), .C1(_03716_ ), .C2(_03719_ ), .ZN(_03720_ ) );
NOR2_X1 _11390_ ( .A1(_03700_ ), .A2(_03720_ ), .ZN(_03721_ ) );
INV_X1 _11391_ ( .A(_03721_ ), .ZN(_03722_ ) );
AND2_X1 _11392_ ( .A1(_03306_ ), .A2(\IF_ID_inst [19] ), .ZN(_03723_ ) );
OAI21_X1 _11393_ ( .A(_03672_ ), .B1(_03723_ ), .B2(_03588_ ), .ZN(_03724_ ) );
XNOR2_X1 _11394_ ( .A(_03724_ ), .B(\IF_ID_pc [19] ), .ZN(_03725_ ) );
XNOR2_X1 _11395_ ( .A(_03592_ ), .B(_02071_ ), .ZN(_03726_ ) );
AND2_X1 _11396_ ( .A1(_03725_ ), .A2(_03726_ ), .ZN(_03727_ ) );
AND2_X1 _11397_ ( .A1(_03306_ ), .A2(\IF_ID_inst [18] ), .ZN(_03728_ ) );
INV_X1 _11398_ ( .A(_03728_ ), .ZN(_03729_ ) );
AOI21_X1 _11399_ ( .A(_03589_ ), .B1(_03729_ ), .B2(_03664_ ), .ZN(_03730_ ) );
XNOR2_X1 _11400_ ( .A(_03730_ ), .B(_01932_ ), .ZN(_03731_ ) );
AND2_X1 _11401_ ( .A1(_03306_ ), .A2(\IF_ID_inst [17] ), .ZN(_03732_ ) );
MUX2_X1 _11402_ ( .A(_03530_ ), .B(_03732_ ), .S(_03606_ ), .Z(_03733_ ) );
XNOR2_X1 _11403_ ( .A(_03733_ ), .B(_01952_ ), .ZN(_03734_ ) );
AND3_X1 _11404_ ( .A1(_03727_ ), .A2(_03731_ ), .A3(_03734_ ), .ZN(_03735_ ) );
AND2_X1 _11405_ ( .A1(_03722_ ), .A2(_03735_ ), .ZN(_03736_ ) );
AND2_X1 _11406_ ( .A1(_03733_ ), .A2(\IF_ID_pc [17] ), .ZN(_03737_ ) );
AOI21_X1 _11407_ ( .A(_03591_ ), .B1(_03729_ ), .B2(_03606_ ), .ZN(_03738_ ) );
AND2_X1 _11408_ ( .A1(_03738_ ), .A2(\IF_ID_pc [18] ), .ZN(_03739_ ) );
OAI221_X1 _11409_ ( .A(_03727_ ), .B1(\IF_ID_pc [18] ), .B2(_03730_ ), .C1(_03737_ ), .C2(_03739_ ), .ZN(_03740_ ) );
NOR2_X1 _11410_ ( .A1(_03724_ ), .A2(_02090_ ), .ZN(_03741_ ) );
AND2_X1 _11411_ ( .A1(_03726_ ), .A2(_03741_ ), .ZN(_03742_ ) );
AOI21_X1 _11412_ ( .A(_03742_ ), .B1(\IF_ID_pc [20] ), .B2(_03592_ ), .ZN(_03743_ ) );
AND2_X1 _11413_ ( .A1(_03740_ ), .A2(_03743_ ), .ZN(_03744_ ) );
INV_X1 _11414_ ( .A(_03744_ ), .ZN(_03745_ ) );
NOR2_X1 _11415_ ( .A1(_03736_ ), .A2(_03745_ ), .ZN(_03746_ ) );
INV_X1 _11416_ ( .A(_03746_ ), .ZN(_03747_ ) );
XNOR2_X1 _11417_ ( .A(_03592_ ), .B(_02028_ ), .ZN(_03748_ ) );
XNOR2_X1 _11418_ ( .A(_03592_ ), .B(_02074_ ), .ZN(_03749_ ) );
AND2_X1 _11419_ ( .A1(_03748_ ), .A2(_03749_ ), .ZN(_03750_ ) );
XNOR2_X1 _11420_ ( .A(_03593_ ), .B(_02031_ ), .ZN(_03751_ ) );
INV_X1 _11421_ ( .A(_03751_ ), .ZN(_03752_ ) );
XNOR2_X1 _11422_ ( .A(_03593_ ), .B(\IF_ID_pc [22] ), .ZN(_03753_ ) );
NOR2_X1 _11423_ ( .A1(_03752_ ), .A2(_03753_ ), .ZN(_03754_ ) );
AND3_X1 _11424_ ( .A1(_03747_ ), .A2(_03750_ ), .A3(_03754_ ), .ZN(_03755_ ) );
AND2_X1 _11425_ ( .A1(_03593_ ), .A2(\IF_ID_pc [22] ), .ZN(_03756_ ) );
AND2_X1 _11426_ ( .A1(_03593_ ), .A2(\IF_ID_pc [21] ), .ZN(_03757_ ) );
OAI21_X1 _11427_ ( .A(_03750_ ), .B1(_03756_ ), .B2(_03757_ ), .ZN(_03758_ ) );
NAND2_X1 _11428_ ( .A1(_03594_ ), .A2(\IF_ID_pc [24] ), .ZN(_03759_ ) );
NAND2_X1 _11429_ ( .A1(_03594_ ), .A2(\IF_ID_pc [23] ), .ZN(_03760_ ) );
NAND3_X1 _11430_ ( .A1(_03758_ ), .A2(_03759_ ), .A3(_03760_ ), .ZN(_03761_ ) );
OAI21_X1 _11431_ ( .A(_03601_ ), .B1(_03755_ ), .B2(_03761_ ), .ZN(_03762_ ) );
OAI21_X1 _11432_ ( .A(_03593_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_03763_ ) );
INV_X1 _11433_ ( .A(_03763_ ), .ZN(_03764_ ) );
AND3_X1 _11434_ ( .A1(_03598_ ), .A2(_03597_ ), .A3(_03764_ ), .ZN(_03765_ ) );
AND2_X1 _11435_ ( .A1(_03594_ ), .A2(\IF_ID_pc [28] ), .ZN(_03766_ ) );
AND2_X1 _11436_ ( .A1(_03594_ ), .A2(\IF_ID_pc [27] ), .ZN(_03767_ ) );
NOR3_X1 _11437_ ( .A1(_03765_ ), .A2(_03766_ ), .A3(_03767_ ), .ZN(_03768_ ) );
AOI21_X1 _11438_ ( .A(_03596_ ), .B1(_03762_ ), .B2(_03768_ ), .ZN(_03769_ ) );
AND2_X1 _11439_ ( .A1(_03594_ ), .A2(\IF_ID_pc [30] ), .ZN(_03770_ ) );
NOR2_X1 _11440_ ( .A1(_03594_ ), .A2(\IF_ID_pc [30] ), .ZN(_03771_ ) );
OR4_X1 _11441_ ( .A1(_03590_ ), .A2(_03769_ ), .A3(_03770_ ), .A4(_03771_ ), .ZN(_03772_ ) );
INV_X1 _11442_ ( .A(_03439_ ), .ZN(_03773_ ) );
BUF_X4 _11443_ ( .A(_03773_ ), .Z(_03774_ ) );
BUF_X4 _11444_ ( .A(_03774_ ), .Z(_03775_ ) );
OAI22_X1 _11445_ ( .A1(_03769_ ), .A2(_03590_ ), .B1(_03770_ ), .B2(_03771_ ), .ZN(_03776_ ) );
NAND3_X1 _11446_ ( .A1(_03772_ ), .A2(_03775_ ), .A3(_03776_ ), .ZN(_03777_ ) );
BUF_X4 _11447_ ( .A(_03581_ ), .Z(_03778_ ) );
BUF_X4 _11448_ ( .A(_03774_ ), .Z(_03779_ ) );
BUF_X4 _11449_ ( .A(_03779_ ), .Z(_03780_ ) );
OAI211_X1 _11450_ ( .A(_03777_ ), .B(_03778_ ), .C1(\myexu.pc_jump [30] ), .C2(_03780_ ), .ZN(_03781_ ) );
NAND2_X1 _11451_ ( .A1(\mtvec [30] ), .A2(\myifu.to_reset ), .ZN(_03782_ ) );
AOI21_X1 _11452_ ( .A(fanout_net_4 ), .B1(_03781_ ), .B2(_03782_ ), .ZN(_00282_ ) );
BUF_X4 _11453_ ( .A(_03581_ ), .Z(_03783_ ) );
INV_X1 _11454_ ( .A(_03410_ ), .ZN(_03784_ ) );
NAND3_X1 _11455_ ( .A1(_03436_ ), .A2(_03415_ ), .A3(_03421_ ), .ZN(_03785_ ) );
OAI211_X1 _11456_ ( .A(check_quest ), .B(_03423_ ), .C1(_03784_ ), .C2(_03785_ ), .ZN(_03786_ ) );
XNOR2_X1 _11457_ ( .A(_03746_ ), .B(_03751_ ), .ZN(_03787_ ) );
BUF_X4 _11458_ ( .A(_03439_ ), .Z(_03788_ ) );
OAI211_X1 _11459_ ( .A(_03783_ ), .B(_03786_ ), .C1(_03787_ ), .C2(_03788_ ), .ZN(_03789_ ) );
NAND2_X1 _11460_ ( .A1(\mtvec [21] ), .A2(\myifu.to_reset ), .ZN(_03790_ ) );
AOI21_X1 _11461_ ( .A(fanout_net_4 ), .B1(_03789_ ), .B2(_03790_ ), .ZN(_00283_ ) );
AND3_X1 _11462_ ( .A1(_03722_ ), .A2(_03731_ ), .A3(_03734_ ), .ZN(_03791_ ) );
AND2_X1 _11463_ ( .A1(_03730_ ), .A2(\IF_ID_pc [18] ), .ZN(_03792_ ) );
AND2_X1 _11464_ ( .A1(_03731_ ), .A2(_03737_ ), .ZN(_03793_ ) );
OR3_X1 _11465_ ( .A1(_03791_ ), .A2(_03792_ ), .A3(_03793_ ), .ZN(_03794_ ) );
AOI21_X1 _11466_ ( .A(_03741_ ), .B1(_03794_ ), .B2(_03725_ ), .ZN(_03795_ ) );
XNOR2_X1 _11467_ ( .A(_03795_ ), .B(_03726_ ), .ZN(_03796_ ) );
MUX2_X1 _11468_ ( .A(\myexu.pc_jump [20] ), .B(_03796_ ), .S(_03774_ ), .Z(_03797_ ) );
MUX2_X1 _11469_ ( .A(\mtvec [20] ), .B(_03797_ ), .S(_03580_ ), .Z(_03798_ ) );
AND2_X1 _11470_ ( .A1(_03798_ ), .A2(_01748_ ), .ZN(_00284_ ) );
INV_X1 _11471_ ( .A(\mtvec [19] ), .ZN(_03799_ ) );
XOR2_X1 _11472_ ( .A(_03794_ ), .B(_03725_ ), .Z(_03800_ ) );
NAND2_X1 _11473_ ( .A1(_03800_ ), .A2(_03779_ ), .ZN(_03801_ ) );
AOI21_X1 _11474_ ( .A(\myifu.to_reset ), .B1(_03439_ ), .B2(\myexu.pc_jump [19] ), .ZN(_03802_ ) );
AOI221_X4 _11475_ ( .A(fanout_net_4 ), .B1(_03799_ ), .B2(\myifu.to_reset ), .C1(_03801_ ), .C2(_03802_ ), .ZN(_00285_ ) );
AOI21_X1 _11476_ ( .A(_03737_ ), .B1(_03722_ ), .B2(_03734_ ), .ZN(_03803_ ) );
XNOR2_X1 _11477_ ( .A(_03803_ ), .B(_03731_ ), .ZN(_03804_ ) );
MUX2_X1 _11478_ ( .A(\myexu.pc_jump [18] ), .B(_03804_ ), .S(_03774_ ), .Z(_03805_ ) );
MUX2_X1 _11479_ ( .A(\mtvec [18] ), .B(_03805_ ), .S(_03580_ ), .Z(_03806_ ) );
AND2_X1 _11480_ ( .A1(_03806_ ), .A2(_01748_ ), .ZN(_00286_ ) );
XOR2_X1 _11481_ ( .A(_03721_ ), .B(_03734_ ), .Z(_03807_ ) );
NAND2_X1 _11482_ ( .A1(_03807_ ), .A2(_03775_ ), .ZN(_03808_ ) );
OAI211_X1 _11483_ ( .A(_03808_ ), .B(_03778_ ), .C1(\myexu.pc_jump [17] ), .C2(_03780_ ), .ZN(_03809_ ) );
NAND2_X1 _11484_ ( .A1(\mtvec [17] ), .A2(\myifu.to_reset ), .ZN(_03810_ ) );
AOI21_X1 _11485_ ( .A(fanout_net_4 ), .B1(_03809_ ), .B2(_03810_ ), .ZN(_00287_ ) );
INV_X1 _11486_ ( .A(_03699_ ), .ZN(_03811_ ) );
AOI21_X1 _11487_ ( .A(_03811_ ), .B1(_03653_ ), .B2(_03656_ ), .ZN(_03812_ ) );
OAI21_X1 _11488_ ( .A(_03676_ ), .B1(_03812_ ), .B2(_03711_ ), .ZN(_03813_ ) );
NAND2_X1 _11489_ ( .A1(_03813_ ), .A2(_03719_ ), .ZN(_03814_ ) );
AOI21_X1 _11490_ ( .A(_03713_ ), .B1(_03814_ ), .B2(_03661_ ), .ZN(_03815_ ) );
XNOR2_X1 _11491_ ( .A(_03815_ ), .B(_03666_ ), .ZN(_03816_ ) );
MUX2_X1 _11492_ ( .A(\myexu.pc_jump [16] ), .B(_03816_ ), .S(_03774_ ), .Z(_03817_ ) );
MUX2_X1 _11493_ ( .A(\mtvec [16] ), .B(_03817_ ), .S(_03580_ ), .Z(_03818_ ) );
AND2_X1 _11494_ ( .A1(_03818_ ), .A2(_01748_ ), .ZN(_00288_ ) );
XNOR2_X1 _11495_ ( .A(_03814_ ), .B(_03661_ ), .ZN(_03819_ ) );
NAND2_X1 _11496_ ( .A1(_03819_ ), .A2(_03775_ ), .ZN(_03820_ ) );
OAI211_X1 _11497_ ( .A(_03820_ ), .B(_03778_ ), .C1(\myexu.pc_jump [15] ), .C2(_03780_ ), .ZN(_03821_ ) );
NAND2_X1 _11498_ ( .A1(\mtvec [15] ), .A2(\myifu.to_reset ), .ZN(_03822_ ) );
AOI21_X1 _11499_ ( .A(fanout_net_4 ), .B1(_03821_ ), .B2(_03822_ ), .ZN(_00289_ ) );
NOR2_X1 _11500_ ( .A1(_03812_ ), .A2(_03711_ ), .ZN(_03823_ ) );
INV_X1 _11501_ ( .A(_03823_ ), .ZN(_03824_ ) );
AOI21_X1 _11502_ ( .A(_03718_ ), .B1(_03824_ ), .B2(_03675_ ), .ZN(_03825_ ) );
XNOR2_X1 _11503_ ( .A(_03825_ ), .B(_03671_ ), .ZN(_03826_ ) );
MUX2_X1 _11504_ ( .A(\myexu.pc_jump [14] ), .B(_03826_ ), .S(_03774_ ), .Z(_03827_ ) );
MUX2_X1 _11505_ ( .A(\mtvec [14] ), .B(_03827_ ), .S(_03580_ ), .Z(_03828_ ) );
AND2_X1 _11506_ ( .A1(_03828_ ), .A2(_01748_ ), .ZN(_00290_ ) );
XOR2_X1 _11507_ ( .A(_03823_ ), .B(_03675_ ), .Z(_03829_ ) );
NAND2_X1 _11508_ ( .A1(_03829_ ), .A2(_03775_ ), .ZN(_03830_ ) );
OAI211_X1 _11509_ ( .A(_03830_ ), .B(_03778_ ), .C1(\myexu.pc_jump [13] ), .C2(_03780_ ), .ZN(_03831_ ) );
NAND2_X1 _11510_ ( .A1(\mtvec [13] ), .A2(\myifu.to_reset ), .ZN(_03832_ ) );
AOI21_X1 _11511_ ( .A(fanout_net_4 ), .B1(_03831_ ), .B2(_03832_ ), .ZN(_00291_ ) );
OR3_X1 _11512_ ( .A1(_03437_ ), .A2(_03438_ ), .A3(\myexu.pc_jump [12] ), .ZN(_03833_ ) );
INV_X1 _11513_ ( .A(_03698_ ), .ZN(_03834_ ) );
AOI21_X1 _11514_ ( .A(_03834_ ), .B1(_03653_ ), .B2(_03656_ ), .ZN(_03835_ ) );
OR3_X1 _11515_ ( .A1(_03835_ ), .A2(_03702_ ), .A3(_03697_ ), .ZN(_03836_ ) );
AND3_X1 _11516_ ( .A1(_03836_ ), .A2(_03681_ ), .A3(_03704_ ), .ZN(_03837_ ) );
NOR2_X1 _11517_ ( .A1(_03837_ ), .A2(_03709_ ), .ZN(_03838_ ) );
AND2_X1 _11518_ ( .A1(_03684_ ), .A2(_03685_ ), .ZN(_03839_ ) );
XNOR2_X1 _11519_ ( .A(_03838_ ), .B(_03839_ ), .ZN(_03840_ ) );
OAI211_X1 _11520_ ( .A(_03783_ ), .B(_03833_ ), .C1(_03840_ ), .C2(_03788_ ), .ZN(_03841_ ) );
NAND2_X1 _11521_ ( .A1(\mtvec [12] ), .A2(\myifu.to_reset ), .ZN(_03842_ ) );
AOI21_X1 _11522_ ( .A(fanout_net_4 ), .B1(_03841_ ), .B2(_03842_ ), .ZN(_00292_ ) );
AND3_X1 _11523_ ( .A1(_03762_ ), .A2(_03768_ ), .A3(_03596_ ), .ZN(_03843_ ) );
OAI21_X1 _11524_ ( .A(_03779_ ), .B1(_03843_ ), .B2(_03769_ ), .ZN(_03844_ ) );
OAI211_X1 _11525_ ( .A(_03844_ ), .B(_03778_ ), .C1(\myexu.pc_jump [29] ), .C2(_03780_ ), .ZN(_03845_ ) );
NAND2_X1 _11526_ ( .A1(\mtvec [29] ), .A2(\myifu.to_reset ), .ZN(_03846_ ) );
AOI21_X1 _11527_ ( .A(fanout_net_4 ), .B1(_03845_ ), .B2(_03846_ ), .ZN(_00293_ ) );
AOI21_X1 _11528_ ( .A(_03681_ ), .B1(_03836_ ), .B2(_03704_ ), .ZN(_03847_ ) );
OAI21_X1 _11529_ ( .A(_03779_ ), .B1(_03837_ ), .B2(_03847_ ), .ZN(_03848_ ) );
OAI211_X1 _11530_ ( .A(_03848_ ), .B(_03778_ ), .C1(\myexu.pc_jump [11] ), .C2(_03780_ ), .ZN(_03849_ ) );
NAND2_X1 _11531_ ( .A1(\mtvec [11] ), .A2(\myifu.to_reset ), .ZN(_03850_ ) );
AOI21_X1 _11532_ ( .A(fanout_net_4 ), .B1(_03849_ ), .B2(_03850_ ), .ZN(_00294_ ) );
NOR2_X1 _11533_ ( .A1(_03835_ ), .A2(_03697_ ), .ZN(_03851_ ) );
INV_X1 _11534_ ( .A(_03851_ ), .ZN(_03852_ ) );
OAI21_X1 _11535_ ( .A(_03774_ ), .B1(_03852_ ), .B2(_03690_ ), .ZN(_03853_ ) );
AOI21_X1 _11536_ ( .A(_03853_ ), .B1(_03852_ ), .B2(_03690_ ), .ZN(_03854_ ) );
AOI211_X1 _11537_ ( .A(\myifu.to_reset ), .B(_03854_ ), .C1(\myexu.pc_jump [10] ), .C2(_03788_ ), .ZN(_03855_ ) );
NOR2_X1 _11538_ ( .A1(_03783_ ), .A2(\mtvec [10] ), .ZN(_03856_ ) );
NOR3_X1 _11539_ ( .A1(_03855_ ), .A2(fanout_net_4 ), .A3(_03856_ ), .ZN(_00295_ ) );
AND3_X1 _11540_ ( .A1(_03653_ ), .A2(_03656_ ), .A3(_03834_ ), .ZN(_03857_ ) );
OAI21_X1 _11541_ ( .A(_03779_ ), .B1(_03857_ ), .B2(_03835_ ), .ZN(_03858_ ) );
OAI211_X1 _11542_ ( .A(_03858_ ), .B(_03778_ ), .C1(\myexu.pc_jump [9] ), .C2(_03780_ ), .ZN(_03859_ ) );
NAND2_X1 _11543_ ( .A1(\mtvec [9] ), .A2(\myifu.to_reset ), .ZN(_03860_ ) );
AOI21_X1 _11544_ ( .A(fanout_net_4 ), .B1(_03859_ ), .B2(_03860_ ), .ZN(_00296_ ) );
NOR2_X1 _11545_ ( .A1(_03647_ ), .A2(_03648_ ), .ZN(_03861_ ) );
INV_X1 _11546_ ( .A(_03861_ ), .ZN(_03862_ ) );
XNOR2_X1 _11547_ ( .A(_03651_ ), .B(\IF_ID_pc [8] ), .ZN(_03863_ ) );
OAI21_X1 _11548_ ( .A(_03774_ ), .B1(_03862_ ), .B2(_03863_ ), .ZN(_03864_ ) );
AOI21_X1 _11549_ ( .A(_03864_ ), .B1(_03862_ ), .B2(_03863_ ), .ZN(_03865_ ) );
AOI211_X1 _11550_ ( .A(\myifu.to_reset ), .B(_03865_ ), .C1(\myexu.pc_jump [8] ), .C2(_03788_ ), .ZN(_03866_ ) );
NOR2_X1 _11551_ ( .A1(_03783_ ), .A2(\mtvec [8] ), .ZN(_03867_ ) );
NOR3_X1 _11552_ ( .A1(_03866_ ), .A2(fanout_net_4 ), .A3(_03867_ ), .ZN(_00297_ ) );
NOR3_X1 _11553_ ( .A1(_03642_ ), .A2(_03605_ ), .A3(_03645_ ), .ZN(_03868_ ) );
OAI21_X1 _11554_ ( .A(_03779_ ), .B1(_03647_ ), .B2(_03868_ ), .ZN(_03869_ ) );
OAI211_X1 _11555_ ( .A(_03869_ ), .B(_03778_ ), .C1(\myexu.pc_jump [7] ), .C2(_03780_ ), .ZN(_03870_ ) );
NAND2_X1 _11556_ ( .A1(\mtvec [7] ), .A2(\myifu.to_reset ), .ZN(_03871_ ) );
AOI21_X1 _11557_ ( .A(fanout_net_4 ), .B1(_03870_ ), .B2(_03871_ ), .ZN(_00298_ ) );
AOI21_X1 _11558_ ( .A(_03611_ ), .B1(_03638_ ), .B2(_03641_ ), .ZN(_03872_ ) );
OR3_X1 _11559_ ( .A1(_03872_ ), .A2(_03643_ ), .A3(_03616_ ), .ZN(_03873_ ) );
OAI21_X1 _11560_ ( .A(_03616_ ), .B1(_03872_ ), .B2(_03643_ ), .ZN(_03874_ ) );
AOI21_X1 _11561_ ( .A(_03439_ ), .B1(_03873_ ), .B2(_03874_ ), .ZN(_03875_ ) );
AOI211_X1 _11562_ ( .A(\myifu.to_reset ), .B(_03875_ ), .C1(\myexu.pc_jump [6] ), .C2(_03788_ ), .ZN(_03876_ ) );
NOR2_X1 _11563_ ( .A1(_03783_ ), .A2(\mtvec [6] ), .ZN(_03877_ ) );
NOR3_X1 _11564_ ( .A1(_03876_ ), .A2(fanout_net_4 ), .A3(_03877_ ), .ZN(_00299_ ) );
AND3_X1 _11565_ ( .A1(_03638_ ), .A2(_03641_ ), .A3(_03611_ ), .ZN(_03878_ ) );
OAI21_X1 _11566_ ( .A(_03779_ ), .B1(_03878_ ), .B2(_03872_ ), .ZN(_03879_ ) );
OAI211_X1 _11567_ ( .A(_03879_ ), .B(_03778_ ), .C1(\myexu.pc_jump [5] ), .C2(_03775_ ), .ZN(_03880_ ) );
NAND2_X1 _11568_ ( .A1(\mtvec [5] ), .A2(\myifu.to_reset ), .ZN(_03881_ ) );
AOI21_X1 _11569_ ( .A(fanout_net_4 ), .B1(_03880_ ), .B2(_03881_ ), .ZN(_00300_ ) );
AND2_X1 _11570_ ( .A1(\mtvec [4] ), .A2(\myifu.to_reset ), .ZN(_03882_ ) );
OR2_X1 _11571_ ( .A1(_03627_ ), .A2(_03632_ ), .ZN(_03883_ ) );
NAND2_X1 _11572_ ( .A1(_03883_ ), .A2(_03639_ ), .ZN(_03884_ ) );
XNOR2_X1 _11573_ ( .A(_03884_ ), .B(_03637_ ), .ZN(_03885_ ) );
MUX2_X1 _11574_ ( .A(\myexu.pc_jump [4] ), .B(_03885_ ), .S(_03774_ ), .Z(_03886_ ) );
AOI21_X1 _11575_ ( .A(_03882_ ), .B1(_03886_ ), .B2(_03581_ ), .ZN(_03887_ ) );
NOR2_X1 _11576_ ( .A1(_03887_ ), .A2(fanout_net_4 ), .ZN(_00301_ ) );
XOR2_X1 _11577_ ( .A(_03627_ ), .B(_03632_ ), .Z(_03888_ ) );
MUX2_X1 _11578_ ( .A(\myexu.pc_jump [3] ), .B(_03888_ ), .S(_03773_ ), .Z(_03889_ ) );
AND2_X1 _11579_ ( .A1(_03889_ ), .A2(_03580_ ), .ZN(_03890_ ) );
AOI21_X1 _11580_ ( .A(_03890_ ), .B1(\mtvec [3] ), .B2(\myifu.to_reset ), .ZN(_03891_ ) );
NOR2_X1 _11581_ ( .A1(_03891_ ), .A2(reset ), .ZN(_00302_ ) );
AND2_X1 _11582_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
OAI21_X1 _11583_ ( .A(_01586_ ), .B1(\myifu.pc_$_SDFFE_PP1P__Q_E ), .B2(fanout_net_13 ), .ZN(_03892_ ) );
AOI21_X1 _11584_ ( .A(_03892_ ), .B1(_03887_ ), .B2(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_00303_ ) );
NOR2_X1 _11585_ ( .A1(_03581_ ), .A2(\mtvec [2] ), .ZN(_03893_ ) );
XNOR2_X1 _11586_ ( .A(_03620_ ), .B(_03624_ ), .ZN(_03894_ ) );
MUX2_X1 _11587_ ( .A(_03894_ ), .B(_03433_ ), .S(_03439_ ), .Z(_03895_ ) );
AOI211_X1 _11588_ ( .A(reset ), .B(_03893_ ), .C1(_03895_ ), .C2(_03783_ ), .ZN(_00304_ ) );
OAI21_X1 _11589_ ( .A(_01586_ ), .B1(\myifu.pc_$_SDFFE_PP1P__Q_E ), .B2(fanout_net_9 ), .ZN(_03896_ ) );
AOI21_X1 _11590_ ( .A(_03896_ ), .B1(_03891_ ), .B2(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_00305_ ) );
NOR2_X1 _11591_ ( .A1(_03755_ ), .A2(_03761_ ), .ZN(_03897_ ) );
INV_X1 _11592_ ( .A(_03599_ ), .ZN(_03898_ ) );
INV_X1 _11593_ ( .A(_03600_ ), .ZN(_03899_ ) );
NOR3_X1 _11594_ ( .A1(_03897_ ), .A2(_03898_ ), .A3(_03899_ ), .ZN(_03900_ ) );
OAI21_X1 _11595_ ( .A(_03598_ ), .B1(_03900_ ), .B2(_03764_ ), .ZN(_03901_ ) );
INV_X1 _11596_ ( .A(_03767_ ), .ZN(_03902_ ) );
AND3_X1 _11597_ ( .A1(_03901_ ), .A2(_03597_ ), .A3(_03902_ ), .ZN(_03903_ ) );
AOI21_X1 _11598_ ( .A(_03597_ ), .B1(_03901_ ), .B2(_03902_ ), .ZN(_03904_ ) );
OR3_X1 _11599_ ( .A1(_03903_ ), .A2(_03904_ ), .A3(_03439_ ), .ZN(_03905_ ) );
OAI211_X1 _11600_ ( .A(_03905_ ), .B(_03778_ ), .C1(\myexu.pc_jump [28] ), .C2(_03775_ ), .ZN(_03906_ ) );
NAND2_X1 _11601_ ( .A1(\mtvec [28] ), .A2(\myifu.to_reset ), .ZN(_03907_ ) );
AOI21_X1 _11602_ ( .A(reset ), .B1(_03906_ ), .B2(_03907_ ), .ZN(_00306_ ) );
NOR2_X1 _11603_ ( .A1(_03581_ ), .A2(\mtvec [1] ), .ZN(_03908_ ) );
XNOR2_X1 _11604_ ( .A(_03623_ ), .B(_03430_ ), .ZN(_03909_ ) );
MUX2_X1 _11605_ ( .A(_03909_ ), .B(_03432_ ), .S(_03439_ ), .Z(_03910_ ) );
AOI211_X1 _11606_ ( .A(reset ), .B(_03908_ ), .C1(_03910_ ), .C2(_03783_ ), .ZN(_00307_ ) );
NOR2_X1 _11607_ ( .A1(_03900_ ), .A2(_03764_ ), .ZN(_03911_ ) );
XOR2_X1 _11608_ ( .A(_03911_ ), .B(_03598_ ), .Z(_03912_ ) );
NAND2_X1 _11609_ ( .A1(_03912_ ), .A2(_03775_ ), .ZN(_03913_ ) );
OAI211_X1 _11610_ ( .A(_03913_ ), .B(_03581_ ), .C1(\myexu.pc_jump [27] ), .C2(_03775_ ), .ZN(_03914_ ) );
NAND2_X1 _11611_ ( .A1(\mtvec [27] ), .A2(\myifu.to_reset ), .ZN(_03915_ ) );
AOI21_X1 _11612_ ( .A(reset ), .B1(_03914_ ), .B2(_03915_ ), .ZN(_00308_ ) );
NOR2_X1 _11613_ ( .A1(_03897_ ), .A2(_03899_ ), .ZN(_03916_ ) );
AND2_X1 _11614_ ( .A1(_03594_ ), .A2(\IF_ID_pc [25] ), .ZN(_03917_ ) );
OR3_X1 _11615_ ( .A1(_03916_ ), .A2(_03917_ ), .A3(_03898_ ), .ZN(_03918_ ) );
OAI21_X1 _11616_ ( .A(_03898_ ), .B1(_03916_ ), .B2(_03917_ ), .ZN(_03919_ ) );
NAND3_X1 _11617_ ( .A1(_03918_ ), .A2(_03779_ ), .A3(_03919_ ), .ZN(_03920_ ) );
OAI211_X1 _11618_ ( .A(_03920_ ), .B(_03581_ ), .C1(\myexu.pc_jump [26] ), .C2(_03775_ ), .ZN(_03921_ ) );
NAND2_X1 _11619_ ( .A1(\mtvec [26] ), .A2(\myifu.to_reset ), .ZN(_03922_ ) );
AOI21_X1 _11620_ ( .A(reset ), .B1(_03921_ ), .B2(_03922_ ), .ZN(_00309_ ) );
AND4_X1 _11621_ ( .A1(_03750_ ), .A2(_03722_ ), .A3(_03754_ ), .A4(_03735_ ), .ZN(_03923_ ) );
AND3_X1 _11622_ ( .A1(_03745_ ), .A2(_03750_ ), .A3(_03754_ ), .ZN(_03924_ ) );
NOR4_X1 _11623_ ( .A1(_03923_ ), .A2(_03761_ ), .A3(_03924_ ), .A4(_03600_ ), .ZN(_03925_ ) );
OAI21_X1 _11624_ ( .A(_03779_ ), .B1(_03916_ ), .B2(_03925_ ), .ZN(_03926_ ) );
OAI211_X1 _11625_ ( .A(_03926_ ), .B(_03581_ ), .C1(\myexu.pc_jump [25] ), .C2(_03775_ ), .ZN(_03927_ ) );
NAND2_X1 _11626_ ( .A1(\mtvec [25] ), .A2(\myifu.to_reset ), .ZN(_03928_ ) );
AOI21_X1 _11627_ ( .A(reset ), .B1(_03927_ ), .B2(_03928_ ), .ZN(_00310_ ) );
OAI21_X1 _11628_ ( .A(_03754_ ), .B1(_03736_ ), .B2(_03745_ ), .ZN(_03929_ ) );
OAI21_X1 _11629_ ( .A(_03594_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_03930_ ) );
NAND2_X1 _11630_ ( .A1(_03929_ ), .A2(_03930_ ), .ZN(_03931_ ) );
NAND2_X1 _11631_ ( .A1(_03931_ ), .A2(_03749_ ), .ZN(_03932_ ) );
AND2_X1 _11632_ ( .A1(_03932_ ), .A2(_03760_ ), .ZN(_03933_ ) );
XNOR2_X1 _11633_ ( .A(_03933_ ), .B(_03748_ ), .ZN(_03934_ ) );
AND2_X1 _11634_ ( .A1(_03934_ ), .A2(_03774_ ), .ZN(_03935_ ) );
AOI211_X1 _11635_ ( .A(\myifu.to_reset ), .B(_03935_ ), .C1(\myexu.pc_jump [24] ), .C2(_03788_ ), .ZN(_03936_ ) );
NOR2_X1 _11636_ ( .A1(_03783_ ), .A2(\mtvec [24] ), .ZN(_03937_ ) );
NOR3_X1 _11637_ ( .A1(_03936_ ), .A2(reset ), .A3(_03937_ ), .ZN(_00311_ ) );
OR3_X1 _11638_ ( .A1(_03437_ ), .A2(_03438_ ), .A3(\myexu.pc_jump [23] ), .ZN(_03938_ ) );
XOR2_X1 _11639_ ( .A(_03931_ ), .B(_03749_ ), .Z(_03939_ ) );
OAI211_X1 _11640_ ( .A(_03783_ ), .B(_03938_ ), .C1(_03939_ ), .C2(_03788_ ), .ZN(_03940_ ) );
NAND2_X1 _11641_ ( .A1(\mtvec [23] ), .A2(\myifu.to_reset ), .ZN(_03941_ ) );
AOI21_X1 _11642_ ( .A(reset ), .B1(_03940_ ), .B2(_03941_ ), .ZN(_00312_ ) );
INV_X1 _11643_ ( .A(_03736_ ), .ZN(_03942_ ) );
AOI21_X1 _11644_ ( .A(_03752_ ), .B1(_03942_ ), .B2(_03744_ ), .ZN(_03943_ ) );
OR3_X1 _11645_ ( .A1(_03943_ ), .A2(_03757_ ), .A3(_03753_ ), .ZN(_03944_ ) );
OAI21_X1 _11646_ ( .A(_03753_ ), .B1(_03943_ ), .B2(_03757_ ), .ZN(_03945_ ) );
AOI21_X1 _11647_ ( .A(_03439_ ), .B1(_03944_ ), .B2(_03945_ ), .ZN(_03946_ ) );
AOI211_X1 _11648_ ( .A(\myifu.to_reset ), .B(_03946_ ), .C1(\myexu.pc_jump [22] ), .C2(_03788_ ), .ZN(_03947_ ) );
NOR2_X1 _11649_ ( .A1(_03783_ ), .A2(\mtvec [22] ), .ZN(_03948_ ) );
NOR3_X1 _11650_ ( .A1(_03947_ ), .A2(reset ), .A3(_03948_ ), .ZN(_00313_ ) );
NAND2_X1 _11651_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_03949_ ) );
NOR3_X1 _11652_ ( .A1(_03769_ ), .A2(_03590_ ), .A3(_03770_ ), .ZN(_03950_ ) );
NOR2_X1 _11653_ ( .A1(_03950_ ), .A2(_03771_ ), .ZN(_03951_ ) );
XNOR2_X1 _11654_ ( .A(_03594_ ), .B(\IF_ID_pc [31] ), .ZN(_03952_ ) );
OAI21_X1 _11655_ ( .A(_03779_ ), .B1(_03951_ ), .B2(_03952_ ), .ZN(_03953_ ) );
AOI21_X1 _11656_ ( .A(_03953_ ), .B1(_03951_ ), .B2(_03952_ ), .ZN(_03954_ ) );
OAI21_X1 _11657_ ( .A(_03581_ ), .B1(_03780_ ), .B2(\myexu.pc_jump [31] ), .ZN(_03955_ ) );
OAI211_X1 _11658_ ( .A(_01748_ ), .B(_03949_ ), .C1(_03954_ ), .C2(_03955_ ), .ZN(_00314_ ) );
INV_X1 _11659_ ( .A(\myifu.tmp_offset [2] ), .ZN(_03956_ ) );
AND3_X1 _11660_ ( .A1(_02170_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .A3(_02173_ ), .ZN(_03957_ ) );
NOR2_X1 _11661_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_03958_ ) );
NAND2_X1 _11662_ ( .A1(_03958_ ), .A2(io_master_rvalid ), .ZN(_03959_ ) );
AOI21_X1 _11663_ ( .A(_03957_ ), .B1(_02175_ ), .B2(_03959_ ), .ZN(_03960_ ) );
INV_X1 _11664_ ( .A(\io_master_rid [3] ), .ZN(_03961_ ) );
INV_X1 _11665_ ( .A(\io_master_rid [2] ), .ZN(_03962_ ) );
INV_X1 _11666_ ( .A(\io_master_rid [1] ), .ZN(_03963_ ) );
NAND4_X1 _11667_ ( .A1(_03961_ ), .A2(_03962_ ), .A3(_03963_ ), .A4(\io_master_rid [0] ), .ZN(_03964_ ) );
AOI21_X1 _11668_ ( .A(_02087_ ), .B1(_02175_ ), .B2(_03964_ ), .ZN(_03965_ ) );
AND2_X1 _11669_ ( .A1(_03960_ ), .A2(_03965_ ), .ZN(_03966_ ) );
INV_X1 _11670_ ( .A(_03966_ ), .ZN(_03967_ ) );
NOR2_X1 _11671_ ( .A1(_02174_ ), .A2(io_master_rlast ), .ZN(_03968_ ) );
OAI211_X1 _11672_ ( .A(_01679_ ), .B(_03956_ ), .C1(_03967_ ), .C2(_03968_ ), .ZN(_03969_ ) );
INV_X1 _11673_ ( .A(_03969_ ), .ZN(_00315_ ) );
NOR3_X1 _11674_ ( .A1(reset ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00316_ ) );
AND3_X1 _11675_ ( .A1(_02221_ ), .A2(_03440_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_03970_ ) );
INV_X1 _11676_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_03971_ ) );
MUX2_X1 _11677_ ( .A(_02221_ ), .B(_03971_ ), .S(\myifu.to_reset ), .Z(_03972_ ) );
AOI211_X1 _11678_ ( .A(reset ), .B(_03970_ ), .C1(_03972_ ), .C2(\myifu.state [1] ), .ZN(_00317_ ) );
NOR2_X1 _11679_ ( .A1(_02159_ ), .A2(_02151_ ), .ZN(_03973_ ) );
INV_X1 _11680_ ( .A(_03973_ ), .ZN(_03974_ ) );
BUF_X2 _11681_ ( .A(_03974_ ), .Z(_03975_ ) );
BUF_X4 _11682_ ( .A(_02233_ ), .Z(_03976_ ) );
MUX2_X1 _11683_ ( .A(\LS_WB_waddr_csreg [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_03976_ ), .Z(_03977_ ) );
BUF_X4 _11684_ ( .A(_02056_ ), .Z(_03978_ ) );
NOR2_X1 _11685_ ( .A1(_03978_ ), .A2(\EX_LS_flag [1] ), .ZN(_03979_ ) );
OR2_X1 _11686_ ( .A1(_03979_ ), .A2(_02130_ ), .ZN(_03980_ ) );
NOR2_X1 _11687_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_03981_ ) );
AND2_X2 _11688_ ( .A1(_03981_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_03982_ ) );
NOR2_X2 _11689_ ( .A1(_03980_ ), .A2(_03982_ ), .ZN(_03983_ ) );
BUF_X4 _11690_ ( .A(_03983_ ), .Z(_03984_ ) );
BUF_X2 _11691_ ( .A(_03984_ ), .Z(_03985_ ) );
AND3_X1 _11692_ ( .A1(_03975_ ), .A2(_03977_ ), .A3(_03985_ ), .ZN(_00320_ ) );
NOR2_X1 _11693_ ( .A1(_03973_ ), .A2(_03982_ ), .ZN(_03986_ ) );
INV_X1 _11694_ ( .A(_03986_ ), .ZN(_03987_ ) );
BUF_X4 _11695_ ( .A(_02149_ ), .Z(_03988_ ) );
NAND3_X1 _11696_ ( .A1(_03988_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_03989_ ) );
BUF_X4 _11697_ ( .A(_03978_ ), .Z(_03990_ ) );
NAND2_X1 _11698_ ( .A1(_03990_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03991_ ) );
AOI211_X1 _11699_ ( .A(_02134_ ), .B(_03987_ ), .C1(_03989_ ), .C2(_03991_ ), .ZN(_00321_ ) );
NAND3_X1 _11700_ ( .A1(_03988_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_03992_ ) );
NAND2_X1 _11701_ ( .A1(_03990_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_03993_ ) );
AOI211_X1 _11702_ ( .A(_02134_ ), .B(_03987_ ), .C1(_03992_ ), .C2(_03993_ ), .ZN(_00322_ ) );
NAND3_X1 _11703_ ( .A1(_03988_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_03994_ ) );
NAND2_X1 _11704_ ( .A1(_03990_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_03995_ ) );
AOI211_X1 _11705_ ( .A(_02134_ ), .B(_03987_ ), .C1(_03994_ ), .C2(_03995_ ), .ZN(_00323_ ) );
NAND3_X1 _11706_ ( .A1(_03988_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_03996_ ) );
NAND2_X1 _11707_ ( .A1(_03990_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03997_ ) );
AOI211_X1 _11708_ ( .A(_02134_ ), .B(_03987_ ), .C1(_03996_ ), .C2(_03997_ ), .ZN(_00324_ ) );
NAND3_X1 _11709_ ( .A1(_03988_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_03998_ ) );
NAND2_X1 _11710_ ( .A1(_03990_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_03999_ ) );
AOI211_X1 _11711_ ( .A(_02134_ ), .B(_03987_ ), .C1(_03998_ ), .C2(_03999_ ), .ZN(_00325_ ) );
NAND3_X1 _11712_ ( .A1(_03988_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_04000_ ) );
NAND2_X1 _11713_ ( .A1(_03990_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_04001_ ) );
AOI211_X1 _11714_ ( .A(_02134_ ), .B(_03987_ ), .C1(_04000_ ), .C2(_04001_ ), .ZN(_00326_ ) );
NAND3_X1 _11715_ ( .A1(_03988_ ), .A2(fanout_net_6 ), .A3(\EX_LS_flag [2] ), .ZN(_04002_ ) );
NAND2_X1 _11716_ ( .A1(_03990_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_04003_ ) );
AOI211_X1 _11717_ ( .A(_02134_ ), .B(_03987_ ), .C1(_04002_ ), .C2(_04003_ ), .ZN(_00327_ ) );
NOR4_X1 _11718_ ( .A1(_03990_ ), .A2(_02148_ ), .A3(\EX_LS_dest_csreg_mem [9] ), .A4(\EX_LS_flag [0] ), .ZN(_04004_ ) );
NOR2_X1 _11719_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_04005_ ) );
OAI211_X1 _11720_ ( .A(_03986_ ), .B(_02132_ ), .C1(_04004_ ), .C2(_04005_ ), .ZN(_00328_ ) );
NOR4_X1 _11721_ ( .A1(_03990_ ), .A2(_02148_ ), .A3(\EX_LS_dest_csreg_mem [8] ), .A4(\EX_LS_flag [0] ), .ZN(_04006_ ) );
NOR2_X1 _11722_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_04007_ ) );
OAI211_X1 _11723_ ( .A(_03986_ ), .B(_02132_ ), .C1(_04006_ ), .C2(_04007_ ), .ZN(_00329_ ) );
NOR4_X1 _11724_ ( .A1(_03990_ ), .A2(_02148_ ), .A3(\EX_LS_dest_csreg_mem [6] ), .A4(\EX_LS_flag [0] ), .ZN(_04008_ ) );
NOR2_X1 _11725_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_04009_ ) );
OAI211_X1 _11726_ ( .A(_03986_ ), .B(_02132_ ), .C1(_04008_ ), .C2(_04009_ ), .ZN(_00330_ ) );
BUF_X4 _11727_ ( .A(_03978_ ), .Z(_04010_ ) );
NOR4_X1 _11728_ ( .A1(_04010_ ), .A2(_02148_ ), .A3(fanout_net_5 ), .A4(\EX_LS_flag [0] ), .ZN(_04011_ ) );
NOR2_X1 _11729_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_04012_ ) );
OAI211_X1 _11730_ ( .A(_03986_ ), .B(_02132_ ), .C1(_04011_ ), .C2(_04012_ ), .ZN(_00331_ ) );
INV_X1 _11731_ ( .A(\mysc.state [2] ), .ZN(_04013_ ) );
NOR2_X1 _11732_ ( .A1(_04013_ ), .A2(reset ), .ZN(_00339_ ) );
INV_X1 _11733_ ( .A(IDU_valid_EXU ), .ZN(_04014_ ) );
NOR2_X1 _11734_ ( .A1(_04014_ ), .A2(EXU_valid_LSU ), .ZN(\myexu.state_$_ANDNOT__B_Y ) );
INV_X1 _11735_ ( .A(\ID_EX_typ [6] ), .ZN(_04015_ ) );
NAND2_X1 _11736_ ( .A1(_04015_ ), .A2(\ID_EX_typ [7] ), .ZN(_04016_ ) );
INV_X1 _11737_ ( .A(\ID_EX_typ [5] ), .ZN(_04017_ ) );
NOR2_X1 _11738_ ( .A1(_04016_ ), .A2(_04017_ ), .ZN(_04018_ ) );
INV_X1 _11739_ ( .A(fanout_net_7 ), .ZN(_04019_ ) );
AND2_X2 _11740_ ( .A1(_04018_ ), .A2(_04019_ ), .ZN(_04020_ ) );
NOR3_X1 _11741_ ( .A1(_04016_ ), .A2(\ID_EX_typ [5] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04021_ ) );
OAI21_X1 _11742_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .B1(_04020_ ), .B2(_04021_ ), .ZN(_04022_ ) );
INV_X1 _11743_ ( .A(\myec.state [1] ), .ZN(_04023_ ) );
NAND2_X1 _11744_ ( .A1(_04023_ ), .A2(\myec.state [0] ), .ZN(_04024_ ) );
AND2_X1 _11745_ ( .A1(_04024_ ), .A2(_03221_ ), .ZN(_04025_ ) );
BUF_X2 _11746_ ( .A(_04025_ ), .Z(_04026_ ) );
INV_X1 _11747_ ( .A(\myexu.state_$_ANDNOT__B_Y ), .ZN(_04027_ ) );
OAI22_X1 _11748_ ( .A1(_04027_ ), .A2(_04016_ ), .B1(_03438_ ), .B2(check_assert ), .ZN(_04028_ ) );
AND3_X1 _11749_ ( .A1(_04022_ ), .A2(_04026_ ), .A3(_04028_ ), .ZN(_00132_ ) );
CLKBUF_X2 _11750_ ( .A(_04024_ ), .Z(_04029_ ) );
CLKBUF_X2 _11751_ ( .A(_04029_ ), .Z(_04030_ ) );
AND3_X1 _11752_ ( .A1(_04030_ ), .A2(\ID_EX_rd [4] ), .A3(_03239_ ), .ZN(_00153_ ) );
AND3_X1 _11753_ ( .A1(_04030_ ), .A2(\ID_EX_rd [3] ), .A3(_03239_ ), .ZN(_00154_ ) );
AND3_X1 _11754_ ( .A1(_04030_ ), .A2(\ID_EX_rd [2] ), .A3(_03239_ ), .ZN(_00155_ ) );
AND3_X1 _11755_ ( .A1(_04030_ ), .A2(\ID_EX_rd [1] ), .A3(_03239_ ), .ZN(_00156_ ) );
AND3_X1 _11756_ ( .A1(_04030_ ), .A2(\ID_EX_rd [0] ), .A3(_03239_ ), .ZN(_00157_ ) );
INV_X2 _11757_ ( .A(_04025_ ), .ZN(_04031_ ) );
BUF_X4 _11758_ ( .A(_04031_ ), .Z(_04032_ ) );
XNOR2_X1 _11759_ ( .A(\EX_LS_dest_csreg_mem [8] ), .B(\ID_EX_csr [8] ), .ZN(_04033_ ) );
INV_X1 _11760_ ( .A(\ID_EX_csr [4] ), .ZN(_04034_ ) );
NAND2_X1 _11761_ ( .A1(_04034_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .ZN(_04035_ ) );
INV_X1 _11762_ ( .A(fanout_net_6 ), .ZN(_04036_ ) );
NAND2_X1 _11763_ ( .A1(_04036_ ), .A2(\ID_EX_csr [1] ), .ZN(_04037_ ) );
INV_X1 _11764_ ( .A(\EX_LS_dest_csreg_mem [4] ), .ZN(_04038_ ) );
NAND2_X1 _11765_ ( .A1(_04038_ ), .A2(\ID_EX_csr [4] ), .ZN(_04039_ ) );
INV_X1 _11766_ ( .A(\ID_EX_csr [3] ), .ZN(_04040_ ) );
NAND2_X1 _11767_ ( .A1(_04040_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .ZN(_04041_ ) );
AND4_X1 _11768_ ( .A1(_04035_ ), .A2(_04037_ ), .A3(_04039_ ), .A4(_04041_ ), .ZN(_04042_ ) );
INV_X1 _11769_ ( .A(fanout_net_5 ), .ZN(_04043_ ) );
INV_X1 _11770_ ( .A(\ID_EX_csr [5] ), .ZN(_04044_ ) );
AOI22_X1 _11771_ ( .A1(_04043_ ), .A2(\ID_EX_csr [0] ), .B1(_04044_ ), .B2(\EX_LS_dest_csreg_mem [5] ), .ZN(_04045_ ) );
OR2_X1 _11772_ ( .A1(_04044_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .ZN(_04046_ ) );
INV_X1 _11773_ ( .A(\ID_EX_csr [1] ), .ZN(_04047_ ) );
NAND2_X1 _11774_ ( .A1(_04047_ ), .A2(fanout_net_6 ), .ZN(_04048_ ) );
AND4_X1 _11775_ ( .A1(_04042_ ), .A2(_04045_ ), .A3(_04046_ ), .A4(_04048_ ), .ZN(_04049_ ) );
INV_X1 _11776_ ( .A(\ID_EX_csr [9] ), .ZN(_04050_ ) );
NAND2_X1 _11777_ ( .A1(_04050_ ), .A2(\EX_LS_dest_csreg_mem [9] ), .ZN(_04051_ ) );
INV_X1 _11778_ ( .A(\EX_LS_dest_csreg_mem [3] ), .ZN(_04052_ ) );
NAND2_X1 _11779_ ( .A1(_04052_ ), .A2(\ID_EX_csr [3] ), .ZN(_04053_ ) );
AND4_X2 _11780_ ( .A1(_04033_ ), .A2(_04049_ ), .A3(_04051_ ), .A4(_04053_ ), .ZN(_04054_ ) );
INV_X1 _11781_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_04055_ ) );
INV_X1 _11782_ ( .A(\EX_LS_dest_csreg_mem [7] ), .ZN(_04056_ ) );
AOI22_X1 _11783_ ( .A1(_04055_ ), .A2(\ID_EX_csr [9] ), .B1(_04056_ ), .B2(\ID_EX_csr [7] ), .ZN(_04057_ ) );
XNOR2_X1 _11784_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_04058_ ) );
INV_X1 _11785_ ( .A(\ID_EX_csr [0] ), .ZN(_04059_ ) );
INV_X1 _11786_ ( .A(\ID_EX_csr [7] ), .ZN(_04060_ ) );
AOI22_X1 _11787_ ( .A1(fanout_net_5 ), .A2(_04059_ ), .B1(_04060_ ), .B2(\EX_LS_dest_csreg_mem [7] ), .ZN(_04061_ ) );
NAND4_X1 _11788_ ( .A1(_02233_ ), .A2(_04057_ ), .A3(_04058_ ), .A4(_04061_ ), .ZN(_04062_ ) );
XOR2_X1 _11789_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .Z(_04063_ ) );
XOR2_X1 _11790_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .Z(_04064_ ) );
XOR2_X1 _11791_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .Z(_04065_ ) );
NOR4_X1 _11792_ ( .A1(_04062_ ), .A2(_04063_ ), .A3(_04064_ ), .A4(_04065_ ), .ZN(_04066_ ) );
AND3_X1 _11793_ ( .A1(_04054_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_04066_ ), .ZN(_04067_ ) );
AND2_X1 _11794_ ( .A1(_04054_ ), .A2(_04066_ ), .ZN(_04068_ ) );
INV_X1 _11795_ ( .A(_04068_ ), .ZN(_04069_ ) );
INV_X1 _11796_ ( .A(\ID_EX_csr [11] ), .ZN(_04070_ ) );
NAND3_X1 _11797_ ( .A1(_04070_ ), .A2(\ID_EX_csr [9] ), .A3(\ID_EX_csr [8] ), .ZN(_04071_ ) );
NOR2_X1 _11798_ ( .A1(_04071_ ), .A2(\ID_EX_csr [10] ), .ZN(_04072_ ) );
INV_X1 _11799_ ( .A(\ID_EX_csr [6] ), .ZN(_04073_ ) );
NOR3_X1 _11800_ ( .A1(_04073_ ), .A2(\ID_EX_csr [5] ), .A3(\ID_EX_csr [4] ), .ZN(_04074_ ) );
AND3_X1 _11801_ ( .A1(_04072_ ), .A2(_04060_ ), .A3(_04074_ ), .ZN(_04075_ ) );
BUF_X4 _11802_ ( .A(_04075_ ), .Z(_04076_ ) );
BUF_X4 _11803_ ( .A(_04076_ ), .Z(_04077_ ) );
INV_X1 _11804_ ( .A(\ID_EX_csr [2] ), .ZN(_04078_ ) );
NAND2_X1 _11805_ ( .A1(_04040_ ), .A2(_04078_ ), .ZN(_04079_ ) );
NAND2_X1 _11806_ ( .A1(_04047_ ), .A2(\ID_EX_csr [0] ), .ZN(_04080_ ) );
NOR2_X1 _11807_ ( .A1(_04079_ ), .A2(_04080_ ), .ZN(_04081_ ) );
BUF_X4 _11808_ ( .A(_04081_ ), .Z(_04082_ ) );
NAND3_X1 _11809_ ( .A1(_04077_ ), .A2(\mepc [30] ), .A3(_04082_ ), .ZN(_04083_ ) );
NAND3_X1 _11810_ ( .A1(_04040_ ), .A2(_04078_ ), .A3(\ID_EX_csr [1] ), .ZN(_04084_ ) );
NOR2_X1 _11811_ ( .A1(_04084_ ), .A2(\ID_EX_csr [0] ), .ZN(_04085_ ) );
BUF_X2 _11812_ ( .A(_04085_ ), .Z(_04086_ ) );
NAND3_X1 _11813_ ( .A1(_04077_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_04086_ ), .ZN(_04087_ ) );
AND2_X1 _11814_ ( .A1(_04083_ ), .A2(_04087_ ), .ZN(_04088_ ) );
NOR2_X1 _11815_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_04089_ ) );
NAND3_X1 _11816_ ( .A1(_04089_ ), .A2(_04044_ ), .A3(_04034_ ), .ZN(_04090_ ) );
NOR3_X1 _11817_ ( .A1(_04090_ ), .A2(\ID_EX_csr [10] ), .A3(_04071_ ), .ZN(_04091_ ) );
BUF_X4 _11818_ ( .A(_04091_ ), .Z(_04092_ ) );
BUF_X4 _11819_ ( .A(_04092_ ), .Z(_04093_ ) );
BUF_X2 _11820_ ( .A(_04093_ ), .Z(_04094_ ) );
NOR3_X1 _11821_ ( .A1(_04080_ ), .A2(\ID_EX_csr [3] ), .A3(_04078_ ), .ZN(_04095_ ) );
BUF_X2 _11822_ ( .A(_04095_ ), .Z(_04096_ ) );
BUF_X2 _11823_ ( .A(_04096_ ), .Z(_04097_ ) );
NAND3_X1 _11824_ ( .A1(_04094_ ), .A2(\mtvec [30] ), .A3(_04097_ ), .ZN(_04098_ ) );
NAND4_X1 _11825_ ( .A1(_04060_ ), .A2(_04073_ ), .A3(\ID_EX_csr [9] ), .A4(\ID_EX_csr [8] ), .ZN(_04099_ ) );
NAND4_X1 _11826_ ( .A1(_04044_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_04100_ ) );
NOR2_X1 _11827_ ( .A1(_04099_ ), .A2(_04100_ ), .ZN(_04101_ ) );
AND2_X1 _11828_ ( .A1(_04101_ ), .A2(_04081_ ), .ZN(_04102_ ) );
INV_X1 _11829_ ( .A(_04102_ ), .ZN(_04103_ ) );
NOR3_X1 _11830_ ( .A1(_04079_ ), .A2(\ID_EX_csr [1] ), .A3(\ID_EX_csr [0] ), .ZN(_04104_ ) );
BUF_X2 _11831_ ( .A(_04104_ ), .Z(_04105_ ) );
BUF_X2 _11832_ ( .A(_04105_ ), .Z(_04106_ ) );
NAND3_X1 _11833_ ( .A1(_04094_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_04106_ ), .ZN(_04107_ ) );
NAND4_X1 _11834_ ( .A1(_04088_ ), .A2(_04098_ ), .A3(_04103_ ), .A4(_04107_ ), .ZN(_04108_ ) );
AOI21_X1 _11835_ ( .A(_04067_ ), .B1(_04069_ ), .B2(_04108_ ), .ZN(_04109_ ) );
INV_X1 _11836_ ( .A(_04109_ ), .ZN(_04110_ ) );
AND2_X1 _11837_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_04111_ ) );
AND2_X1 _11838_ ( .A1(_04111_ ), .A2(\ID_EX_pc [4] ), .ZN(_04112_ ) );
AND2_X1 _11839_ ( .A1(_04112_ ), .A2(\ID_EX_pc [5] ), .ZN(_04113_ ) );
AND2_X1 _11840_ ( .A1(_04113_ ), .A2(\ID_EX_pc [6] ), .ZN(_04114_ ) );
AND2_X1 _11841_ ( .A1(_04114_ ), .A2(\ID_EX_pc [7] ), .ZN(_04115_ ) );
AND2_X1 _11842_ ( .A1(_04115_ ), .A2(\ID_EX_pc [8] ), .ZN(_04116_ ) );
AND2_X1 _11843_ ( .A1(_04116_ ), .A2(\ID_EX_pc [9] ), .ZN(_04117_ ) );
AND2_X1 _11844_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_04118_ ) );
AND2_X1 _11845_ ( .A1(_04117_ ), .A2(_04118_ ), .ZN(_04119_ ) );
AND2_X1 _11846_ ( .A1(_04119_ ), .A2(\ID_EX_pc [12] ), .ZN(_04120_ ) );
AND2_X1 _11847_ ( .A1(_04120_ ), .A2(\ID_EX_pc [13] ), .ZN(_04121_ ) );
AND3_X1 _11848_ ( .A1(_04121_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_04122_ ) );
AND3_X1 _11849_ ( .A1(_04122_ ), .A2(\ID_EX_pc [17] ), .A3(\ID_EX_pc [16] ), .ZN(_04123_ ) );
AND3_X1 _11850_ ( .A1(_04123_ ), .A2(\ID_EX_pc [19] ), .A3(\ID_EX_pc [18] ), .ZN(_04124_ ) );
AND3_X1 _11851_ ( .A1(_04124_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_04125_ ) );
AND3_X1 _11852_ ( .A1(_04125_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_04126_ ) );
AND3_X1 _11853_ ( .A1(_04126_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_pc [24] ), .ZN(_04127_ ) );
AND3_X1 _11854_ ( .A1(_04127_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_04128_ ) );
NAND3_X1 _11855_ ( .A1(_04128_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_04129_ ) );
XNOR2_X1 _11856_ ( .A(_04129_ ), .B(\ID_EX_pc [30] ), .ZN(_04130_ ) );
XOR2_X1 _11857_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_04131_ ) );
XOR2_X1 _11858_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_04132_ ) );
AND2_X1 _11859_ ( .A1(_04131_ ), .A2(_04132_ ), .ZN(_04133_ ) );
XOR2_X1 _11860_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_04134_ ) );
XOR2_X1 _11861_ ( .A(\ID_EX_pc [21] ), .B(\ID_EX_imm [21] ), .Z(_04135_ ) );
AND2_X1 _11862_ ( .A1(_04134_ ), .A2(_04135_ ), .ZN(_04136_ ) );
AND2_X1 _11863_ ( .A1(_04133_ ), .A2(_04136_ ), .ZN(_04137_ ) );
XOR2_X1 _11864_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_04138_ ) );
XOR2_X1 _11865_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_04139_ ) );
AND2_X1 _11866_ ( .A1(_04138_ ), .A2(_04139_ ), .ZN(_04140_ ) );
XOR2_X1 _11867_ ( .A(\ID_EX_pc [17] ), .B(\ID_EX_imm [17] ), .Z(_04141_ ) );
XOR2_X1 _11868_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_04142_ ) );
AND3_X1 _11869_ ( .A1(_04140_ ), .A2(_04141_ ), .A3(_04142_ ), .ZN(_04143_ ) );
XOR2_X1 _11870_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_04144_ ) );
XOR2_X1 _11871_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_04145_ ) );
AND2_X1 _11872_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_04146_ ) );
AND2_X1 _11873_ ( .A1(_04145_ ), .A2(_04146_ ), .ZN(_04147_ ) );
AND2_X1 _11874_ ( .A1(\ID_EX_pc [1] ), .A2(\ID_EX_imm [1] ), .ZN(_04148_ ) );
OAI21_X1 _11875_ ( .A(_04144_ ), .B1(_04147_ ), .B2(_04148_ ), .ZN(_04149_ ) );
INV_X1 _11876_ ( .A(_04149_ ), .ZN(_04150_ ) );
AND2_X1 _11877_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_04151_ ) );
NOR2_X1 _11878_ ( .A1(_04150_ ), .A2(_04151_ ), .ZN(_04152_ ) );
NOR2_X1 _11879_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_04153_ ) );
NOR2_X1 _11880_ ( .A1(_04152_ ), .A2(_04153_ ), .ZN(_04154_ ) );
AND2_X1 _11881_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_04155_ ) );
NOR2_X1 _11882_ ( .A1(_04154_ ), .A2(_04155_ ), .ZN(_04156_ ) );
AND2_X1 _11883_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_04157_ ) );
NOR2_X1 _11884_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_04158_ ) );
NOR3_X1 _11885_ ( .A1(_04156_ ), .A2(_04157_ ), .A3(_04158_ ), .ZN(_04159_ ) );
NOR2_X1 _11886_ ( .A1(_04159_ ), .A2(_04157_ ), .ZN(_04160_ ) );
NOR2_X1 _11887_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_04161_ ) );
NOR2_X1 _11888_ ( .A1(_04160_ ), .A2(_04161_ ), .ZN(_04162_ ) );
AND2_X1 _11889_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_04163_ ) );
NOR2_X1 _11890_ ( .A1(_04162_ ), .A2(_04163_ ), .ZN(_04164_ ) );
AND2_X1 _11891_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_04165_ ) );
NOR2_X1 _11892_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_04166_ ) );
NOR3_X1 _11893_ ( .A1(_04164_ ), .A2(_04165_ ), .A3(_04166_ ), .ZN(_04167_ ) );
NOR2_X1 _11894_ ( .A1(_04167_ ), .A2(_04165_ ), .ZN(_04168_ ) );
NOR2_X1 _11895_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04169_ ) );
NOR2_X1 _11896_ ( .A1(_04168_ ), .A2(_04169_ ), .ZN(_04170_ ) );
AND2_X1 _11897_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04171_ ) );
NOR2_X1 _11898_ ( .A1(_04170_ ), .A2(_04171_ ), .ZN(_04172_ ) );
INV_X1 _11899_ ( .A(_04172_ ), .ZN(_04173_ ) );
XOR2_X1 _11900_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_04174_ ) );
INV_X1 _11901_ ( .A(_04174_ ), .ZN(_04175_ ) );
XNOR2_X1 _11902_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .ZN(_04176_ ) );
NOR2_X1 _11903_ ( .A1(_04175_ ), .A2(_04176_ ), .ZN(_04177_ ) );
XOR2_X1 _11904_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_04178_ ) );
XOR2_X1 _11905_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_04179_ ) );
AND2_X1 _11906_ ( .A1(_04178_ ), .A2(_04179_ ), .ZN(_04180_ ) );
AND2_X1 _11907_ ( .A1(_04177_ ), .A2(_04180_ ), .ZN(_04181_ ) );
XOR2_X1 _11908_ ( .A(\ID_EX_pc [11] ), .B(\ID_EX_imm [11] ), .Z(_04182_ ) );
XOR2_X1 _11909_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_04183_ ) );
AND2_X1 _11910_ ( .A1(_04182_ ), .A2(_04183_ ), .ZN(_04184_ ) );
XOR2_X1 _11911_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_04185_ ) );
XOR2_X1 _11912_ ( .A(\ID_EX_pc [9] ), .B(\ID_EX_imm [9] ), .Z(_04186_ ) );
AND2_X1 _11913_ ( .A1(_04185_ ), .A2(_04186_ ), .ZN(_04187_ ) );
AND2_X1 _11914_ ( .A1(_04184_ ), .A2(_04187_ ), .ZN(_04188_ ) );
AND3_X1 _11915_ ( .A1(_04173_ ), .A2(_04181_ ), .A3(_04188_ ), .ZN(_04189_ ) );
AND2_X1 _11916_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_04190_ ) );
AND2_X1 _11917_ ( .A1(_04182_ ), .A2(_04190_ ), .ZN(_04191_ ) );
AOI21_X1 _11918_ ( .A(_04191_ ), .B1(\ID_EX_pc [11] ), .B2(\ID_EX_imm [11] ), .ZN(_04192_ ) );
AND2_X1 _11919_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_04193_ ) );
AND2_X1 _11920_ ( .A1(_04186_ ), .A2(_04193_ ), .ZN(_04194_ ) );
AOI21_X1 _11921_ ( .A(_04194_ ), .B1(\ID_EX_pc [9] ), .B2(\ID_EX_imm [9] ), .ZN(_04195_ ) );
INV_X1 _11922_ ( .A(_04184_ ), .ZN(_04196_ ) );
OAI21_X1 _11923_ ( .A(_04192_ ), .B1(_04195_ ), .B2(_04196_ ), .ZN(_04197_ ) );
NAND2_X1 _11924_ ( .A1(_04197_ ), .A2(_04181_ ), .ZN(_04198_ ) );
NAND2_X1 _11925_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_04199_ ) );
NOR2_X1 _11926_ ( .A1(_04176_ ), .A2(_04199_ ), .ZN(_04200_ ) );
AOI21_X1 _11927_ ( .A(_04200_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_04201_ ) );
INV_X1 _11928_ ( .A(_04180_ ), .ZN(_04202_ ) );
OR2_X1 _11929_ ( .A1(_04201_ ), .A2(_04202_ ), .ZN(_04203_ ) );
AND2_X1 _11930_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04204_ ) );
AND2_X1 _11931_ ( .A1(_04178_ ), .A2(_04204_ ), .ZN(_04205_ ) );
AOI21_X1 _11932_ ( .A(_04205_ ), .B1(\ID_EX_pc [15] ), .B2(\ID_EX_imm [15] ), .ZN(_04206_ ) );
AND3_X1 _11933_ ( .A1(_04198_ ), .A2(_04203_ ), .A3(_04206_ ), .ZN(_04207_ ) );
INV_X1 _11934_ ( .A(_04207_ ), .ZN(_04208_ ) );
OAI211_X1 _11935_ ( .A(_04137_ ), .B(_04143_ ), .C1(_04189_ ), .C2(_04208_ ), .ZN(_04209_ ) );
NAND3_X1 _11936_ ( .A1(_04131_ ), .A2(\ID_EX_pc [22] ), .A3(\ID_EX_imm [22] ), .ZN(_04210_ ) );
INV_X1 _11937_ ( .A(\ID_EX_pc [23] ), .ZN(_04211_ ) );
NAND3_X1 _11938_ ( .A1(_04138_ ), .A2(\ID_EX_pc [18] ), .A3(\ID_EX_imm [18] ), .ZN(_04212_ ) );
INV_X1 _11939_ ( .A(\ID_EX_pc [19] ), .ZN(_04213_ ) );
OAI21_X1 _11940_ ( .A(_04212_ ), .B1(_04213_ ), .B2(_02941_ ), .ZN(_04214_ ) );
AND2_X1 _11941_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_04215_ ) );
AND2_X1 _11942_ ( .A1(_04141_ ), .A2(_04215_ ), .ZN(_04216_ ) );
AOI21_X1 _11943_ ( .A(_04216_ ), .B1(\ID_EX_pc [17] ), .B2(\ID_EX_imm [17] ), .ZN(_04217_ ) );
INV_X1 _11944_ ( .A(_04217_ ), .ZN(_04218_ ) );
AOI21_X1 _11945_ ( .A(_04214_ ), .B1(_04218_ ), .B2(_04140_ ), .ZN(_04219_ ) );
INV_X1 _11946_ ( .A(_04137_ ), .ZN(_04220_ ) );
OAI221_X1 _11947_ ( .A(_04210_ ), .B1(_04211_ ), .B2(_02397_ ), .C1(_04219_ ), .C2(_04220_ ), .ZN(_04221_ ) );
AND2_X1 _11948_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_04222_ ) );
AND2_X1 _11949_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_04223_ ) );
AOI21_X1 _11950_ ( .A(_04222_ ), .B1(_04135_ ), .B2(_04223_ ), .ZN(_04224_ ) );
INV_X1 _11951_ ( .A(_04224_ ), .ZN(_04225_ ) );
AOI21_X1 _11952_ ( .A(_04221_ ), .B1(_04133_ ), .B2(_04225_ ), .ZN(_04226_ ) );
NAND2_X1 _11953_ ( .A1(_04209_ ), .A2(_04226_ ), .ZN(_04227_ ) );
XOR2_X1 _11954_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_04228_ ) );
XOR2_X1 _11955_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_04229_ ) );
AND2_X1 _11956_ ( .A1(_04228_ ), .A2(_04229_ ), .ZN(_04230_ ) );
XOR2_X1 _11957_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_04231_ ) );
AND2_X1 _11958_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_04232_ ) );
NOR2_X1 _11959_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_04233_ ) );
NOR2_X1 _11960_ ( .A1(_04232_ ), .A2(_04233_ ), .ZN(_04234_ ) );
AND2_X1 _11961_ ( .A1(_04231_ ), .A2(_04234_ ), .ZN(_04235_ ) );
NAND3_X1 _11962_ ( .A1(_04227_ ), .A2(_04230_ ), .A3(_04235_ ), .ZN(_04236_ ) );
AND3_X1 _11963_ ( .A1(_04228_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_imm [26] ), .ZN(_04237_ ) );
NAND2_X1 _11964_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_04238_ ) );
OR3_X1 _11965_ ( .A1(_04232_ ), .A2(_04233_ ), .A3(_04238_ ), .ZN(_04239_ ) );
INV_X1 _11966_ ( .A(\ID_EX_pc [25] ), .ZN(_04240_ ) );
OAI21_X1 _11967_ ( .A(_04239_ ), .B1(_04240_ ), .B2(_03016_ ), .ZN(_04241_ ) );
AOI221_X4 _11968_ ( .A(_04237_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .C1(_04230_ ), .C2(_04241_ ), .ZN(_04242_ ) );
NAND2_X1 _11969_ ( .A1(_04236_ ), .A2(_04242_ ), .ZN(_04243_ ) );
XOR2_X1 _11970_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_04244_ ) );
NAND2_X1 _11971_ ( .A1(_04243_ ), .A2(_04244_ ), .ZN(_04245_ ) );
NAND2_X1 _11972_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_04246_ ) );
INV_X1 _11973_ ( .A(\ID_EX_pc [29] ), .ZN(_04247_ ) );
AOI22_X1 _11974_ ( .A1(_04245_ ), .A2(_04246_ ), .B1(_04247_ ), .B2(_03119_ ), .ZN(_04248_ ) );
AND2_X1 _11975_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_04249_ ) );
OR2_X1 _11976_ ( .A1(_04248_ ), .A2(_04249_ ), .ZN(_04250_ ) );
XOR2_X1 _11977_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .Z(_04251_ ) );
XOR2_X1 _11978_ ( .A(_04250_ ), .B(_04251_ ), .Z(_04252_ ) );
NOR2_X1 _11979_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_7 ), .ZN(_04253_ ) );
AND2_X1 _11980_ ( .A1(_04253_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04254_ ) );
INV_X1 _11981_ ( .A(_04254_ ), .ZN(_04255_ ) );
INV_X1 _11982_ ( .A(_02940_ ), .ZN(_04256_ ) );
INV_X1 _11983_ ( .A(_02335_ ), .ZN(_04257_ ) );
XNOR2_X1 _11984_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .ZN(_04258_ ) );
NAND2_X1 _11985_ ( .A1(_02239_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_04259_ ) );
NAND4_X4 _11986_ ( .A1(_02235_ ), .A2(_04257_ ), .A3(_04258_ ), .A4(_04259_ ), .ZN(_04260_ ) );
BUF_X8 _11987_ ( .A(_04260_ ), .Z(_04261_ ) );
BUF_X4 _11988_ ( .A(_04261_ ), .Z(_04262_ ) );
CLKBUF_X2 _11989_ ( .A(_04262_ ), .Z(_04263_ ) );
NOR2_X1 _11990_ ( .A1(_02239_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_04264_ ) );
AOI21_X1 _11991_ ( .A(_04264_ ), .B1(_02237_ ), .B2(\ID_EX_rs2 [3] ), .ZN(_04265_ ) );
XNOR2_X1 _11992_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_04266_ ) );
XNOR2_X1 _11993_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_04267_ ) );
AOI21_X1 _11994_ ( .A(_02243_ ), .B1(\EX_LS_dest_reg [3] ), .B2(_03479_ ), .ZN(_04268_ ) );
NAND4_X1 _11995_ ( .A1(_04265_ ), .A2(_04266_ ), .A3(_04267_ ), .A4(_04268_ ), .ZN(_04269_ ) );
CLKBUF_X2 _11996_ ( .A(_04269_ ), .Z(_04270_ ) );
BUF_X2 _11997_ ( .A(_04270_ ), .Z(_04271_ ) );
CLKBUF_X2 _11998_ ( .A(_04271_ ), .Z(_04272_ ) );
OR3_X1 _11999_ ( .A1(_04263_ ), .A2(\EX_LS_result_reg [19] ), .A3(_04272_ ), .ZN(_04273_ ) );
INV_X1 _12000_ ( .A(fanout_net_43 ), .ZN(_04274_ ) );
BUF_X4 _12001_ ( .A(_04274_ ), .Z(_04275_ ) );
INV_X1 _12002_ ( .A(fanout_net_31 ), .ZN(_04276_ ) );
CLKBUF_X2 _12003_ ( .A(_04276_ ), .Z(_04277_ ) );
BUF_X2 _12004_ ( .A(_04277_ ), .Z(_04278_ ) );
CLKBUF_X2 _12005_ ( .A(_04278_ ), .Z(_04279_ ) );
OR2_X1 _12006_ ( .A1(_04279_ ), .A2(\myreg.Reg[3][19] ), .ZN(_04280_ ) );
OAI211_X1 _12007_ ( .A(_04280_ ), .B(fanout_net_40 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[2][19] ), .ZN(_04281_ ) );
INV_X1 _12008_ ( .A(fanout_net_42 ), .ZN(_04282_ ) );
BUF_X4 _12009_ ( .A(_04282_ ), .Z(_04283_ ) );
BUF_X4 _12010_ ( .A(_04283_ ), .Z(_04284_ ) );
BUF_X4 _12011_ ( .A(_04284_ ), .Z(_04285_ ) );
OR2_X1 _12012_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[0][19] ), .ZN(_04286_ ) );
INV_X1 _12013_ ( .A(fanout_net_40 ), .ZN(_04287_ ) );
BUF_X4 _12014_ ( .A(_04287_ ), .Z(_04288_ ) );
BUF_X4 _12015_ ( .A(_04288_ ), .Z(_04289_ ) );
BUF_X4 _12016_ ( .A(_04289_ ), .Z(_04290_ ) );
BUF_X4 _12017_ ( .A(_04290_ ), .Z(_04291_ ) );
BUF_X2 _12018_ ( .A(_04276_ ), .Z(_04292_ ) );
BUF_X2 _12019_ ( .A(_04292_ ), .Z(_04293_ ) );
BUF_X4 _12020_ ( .A(_04293_ ), .Z(_04294_ ) );
OAI211_X1 _12021_ ( .A(_04286_ ), .B(_04291_ ), .C1(_04294_ ), .C2(\myreg.Reg[1][19] ), .ZN(_04295_ ) );
NAND3_X1 _12022_ ( .A1(_04281_ ), .A2(_04285_ ), .A3(_04295_ ), .ZN(_04296_ ) );
MUX2_X1 _12023_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_31 ), .Z(_04297_ ) );
MUX2_X1 _12024_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_31 ), .Z(_04298_ ) );
MUX2_X1 _12025_ ( .A(_04297_ ), .B(_04298_ ), .S(_04290_ ), .Z(_04299_ ) );
BUF_X4 _12026_ ( .A(_04285_ ), .Z(_04300_ ) );
OAI211_X1 _12027_ ( .A(_04275_ ), .B(_04296_ ), .C1(_04299_ ), .C2(_04300_ ), .ZN(_04301_ ) );
OR2_X1 _12028_ ( .A1(_04293_ ), .A2(\myreg.Reg[13][19] ), .ZN(_04302_ ) );
OAI211_X1 _12029_ ( .A(_04302_ ), .B(_04291_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[12][19] ), .ZN(_04303_ ) );
OR2_X1 _12030_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[14][19] ), .ZN(_04304_ ) );
OAI211_X1 _12031_ ( .A(_04304_ ), .B(fanout_net_40 ), .C1(_04294_ ), .C2(\myreg.Reg[15][19] ), .ZN(_04305_ ) );
NAND3_X1 _12032_ ( .A1(_04303_ ), .A2(fanout_net_42 ), .A3(_04305_ ), .ZN(_04306_ ) );
MUX2_X1 _12033_ ( .A(\myreg.Reg[8][19] ), .B(\myreg.Reg[9][19] ), .S(fanout_net_31 ), .Z(_04307_ ) );
MUX2_X1 _12034_ ( .A(\myreg.Reg[10][19] ), .B(\myreg.Reg[11][19] ), .S(fanout_net_31 ), .Z(_04308_ ) );
MUX2_X1 _12035_ ( .A(_04307_ ), .B(_04308_ ), .S(fanout_net_40 ), .Z(_04309_ ) );
OAI211_X1 _12036_ ( .A(fanout_net_43 ), .B(_04306_ ), .C1(_04309_ ), .C2(fanout_net_42 ), .ZN(_04310_ ) );
OAI211_X1 _12037_ ( .A(_04301_ ), .B(_04310_ ), .C1(_04263_ ), .C2(_04272_ ), .ZN(_04311_ ) );
NAND2_X1 _12038_ ( .A1(_04273_ ), .A2(_04311_ ), .ZN(_04312_ ) );
XNOR2_X2 _12039_ ( .A(_04256_ ), .B(_04312_ ), .ZN(_04313_ ) );
OR2_X1 _12040_ ( .A1(_04279_ ), .A2(\myreg.Reg[9][18] ), .ZN(_04314_ ) );
BUF_X4 _12041_ ( .A(_04290_ ), .Z(_04315_ ) );
OAI211_X1 _12042_ ( .A(_04314_ ), .B(_04315_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[8][18] ), .ZN(_04316_ ) );
OR2_X1 _12043_ ( .A1(_04279_ ), .A2(\myreg.Reg[11][18] ), .ZN(_04317_ ) );
OAI211_X1 _12044_ ( .A(_04317_ ), .B(fanout_net_40 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[10][18] ), .ZN(_04318_ ) );
NAND3_X1 _12045_ ( .A1(_04316_ ), .A2(_04318_ ), .A3(_04300_ ), .ZN(_04319_ ) );
MUX2_X1 _12046_ ( .A(\myreg.Reg[14][18] ), .B(\myreg.Reg[15][18] ), .S(fanout_net_31 ), .Z(_04320_ ) );
MUX2_X1 _12047_ ( .A(\myreg.Reg[12][18] ), .B(\myreg.Reg[13][18] ), .S(fanout_net_31 ), .Z(_04321_ ) );
MUX2_X1 _12048_ ( .A(_04320_ ), .B(_04321_ ), .S(_04291_ ), .Z(_04322_ ) );
BUF_X4 _12049_ ( .A(_04285_ ), .Z(_04323_ ) );
OAI211_X1 _12050_ ( .A(fanout_net_43 ), .B(_04319_ ), .C1(_04322_ ), .C2(_04323_ ), .ZN(_04324_ ) );
MUX2_X1 _12051_ ( .A(\myreg.Reg[2][18] ), .B(\myreg.Reg[3][18] ), .S(fanout_net_31 ), .Z(_04325_ ) );
AND2_X1 _12052_ ( .A1(_04325_ ), .A2(fanout_net_40 ), .ZN(_04326_ ) );
BUF_X4 _12053_ ( .A(_04291_ ), .Z(_04327_ ) );
MUX2_X1 _12054_ ( .A(\myreg.Reg[0][18] ), .B(\myreg.Reg[1][18] ), .S(fanout_net_31 ), .Z(_04328_ ) );
AOI211_X1 _12055_ ( .A(fanout_net_42 ), .B(_04326_ ), .C1(_04327_ ), .C2(_04328_ ), .ZN(_04329_ ) );
MUX2_X1 _12056_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_31 ), .Z(_04330_ ) );
MUX2_X1 _12057_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_31 ), .Z(_04331_ ) );
MUX2_X1 _12058_ ( .A(_04330_ ), .B(_04331_ ), .S(_04290_ ), .Z(_04332_ ) );
OAI21_X1 _12059_ ( .A(_04275_ ), .B1(_04332_ ), .B2(_04300_ ), .ZN(_04333_ ) );
CLKBUF_X3 _12060_ ( .A(_04262_ ), .Z(_04334_ ) );
BUF_X2 _12061_ ( .A(_04271_ ), .Z(_04335_ ) );
OAI221_X1 _12062_ ( .A(_04324_ ), .B1(_04329_ ), .B2(_04333_ ), .C1(_04334_ ), .C2(_04335_ ), .ZN(_04336_ ) );
OR3_X1 _12063_ ( .A1(_04263_ ), .A2(\EX_LS_result_reg [18] ), .A3(_04272_ ), .ZN(_04337_ ) );
NAND2_X1 _12064_ ( .A1(_04336_ ), .A2(_04337_ ), .ZN(_04338_ ) );
NAND2_X1 _12065_ ( .A1(_04338_ ), .A2(_02917_ ), .ZN(_04339_ ) );
NAND4_X1 _12066_ ( .A1(_04336_ ), .A2(_04337_ ), .A3(_02897_ ), .A4(_02916_ ), .ZN(_04340_ ) );
AND3_X1 _12067_ ( .A1(_04313_ ), .A2(_04339_ ), .A3(_04340_ ), .ZN(_04341_ ) );
INV_X1 _12068_ ( .A(_02472_ ), .ZN(_04342_ ) );
OR2_X1 _12069_ ( .A1(_04294_ ), .A2(\myreg.Reg[9][16] ), .ZN(_04343_ ) );
OAI211_X1 _12070_ ( .A(_04343_ ), .B(_04327_ ), .C1(fanout_net_31 ), .C2(\myreg.Reg[8][16] ), .ZN(_04344_ ) );
BUF_X4 _12071_ ( .A(_04300_ ), .Z(_04345_ ) );
OR2_X1 _12072_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[10][16] ), .ZN(_04346_ ) );
BUF_X4 _12073_ ( .A(_04294_ ), .Z(_04347_ ) );
OAI211_X1 _12074_ ( .A(_04346_ ), .B(fanout_net_40 ), .C1(_04347_ ), .C2(\myreg.Reg[11][16] ), .ZN(_04348_ ) );
NAND3_X1 _12075_ ( .A1(_04344_ ), .A2(_04345_ ), .A3(_04348_ ), .ZN(_04349_ ) );
MUX2_X1 _12076_ ( .A(\myreg.Reg[14][16] ), .B(\myreg.Reg[15][16] ), .S(fanout_net_31 ), .Z(_04350_ ) );
MUX2_X1 _12077_ ( .A(\myreg.Reg[12][16] ), .B(\myreg.Reg[13][16] ), .S(fanout_net_31 ), .Z(_04351_ ) );
MUX2_X1 _12078_ ( .A(_04350_ ), .B(_04351_ ), .S(_04327_ ), .Z(_04352_ ) );
BUF_X4 _12079_ ( .A(_04300_ ), .Z(_04353_ ) );
OAI211_X1 _12080_ ( .A(fanout_net_43 ), .B(_04349_ ), .C1(_04352_ ), .C2(_04353_ ), .ZN(_04354_ ) );
MUX2_X1 _12081_ ( .A(\myreg.Reg[2][16] ), .B(\myreg.Reg[3][16] ), .S(fanout_net_31 ), .Z(_04355_ ) );
AND2_X1 _12082_ ( .A1(_04355_ ), .A2(fanout_net_40 ), .ZN(_04356_ ) );
BUF_X4 _12083_ ( .A(_04315_ ), .Z(_04357_ ) );
MUX2_X1 _12084_ ( .A(\myreg.Reg[0][16] ), .B(\myreg.Reg[1][16] ), .S(fanout_net_31 ), .Z(_04358_ ) );
AOI211_X1 _12085_ ( .A(fanout_net_42 ), .B(_04356_ ), .C1(_04357_ ), .C2(_04358_ ), .ZN(_04359_ ) );
BUF_X4 _12086_ ( .A(_04275_ ), .Z(_04360_ ) );
MUX2_X1 _12087_ ( .A(\myreg.Reg[6][16] ), .B(\myreg.Reg[7][16] ), .S(fanout_net_31 ), .Z(_04361_ ) );
MUX2_X1 _12088_ ( .A(\myreg.Reg[4][16] ), .B(\myreg.Reg[5][16] ), .S(fanout_net_31 ), .Z(_04362_ ) );
BUF_X4 _12089_ ( .A(_04290_ ), .Z(_04363_ ) );
MUX2_X1 _12090_ ( .A(_04361_ ), .B(_04362_ ), .S(_04363_ ), .Z(_04364_ ) );
OAI21_X1 _12091_ ( .A(_04360_ ), .B1(_04364_ ), .B2(_04345_ ), .ZN(_04365_ ) );
BUF_X2 _12092_ ( .A(_04263_ ), .Z(_04366_ ) );
BUF_X2 _12093_ ( .A(_04272_ ), .Z(_04367_ ) );
OAI221_X1 _12094_ ( .A(_04354_ ), .B1(_04359_ ), .B2(_04365_ ), .C1(_04366_ ), .C2(_04367_ ), .ZN(_04368_ ) );
OR3_X1 _12095_ ( .A1(_04334_ ), .A2(\EX_LS_result_reg [16] ), .A3(_04335_ ), .ZN(_04369_ ) );
NAND2_X1 _12096_ ( .A1(_04368_ ), .A2(_04369_ ), .ZN(_04370_ ) );
XNOR2_X1 _12097_ ( .A(_04342_ ), .B(_04370_ ), .ZN(_04371_ ) );
INV_X1 _12098_ ( .A(_02965_ ), .ZN(_04372_ ) );
OR3_X1 _12099_ ( .A1(_04263_ ), .A2(\EX_LS_result_reg [17] ), .A3(_04272_ ), .ZN(_04373_ ) );
OR2_X1 _12100_ ( .A1(_04279_ ), .A2(\myreg.Reg[7][17] ), .ZN(_04374_ ) );
OAI211_X1 _12101_ ( .A(_04374_ ), .B(fanout_net_40 ), .C1(fanout_net_31 ), .C2(\myreg.Reg[6][17] ), .ZN(_04375_ ) );
OR2_X1 _12102_ ( .A1(fanout_net_31 ), .A2(\myreg.Reg[4][17] ), .ZN(_04376_ ) );
OAI211_X1 _12103_ ( .A(_04376_ ), .B(_04291_ ), .C1(_04294_ ), .C2(\myreg.Reg[5][17] ), .ZN(_04377_ ) );
NAND3_X1 _12104_ ( .A1(_04375_ ), .A2(fanout_net_42 ), .A3(_04377_ ), .ZN(_04378_ ) );
MUX2_X1 _12105_ ( .A(\myreg.Reg[2][17] ), .B(\myreg.Reg[3][17] ), .S(fanout_net_31 ), .Z(_04379_ ) );
MUX2_X1 _12106_ ( .A(\myreg.Reg[0][17] ), .B(\myreg.Reg[1][17] ), .S(fanout_net_31 ), .Z(_04380_ ) );
MUX2_X1 _12107_ ( .A(_04379_ ), .B(_04380_ ), .S(_04291_ ), .Z(_04381_ ) );
OAI211_X1 _12108_ ( .A(_04275_ ), .B(_04378_ ), .C1(_04381_ ), .C2(fanout_net_42 ), .ZN(_04382_ ) );
NOR2_X1 _12109_ ( .A1(_04294_ ), .A2(\myreg.Reg[11][17] ), .ZN(_04383_ ) );
OAI21_X1 _12110_ ( .A(fanout_net_40 ), .B1(fanout_net_31 ), .B2(\myreg.Reg[10][17] ), .ZN(_04384_ ) );
NOR2_X1 _12111_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[8][17] ), .ZN(_04385_ ) );
OAI21_X1 _12112_ ( .A(_04291_ ), .B1(_04294_ ), .B2(\myreg.Reg[9][17] ), .ZN(_04386_ ) );
OAI221_X1 _12113_ ( .A(_04285_ ), .B1(_04383_ ), .B2(_04384_ ), .C1(_04385_ ), .C2(_04386_ ), .ZN(_04387_ ) );
MUX2_X1 _12114_ ( .A(\myreg.Reg[12][17] ), .B(\myreg.Reg[13][17] ), .S(fanout_net_32 ), .Z(_04388_ ) );
MUX2_X1 _12115_ ( .A(\myreg.Reg[14][17] ), .B(\myreg.Reg[15][17] ), .S(fanout_net_32 ), .Z(_04389_ ) );
MUX2_X1 _12116_ ( .A(_04388_ ), .B(_04389_ ), .S(fanout_net_40 ), .Z(_04390_ ) );
OAI211_X1 _12117_ ( .A(fanout_net_43 ), .B(_04387_ ), .C1(_04390_ ), .C2(_04323_ ), .ZN(_04391_ ) );
OAI211_X1 _12118_ ( .A(_04382_ ), .B(_04391_ ), .C1(_04334_ ), .C2(_04335_ ), .ZN(_04392_ ) );
NAND2_X1 _12119_ ( .A1(_04373_ ), .A2(_04392_ ), .ZN(_04393_ ) );
XNOR2_X1 _12120_ ( .A(_04372_ ), .B(_04393_ ), .ZN(_04394_ ) );
AND3_X1 _12121_ ( .A1(_04341_ ), .A2(_04371_ ), .A3(_04394_ ), .ZN(_04395_ ) );
INV_X1 _12122_ ( .A(_02373_ ), .ZN(_04396_ ) );
OR3_X1 _12123_ ( .A1(_04263_ ), .A2(\EX_LS_result_reg [22] ), .A3(_04272_ ), .ZN(_04397_ ) );
OR2_X1 _12124_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[0][22] ), .ZN(_04398_ ) );
BUF_X2 _12125_ ( .A(_04279_ ), .Z(_04399_ ) );
OAI211_X1 _12126_ ( .A(_04398_ ), .B(_04315_ ), .C1(_04399_ ), .C2(\myreg.Reg[1][22] ), .ZN(_04400_ ) );
OR2_X1 _12127_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][22] ), .ZN(_04401_ ) );
OAI211_X1 _12128_ ( .A(_04401_ ), .B(fanout_net_40 ), .C1(_04399_ ), .C2(\myreg.Reg[3][22] ), .ZN(_04402_ ) );
NAND3_X1 _12129_ ( .A1(_04400_ ), .A2(_04402_ ), .A3(_04300_ ), .ZN(_04403_ ) );
MUX2_X1 _12130_ ( .A(\myreg.Reg[6][22] ), .B(\myreg.Reg[7][22] ), .S(fanout_net_32 ), .Z(_04404_ ) );
MUX2_X1 _12131_ ( .A(\myreg.Reg[4][22] ), .B(\myreg.Reg[5][22] ), .S(fanout_net_32 ), .Z(_04405_ ) );
MUX2_X1 _12132_ ( .A(_04404_ ), .B(_04405_ ), .S(_04315_ ), .Z(_04406_ ) );
OAI211_X1 _12133_ ( .A(_04275_ ), .B(_04403_ ), .C1(_04406_ ), .C2(_04323_ ), .ZN(_04407_ ) );
OR2_X1 _12134_ ( .A1(_04279_ ), .A2(\myreg.Reg[15][22] ), .ZN(_04408_ ) );
OAI211_X1 _12135_ ( .A(_04408_ ), .B(fanout_net_40 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[14][22] ), .ZN(_04409_ ) );
OR2_X1 _12136_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][22] ), .ZN(_04410_ ) );
OAI211_X1 _12137_ ( .A(_04410_ ), .B(_04315_ ), .C1(_04399_ ), .C2(\myreg.Reg[13][22] ), .ZN(_04411_ ) );
NAND3_X1 _12138_ ( .A1(_04409_ ), .A2(fanout_net_42 ), .A3(_04411_ ), .ZN(_04412_ ) );
MUX2_X1 _12139_ ( .A(\myreg.Reg[8][22] ), .B(\myreg.Reg[9][22] ), .S(fanout_net_32 ), .Z(_04413_ ) );
MUX2_X1 _12140_ ( .A(\myreg.Reg[10][22] ), .B(\myreg.Reg[11][22] ), .S(fanout_net_32 ), .Z(_04414_ ) );
MUX2_X1 _12141_ ( .A(_04413_ ), .B(_04414_ ), .S(fanout_net_40 ), .Z(_04415_ ) );
OAI211_X1 _12142_ ( .A(fanout_net_43 ), .B(_04412_ ), .C1(_04415_ ), .C2(fanout_net_42 ), .ZN(_04416_ ) );
OAI211_X1 _12143_ ( .A(_04407_ ), .B(_04416_ ), .C1(_04334_ ), .C2(_04335_ ), .ZN(_04417_ ) );
NAND2_X1 _12144_ ( .A1(_04397_ ), .A2(_04417_ ), .ZN(_04418_ ) );
XNOR2_X1 _12145_ ( .A(_04396_ ), .B(_04418_ ), .ZN(_04419_ ) );
INV_X1 _12146_ ( .A(_02396_ ), .ZN(_04420_ ) );
OR3_X1 _12147_ ( .A1(_04263_ ), .A2(\EX_LS_result_reg [23] ), .A3(_04272_ ), .ZN(_04421_ ) );
OR2_X1 _12148_ ( .A1(_04279_ ), .A2(\myreg.Reg[1][23] ), .ZN(_04422_ ) );
OAI211_X1 _12149_ ( .A(_04422_ ), .B(_04291_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[0][23] ), .ZN(_04423_ ) );
OR2_X1 _12150_ ( .A1(_04293_ ), .A2(\myreg.Reg[3][23] ), .ZN(_04424_ ) );
OAI211_X1 _12151_ ( .A(_04424_ ), .B(fanout_net_40 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[2][23] ), .ZN(_04425_ ) );
NAND3_X1 _12152_ ( .A1(_04423_ ), .A2(_04425_ ), .A3(_04285_ ), .ZN(_04426_ ) );
MUX2_X1 _12153_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_32 ), .Z(_04427_ ) );
MUX2_X1 _12154_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_32 ), .Z(_04428_ ) );
MUX2_X1 _12155_ ( .A(_04427_ ), .B(_04428_ ), .S(_04290_ ), .Z(_04429_ ) );
OAI211_X1 _12156_ ( .A(_04275_ ), .B(_04426_ ), .C1(_04429_ ), .C2(_04323_ ), .ZN(_04430_ ) );
OR2_X1 _12157_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[14][23] ), .ZN(_04431_ ) );
OAI211_X1 _12158_ ( .A(_04431_ ), .B(fanout_net_40 ), .C1(_04294_ ), .C2(\myreg.Reg[15][23] ), .ZN(_04432_ ) );
OR2_X1 _12159_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[12][23] ), .ZN(_04433_ ) );
OAI211_X1 _12160_ ( .A(_04433_ ), .B(_04291_ ), .C1(_04294_ ), .C2(\myreg.Reg[13][23] ), .ZN(_04434_ ) );
NAND3_X1 _12161_ ( .A1(_04432_ ), .A2(_04434_ ), .A3(fanout_net_42 ), .ZN(_04435_ ) );
MUX2_X1 _12162_ ( .A(\myreg.Reg[8][23] ), .B(\myreg.Reg[9][23] ), .S(fanout_net_32 ), .Z(_04436_ ) );
MUX2_X1 _12163_ ( .A(\myreg.Reg[10][23] ), .B(\myreg.Reg[11][23] ), .S(fanout_net_32 ), .Z(_04437_ ) );
MUX2_X1 _12164_ ( .A(_04436_ ), .B(_04437_ ), .S(fanout_net_40 ), .Z(_04438_ ) );
OAI211_X1 _12165_ ( .A(fanout_net_43 ), .B(_04435_ ), .C1(_04438_ ), .C2(fanout_net_42 ), .ZN(_04439_ ) );
OAI211_X1 _12166_ ( .A(_04430_ ), .B(_04439_ ), .C1(_04263_ ), .C2(_04272_ ), .ZN(_04440_ ) );
NAND2_X1 _12167_ ( .A1(_04421_ ), .A2(_04440_ ), .ZN(_04441_ ) );
XNOR2_X1 _12168_ ( .A(_04420_ ), .B(_04441_ ), .ZN(_04442_ ) );
AND2_X1 _12169_ ( .A1(_04419_ ), .A2(_04442_ ), .ZN(_04443_ ) );
INV_X1 _12170_ ( .A(_02422_ ), .ZN(_04444_ ) );
OR3_X1 _12171_ ( .A1(_04334_ ), .A2(\EX_LS_result_reg [20] ), .A3(_04335_ ), .ZN(_04445_ ) );
OR2_X1 _12172_ ( .A1(_04294_ ), .A2(\myreg.Reg[1][20] ), .ZN(_04446_ ) );
OAI211_X1 _12173_ ( .A(_04446_ ), .B(_04327_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[0][20] ), .ZN(_04447_ ) );
OR2_X1 _12174_ ( .A1(fanout_net_32 ), .A2(\myreg.Reg[2][20] ), .ZN(_04448_ ) );
BUF_X2 _12175_ ( .A(_04279_ ), .Z(_04449_ ) );
OAI211_X1 _12176_ ( .A(_04448_ ), .B(fanout_net_40 ), .C1(_04449_ ), .C2(\myreg.Reg[3][20] ), .ZN(_04450_ ) );
NAND3_X1 _12177_ ( .A1(_04447_ ), .A2(_04323_ ), .A3(_04450_ ), .ZN(_04451_ ) );
MUX2_X1 _12178_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_32 ), .Z(_04452_ ) );
MUX2_X1 _12179_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_32 ), .Z(_04453_ ) );
MUX2_X1 _12180_ ( .A(_04452_ ), .B(_04453_ ), .S(_04363_ ), .Z(_04454_ ) );
OAI211_X1 _12181_ ( .A(_04360_ ), .B(_04451_ ), .C1(_04454_ ), .C2(_04345_ ), .ZN(_04455_ ) );
OR2_X1 _12182_ ( .A1(_04279_ ), .A2(\myreg.Reg[15][20] ), .ZN(_04456_ ) );
OAI211_X1 _12183_ ( .A(_04456_ ), .B(fanout_net_40 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[14][20] ), .ZN(_04457_ ) );
OR2_X1 _12184_ ( .A1(_04279_ ), .A2(\myreg.Reg[13][20] ), .ZN(_04458_ ) );
OAI211_X1 _12185_ ( .A(_04458_ ), .B(_04363_ ), .C1(fanout_net_32 ), .C2(\myreg.Reg[12][20] ), .ZN(_04459_ ) );
NAND3_X1 _12186_ ( .A1(_04457_ ), .A2(_04459_ ), .A3(fanout_net_42 ), .ZN(_04460_ ) );
MUX2_X1 _12187_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_32 ), .Z(_04461_ ) );
MUX2_X1 _12188_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_32 ), .Z(_04462_ ) );
MUX2_X1 _12189_ ( .A(_04461_ ), .B(_04462_ ), .S(fanout_net_40 ), .Z(_04463_ ) );
OAI211_X1 _12190_ ( .A(fanout_net_43 ), .B(_04460_ ), .C1(_04463_ ), .C2(fanout_net_42 ), .ZN(_04464_ ) );
OAI211_X1 _12191_ ( .A(_04455_ ), .B(_04464_ ), .C1(_04366_ ), .C2(_04367_ ), .ZN(_04465_ ) );
NAND2_X1 _12192_ ( .A1(_04445_ ), .A2(_04465_ ), .ZN(_04466_ ) );
XNOR2_X1 _12193_ ( .A(_04444_ ), .B(_04466_ ), .ZN(_04467_ ) );
AND2_X2 _12194_ ( .A1(_02443_ ), .A2(_02444_ ), .ZN(_04468_ ) );
INV_X1 _12195_ ( .A(_04468_ ), .ZN(_04469_ ) );
OR3_X1 _12196_ ( .A1(_04262_ ), .A2(\EX_LS_result_reg [21] ), .A3(_04271_ ), .ZN(_04470_ ) );
OR2_X1 _12197_ ( .A1(_04293_ ), .A2(\myreg.Reg[1][21] ), .ZN(_04471_ ) );
OAI211_X1 _12198_ ( .A(_04471_ ), .B(_04291_ ), .C1(\myreg.Reg[0][21] ), .C2(fanout_net_32 ), .ZN(_04472_ ) );
OR2_X1 _12199_ ( .A1(_04293_ ), .A2(\myreg.Reg[3][21] ), .ZN(_04473_ ) );
OAI211_X1 _12200_ ( .A(_04473_ ), .B(fanout_net_40 ), .C1(fanout_net_32 ), .C2(\myreg.Reg[2][21] ), .ZN(_04474_ ) );
NAND3_X1 _12201_ ( .A1(_04472_ ), .A2(_04474_ ), .A3(_04285_ ), .ZN(_04475_ ) );
MUX2_X1 _12202_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_32 ), .Z(_04476_ ) );
MUX2_X1 _12203_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_33 ), .Z(_04477_ ) );
MUX2_X1 _12204_ ( .A(_04476_ ), .B(_04477_ ), .S(_04290_ ), .Z(_04478_ ) );
OAI211_X1 _12205_ ( .A(_04275_ ), .B(_04475_ ), .C1(_04478_ ), .C2(_04300_ ), .ZN(_04479_ ) );
OR2_X1 _12206_ ( .A1(_04293_ ), .A2(\myreg.Reg[15][21] ), .ZN(_04480_ ) );
OAI211_X1 _12207_ ( .A(_04480_ ), .B(fanout_net_40 ), .C1(fanout_net_33 ), .C2(\myreg.Reg[14][21] ), .ZN(_04481_ ) );
OR2_X1 _12208_ ( .A1(_04293_ ), .A2(\myreg.Reg[13][21] ), .ZN(_04482_ ) );
OAI211_X1 _12209_ ( .A(_04482_ ), .B(_04290_ ), .C1(fanout_net_33 ), .C2(\myreg.Reg[12][21] ), .ZN(_04483_ ) );
NAND3_X1 _12210_ ( .A1(_04481_ ), .A2(_04483_ ), .A3(fanout_net_42 ), .ZN(_04484_ ) );
MUX2_X1 _12211_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_33 ), .Z(_04485_ ) );
MUX2_X1 _12212_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_33 ), .Z(_04486_ ) );
MUX2_X1 _12213_ ( .A(_04485_ ), .B(_04486_ ), .S(fanout_net_40 ), .Z(_04487_ ) );
OAI211_X1 _12214_ ( .A(fanout_net_43 ), .B(_04484_ ), .C1(_04487_ ), .C2(fanout_net_42 ), .ZN(_04488_ ) );
OAI211_X1 _12215_ ( .A(_04479_ ), .B(_04488_ ), .C1(_04263_ ), .C2(_04272_ ), .ZN(_04489_ ) );
NAND2_X1 _12216_ ( .A1(_04470_ ), .A2(_04489_ ), .ZN(_04490_ ) );
XNOR2_X1 _12217_ ( .A(_04469_ ), .B(_04490_ ), .ZN(_04491_ ) );
AND3_X1 _12218_ ( .A1(_04443_ ), .A2(_04467_ ), .A3(_04491_ ), .ZN(_04492_ ) );
AND2_X1 _12219_ ( .A1(_04395_ ), .A2(_04492_ ), .ZN(_04493_ ) );
OR3_X1 _12220_ ( .A1(_04334_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_04335_ ), .ZN(_04494_ ) );
NAND2_X1 _12221_ ( .A1(_03074_ ), .A2(fanout_net_33 ), .ZN(_04495_ ) );
OAI211_X1 _12222_ ( .A(_04495_ ), .B(_04327_ ), .C1(fanout_net_33 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04496_ ) );
NAND2_X1 _12223_ ( .A1(_03077_ ), .A2(fanout_net_33 ), .ZN(_04497_ ) );
OAI211_X1 _12224_ ( .A(_04497_ ), .B(fanout_net_40 ), .C1(fanout_net_33 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04498_ ) );
NAND3_X1 _12225_ ( .A1(_04496_ ), .A2(_04498_ ), .A3(_04323_ ), .ZN(_04499_ ) );
MUX2_X1 _12226_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04500_ ) );
MUX2_X1 _12227_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04501_ ) );
MUX2_X1 _12228_ ( .A(_04500_ ), .B(_04501_ ), .S(_04363_ ), .Z(_04502_ ) );
OAI211_X1 _12229_ ( .A(_04360_ ), .B(_04499_ ), .C1(_04502_ ), .C2(_04353_ ), .ZN(_04503_ ) );
OR2_X1 _12230_ ( .A1(fanout_net_33 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04504_ ) );
OAI211_X1 _12231_ ( .A(_04504_ ), .B(fanout_net_40 ), .C1(_04347_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04505_ ) );
OR2_X1 _12232_ ( .A1(fanout_net_33 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04506_ ) );
OAI211_X1 _12233_ ( .A(_04506_ ), .B(_04327_ ), .C1(_04449_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04507_ ) );
NAND3_X1 _12234_ ( .A1(_04505_ ), .A2(_04507_ ), .A3(fanout_net_42 ), .ZN(_04508_ ) );
MUX2_X1 _12235_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04509_ ) );
MUX2_X1 _12236_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04510_ ) );
MUX2_X1 _12237_ ( .A(_04509_ ), .B(_04510_ ), .S(fanout_net_40 ), .Z(_04511_ ) );
OAI211_X1 _12238_ ( .A(fanout_net_43 ), .B(_04508_ ), .C1(_04511_ ), .C2(fanout_net_42 ), .ZN(_04512_ ) );
OAI211_X1 _12239_ ( .A(_04503_ ), .B(_04512_ ), .C1(_04366_ ), .C2(_04367_ ), .ZN(_04513_ ) );
NAND2_X1 _12240_ ( .A1(_04494_ ), .A2(_04513_ ), .ZN(_04514_ ) );
XNOR2_X1 _12241_ ( .A(_04514_ ), .B(_03095_ ), .ZN(_04515_ ) );
OR3_X1 _12242_ ( .A1(_04334_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04335_ ), .ZN(_04516_ ) );
OR2_X1 _12243_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04517_ ) );
OAI211_X1 _12244_ ( .A(_04517_ ), .B(_04327_ ), .C1(_04449_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04518_ ) );
OR2_X1 _12245_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04519_ ) );
OAI211_X1 _12246_ ( .A(_04519_ ), .B(fanout_net_40 ), .C1(_04449_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04520_ ) );
NAND3_X1 _12247_ ( .A1(_04518_ ), .A2(_04520_ ), .A3(fanout_net_42 ), .ZN(_04521_ ) );
MUX2_X1 _12248_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04522_ ) );
MUX2_X1 _12249_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04523_ ) );
MUX2_X1 _12250_ ( .A(_04522_ ), .B(_04523_ ), .S(_04363_ ), .Z(_04524_ ) );
OAI211_X1 _12251_ ( .A(_04360_ ), .B(_04521_ ), .C1(_04524_ ), .C2(fanout_net_42 ), .ZN(_04525_ ) );
NOR2_X1 _12252_ ( .A1(_04399_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04526_ ) );
OAI21_X1 _12253_ ( .A(fanout_net_40 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04527_ ) );
NOR2_X1 _12254_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04528_ ) );
OAI21_X1 _12255_ ( .A(_04363_ ), .B1(_04449_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04529_ ) );
OAI221_X1 _12256_ ( .A(_04323_ ), .B1(_04526_ ), .B2(_04527_ ), .C1(_04528_ ), .C2(_04529_ ), .ZN(_04530_ ) );
MUX2_X1 _12257_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04531_ ) );
MUX2_X1 _12258_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04532_ ) );
MUX2_X1 _12259_ ( .A(_04531_ ), .B(_04532_ ), .S(fanout_net_40 ), .Z(_04533_ ) );
OAI211_X1 _12260_ ( .A(fanout_net_43 ), .B(_04530_ ), .C1(_04533_ ), .C2(_04345_ ), .ZN(_04534_ ) );
OAI211_X1 _12261_ ( .A(_04525_ ), .B(_04534_ ), .C1(_04366_ ), .C2(_04367_ ), .ZN(_04535_ ) );
NAND2_X1 _12262_ ( .A1(_04516_ ), .A2(_04535_ ), .ZN(_04536_ ) );
XNOR2_X1 _12263_ ( .A(_04536_ ), .B(_03118_ ), .ZN(_04537_ ) );
AND2_X1 _12264_ ( .A1(_04515_ ), .A2(_04537_ ), .ZN(_04538_ ) );
OR3_X1 _12265_ ( .A1(_04366_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04367_ ), .ZN(_04539_ ) );
OR2_X1 _12266_ ( .A1(_04399_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04540_ ) );
OAI211_X1 _12267_ ( .A(_04540_ ), .B(fanout_net_40 ), .C1(fanout_net_33 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04541_ ) );
OR2_X1 _12268_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04542_ ) );
OAI211_X1 _12269_ ( .A(_04542_ ), .B(_04357_ ), .C1(_04347_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04543_ ) );
NAND3_X1 _12270_ ( .A1(_04541_ ), .A2(fanout_net_42 ), .A3(_04543_ ), .ZN(_04544_ ) );
MUX2_X1 _12271_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04545_ ) );
MUX2_X1 _12272_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04546_ ) );
MUX2_X1 _12273_ ( .A(_04545_ ), .B(_04546_ ), .S(_04357_ ), .Z(_04547_ ) );
OAI211_X1 _12274_ ( .A(_04360_ ), .B(_04544_ ), .C1(_04547_ ), .C2(fanout_net_42 ), .ZN(_04548_ ) );
NOR2_X1 _12275_ ( .A1(_04347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04549_ ) );
OAI21_X1 _12276_ ( .A(fanout_net_41 ), .B1(fanout_net_33 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04550_ ) );
NOR2_X1 _12277_ ( .A1(fanout_net_33 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04551_ ) );
OAI21_X1 _12278_ ( .A(_04357_ ), .B1(_04347_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04552_ ) );
OAI221_X1 _12279_ ( .A(_04345_ ), .B1(_04549_ ), .B2(_04550_ ), .C1(_04551_ ), .C2(_04552_ ), .ZN(_04553_ ) );
MUX2_X1 _12280_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_33 ), .Z(_04554_ ) );
MUX2_X1 _12281_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04555_ ) );
MUX2_X1 _12282_ ( .A(_04554_ ), .B(_04555_ ), .S(fanout_net_41 ), .Z(_04556_ ) );
OAI211_X1 _12283_ ( .A(fanout_net_43 ), .B(_04553_ ), .C1(_04556_ ), .C2(_04353_ ), .ZN(_04557_ ) );
OAI211_X1 _12284_ ( .A(_04548_ ), .B(_04557_ ), .C1(_04366_ ), .C2(_04367_ ), .ZN(_04558_ ) );
NAND2_X1 _12285_ ( .A1(_04539_ ), .A2(_04558_ ), .ZN(_04559_ ) );
XNOR2_X1 _12286_ ( .A(_04559_ ), .B(_03149_ ), .ZN(_04560_ ) );
OR3_X1 _12287_ ( .A1(_04334_ ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_04335_ ), .ZN(_04561_ ) );
OR2_X1 _12288_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04562_ ) );
OAI211_X1 _12289_ ( .A(_04562_ ), .B(_04327_ ), .C1(_04347_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04563_ ) );
OR2_X1 _12290_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04564_ ) );
OAI211_X1 _12291_ ( .A(_04564_ ), .B(fanout_net_41 ), .C1(_04449_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04565_ ) );
NAND3_X1 _12292_ ( .A1(_04563_ ), .A2(_04565_ ), .A3(_04323_ ), .ZN(_04566_ ) );
MUX2_X1 _12293_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04567_ ) );
MUX2_X1 _12294_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04568_ ) );
MUX2_X1 _12295_ ( .A(_04567_ ), .B(_04568_ ), .S(_04363_ ), .Z(_04569_ ) );
OAI211_X1 _12296_ ( .A(fanout_net_43 ), .B(_04566_ ), .C1(_04569_ ), .C2(_04353_ ), .ZN(_04570_ ) );
OR2_X1 _12297_ ( .A1(fanout_net_34 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04571_ ) );
OAI211_X1 _12298_ ( .A(_04571_ ), .B(_04327_ ), .C1(_04347_ ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04572_ ) );
NAND2_X1 _12299_ ( .A1(_02266_ ), .A2(fanout_net_34 ), .ZN(_04573_ ) );
OAI211_X1 _12300_ ( .A(_04573_ ), .B(fanout_net_41 ), .C1(fanout_net_34 ), .C2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04574_ ) );
NAND3_X1 _12301_ ( .A1(_04572_ ), .A2(_04574_ ), .A3(_04323_ ), .ZN(_04575_ ) );
MUX2_X1 _12302_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04576_ ) );
MUX2_X1 _12303_ ( .A(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04577_ ) );
MUX2_X1 _12304_ ( .A(_04576_ ), .B(_04577_ ), .S(_04363_ ), .Z(_04578_ ) );
OAI211_X1 _12305_ ( .A(_04360_ ), .B(_04575_ ), .C1(_04578_ ), .C2(_04353_ ), .ZN(_04579_ ) );
OAI211_X1 _12306_ ( .A(_04570_ ), .B(_04579_ ), .C1(_04366_ ), .C2(_04367_ ), .ZN(_04580_ ) );
NAND2_X1 _12307_ ( .A1(_04561_ ), .A2(_04580_ ), .ZN(_04581_ ) );
INV_X1 _12308_ ( .A(_04581_ ), .ZN(_04582_ ) );
XNOR2_X1 _12309_ ( .A(_02297_ ), .B(_04582_ ), .ZN(_04583_ ) );
AND3_X1 _12310_ ( .A1(_04538_ ), .A2(_04560_ ), .A3(_04583_ ), .ZN(_04584_ ) );
NOR2_X2 _12311_ ( .A1(_04260_ ), .A2(_04269_ ), .ZN(_04585_ ) );
NAND2_X1 _12312_ ( .A1(_04585_ ), .A2(\EX_LS_result_reg [26] ), .ZN(_04586_ ) );
OR2_X1 _12313_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04587_ ) );
OAI211_X1 _12314_ ( .A(_04587_ ), .B(fanout_net_41 ), .C1(_04399_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04588_ ) );
MUX2_X1 _12315_ ( .A(_03054_ ), .B(_03055_ ), .S(fanout_net_34 ), .Z(_04589_ ) );
OAI211_X1 _12316_ ( .A(_04588_ ), .B(_04300_ ), .C1(_04589_ ), .C2(fanout_net_41 ), .ZN(_04590_ ) );
MUX2_X1 _12317_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04591_ ) );
MUX2_X1 _12318_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04592_ ) );
MUX2_X1 _12319_ ( .A(_04591_ ), .B(_04592_ ), .S(_04315_ ), .Z(_04593_ ) );
OAI211_X1 _12320_ ( .A(fanout_net_43 ), .B(_04590_ ), .C1(_04593_ ), .C2(_04345_ ), .ZN(_04594_ ) );
OR2_X1 _12321_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04595_ ) );
OAI211_X1 _12322_ ( .A(_04595_ ), .B(_04315_ ), .C1(_04399_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04596_ ) );
NOR2_X1 _12323_ ( .A1(_04449_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04597_ ) );
OAI21_X1 _12324_ ( .A(fanout_net_41 ), .B1(fanout_net_34 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04598_ ) );
OAI211_X1 _12325_ ( .A(_04596_ ), .B(_04300_ ), .C1(_04597_ ), .C2(_04598_ ), .ZN(_04599_ ) );
MUX2_X1 _12326_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04600_ ) );
MUX2_X1 _12327_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04601_ ) );
MUX2_X1 _12328_ ( .A(_04600_ ), .B(_04601_ ), .S(_04315_ ), .Z(_04602_ ) );
OAI211_X1 _12329_ ( .A(_04360_ ), .B(_04599_ ), .C1(_04602_ ), .C2(_04345_ ), .ZN(_04603_ ) );
OAI211_X1 _12330_ ( .A(_04594_ ), .B(_04603_ ), .C1(_04334_ ), .C2(_04335_ ), .ZN(_04604_ ) );
NAND2_X1 _12331_ ( .A1(_04586_ ), .A2(_04604_ ), .ZN(_04605_ ) );
XNOR2_X1 _12332_ ( .A(_04605_ ), .B(_03063_ ), .ZN(_04606_ ) );
INV_X1 _12333_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04607_ ) );
OR3_X1 _12334_ ( .A1(_04263_ ), .A2(_04607_ ), .A3(_04272_ ), .ZN(_04608_ ) );
OR2_X1 _12335_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04609_ ) );
OAI211_X1 _12336_ ( .A(_04609_ ), .B(_04363_ ), .C1(_04449_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04610_ ) );
NAND2_X1 _12337_ ( .A1(_02308_ ), .A2(fanout_net_34 ), .ZN(_04611_ ) );
OAI211_X1 _12338_ ( .A(_04611_ ), .B(fanout_net_41 ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04612_ ) );
NAND3_X1 _12339_ ( .A1(_04610_ ), .A2(_04612_ ), .A3(_04323_ ), .ZN(_04613_ ) );
MUX2_X1 _12340_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04614_ ) );
MUX2_X1 _12341_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04615_ ) );
MUX2_X1 _12342_ ( .A(_04614_ ), .B(_04615_ ), .S(_04315_ ), .Z(_04616_ ) );
OAI211_X1 _12343_ ( .A(fanout_net_43 ), .B(_04613_ ), .C1(_04616_ ), .C2(_04345_ ), .ZN(_04617_ ) );
OR2_X1 _12344_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04618_ ) );
OAI211_X1 _12345_ ( .A(_04618_ ), .B(_04363_ ), .C1(_04449_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04619_ ) );
NAND2_X1 _12346_ ( .A1(_02323_ ), .A2(fanout_net_34 ), .ZN(_04620_ ) );
OAI211_X1 _12347_ ( .A(_04620_ ), .B(fanout_net_41 ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04621_ ) );
NAND3_X1 _12348_ ( .A1(_04619_ ), .A2(_04621_ ), .A3(_04300_ ), .ZN(_04622_ ) );
MUX2_X1 _12349_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04623_ ) );
MUX2_X1 _12350_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_34 ), .Z(_04624_ ) );
MUX2_X1 _12351_ ( .A(_04623_ ), .B(_04624_ ), .S(_04315_ ), .Z(_04625_ ) );
OAI211_X1 _12352_ ( .A(_04360_ ), .B(_04622_ ), .C1(_04625_ ), .C2(_04345_ ), .ZN(_04626_ ) );
OAI211_X1 _12353_ ( .A(_04617_ ), .B(_04626_ ), .C1(_04334_ ), .C2(_04335_ ), .ZN(_04627_ ) );
NAND2_X1 _12354_ ( .A1(_04608_ ), .A2(_04627_ ), .ZN(_04628_ ) );
XNOR2_X1 _12355_ ( .A(_04628_ ), .B(_02348_ ), .ZN(_04629_ ) );
AND2_X1 _12356_ ( .A1(_04606_ ), .A2(_04629_ ), .ZN(_04630_ ) );
INV_X1 _12357_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04631_ ) );
OR3_X1 _12358_ ( .A1(_04366_ ), .A2(_04631_ ), .A3(_04367_ ), .ZN(_04632_ ) );
OR2_X1 _12359_ ( .A1(_04399_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04633_ ) );
OAI211_X1 _12360_ ( .A(_04633_ ), .B(fanout_net_41 ), .C1(fanout_net_34 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04634_ ) );
OR2_X1 _12361_ ( .A1(fanout_net_34 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04635_ ) );
OAI211_X1 _12362_ ( .A(_04635_ ), .B(_04357_ ), .C1(_04347_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04636_ ) );
NAND3_X1 _12363_ ( .A1(_04634_ ), .A2(_04353_ ), .A3(_04636_ ), .ZN(_04637_ ) );
MUX2_X1 _12364_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04638_ ) );
MUX2_X1 _12365_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04639_ ) );
MUX2_X1 _12366_ ( .A(_04638_ ), .B(_04639_ ), .S(_04357_ ), .Z(_04640_ ) );
OAI211_X1 _12367_ ( .A(fanout_net_43 ), .B(_04637_ ), .C1(_04640_ ), .C2(_04353_ ), .ZN(_04641_ ) );
OR2_X1 _12368_ ( .A1(_04399_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04642_ ) );
OAI211_X1 _12369_ ( .A(_04642_ ), .B(_04357_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04643_ ) );
NAND2_X1 _12370_ ( .A1(_03019_ ), .A2(fanout_net_35 ), .ZN(_04644_ ) );
OAI211_X1 _12371_ ( .A(_04644_ ), .B(fanout_net_41 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04645_ ) );
NAND3_X1 _12372_ ( .A1(_04643_ ), .A2(_04645_ ), .A3(_04353_ ), .ZN(_04646_ ) );
MUX2_X1 _12373_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04647_ ) );
MUX2_X1 _12374_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04648_ ) );
MUX2_X1 _12375_ ( .A(_04647_ ), .B(_04648_ ), .S(_04327_ ), .Z(_04649_ ) );
OAI211_X1 _12376_ ( .A(_04360_ ), .B(_04646_ ), .C1(_04649_ ), .C2(_04353_ ), .ZN(_04650_ ) );
OAI211_X1 _12377_ ( .A(_04641_ ), .B(_04650_ ), .C1(_04366_ ), .C2(_04367_ ), .ZN(_04651_ ) );
NAND2_X1 _12378_ ( .A1(_04632_ ), .A2(_04651_ ), .ZN(_04652_ ) );
XNOR2_X1 _12379_ ( .A(_04652_ ), .B(_03039_ ), .ZN(_04653_ ) );
OR2_X1 _12380_ ( .A1(_04449_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04654_ ) );
OAI211_X1 _12381_ ( .A(_04654_ ), .B(_04357_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04655_ ) );
OR2_X1 _12382_ ( .A1(_04399_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04656_ ) );
OAI211_X1 _12383_ ( .A(_04656_ ), .B(fanout_net_41 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04657_ ) );
NAND3_X1 _12384_ ( .A1(_04655_ ), .A2(_04657_ ), .A3(fanout_net_42 ), .ZN(_04658_ ) );
MUX2_X1 _12385_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04659_ ) );
MUX2_X1 _12386_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04660_ ) );
MUX2_X1 _12387_ ( .A(_04659_ ), .B(_04660_ ), .S(_04357_ ), .Z(_04661_ ) );
OAI211_X1 _12388_ ( .A(_04360_ ), .B(_04658_ ), .C1(_04661_ ), .C2(fanout_net_42 ), .ZN(_04662_ ) );
NOR2_X1 _12389_ ( .A1(_04347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04663_ ) );
OAI21_X1 _12390_ ( .A(fanout_net_41 ), .B1(fanout_net_35 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04664_ ) );
NOR2_X1 _12391_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04665_ ) );
OAI21_X1 _12392_ ( .A(_04357_ ), .B1(_04347_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04666_ ) );
OAI221_X1 _12393_ ( .A(_04345_ ), .B1(_04663_ ), .B2(_04664_ ), .C1(_04665_ ), .C2(_04666_ ), .ZN(_04667_ ) );
MUX2_X1 _12394_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04668_ ) );
MUX2_X1 _12395_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04669_ ) );
MUX2_X1 _12396_ ( .A(_04668_ ), .B(_04669_ ), .S(fanout_net_41 ), .Z(_04670_ ) );
OAI211_X1 _12397_ ( .A(fanout_net_43 ), .B(_04667_ ), .C1(_04670_ ), .C2(_04353_ ), .ZN(_04671_ ) );
AOI21_X1 _12398_ ( .A(_04585_ ), .B1(_04662_ ), .B2(_04671_ ), .ZN(_04672_ ) );
NOR3_X1 _12399_ ( .A1(_04366_ ), .A2(\EX_LS_result_reg [24] ), .A3(_04367_ ), .ZN(_04673_ ) );
NOR2_X1 _12400_ ( .A1(_04672_ ), .A2(_04673_ ), .ZN(_04674_ ) );
XNOR2_X1 _12401_ ( .A(_04674_ ), .B(_03196_ ), .ZN(_04675_ ) );
AND3_X1 _12402_ ( .A1(_04630_ ), .A2(_04653_ ), .A3(_04675_ ), .ZN(_04676_ ) );
AND2_X1 _12403_ ( .A1(_04584_ ), .A2(_04676_ ), .ZN(_04677_ ) );
INV_X1 _12404_ ( .A(_02815_ ), .ZN(_04678_ ) );
OR3_X1 _12405_ ( .A1(_04261_ ), .A2(\EX_LS_result_reg [15] ), .A3(_04270_ ), .ZN(_04679_ ) );
OR2_X1 _12406_ ( .A1(_04277_ ), .A2(\myreg.Reg[9][15] ), .ZN(_04680_ ) );
BUF_X4 _12407_ ( .A(_04288_ ), .Z(_04681_ ) );
OAI211_X1 _12408_ ( .A(_04680_ ), .B(_04681_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[8][15] ), .ZN(_04682_ ) );
OR2_X1 _12409_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[10][15] ), .ZN(_04683_ ) );
BUF_X4 _12410_ ( .A(_04277_ ), .Z(_04684_ ) );
OAI211_X1 _12411_ ( .A(_04683_ ), .B(fanout_net_41 ), .C1(_04684_ ), .C2(\myreg.Reg[11][15] ), .ZN(_04685_ ) );
NAND3_X1 _12412_ ( .A1(_04682_ ), .A2(_04284_ ), .A3(_04685_ ), .ZN(_04686_ ) );
MUX2_X1 _12413_ ( .A(\myreg.Reg[14][15] ), .B(\myreg.Reg[15][15] ), .S(fanout_net_35 ), .Z(_04687_ ) );
MUX2_X1 _12414_ ( .A(\myreg.Reg[12][15] ), .B(\myreg.Reg[13][15] ), .S(fanout_net_35 ), .Z(_04688_ ) );
BUF_X4 _12415_ ( .A(_04288_ ), .Z(_04689_ ) );
MUX2_X1 _12416_ ( .A(_04687_ ), .B(_04688_ ), .S(_04689_ ), .Z(_04690_ ) );
BUF_X4 _12417_ ( .A(_04283_ ), .Z(_04691_ ) );
OAI211_X1 _12418_ ( .A(fanout_net_43 ), .B(_04686_ ), .C1(_04690_ ), .C2(_04691_ ), .ZN(_04692_ ) );
BUF_X4 _12419_ ( .A(_04274_ ), .Z(_04693_ ) );
NOR2_X1 _12420_ ( .A1(_04684_ ), .A2(\myreg.Reg[3][15] ), .ZN(_04694_ ) );
OAI21_X1 _12421_ ( .A(fanout_net_41 ), .B1(fanout_net_35 ), .B2(\myreg.Reg[2][15] ), .ZN(_04695_ ) );
NOR2_X1 _12422_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[0][15] ), .ZN(_04696_ ) );
OAI21_X1 _12423_ ( .A(_04689_ ), .B1(_04684_ ), .B2(\myreg.Reg[1][15] ), .ZN(_04697_ ) );
OAI221_X1 _12424_ ( .A(_04284_ ), .B1(_04694_ ), .B2(_04695_ ), .C1(_04696_ ), .C2(_04697_ ), .ZN(_04698_ ) );
MUX2_X1 _12425_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_35 ), .Z(_04699_ ) );
MUX2_X1 _12426_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_35 ), .Z(_04700_ ) );
MUX2_X1 _12427_ ( .A(_04699_ ), .B(_04700_ ), .S(_04689_ ), .Z(_04701_ ) );
OAI211_X1 _12428_ ( .A(_04693_ ), .B(_04698_ ), .C1(_04701_ ), .C2(_04691_ ), .ZN(_04702_ ) );
BUF_X4 _12429_ ( .A(_04260_ ), .Z(_04703_ ) );
BUF_X2 _12430_ ( .A(_04269_ ), .Z(_04704_ ) );
OAI211_X1 _12431_ ( .A(_04692_ ), .B(_04702_ ), .C1(_04703_ ), .C2(_04704_ ), .ZN(_04705_ ) );
NAND2_X1 _12432_ ( .A1(_04679_ ), .A2(_04705_ ), .ZN(_04706_ ) );
XNOR2_X1 _12433_ ( .A(_04678_ ), .B(_04706_ ), .ZN(_04707_ ) );
INV_X1 _12434_ ( .A(_02838_ ), .ZN(_04708_ ) );
OR3_X1 _12435_ ( .A1(_04703_ ), .A2(\EX_LS_result_reg [14] ), .A3(_04704_ ), .ZN(_04709_ ) );
BUF_X2 _12436_ ( .A(_04276_ ), .Z(_04710_ ) );
OR2_X1 _12437_ ( .A1(_04710_ ), .A2(\myreg.Reg[1][14] ), .ZN(_04711_ ) );
OAI211_X1 _12438_ ( .A(_04711_ ), .B(_04290_ ), .C1(fanout_net_35 ), .C2(\myreg.Reg[0][14] ), .ZN(_04712_ ) );
OR2_X1 _12439_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[2][14] ), .ZN(_04713_ ) );
OAI211_X1 _12440_ ( .A(_04713_ ), .B(fanout_net_41 ), .C1(_04293_ ), .C2(\myreg.Reg[3][14] ), .ZN(_04714_ ) );
NAND3_X1 _12441_ ( .A1(_04712_ ), .A2(_04691_ ), .A3(_04714_ ), .ZN(_04715_ ) );
MUX2_X1 _12442_ ( .A(\myreg.Reg[6][14] ), .B(\myreg.Reg[7][14] ), .S(fanout_net_35 ), .Z(_04716_ ) );
MUX2_X1 _12443_ ( .A(\myreg.Reg[4][14] ), .B(\myreg.Reg[5][14] ), .S(fanout_net_35 ), .Z(_04717_ ) );
BUF_X4 _12444_ ( .A(_04288_ ), .Z(_04718_ ) );
MUX2_X1 _12445_ ( .A(_04716_ ), .B(_04717_ ), .S(_04718_ ), .Z(_04719_ ) );
OAI211_X1 _12446_ ( .A(_04275_ ), .B(_04715_ ), .C1(_04719_ ), .C2(_04285_ ), .ZN(_04720_ ) );
OR2_X1 _12447_ ( .A1(_04292_ ), .A2(\myreg.Reg[15][14] ), .ZN(_04721_ ) );
OAI211_X1 _12448_ ( .A(_04721_ ), .B(fanout_net_41 ), .C1(fanout_net_35 ), .C2(\myreg.Reg[14][14] ), .ZN(_04722_ ) );
OR2_X1 _12449_ ( .A1(fanout_net_35 ), .A2(\myreg.Reg[12][14] ), .ZN(_04723_ ) );
OAI211_X1 _12450_ ( .A(_04723_ ), .B(_04718_ ), .C1(_04278_ ), .C2(\myreg.Reg[13][14] ), .ZN(_04724_ ) );
NAND3_X1 _12451_ ( .A1(_04722_ ), .A2(fanout_net_42 ), .A3(_04724_ ), .ZN(_04725_ ) );
MUX2_X1 _12452_ ( .A(\myreg.Reg[8][14] ), .B(\myreg.Reg[9][14] ), .S(fanout_net_35 ), .Z(_04726_ ) );
MUX2_X1 _12453_ ( .A(\myreg.Reg[10][14] ), .B(\myreg.Reg[11][14] ), .S(fanout_net_36 ), .Z(_04727_ ) );
MUX2_X1 _12454_ ( .A(_04726_ ), .B(_04727_ ), .S(fanout_net_41 ), .Z(_04728_ ) );
OAI211_X1 _12455_ ( .A(fanout_net_43 ), .B(_04725_ ), .C1(_04728_ ), .C2(fanout_net_42 ), .ZN(_04729_ ) );
OAI211_X1 _12456_ ( .A(_04720_ ), .B(_04729_ ), .C1(_04262_ ), .C2(_04271_ ), .ZN(_04730_ ) );
NAND2_X1 _12457_ ( .A1(_04709_ ), .A2(_04730_ ), .ZN(_04731_ ) );
XNOR2_X1 _12458_ ( .A(_04708_ ), .B(_04731_ ), .ZN(_04732_ ) );
AND2_X1 _12459_ ( .A1(_04707_ ), .A2(_04732_ ), .ZN(_04733_ ) );
INV_X1 _12460_ ( .A(_02886_ ), .ZN(_04734_ ) );
OR3_X1 _12461_ ( .A1(_04261_ ), .A2(\EX_LS_result_reg [12] ), .A3(_04270_ ), .ZN(_04735_ ) );
OR2_X1 _12462_ ( .A1(_04277_ ), .A2(\myreg.Reg[9][12] ), .ZN(_04736_ ) );
OAI211_X1 _12463_ ( .A(_04736_ ), .B(_04681_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[8][12] ), .ZN(_04737_ ) );
OR2_X1 _12464_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[10][12] ), .ZN(_04738_ ) );
OAI211_X1 _12465_ ( .A(_04738_ ), .B(fanout_net_41 ), .C1(_04684_ ), .C2(\myreg.Reg[11][12] ), .ZN(_04739_ ) );
NAND3_X1 _12466_ ( .A1(_04737_ ), .A2(_04284_ ), .A3(_04739_ ), .ZN(_04740_ ) );
MUX2_X1 _12467_ ( .A(\myreg.Reg[14][12] ), .B(\myreg.Reg[15][12] ), .S(fanout_net_36 ), .Z(_04741_ ) );
MUX2_X1 _12468_ ( .A(\myreg.Reg[12][12] ), .B(\myreg.Reg[13][12] ), .S(fanout_net_36 ), .Z(_04742_ ) );
MUX2_X1 _12469_ ( .A(_04741_ ), .B(_04742_ ), .S(_04689_ ), .Z(_04743_ ) );
OAI211_X1 _12470_ ( .A(fanout_net_43 ), .B(_04740_ ), .C1(_04743_ ), .C2(_04691_ ), .ZN(_04744_ ) );
NOR2_X1 _12471_ ( .A1(_04710_ ), .A2(\myreg.Reg[3][12] ), .ZN(_04745_ ) );
OAI21_X1 _12472_ ( .A(fanout_net_41 ), .B1(fanout_net_36 ), .B2(\myreg.Reg[2][12] ), .ZN(_04746_ ) );
NOR2_X1 _12473_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[0][12] ), .ZN(_04747_ ) );
OAI21_X1 _12474_ ( .A(_04289_ ), .B1(_04710_ ), .B2(\myreg.Reg[1][12] ), .ZN(_04748_ ) );
OAI221_X1 _12475_ ( .A(_04284_ ), .B1(_04745_ ), .B2(_04746_ ), .C1(_04747_ ), .C2(_04748_ ), .ZN(_04749_ ) );
MUX2_X1 _12476_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_36 ), .Z(_04750_ ) );
MUX2_X1 _12477_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_36 ), .Z(_04751_ ) );
MUX2_X1 _12478_ ( .A(_04750_ ), .B(_04751_ ), .S(_04289_ ), .Z(_04752_ ) );
BUF_X4 _12479_ ( .A(_04283_ ), .Z(_04753_ ) );
OAI211_X1 _12480_ ( .A(_04693_ ), .B(_04749_ ), .C1(_04752_ ), .C2(_04753_ ), .ZN(_04754_ ) );
OAI211_X1 _12481_ ( .A(_04744_ ), .B(_04754_ ), .C1(_04703_ ), .C2(_04704_ ), .ZN(_04755_ ) );
NAND2_X1 _12482_ ( .A1(_04735_ ), .A2(_04755_ ), .ZN(_04756_ ) );
XNOR2_X1 _12483_ ( .A(_04734_ ), .B(_04756_ ), .ZN(_04757_ ) );
AND2_X2 _12484_ ( .A1(_02860_ ), .A2(_02861_ ), .ZN(_04758_ ) );
INV_X1 _12485_ ( .A(_04758_ ), .ZN(_04759_ ) );
OR3_X1 _12486_ ( .A1(_04703_ ), .A2(\EX_LS_result_reg [13] ), .A3(_04704_ ), .ZN(_04760_ ) );
OR2_X1 _12487_ ( .A1(_04292_ ), .A2(\myreg.Reg[3][13] ), .ZN(_04761_ ) );
OAI211_X1 _12488_ ( .A(_04761_ ), .B(fanout_net_41 ), .C1(fanout_net_36 ), .C2(\myreg.Reg[2][13] ), .ZN(_04762_ ) );
OR2_X1 _12489_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[0][13] ), .ZN(_04763_ ) );
OAI211_X1 _12490_ ( .A(_04763_ ), .B(_04718_ ), .C1(_04278_ ), .C2(\myreg.Reg[1][13] ), .ZN(_04764_ ) );
NAND3_X1 _12491_ ( .A1(_04762_ ), .A2(_04753_ ), .A3(_04764_ ), .ZN(_04765_ ) );
MUX2_X1 _12492_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(fanout_net_36 ), .Z(_04766_ ) );
MUX2_X1 _12493_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(fanout_net_36 ), .Z(_04767_ ) );
MUX2_X1 _12494_ ( .A(_04766_ ), .B(_04767_ ), .S(_04681_ ), .Z(_04768_ ) );
OAI211_X1 _12495_ ( .A(_04693_ ), .B(_04765_ ), .C1(_04768_ ), .C2(_04285_ ), .ZN(_04769_ ) );
OR2_X1 _12496_ ( .A1(_04292_ ), .A2(\myreg.Reg[13][13] ), .ZN(_04770_ ) );
OAI211_X1 _12497_ ( .A(_04770_ ), .B(_04718_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[12][13] ), .ZN(_04771_ ) );
OR2_X1 _12498_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][13] ), .ZN(_04772_ ) );
OAI211_X1 _12499_ ( .A(_04772_ ), .B(fanout_net_41 ), .C1(_04278_ ), .C2(\myreg.Reg[15][13] ), .ZN(_04773_ ) );
NAND3_X1 _12500_ ( .A1(_04771_ ), .A2(fanout_net_42 ), .A3(_04773_ ), .ZN(_04774_ ) );
MUX2_X1 _12501_ ( .A(\myreg.Reg[8][13] ), .B(\myreg.Reg[9][13] ), .S(fanout_net_36 ), .Z(_04775_ ) );
MUX2_X1 _12502_ ( .A(\myreg.Reg[10][13] ), .B(\myreg.Reg[11][13] ), .S(fanout_net_36 ), .Z(_04776_ ) );
MUX2_X1 _12503_ ( .A(_04775_ ), .B(_04776_ ), .S(fanout_net_41 ), .Z(_04777_ ) );
OAI211_X1 _12504_ ( .A(fanout_net_43 ), .B(_04774_ ), .C1(_04777_ ), .C2(fanout_net_42 ), .ZN(_04778_ ) );
OAI211_X1 _12505_ ( .A(_04769_ ), .B(_04778_ ), .C1(_04262_ ), .C2(_04271_ ), .ZN(_04779_ ) );
NAND2_X1 _12506_ ( .A1(_04760_ ), .A2(_04779_ ), .ZN(_04780_ ) );
XNOR2_X1 _12507_ ( .A(_04759_ ), .B(_04780_ ), .ZN(_04781_ ) );
AND3_X1 _12508_ ( .A1(_04733_ ), .A2(_04757_ ), .A3(_04781_ ), .ZN(_04782_ ) );
AND2_X2 _12509_ ( .A1(_02545_ ), .A2(_02546_ ), .ZN(_04783_ ) );
INV_X1 _12510_ ( .A(_04783_ ), .ZN(_04784_ ) );
OR3_X1 _12511_ ( .A1(_04261_ ), .A2(\EX_LS_result_reg [11] ), .A3(_04270_ ), .ZN(_04785_ ) );
OR2_X1 _12512_ ( .A1(_04277_ ), .A2(\myreg.Reg[1][11] ), .ZN(_04786_ ) );
OAI211_X1 _12513_ ( .A(_04786_ ), .B(_04689_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[0][11] ), .ZN(_04787_ ) );
BUF_X2 _12514_ ( .A(_04276_ ), .Z(_04788_ ) );
OR2_X1 _12515_ ( .A1(_04788_ ), .A2(\myreg.Reg[3][11] ), .ZN(_04789_ ) );
OAI211_X1 _12516_ ( .A(_04789_ ), .B(fanout_net_41 ), .C1(fanout_net_36 ), .C2(\myreg.Reg[2][11] ), .ZN(_04790_ ) );
NAND3_X1 _12517_ ( .A1(_04787_ ), .A2(_04790_ ), .A3(_04284_ ), .ZN(_04791_ ) );
MUX2_X1 _12518_ ( .A(\myreg.Reg[6][11] ), .B(\myreg.Reg[7][11] ), .S(fanout_net_36 ), .Z(_04792_ ) );
MUX2_X1 _12519_ ( .A(\myreg.Reg[4][11] ), .B(\myreg.Reg[5][11] ), .S(fanout_net_36 ), .Z(_04793_ ) );
MUX2_X1 _12520_ ( .A(_04792_ ), .B(_04793_ ), .S(_04289_ ), .Z(_04794_ ) );
OAI211_X1 _12521_ ( .A(_04693_ ), .B(_04791_ ), .C1(_04794_ ), .C2(_04753_ ), .ZN(_04795_ ) );
OR2_X1 _12522_ ( .A1(_04277_ ), .A2(\myreg.Reg[13][11] ), .ZN(_04796_ ) );
OAI211_X1 _12523_ ( .A(_04796_ ), .B(_04689_ ), .C1(fanout_net_36 ), .C2(\myreg.Reg[12][11] ), .ZN(_04797_ ) );
OR2_X1 _12524_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][11] ), .ZN(_04798_ ) );
OAI211_X1 _12525_ ( .A(_04798_ ), .B(fanout_net_41 ), .C1(_04710_ ), .C2(\myreg.Reg[15][11] ), .ZN(_04799_ ) );
NAND3_X1 _12526_ ( .A1(_04797_ ), .A2(fanout_net_42 ), .A3(_04799_ ), .ZN(_04800_ ) );
MUX2_X1 _12527_ ( .A(\myreg.Reg[8][11] ), .B(\myreg.Reg[9][11] ), .S(fanout_net_36 ), .Z(_04801_ ) );
MUX2_X1 _12528_ ( .A(\myreg.Reg[10][11] ), .B(\myreg.Reg[11][11] ), .S(fanout_net_36 ), .Z(_04802_ ) );
MUX2_X1 _12529_ ( .A(_04801_ ), .B(_04802_ ), .S(fanout_net_41 ), .Z(_04803_ ) );
OAI211_X1 _12530_ ( .A(fanout_net_43 ), .B(_04800_ ), .C1(_04803_ ), .C2(fanout_net_42 ), .ZN(_04804_ ) );
OAI211_X1 _12531_ ( .A(_04795_ ), .B(_04804_ ), .C1(_04703_ ), .C2(_04704_ ), .ZN(_04805_ ) );
NAND2_X1 _12532_ ( .A1(_04785_ ), .A2(_04805_ ), .ZN(_04806_ ) );
XNOR2_X1 _12533_ ( .A(_04784_ ), .B(_04806_ ), .ZN(_04807_ ) );
INV_X1 _12534_ ( .A(_02571_ ), .ZN(_04808_ ) );
OR3_X1 _12535_ ( .A1(_04703_ ), .A2(\EX_LS_result_reg [10] ), .A3(_04704_ ), .ZN(_04809_ ) );
OR2_X1 _12536_ ( .A1(_04292_ ), .A2(\myreg.Reg[3][10] ), .ZN(_04810_ ) );
OAI211_X1 _12537_ ( .A(_04810_ ), .B(fanout_net_41 ), .C1(fanout_net_36 ), .C2(\myreg.Reg[2][10] ), .ZN(_04811_ ) );
OR2_X1 _12538_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[0][10] ), .ZN(_04812_ ) );
OAI211_X1 _12539_ ( .A(_04812_ ), .B(_04718_ ), .C1(_04278_ ), .C2(\myreg.Reg[1][10] ), .ZN(_04813_ ) );
NAND3_X1 _12540_ ( .A1(_04811_ ), .A2(_04753_ ), .A3(_04813_ ), .ZN(_04814_ ) );
MUX2_X1 _12541_ ( .A(\myreg.Reg[6][10] ), .B(\myreg.Reg[7][10] ), .S(fanout_net_36 ), .Z(_04815_ ) );
MUX2_X1 _12542_ ( .A(\myreg.Reg[4][10] ), .B(\myreg.Reg[5][10] ), .S(fanout_net_36 ), .Z(_04816_ ) );
MUX2_X1 _12543_ ( .A(_04815_ ), .B(_04816_ ), .S(_04681_ ), .Z(_04817_ ) );
OAI211_X1 _12544_ ( .A(_04275_ ), .B(_04814_ ), .C1(_04817_ ), .C2(_04285_ ), .ZN(_04818_ ) );
OR2_X1 _12545_ ( .A1(fanout_net_36 ), .A2(\myreg.Reg[14][10] ), .ZN(_04819_ ) );
OAI211_X1 _12546_ ( .A(_04819_ ), .B(fanout_net_41 ), .C1(_04278_ ), .C2(\myreg.Reg[15][10] ), .ZN(_04820_ ) );
OR2_X1 _12547_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][10] ), .ZN(_04821_ ) );
OAI211_X1 _12548_ ( .A(_04821_ ), .B(_04718_ ), .C1(_04278_ ), .C2(\myreg.Reg[13][10] ), .ZN(_04822_ ) );
NAND3_X1 _12549_ ( .A1(_04820_ ), .A2(_04822_ ), .A3(fanout_net_42 ), .ZN(_04823_ ) );
MUX2_X1 _12550_ ( .A(\myreg.Reg[8][10] ), .B(\myreg.Reg[9][10] ), .S(fanout_net_37 ), .Z(_04824_ ) );
MUX2_X1 _12551_ ( .A(\myreg.Reg[10][10] ), .B(\myreg.Reg[11][10] ), .S(fanout_net_37 ), .Z(_04825_ ) );
MUX2_X1 _12552_ ( .A(_04824_ ), .B(_04825_ ), .S(fanout_net_41 ), .Z(_04826_ ) );
OAI211_X1 _12553_ ( .A(fanout_net_43 ), .B(_04823_ ), .C1(_04826_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04827_ ) );
OAI211_X1 _12554_ ( .A(_04818_ ), .B(_04827_ ), .C1(_04262_ ), .C2(_04271_ ), .ZN(_04828_ ) );
NAND2_X1 _12555_ ( .A1(_04809_ ), .A2(_04828_ ), .ZN(_04829_ ) );
XNOR2_X1 _12556_ ( .A(_04808_ ), .B(_04829_ ), .ZN(_04830_ ) );
AND2_X1 _12557_ ( .A1(_04807_ ), .A2(_04830_ ), .ZN(_04831_ ) );
AND2_X2 _12558_ ( .A1(_02520_ ), .A2(_02521_ ), .ZN(_04832_ ) );
INV_X1 _12559_ ( .A(_04832_ ), .ZN(_04833_ ) );
OR3_X1 _12560_ ( .A1(_04261_ ), .A2(\EX_LS_result_reg [9] ), .A3(_04270_ ), .ZN(_04834_ ) );
OR2_X1 _12561_ ( .A1(_04788_ ), .A2(\myreg.Reg[1][9] ), .ZN(_04835_ ) );
OAI211_X1 _12562_ ( .A(_04835_ ), .B(_04689_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[0][9] ), .ZN(_04836_ ) );
OR2_X1 _12563_ ( .A1(_04788_ ), .A2(\myreg.Reg[3][9] ), .ZN(_04837_ ) );
OAI211_X1 _12564_ ( .A(_04837_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[2][9] ), .ZN(_04838_ ) );
NAND3_X1 _12565_ ( .A1(_04836_ ), .A2(_04838_ ), .A3(_04283_ ), .ZN(_04839_ ) );
MUX2_X1 _12566_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_37 ), .Z(_04840_ ) );
MUX2_X1 _12567_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_37 ), .Z(_04841_ ) );
MUX2_X1 _12568_ ( .A(_04840_ ), .B(_04841_ ), .S(_04289_ ), .Z(_04842_ ) );
OAI211_X1 _12569_ ( .A(_04693_ ), .B(_04839_ ), .C1(_04842_ ), .C2(_04753_ ), .ZN(_04843_ ) );
OR2_X1 _12570_ ( .A1(_04788_ ), .A2(\myreg.Reg[13][9] ), .ZN(_04844_ ) );
OAI211_X1 _12571_ ( .A(_04844_ ), .B(_04289_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[12][9] ), .ZN(_04845_ ) );
OR2_X1 _12572_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[14][9] ), .ZN(_04846_ ) );
OAI211_X1 _12573_ ( .A(_04846_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04710_ ), .C2(\myreg.Reg[15][9] ), .ZN(_04847_ ) );
NAND3_X1 _12574_ ( .A1(_04845_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04847_ ), .ZN(_04848_ ) );
MUX2_X1 _12575_ ( .A(\myreg.Reg[8][9] ), .B(\myreg.Reg[9][9] ), .S(fanout_net_37 ), .Z(_04849_ ) );
MUX2_X1 _12576_ ( .A(\myreg.Reg[10][9] ), .B(\myreg.Reg[11][9] ), .S(fanout_net_37 ), .Z(_04850_ ) );
MUX2_X1 _12577_ ( .A(_04849_ ), .B(_04850_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04851_ ) );
OAI211_X1 _12578_ ( .A(fanout_net_43 ), .B(_04848_ ), .C1(_04851_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04852_ ) );
OAI211_X1 _12579_ ( .A(_04843_ ), .B(_04852_ ), .C1(_04703_ ), .C2(_04704_ ), .ZN(_04853_ ) );
NAND2_X2 _12580_ ( .A1(_04834_ ), .A2(_04853_ ), .ZN(_04854_ ) );
XNOR2_X1 _12581_ ( .A(_04833_ ), .B(_04854_ ), .ZN(_04855_ ) );
INV_X1 _12582_ ( .A(_02498_ ), .ZN(_04856_ ) );
OR3_X1 _12583_ ( .A1(_04262_ ), .A2(\EX_LS_result_reg [8] ), .A3(_04704_ ), .ZN(_04857_ ) );
OR2_X1 _12584_ ( .A1(_04710_ ), .A2(\myreg.Reg[3][8] ), .ZN(_04858_ ) );
OAI211_X1 _12585_ ( .A(_04858_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[2][8] ), .ZN(_04859_ ) );
OR2_X1 _12586_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][8] ), .ZN(_04860_ ) );
OAI211_X1 _12587_ ( .A(_04860_ ), .B(_04290_ ), .C1(_04293_ ), .C2(\myreg.Reg[1][8] ), .ZN(_04861_ ) );
NAND3_X1 _12588_ ( .A1(_04859_ ), .A2(_04691_ ), .A3(_04861_ ), .ZN(_04862_ ) );
MUX2_X1 _12589_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_37 ), .Z(_04863_ ) );
MUX2_X1 _12590_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_37 ), .Z(_04864_ ) );
MUX2_X1 _12591_ ( .A(_04863_ ), .B(_04864_ ), .S(_04718_ ), .Z(_04865_ ) );
OAI211_X1 _12592_ ( .A(_04275_ ), .B(_04862_ ), .C1(_04865_ ), .C2(_04285_ ), .ZN(_04866_ ) );
OR2_X1 _12593_ ( .A1(_04710_ ), .A2(\myreg.Reg[15][8] ), .ZN(_04867_ ) );
OAI211_X1 _12594_ ( .A(_04867_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][8] ), .ZN(_04868_ ) );
OR2_X1 _12595_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][8] ), .ZN(_04869_ ) );
OAI211_X1 _12596_ ( .A(_04869_ ), .B(_04718_ ), .C1(_04293_ ), .C2(\myreg.Reg[13][8] ), .ZN(_04870_ ) );
NAND3_X1 _12597_ ( .A1(_04868_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04870_ ), .ZN(_04871_ ) );
MUX2_X1 _12598_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_37 ), .Z(_04872_ ) );
MUX2_X1 _12599_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_37 ), .Z(_04873_ ) );
MUX2_X1 _12600_ ( .A(_04872_ ), .B(_04873_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04874_ ) );
OAI211_X1 _12601_ ( .A(fanout_net_43 ), .B(_04871_ ), .C1(_04874_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04875_ ) );
OAI211_X1 _12602_ ( .A(_04866_ ), .B(_04875_ ), .C1(_04262_ ), .C2(_04271_ ), .ZN(_04876_ ) );
NAND2_X1 _12603_ ( .A1(_04857_ ), .A2(_04876_ ), .ZN(_04877_ ) );
XNOR2_X1 _12604_ ( .A(_04856_ ), .B(_04877_ ), .ZN(_04878_ ) );
AND2_X1 _12605_ ( .A1(_04855_ ), .A2(_04878_ ), .ZN(_04879_ ) );
AND2_X1 _12606_ ( .A1(_04831_ ), .A2(_04879_ ), .ZN(_04880_ ) );
AND2_X1 _12607_ ( .A1(_04782_ ), .A2(_04880_ ), .ZN(_04881_ ) );
AND3_X1 _12608_ ( .A1(_04493_ ), .A2(_04677_ ), .A3(_04881_ ), .ZN(_04882_ ) );
INV_X1 _12609_ ( .A(_02670_ ), .ZN(_04883_ ) );
OR3_X1 _12610_ ( .A1(_04261_ ), .A2(\EX_LS_result_reg [6] ), .A3(_04270_ ), .ZN(_04884_ ) );
OR2_X1 _12611_ ( .A1(_04788_ ), .A2(\myreg.Reg[7][6] ), .ZN(_04885_ ) );
OAI211_X1 _12612_ ( .A(_04885_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_37 ), .C2(\myreg.Reg[6][6] ), .ZN(_04886_ ) );
OR2_X1 _12613_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[4][6] ), .ZN(_04887_ ) );
OAI211_X1 _12614_ ( .A(_04887_ ), .B(_04289_ ), .C1(_04710_ ), .C2(\myreg.Reg[5][6] ), .ZN(_04888_ ) );
NAND3_X1 _12615_ ( .A1(_04886_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04888_ ), .ZN(_04889_ ) );
MUX2_X1 _12616_ ( .A(\myreg.Reg[2][6] ), .B(\myreg.Reg[3][6] ), .S(fanout_net_37 ), .Z(_04890_ ) );
MUX2_X1 _12617_ ( .A(\myreg.Reg[0][6] ), .B(\myreg.Reg[1][6] ), .S(fanout_net_37 ), .Z(_04891_ ) );
MUX2_X1 _12618_ ( .A(_04890_ ), .B(_04891_ ), .S(_04288_ ), .Z(_04892_ ) );
OAI211_X1 _12619_ ( .A(_04274_ ), .B(_04889_ ), .C1(_04892_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04893_ ) );
NOR2_X1 _12620_ ( .A1(_04292_ ), .A2(\myreg.Reg[11][6] ), .ZN(_04894_ ) );
OAI21_X1 _12621_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_37 ), .B2(\myreg.Reg[10][6] ), .ZN(_04895_ ) );
NOR2_X1 _12622_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][6] ), .ZN(_04896_ ) );
OAI21_X1 _12623_ ( .A(_04288_ ), .B1(_04292_ ), .B2(\myreg.Reg[9][6] ), .ZN(_04897_ ) );
OAI221_X1 _12624_ ( .A(_04283_ ), .B1(_04894_ ), .B2(_04895_ ), .C1(_04896_ ), .C2(_04897_ ), .ZN(_04898_ ) );
MUX2_X1 _12625_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(fanout_net_37 ), .Z(_04899_ ) );
MUX2_X1 _12626_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(fanout_net_37 ), .Z(_04900_ ) );
MUX2_X1 _12627_ ( .A(_04899_ ), .B(_04900_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04901_ ) );
OAI211_X1 _12628_ ( .A(fanout_net_43 ), .B(_04898_ ), .C1(_04901_ ), .C2(_04753_ ), .ZN(_04902_ ) );
OAI211_X1 _12629_ ( .A(_04893_ ), .B(_04902_ ), .C1(_04261_ ), .C2(_04270_ ), .ZN(_04903_ ) );
NAND2_X1 _12630_ ( .A1(_04884_ ), .A2(_04903_ ), .ZN(_04904_ ) );
XNOR2_X1 _12631_ ( .A(_04883_ ), .B(_04904_ ), .ZN(_04905_ ) );
AND2_X2 _12632_ ( .A1(_02646_ ), .A2(_02647_ ), .ZN(_04906_ ) );
INV_X1 _12633_ ( .A(_04906_ ), .ZN(_04907_ ) );
OR3_X1 _12634_ ( .A1(_04261_ ), .A2(\EX_LS_result_reg [7] ), .A3(_04270_ ), .ZN(_04908_ ) );
OR2_X1 _12635_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[4][7] ), .ZN(_04909_ ) );
OAI211_X1 _12636_ ( .A(_04909_ ), .B(_04289_ ), .C1(_04710_ ), .C2(\myreg.Reg[5][7] ), .ZN(_04910_ ) );
OR2_X1 _12637_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[6][7] ), .ZN(_04911_ ) );
OAI211_X1 _12638_ ( .A(_04911_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04710_ ), .C2(\myreg.Reg[7][7] ), .ZN(_04912_ ) );
NAND3_X1 _12639_ ( .A1(_04910_ ), .A2(_04912_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04913_ ) );
MUX2_X1 _12640_ ( .A(\myreg.Reg[2][7] ), .B(\myreg.Reg[3][7] ), .S(fanout_net_37 ), .Z(_04914_ ) );
MUX2_X1 _12641_ ( .A(\myreg.Reg[0][7] ), .B(\myreg.Reg[1][7] ), .S(fanout_net_38 ), .Z(_04915_ ) );
MUX2_X1 _12642_ ( .A(_04914_ ), .B(_04915_ ), .S(_04288_ ), .Z(_04916_ ) );
OAI211_X1 _12643_ ( .A(_04693_ ), .B(_04913_ ), .C1(_04916_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04917_ ) );
NOR2_X1 _12644_ ( .A1(_04292_ ), .A2(\myreg.Reg[11][7] ), .ZN(_04918_ ) );
OAI21_X1 _12645_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_38 ), .B2(\myreg.Reg[10][7] ), .ZN(_04919_ ) );
NOR2_X1 _12646_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[8][7] ), .ZN(_04920_ ) );
OAI21_X1 _12647_ ( .A(_04288_ ), .B1(_04292_ ), .B2(\myreg.Reg[9][7] ), .ZN(_04921_ ) );
OAI221_X1 _12648_ ( .A(_04283_ ), .B1(_04918_ ), .B2(_04919_ ), .C1(_04920_ ), .C2(_04921_ ), .ZN(_04922_ ) );
MUX2_X1 _12649_ ( .A(\myreg.Reg[12][7] ), .B(\myreg.Reg[13][7] ), .S(fanout_net_38 ), .Z(_04923_ ) );
MUX2_X1 _12650_ ( .A(\myreg.Reg[14][7] ), .B(\myreg.Reg[15][7] ), .S(fanout_net_38 ), .Z(_04924_ ) );
MUX2_X1 _12651_ ( .A(_04923_ ), .B(_04924_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_04925_ ) );
OAI211_X1 _12652_ ( .A(fanout_net_43 ), .B(_04922_ ), .C1(_04925_ ), .C2(_04753_ ), .ZN(_04926_ ) );
OAI211_X1 _12653_ ( .A(_04917_ ), .B(_04926_ ), .C1(_04261_ ), .C2(_04704_ ), .ZN(_04927_ ) );
NAND2_X1 _12654_ ( .A1(_04908_ ), .A2(_04927_ ), .ZN(_04928_ ) );
XNOR2_X1 _12655_ ( .A(_04907_ ), .B(_04928_ ), .ZN(_04929_ ) );
AND2_X1 _12656_ ( .A1(_04905_ ), .A2(_04929_ ), .ZN(_04930_ ) );
OR3_X1 _12657_ ( .A1(_04703_ ), .A2(\EX_LS_result_reg [4] ), .A3(_04270_ ), .ZN(_04931_ ) );
OR2_X1 _12658_ ( .A1(_04277_ ), .A2(\myreg.Reg[9][4] ), .ZN(_04932_ ) );
OAI211_X1 _12659_ ( .A(_04932_ ), .B(_04681_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[8][4] ), .ZN(_04933_ ) );
OR2_X1 _12660_ ( .A1(_04277_ ), .A2(\myreg.Reg[11][4] ), .ZN(_04934_ ) );
OAI211_X1 _12661_ ( .A(_04934_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_38 ), .C2(\myreg.Reg[10][4] ), .ZN(_04935_ ) );
NAND3_X1 _12662_ ( .A1(_04933_ ), .A2(_04935_ ), .A3(_04753_ ), .ZN(_04936_ ) );
MUX2_X1 _12663_ ( .A(\myreg.Reg[14][4] ), .B(\myreg.Reg[15][4] ), .S(fanout_net_38 ), .Z(_04937_ ) );
MUX2_X1 _12664_ ( .A(\myreg.Reg[12][4] ), .B(\myreg.Reg[13][4] ), .S(fanout_net_38 ), .Z(_04938_ ) );
MUX2_X1 _12665_ ( .A(_04937_ ), .B(_04938_ ), .S(_04681_ ), .Z(_04939_ ) );
OAI211_X1 _12666_ ( .A(fanout_net_43 ), .B(_04936_ ), .C1(_04939_ ), .C2(_04691_ ), .ZN(_04940_ ) );
OR2_X1 _12667_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][4] ), .ZN(_04941_ ) );
OAI211_X1 _12668_ ( .A(_04941_ ), .B(_04681_ ), .C1(_04684_ ), .C2(\myreg.Reg[1][4] ), .ZN(_04942_ ) );
NOR2_X1 _12669_ ( .A1(_04278_ ), .A2(\myreg.Reg[3][4] ), .ZN(_04943_ ) );
OAI21_X1 _12670_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_38 ), .B2(\myreg.Reg[2][4] ), .ZN(_04944_ ) );
OAI211_X1 _12671_ ( .A(_04942_ ), .B(_04284_ ), .C1(_04943_ ), .C2(_04944_ ), .ZN(_04945_ ) );
MUX2_X1 _12672_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_38 ), .Z(_04946_ ) );
MUX2_X1 _12673_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_38 ), .Z(_04947_ ) );
MUX2_X1 _12674_ ( .A(_04946_ ), .B(_04947_ ), .S(_04689_ ), .Z(_04948_ ) );
OAI211_X1 _12675_ ( .A(_04693_ ), .B(_04945_ ), .C1(_04948_ ), .C2(_04691_ ), .ZN(_04949_ ) );
OAI211_X1 _12676_ ( .A(_04940_ ), .B(_04949_ ), .C1(_04262_ ), .C2(_04271_ ), .ZN(_04950_ ) );
NAND2_X1 _12677_ ( .A1(_04931_ ), .A2(_04950_ ), .ZN(_04951_ ) );
XNOR2_X1 _12678_ ( .A(_02623_ ), .B(_04951_ ), .ZN(_04952_ ) );
OR2_X1 _12679_ ( .A1(fanout_net_38 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04953_ ) );
OAI211_X1 _12680_ ( .A(_04953_ ), .B(_04681_ ), .C1(_04684_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04954_ ) );
OR2_X1 _12681_ ( .A1(fanout_net_38 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04955_ ) );
OAI211_X1 _12682_ ( .A(_04955_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04684_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04956_ ) );
NAND3_X1 _12683_ ( .A1(_04954_ ), .A2(_04956_ ), .A3(_04284_ ), .ZN(_04957_ ) );
MUX2_X1 _12684_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_38 ), .Z(_04958_ ) );
MUX2_X1 _12685_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_38 ), .Z(_04959_ ) );
MUX2_X1 _12686_ ( .A(_04958_ ), .B(_04959_ ), .S(_04689_ ), .Z(_04960_ ) );
OAI211_X1 _12687_ ( .A(fanout_net_43 ), .B(_04957_ ), .C1(_04960_ ), .C2(_04691_ ), .ZN(_04961_ ) );
NAND2_X1 _12688_ ( .A1(_02578_ ), .A2(fanout_net_38 ), .ZN(_04962_ ) );
OAI211_X1 _12689_ ( .A(_04962_ ), .B(_04289_ ), .C1(fanout_net_38 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04963_ ) );
NOR2_X1 _12690_ ( .A1(_04684_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04964_ ) );
OAI21_X1 _12691_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_38 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04965_ ) );
OAI211_X1 _12692_ ( .A(_04963_ ), .B(_04284_ ), .C1(_04964_ ), .C2(_04965_ ), .ZN(_04966_ ) );
MUX2_X1 _12693_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_38 ), .Z(_04967_ ) );
MUX2_X1 _12694_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_38 ), .Z(_04968_ ) );
MUX2_X1 _12695_ ( .A(_04967_ ), .B(_04968_ ), .S(_04289_ ), .Z(_04969_ ) );
OAI211_X1 _12696_ ( .A(_04693_ ), .B(_04966_ ), .C1(_04969_ ), .C2(_04753_ ), .ZN(_04970_ ) );
AOI21_X1 _12697_ ( .A(_04585_ ), .B1(_04961_ ), .B2(_04970_ ), .ZN(_04971_ ) );
AND2_X1 _12698_ ( .A1(_04585_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04972_ ) );
NOR2_X1 _12699_ ( .A1(_04971_ ), .A2(_04972_ ), .ZN(_04973_ ) );
XNOR2_X1 _12700_ ( .A(_04973_ ), .B(_02598_ ), .ZN(_04974_ ) );
AND3_X1 _12701_ ( .A1(_04930_ ), .A2(_04952_ ), .A3(_04974_ ), .ZN(_04975_ ) );
INV_X1 _12702_ ( .A(_02704_ ), .ZN(_04976_ ) );
OR3_X1 _12703_ ( .A1(_04260_ ), .A2(\EX_LS_result_reg [1] ), .A3(_04269_ ), .ZN(_04977_ ) );
OR2_X1 _12704_ ( .A1(_04276_ ), .A2(\myreg.Reg[9][1] ), .ZN(_04978_ ) );
OAI211_X1 _12705_ ( .A(_04978_ ), .B(_04288_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[8][1] ), .ZN(_04979_ ) );
OR2_X1 _12706_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[10][1] ), .ZN(_04980_ ) );
OAI211_X1 _12707_ ( .A(_04980_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04788_ ), .C2(\myreg.Reg[11][1] ), .ZN(_04981_ ) );
NAND3_X1 _12708_ ( .A1(_04979_ ), .A2(_04283_ ), .A3(_04981_ ), .ZN(_04982_ ) );
MUX2_X1 _12709_ ( .A(\myreg.Reg[14][1] ), .B(\myreg.Reg[15][1] ), .S(fanout_net_38 ), .Z(_04983_ ) );
MUX2_X1 _12710_ ( .A(\myreg.Reg[12][1] ), .B(\myreg.Reg[13][1] ), .S(fanout_net_38 ), .Z(_04984_ ) );
MUX2_X1 _12711_ ( .A(_04983_ ), .B(_04984_ ), .S(_04287_ ), .Z(_04985_ ) );
OAI211_X1 _12712_ ( .A(fanout_net_43 ), .B(_04982_ ), .C1(_04985_ ), .C2(_04283_ ), .ZN(_04986_ ) );
NOR2_X1 _12713_ ( .A1(_04788_ ), .A2(\myreg.Reg[3][1] ), .ZN(_04987_ ) );
OAI21_X1 _12714_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_38 ), .B2(\myreg.Reg[2][1] ), .ZN(_04988_ ) );
NOR2_X1 _12715_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][1] ), .ZN(_04989_ ) );
OAI21_X1 _12716_ ( .A(_04287_ ), .B1(_04788_ ), .B2(\myreg.Reg[1][1] ), .ZN(_04990_ ) );
OAI221_X1 _12717_ ( .A(_04282_ ), .B1(_04987_ ), .B2(_04988_ ), .C1(_04989_ ), .C2(_04990_ ), .ZN(_04991_ ) );
MUX2_X1 _12718_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(fanout_net_38 ), .Z(_04992_ ) );
MUX2_X1 _12719_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(fanout_net_38 ), .Z(_04993_ ) );
MUX2_X1 _12720_ ( .A(_04992_ ), .B(_04993_ ), .S(_04287_ ), .Z(_04994_ ) );
OAI211_X1 _12721_ ( .A(_04274_ ), .B(_04991_ ), .C1(_04994_ ), .C2(_04283_ ), .ZN(_04995_ ) );
OAI211_X1 _12722_ ( .A(_04986_ ), .B(_04995_ ), .C1(_04260_ ), .C2(_04269_ ), .ZN(_04996_ ) );
NAND2_X1 _12723_ ( .A1(_04977_ ), .A2(_04996_ ), .ZN(_04997_ ) );
XNOR2_X1 _12724_ ( .A(_04976_ ), .B(_04997_ ), .ZN(_04998_ ) );
INV_X1 _12725_ ( .A(_02774_ ), .ZN(_04999_ ) );
OR3_X1 _12726_ ( .A1(_04703_ ), .A2(\EX_LS_result_reg [2] ), .A3(_04704_ ), .ZN(_05000_ ) );
OR2_X1 _12727_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[0][2] ), .ZN(_05001_ ) );
OAI211_X1 _12728_ ( .A(_05001_ ), .B(_04718_ ), .C1(_04278_ ), .C2(\myreg.Reg[1][2] ), .ZN(_05002_ ) );
OR2_X1 _12729_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[2][2] ), .ZN(_05003_ ) );
OAI211_X1 _12730_ ( .A(_05003_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04278_ ), .C2(\myreg.Reg[3][2] ), .ZN(_05004_ ) );
NAND3_X1 _12731_ ( .A1(_05002_ ), .A2(_05004_ ), .A3(_04753_ ), .ZN(_05005_ ) );
MUX2_X1 _12732_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_39 ), .Z(_05006_ ) );
MUX2_X1 _12733_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_39 ), .Z(_05007_ ) );
MUX2_X1 _12734_ ( .A(_05006_ ), .B(_05007_ ), .S(_04681_ ), .Z(_05008_ ) );
OAI211_X1 _12735_ ( .A(_04693_ ), .B(_05005_ ), .C1(_05008_ ), .C2(_04691_ ), .ZN(_05009_ ) );
OR2_X1 _12736_ ( .A1(_04292_ ), .A2(\myreg.Reg[15][2] ), .ZN(_05010_ ) );
OAI211_X1 _12737_ ( .A(_05010_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_39 ), .C2(\myreg.Reg[14][2] ), .ZN(_05011_ ) );
OR2_X1 _12738_ ( .A1(_04277_ ), .A2(\myreg.Reg[13][2] ), .ZN(_05012_ ) );
OAI211_X1 _12739_ ( .A(_05012_ ), .B(_04718_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[12][2] ), .ZN(_05013_ ) );
NAND3_X1 _12740_ ( .A1(_05011_ ), .A2(_05013_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05014_ ) );
MUX2_X1 _12741_ ( .A(\myreg.Reg[8][2] ), .B(\myreg.Reg[9][2] ), .S(fanout_net_39 ), .Z(_05015_ ) );
MUX2_X1 _12742_ ( .A(\myreg.Reg[10][2] ), .B(\myreg.Reg[11][2] ), .S(fanout_net_39 ), .Z(_05016_ ) );
MUX2_X1 _12743_ ( .A(_05015_ ), .B(_05016_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_05017_ ) );
OAI211_X1 _12744_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05014_ ), .C1(_05017_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05018_ ) );
OAI211_X1 _12745_ ( .A(_05009_ ), .B(_05018_ ), .C1(_04262_ ), .C2(_04271_ ), .ZN(_05019_ ) );
NAND2_X1 _12746_ ( .A1(_05000_ ), .A2(_05019_ ), .ZN(_05020_ ) );
XNOR2_X1 _12747_ ( .A(_04999_ ), .B(_05020_ ), .ZN(_05021_ ) );
OR3_X1 _12748_ ( .A1(_04261_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04270_ ), .ZN(_05022_ ) );
OR2_X1 _12749_ ( .A1(_04277_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05023_ ) );
OAI211_X1 _12750_ ( .A(_05023_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_39 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_05024_ ) );
OR2_X1 _12751_ ( .A1(fanout_net_39 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_05025_ ) );
OAI211_X1 _12752_ ( .A(_05025_ ), .B(_04681_ ), .C1(_04684_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05026_ ) );
NAND3_X1 _12753_ ( .A1(_05024_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_05026_ ), .ZN(_05027_ ) );
MUX2_X1 _12754_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_39 ), .Z(_05028_ ) );
MUX2_X1 _12755_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_39 ), .Z(_05029_ ) );
MUX2_X1 _12756_ ( .A(_05028_ ), .B(_05029_ ), .S(_04689_ ), .Z(_05030_ ) );
OAI211_X1 _12757_ ( .A(_04693_ ), .B(_05027_ ), .C1(_05030_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05031_ ) );
NOR2_X1 _12758_ ( .A1(_04684_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_05032_ ) );
OAI21_X1 _12759_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_39 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_05033_ ) );
MUX2_X1 _12760_ ( .A(_02743_ ), .B(_02744_ ), .S(fanout_net_39 ), .Z(_05034_ ) );
OAI221_X1 _12761_ ( .A(_04284_ ), .B1(_05032_ ), .B2(_05033_ ), .C1(_05034_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_05035_ ) );
MUX2_X1 _12762_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_39 ), .Z(_05036_ ) );
MUX2_X1 _12763_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_39 ), .Z(_05037_ ) );
MUX2_X1 _12764_ ( .A(_05036_ ), .B(_05037_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_05038_ ) );
OAI211_X1 _12765_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05035_ ), .C1(_05038_ ), .C2(_04691_ ), .ZN(_05039_ ) );
OAI211_X1 _12766_ ( .A(_05031_ ), .B(_05039_ ), .C1(_04703_ ), .C2(_04271_ ), .ZN(_05040_ ) );
NAND2_X1 _12767_ ( .A1(_05022_ ), .A2(_05040_ ), .ZN(_05041_ ) );
XNOR2_X1 _12768_ ( .A(_05041_ ), .B(_02752_ ), .ZN(_05042_ ) );
AND2_X1 _12769_ ( .A1(_05021_ ), .A2(_05042_ ), .ZN(_05043_ ) );
AND2_X2 _12770_ ( .A1(_02726_ ), .A2(_02727_ ), .ZN(_05044_ ) );
OR2_X1 _12771_ ( .A1(_04276_ ), .A2(\myreg.Reg[5][0] ), .ZN(_05045_ ) );
OAI211_X1 _12772_ ( .A(_05045_ ), .B(_04288_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[4][0] ), .ZN(_05046_ ) );
OR2_X1 _12773_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[6][0] ), .ZN(_05047_ ) );
OAI211_X1 _12774_ ( .A(_05047_ ), .B(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_04788_ ), .C2(\myreg.Reg[7][0] ), .ZN(_05048_ ) );
NAND3_X1 _12775_ ( .A1(_05046_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_05048_ ), .ZN(_05049_ ) );
MUX2_X1 _12776_ ( .A(\myreg.Reg[2][0] ), .B(\myreg.Reg[3][0] ), .S(fanout_net_39 ), .Z(_05050_ ) );
MUX2_X1 _12777_ ( .A(\myreg.Reg[0][0] ), .B(\myreg.Reg[1][0] ), .S(fanout_net_39 ), .Z(_05051_ ) );
MUX2_X1 _12778_ ( .A(_05050_ ), .B(_05051_ ), .S(_04287_ ), .Z(_05052_ ) );
OAI211_X1 _12779_ ( .A(_04274_ ), .B(_05049_ ), .C1(_05052_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05053_ ) );
NOR2_X1 _12780_ ( .A1(_04276_ ), .A2(\myreg.Reg[11][0] ), .ZN(_05054_ ) );
OAI21_X1 _12781_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(fanout_net_39 ), .B2(\myreg.Reg[10][0] ), .ZN(_05055_ ) );
NOR2_X1 _12782_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[8][0] ), .ZN(_05056_ ) );
OAI21_X1 _12783_ ( .A(_04287_ ), .B1(_04788_ ), .B2(\myreg.Reg[9][0] ), .ZN(_05057_ ) );
OAI221_X1 _12784_ ( .A(_04282_ ), .B1(_05054_ ), .B2(_05055_ ), .C1(_05056_ ), .C2(_05057_ ), .ZN(_05058_ ) );
MUX2_X1 _12785_ ( .A(\myreg.Reg[12][0] ), .B(\myreg.Reg[13][0] ), .S(fanout_net_39 ), .Z(_05059_ ) );
MUX2_X1 _12786_ ( .A(\myreg.Reg[14][0] ), .B(\myreg.Reg[15][0] ), .S(fanout_net_39 ), .Z(_05060_ ) );
MUX2_X1 _12787_ ( .A(_05059_ ), .B(_05060_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_05061_ ) );
OAI211_X1 _12788_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05058_ ), .C1(_05061_ ), .C2(_04283_ ), .ZN(_05062_ ) );
AOI21_X1 _12789_ ( .A(_04585_ ), .B1(_05053_ ), .B2(_05062_ ), .ZN(_05063_ ) );
AND2_X1 _12790_ ( .A1(_04585_ ), .A2(\EX_LS_result_reg [0] ), .ZN(_05064_ ) );
NOR2_X1 _12791_ ( .A1(_05063_ ), .A2(_05064_ ), .ZN(_05065_ ) );
NOR2_X1 _12792_ ( .A1(_05044_ ), .A2(_05065_ ), .ZN(_05066_ ) );
INV_X1 _12793_ ( .A(_05066_ ), .ZN(_05067_ ) );
NAND2_X1 _12794_ ( .A1(_05044_ ), .A2(_05065_ ), .ZN(_05068_ ) );
AND4_X1 _12795_ ( .A1(_04998_ ), .A2(_05043_ ), .A3(_05067_ ), .A4(_05068_ ), .ZN(_05069_ ) );
AND3_X1 _12796_ ( .A1(_04882_ ), .A2(_04975_ ), .A3(_05069_ ), .ZN(_05070_ ) );
NOR2_X1 _12797_ ( .A1(_04019_ ), .A2(\ID_EX_typ [1] ), .ZN(_05071_ ) );
AND2_X1 _12798_ ( .A1(_05071_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05072_ ) );
BUF_X4 _12799_ ( .A(_05072_ ), .Z(_05073_ ) );
INV_X1 _12800_ ( .A(_05073_ ), .ZN(_05074_ ) );
INV_X2 _12801_ ( .A(fanout_net_8 ), .ZN(_05075_ ) );
BUF_X4 _12802_ ( .A(_05075_ ), .Z(_05076_ ) );
BUF_X2 _12803_ ( .A(_05076_ ), .Z(_05077_ ) );
NAND3_X1 _12804_ ( .A1(_04561_ ), .A2(_05077_ ), .A3(_04580_ ), .ZN(_05078_ ) );
NAND2_X1 _12805_ ( .A1(fanout_net_8 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05079_ ) );
AND2_X2 _12806_ ( .A1(_05078_ ), .A2(_05079_ ), .ZN(_05080_ ) );
XNOR2_X1 _12807_ ( .A(_05080_ ), .B(_02297_ ), .ZN(_05081_ ) );
NAND3_X1 _12808_ ( .A1(_04539_ ), .A2(_05077_ ), .A3(_04558_ ), .ZN(_05082_ ) );
OR2_X1 _12809_ ( .A1(_05077_ ), .A2(\ID_EX_imm [31] ), .ZN(_05083_ ) );
NAND2_X1 _12810_ ( .A1(_05082_ ), .A2(_05083_ ), .ZN(_05084_ ) );
INV_X1 _12811_ ( .A(_03150_ ), .ZN(_05085_ ) );
NAND2_X1 _12812_ ( .A1(_05084_ ), .A2(_05085_ ), .ZN(_05086_ ) );
NAND3_X1 _12813_ ( .A1(_05082_ ), .A2(_03150_ ), .A3(_05083_ ), .ZN(_05087_ ) );
NAND2_X1 _12814_ ( .A1(_05086_ ), .A2(_05087_ ), .ZN(_05088_ ) );
INV_X1 _12815_ ( .A(_05088_ ), .ZN(_05089_ ) );
NOR2_X1 _12816_ ( .A1(_05081_ ), .A2(_05089_ ), .ZN(_05090_ ) );
NAND3_X1 _12817_ ( .A1(_04516_ ), .A2(_05077_ ), .A3(_04535_ ), .ZN(_05091_ ) );
NAND2_X1 _12818_ ( .A1(fanout_net_8 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05092_ ) );
AND2_X2 _12819_ ( .A1(_05091_ ), .A2(_05092_ ), .ZN(_05093_ ) );
INV_X1 _12820_ ( .A(_03118_ ), .ZN(_05094_ ) );
XNOR2_X1 _12821_ ( .A(_05093_ ), .B(_05094_ ), .ZN(_05095_ ) );
INV_X1 _12822_ ( .A(_05095_ ), .ZN(_05096_ ) );
NAND3_X1 _12823_ ( .A1(_04494_ ), .A2(_05077_ ), .A3(_04513_ ), .ZN(_05097_ ) );
NAND2_X1 _12824_ ( .A1(fanout_net_8 ), .A2(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05098_ ) );
AND2_X2 _12825_ ( .A1(_05097_ ), .A2(_05098_ ), .ZN(_05099_ ) );
INV_X1 _12826_ ( .A(_03095_ ), .ZN(_05100_ ) );
XNOR2_X1 _12827_ ( .A(_05099_ ), .B(_05100_ ), .ZN(_05101_ ) );
INV_X1 _12828_ ( .A(_05101_ ), .ZN(_05102_ ) );
AND3_X1 _12829_ ( .A1(_05090_ ), .A2(_05096_ ), .A3(_05102_ ), .ZN(_05103_ ) );
BUF_X4 _12830_ ( .A(_05075_ ), .Z(_05104_ ) );
NAND3_X1 _12831_ ( .A1(_04709_ ), .A2(_04730_ ), .A3(_05104_ ), .ZN(_05105_ ) );
NAND2_X1 _12832_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [14] ), .ZN(_05106_ ) );
AND2_X2 _12833_ ( .A1(_05105_ ), .A2(_05106_ ), .ZN(_05107_ ) );
XNOR2_X1 _12834_ ( .A(_05107_ ), .B(_02838_ ), .ZN(_05108_ ) );
NAND3_X1 _12835_ ( .A1(_04679_ ), .A2(_05104_ ), .A3(_04705_ ), .ZN(_05109_ ) );
NAND2_X1 _12836_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [15] ), .ZN(_05110_ ) );
AND2_X1 _12837_ ( .A1(_05109_ ), .A2(_05110_ ), .ZN(_05111_ ) );
XNOR2_X1 _12838_ ( .A(_05111_ ), .B(_02815_ ), .ZN(_05112_ ) );
NOR2_X1 _12839_ ( .A1(_05108_ ), .A2(_05112_ ), .ZN(_05113_ ) );
NAND3_X1 _12840_ ( .A1(_04760_ ), .A2(_05104_ ), .A3(_04779_ ), .ZN(_05114_ ) );
NAND2_X1 _12841_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [13] ), .ZN(_05115_ ) );
AND2_X2 _12842_ ( .A1(_05114_ ), .A2(_05115_ ), .ZN(_05116_ ) );
XNOR2_X1 _12843_ ( .A(_05116_ ), .B(_04758_ ), .ZN(_05117_ ) );
INV_X1 _12844_ ( .A(_05117_ ), .ZN(_05118_ ) );
NAND2_X1 _12845_ ( .A1(_04756_ ), .A2(_05104_ ), .ZN(_05119_ ) );
OR2_X1 _12846_ ( .A1(_05075_ ), .A2(\ID_EX_imm [12] ), .ZN(_05120_ ) );
NAND2_X1 _12847_ ( .A1(_05119_ ), .A2(_05120_ ), .ZN(_05121_ ) );
XNOR2_X1 _12848_ ( .A(_05121_ ), .B(_02886_ ), .ZN(_05122_ ) );
INV_X1 _12849_ ( .A(_05122_ ), .ZN(_05123_ ) );
AND3_X1 _12850_ ( .A1(_05113_ ), .A2(_05118_ ), .A3(_05123_ ), .ZN(_05124_ ) );
NAND3_X1 _12851_ ( .A1(_04809_ ), .A2(_04828_ ), .A3(_05104_ ), .ZN(_05125_ ) );
NAND2_X1 _12852_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [10] ), .ZN(_05126_ ) );
AND2_X2 _12853_ ( .A1(_05125_ ), .A2(_05126_ ), .ZN(_05127_ ) );
XNOR2_X1 _12854_ ( .A(_05127_ ), .B(_02571_ ), .ZN(_05128_ ) );
NAND3_X1 _12855_ ( .A1(_04785_ ), .A2(_05075_ ), .A3(_04805_ ), .ZN(_05129_ ) );
NAND2_X1 _12856_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [11] ), .ZN(_05130_ ) );
AND2_X1 _12857_ ( .A1(_05129_ ), .A2(_05130_ ), .ZN(_05131_ ) );
XNOR2_X1 _12858_ ( .A(_05131_ ), .B(_04783_ ), .ZN(_05132_ ) );
NOR2_X1 _12859_ ( .A1(_05128_ ), .A2(_05132_ ), .ZN(_05133_ ) );
NAND2_X1 _12860_ ( .A1(_04854_ ), .A2(_05104_ ), .ZN(_05134_ ) );
OR2_X1 _12861_ ( .A1(_05075_ ), .A2(\ID_EX_imm [9] ), .ZN(_05135_ ) );
NAND2_X2 _12862_ ( .A1(_05134_ ), .A2(_05135_ ), .ZN(_05136_ ) );
XNOR2_X1 _12863_ ( .A(_05136_ ), .B(_04832_ ), .ZN(_05137_ ) );
INV_X1 _12864_ ( .A(_05137_ ), .ZN(_05138_ ) );
NAND3_X1 _12865_ ( .A1(_04857_ ), .A2(_04876_ ), .A3(_05104_ ), .ZN(_05139_ ) );
NAND2_X1 _12866_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [8] ), .ZN(_05140_ ) );
AND2_X1 _12867_ ( .A1(_05139_ ), .A2(_05140_ ), .ZN(_05141_ ) );
XNOR2_X1 _12868_ ( .A(_05141_ ), .B(_02498_ ), .ZN(_05142_ ) );
INV_X1 _12869_ ( .A(_05142_ ), .ZN(_05143_ ) );
NAND4_X1 _12870_ ( .A1(_05124_ ), .A2(_05133_ ), .A3(_05138_ ), .A4(_05143_ ), .ZN(_05144_ ) );
NAND3_X1 _12871_ ( .A1(_05022_ ), .A2(_05104_ ), .A3(_05040_ ), .ZN(_05145_ ) );
NAND2_X1 _12872_ ( .A1(fanout_net_8 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_05146_ ) );
AND2_X2 _12873_ ( .A1(_05145_ ), .A2(_05146_ ), .ZN(_05147_ ) );
XNOR2_X1 _12874_ ( .A(_05147_ ), .B(_02781_ ), .ZN(_05148_ ) );
NAND3_X1 _12875_ ( .A1(_05000_ ), .A2(_05019_ ), .A3(_05104_ ), .ZN(_05149_ ) );
NAND2_X1 _12876_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [2] ), .ZN(_05150_ ) );
AND2_X4 _12877_ ( .A1(_05149_ ), .A2(_05150_ ), .ZN(_05151_ ) );
XNOR2_X1 _12878_ ( .A(_05151_ ), .B(_02774_ ), .ZN(_05152_ ) );
NAND2_X1 _12879_ ( .A1(_04997_ ), .A2(_05075_ ), .ZN(_05153_ ) );
NAND2_X1 _12880_ ( .A1(_02705_ ), .A2(fanout_net_8 ), .ZN(_05154_ ) );
NAND2_X1 _12881_ ( .A1(_05153_ ), .A2(_05154_ ), .ZN(_05155_ ) );
BUF_X2 _12882_ ( .A(_05155_ ), .Z(_05156_ ) );
XNOR2_X1 _12883_ ( .A(_05156_ ), .B(_02704_ ), .ZN(_05157_ ) );
INV_X1 _12884_ ( .A(_05044_ ), .ZN(_05158_ ) );
NAND2_X4 _12885_ ( .A1(_05065_ ), .A2(_05075_ ), .ZN(_05159_ ) );
OR2_X2 _12886_ ( .A1(_05075_ ), .A2(\ID_EX_imm [0] ), .ZN(_05160_ ) );
AND3_X1 _12887_ ( .A1(_05158_ ), .A2(_05159_ ), .A3(_05160_ ), .ZN(_05161_ ) );
OR2_X1 _12888_ ( .A1(_05157_ ), .A2(_05161_ ), .ZN(_05162_ ) );
NAND2_X1 _12889_ ( .A1(_05156_ ), .A2(_02704_ ), .ZN(_05163_ ) );
AOI211_X1 _12890_ ( .A(_05148_ ), .B(_05152_ ), .C1(_05162_ ), .C2(_05163_ ), .ZN(_05164_ ) );
AOI21_X1 _12891_ ( .A(_02781_ ), .B1(_05146_ ), .B2(_05145_ ), .ZN(_05165_ ) );
INV_X1 _12892_ ( .A(_05151_ ), .ZN(_05166_ ) );
NOR3_X1 _12893_ ( .A1(_05148_ ), .A2(_04999_ ), .A3(_05166_ ), .ZN(_05167_ ) );
OR3_X1 _12894_ ( .A1(_05164_ ), .A2(_05165_ ), .A3(_05167_ ), .ZN(_05168_ ) );
NAND2_X1 _12895_ ( .A1(_04973_ ), .A2(_05076_ ), .ZN(_05169_ ) );
NAND2_X1 _12896_ ( .A1(_02625_ ), .A2(fanout_net_8 ), .ZN(_05170_ ) );
NAND2_X2 _12897_ ( .A1(_05169_ ), .A2(_05170_ ), .ZN(_05171_ ) );
INV_X1 _12898_ ( .A(_02598_ ), .ZN(_05172_ ) );
XNOR2_X1 _12899_ ( .A(_05171_ ), .B(_05172_ ), .ZN(_05173_ ) );
NAND3_X1 _12900_ ( .A1(_04908_ ), .A2(_05075_ ), .A3(_04927_ ), .ZN(_05174_ ) );
NAND2_X1 _12901_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [7] ), .ZN(_05175_ ) );
AND2_X1 _12902_ ( .A1(_05174_ ), .A2(_05175_ ), .ZN(_05176_ ) );
XNOR2_X1 _12903_ ( .A(_05176_ ), .B(_04906_ ), .ZN(_05177_ ) );
NAND3_X1 _12904_ ( .A1(_04884_ ), .A2(_04903_ ), .A3(_05075_ ), .ZN(_05178_ ) );
NAND2_X1 _12905_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [6] ), .ZN(_05179_ ) );
AND2_X1 _12906_ ( .A1(_05178_ ), .A2(_05179_ ), .ZN(_05180_ ) );
BUF_X2 _12907_ ( .A(_05180_ ), .Z(_05181_ ) );
XNOR2_X1 _12908_ ( .A(_05181_ ), .B(_02670_ ), .ZN(_05182_ ) );
NAND3_X1 _12909_ ( .A1(_04931_ ), .A2(_05104_ ), .A3(_04950_ ), .ZN(_05183_ ) );
NAND2_X1 _12910_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [4] ), .ZN(_05184_ ) );
AND2_X2 _12911_ ( .A1(_05183_ ), .A2(_05184_ ), .ZN(_05185_ ) );
BUF_X4 _12912_ ( .A(_05185_ ), .Z(_05186_ ) );
XNOR2_X2 _12913_ ( .A(_05186_ ), .B(_02622_ ), .ZN(_05187_ ) );
NOR4_X1 _12914_ ( .A1(_05173_ ), .A2(_05177_ ), .A3(_05182_ ), .A4(_05187_ ), .ZN(_05188_ ) );
NAND2_X1 _12915_ ( .A1(_05168_ ), .A2(_05188_ ), .ZN(_05189_ ) );
INV_X1 _12916_ ( .A(_05177_ ), .ZN(_05190_ ) );
INV_X1 _12917_ ( .A(_05182_ ), .ZN(_05191_ ) );
INV_X1 _12918_ ( .A(_05186_ ), .ZN(_05192_ ) );
NOR3_X1 _12919_ ( .A1(_05173_ ), .A2(_02623_ ), .A3(_05192_ ), .ZN(_05193_ ) );
AND3_X1 _12920_ ( .A1(_05169_ ), .A2(_02598_ ), .A3(_05170_ ), .ZN(_05194_ ) );
OAI211_X1 _12921_ ( .A(_05190_ ), .B(_05191_ ), .C1(_05193_ ), .C2(_05194_ ), .ZN(_05195_ ) );
NAND3_X1 _12922_ ( .A1(_05174_ ), .A2(_04906_ ), .A3(_05175_ ), .ZN(_05196_ ) );
NAND3_X1 _12923_ ( .A1(_05190_ ), .A2(_02670_ ), .A3(_05181_ ), .ZN(_05197_ ) );
AND3_X1 _12924_ ( .A1(_05195_ ), .A2(_05196_ ), .A3(_05197_ ), .ZN(_05198_ ) );
AOI21_X1 _12925_ ( .A(_05144_ ), .B1(_05189_ ), .B2(_05198_ ), .ZN(_05199_ ) );
INV_X1 _12926_ ( .A(_05107_ ), .ZN(_05200_ ) );
NOR3_X1 _12927_ ( .A1(_05112_ ), .A2(_04708_ ), .A3(_05200_ ), .ZN(_05201_ ) );
INV_X1 _12928_ ( .A(_05141_ ), .ZN(_05202_ ) );
NOR3_X1 _12929_ ( .A1(_05137_ ), .A2(_04856_ ), .A3(_05202_ ), .ZN(_05203_ ) );
AOI21_X1 _12930_ ( .A(_05203_ ), .B1(_04832_ ), .B2(_05136_ ), .ZN(_05204_ ) );
INV_X1 _12931_ ( .A(_05133_ ), .ZN(_05205_ ) );
INV_X1 _12932_ ( .A(_05131_ ), .ZN(_05206_ ) );
OAI22_X1 _12933_ ( .A1(_05204_ ), .A2(_05205_ ), .B1(_04784_ ), .B2(_05206_ ), .ZN(_05207_ ) );
INV_X1 _12934_ ( .A(_05127_ ), .ZN(_05208_ ) );
NOR3_X1 _12935_ ( .A1(_05132_ ), .A2(_04808_ ), .A3(_05208_ ), .ZN(_05209_ ) );
OAI21_X1 _12936_ ( .A(_05124_ ), .B1(_05207_ ), .B2(_05209_ ), .ZN(_05210_ ) );
AND3_X1 _12937_ ( .A1(_05118_ ), .A2(_02886_ ), .A3(_05121_ ), .ZN(_05211_ ) );
AND3_X1 _12938_ ( .A1(_04758_ ), .A2(_05115_ ), .A3(_05114_ ), .ZN(_05212_ ) );
OAI21_X1 _12939_ ( .A(_05113_ ), .B1(_05211_ ), .B2(_05212_ ), .ZN(_05213_ ) );
INV_X1 _12940_ ( .A(_05111_ ), .ZN(_05214_ ) );
OAI211_X1 _12941_ ( .A(_05210_ ), .B(_05213_ ), .C1(_04678_ ), .C2(_05214_ ), .ZN(_05215_ ) );
OR3_X1 _12942_ ( .A1(_05199_ ), .A2(_05201_ ), .A3(_05215_ ), .ZN(_05216_ ) );
NAND3_X1 _12943_ ( .A1(_04373_ ), .A2(_05076_ ), .A3(_04392_ ), .ZN(_05217_ ) );
NAND2_X1 _12944_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [17] ), .ZN(_05218_ ) );
AND2_X2 _12945_ ( .A1(_05217_ ), .A2(_05218_ ), .ZN(_05219_ ) );
XNOR2_X1 _12946_ ( .A(_05219_ ), .B(_02965_ ), .ZN(_05220_ ) );
INV_X1 _12947_ ( .A(_05220_ ), .ZN(_05221_ ) );
NAND3_X1 _12948_ ( .A1(_04368_ ), .A2(_04369_ ), .A3(_05076_ ), .ZN(_05222_ ) );
NAND2_X1 _12949_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [16] ), .ZN(_05223_ ) );
AND2_X1 _12950_ ( .A1(_05222_ ), .A2(_05223_ ), .ZN(_05224_ ) );
XNOR2_X1 _12951_ ( .A(_05224_ ), .B(_02472_ ), .ZN(_05225_ ) );
INV_X1 _12952_ ( .A(_05225_ ), .ZN(_05226_ ) );
NAND3_X1 _12953_ ( .A1(_04421_ ), .A2(_05076_ ), .A3(_04440_ ), .ZN(_05227_ ) );
NAND2_X1 _12954_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [23] ), .ZN(_05228_ ) );
AND2_X1 _12955_ ( .A1(_05227_ ), .A2(_05228_ ), .ZN(_05229_ ) );
XNOR2_X1 _12956_ ( .A(_05229_ ), .B(_02396_ ), .ZN(_05230_ ) );
NAND3_X1 _12957_ ( .A1(_04397_ ), .A2(_04417_ ), .A3(_05076_ ), .ZN(_05231_ ) );
NAND2_X1 _12958_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [22] ), .ZN(_05232_ ) );
NAND2_X1 _12959_ ( .A1(_05231_ ), .A2(_05232_ ), .ZN(_05233_ ) );
XNOR2_X1 _12960_ ( .A(_05233_ ), .B(_04396_ ), .ZN(_05234_ ) );
NOR2_X1 _12961_ ( .A1(_05230_ ), .A2(_05234_ ), .ZN(_05235_ ) );
NAND3_X1 _12962_ ( .A1(_04445_ ), .A2(_04465_ ), .A3(_05076_ ), .ZN(_05236_ ) );
NAND2_X1 _12963_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [20] ), .ZN(_05237_ ) );
AND2_X2 _12964_ ( .A1(_05236_ ), .A2(_05237_ ), .ZN(_05238_ ) );
XNOR2_X1 _12965_ ( .A(_05238_ ), .B(_02422_ ), .ZN(_05239_ ) );
NAND3_X1 _12966_ ( .A1(_04470_ ), .A2(_05076_ ), .A3(_04489_ ), .ZN(_05240_ ) );
NAND2_X1 _12967_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [21] ), .ZN(_05241_ ) );
AND2_X1 _12968_ ( .A1(_05240_ ), .A2(_05241_ ), .ZN(_05242_ ) );
XNOR2_X1 _12969_ ( .A(_05242_ ), .B(_04468_ ), .ZN(_05243_ ) );
NOR2_X1 _12970_ ( .A1(_05239_ ), .A2(_05243_ ), .ZN(_05244_ ) );
NAND3_X1 _12971_ ( .A1(_04336_ ), .A2(_04337_ ), .A3(_05076_ ), .ZN(_05245_ ) );
NAND2_X1 _12972_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [18] ), .ZN(_05246_ ) );
AND2_X1 _12973_ ( .A1(_05245_ ), .A2(_05246_ ), .ZN(_05247_ ) );
XNOR2_X1 _12974_ ( .A(_05247_ ), .B(_02917_ ), .ZN(_05248_ ) );
INV_X1 _12975_ ( .A(_05248_ ), .ZN(_05249_ ) );
NAND3_X1 _12976_ ( .A1(_04273_ ), .A2(_05076_ ), .A3(_04311_ ), .ZN(_05250_ ) );
NAND2_X1 _12977_ ( .A1(fanout_net_8 ), .A2(\ID_EX_imm [19] ), .ZN(_05251_ ) );
AND2_X1 _12978_ ( .A1(_05250_ ), .A2(_05251_ ), .ZN(_05252_ ) );
XNOR2_X1 _12979_ ( .A(_05252_ ), .B(_02940_ ), .ZN(_05253_ ) );
INV_X1 _12980_ ( .A(_05253_ ), .ZN(_05254_ ) );
AND4_X1 _12981_ ( .A1(_05235_ ), .A2(_05244_ ), .A3(_05249_ ), .A4(_05254_ ), .ZN(_05255_ ) );
AND4_X1 _12982_ ( .A1(_05216_ ), .A2(_05221_ ), .A3(_05226_ ), .A4(_05255_ ), .ZN(_05256_ ) );
NOR3_X1 _12983_ ( .A1(_05230_ ), .A2(_04396_ ), .A3(_05233_ ), .ZN(_05257_ ) );
AND2_X1 _12984_ ( .A1(_05219_ ), .A2(_04372_ ), .ZN(_05258_ ) );
NOR2_X1 _12985_ ( .A1(_05219_ ), .A2(_04372_ ), .ZN(_05259_ ) );
OAI211_X1 _12986_ ( .A(_02472_ ), .B(_05224_ ), .C1(_05258_ ), .C2(_05259_ ), .ZN(_05260_ ) );
INV_X1 _12987_ ( .A(_05219_ ), .ZN(_05261_ ) );
OAI21_X1 _12988_ ( .A(_05260_ ), .B1(_04372_ ), .B2(_05261_ ), .ZN(_05262_ ) );
NAND3_X1 _12989_ ( .A1(_05262_ ), .A2(_05254_ ), .A3(_05249_ ), .ZN(_05263_ ) );
NAND3_X1 _12990_ ( .A1(_05254_ ), .A2(_02917_ ), .A3(_05247_ ), .ZN(_05264_ ) );
NAND3_X1 _12991_ ( .A1(_05250_ ), .A2(_02940_ ), .A3(_05251_ ), .ZN(_05265_ ) );
NAND3_X1 _12992_ ( .A1(_05263_ ), .A2(_05264_ ), .A3(_05265_ ), .ZN(_05266_ ) );
AND3_X1 _12993_ ( .A1(_05266_ ), .A2(_05235_ ), .A3(_05244_ ), .ZN(_05267_ ) );
INV_X1 _12994_ ( .A(_05243_ ), .ZN(_05268_ ) );
AND3_X1 _12995_ ( .A1(_05268_ ), .A2(_02422_ ), .A3(_05238_ ), .ZN(_05269_ ) );
AND3_X1 _12996_ ( .A1(_04468_ ), .A2(_05241_ ), .A3(_05240_ ), .ZN(_05270_ ) );
OAI21_X1 _12997_ ( .A(_05235_ ), .B1(_05269_ ), .B2(_05270_ ), .ZN(_05271_ ) );
INV_X1 _12998_ ( .A(_05229_ ), .ZN(_05272_ ) );
OAI21_X1 _12999_ ( .A(_05271_ ), .B1(_04420_ ), .B2(_05272_ ), .ZN(_05273_ ) );
NOR4_X1 _13000_ ( .A1(_05256_ ), .A2(_05257_ ), .A3(_05267_ ), .A4(_05273_ ), .ZN(_05274_ ) );
NAND3_X1 _13001_ ( .A1(_04608_ ), .A2(_05077_ ), .A3(_04627_ ), .ZN(_05275_ ) );
NAND2_X1 _13002_ ( .A1(_02349_ ), .A2(fanout_net_8 ), .ZN(_05276_ ) );
NAND2_X1 _13003_ ( .A1(_05275_ ), .A2(_05276_ ), .ZN(_05277_ ) );
XNOR2_X1 _13004_ ( .A(_05277_ ), .B(_02348_ ), .ZN(_05278_ ) );
NAND3_X1 _13005_ ( .A1(_04586_ ), .A2(_05077_ ), .A3(_04604_ ), .ZN(_05279_ ) );
NAND2_X1 _13006_ ( .A1(_03064_ ), .A2(fanout_net_8 ), .ZN(_05280_ ) );
NAND2_X1 _13007_ ( .A1(_05279_ ), .A2(_05280_ ), .ZN(_05281_ ) );
INV_X1 _13008_ ( .A(_03063_ ), .ZN(_05282_ ) );
NOR2_X1 _13009_ ( .A1(_05281_ ), .A2(_05282_ ), .ZN(_05283_ ) );
AOI21_X1 _13010_ ( .A(_03063_ ), .B1(_05279_ ), .B2(_05280_ ), .ZN(_05284_ ) );
NOR2_X1 _13011_ ( .A1(_05283_ ), .A2(_05284_ ), .ZN(_05285_ ) );
NOR2_X1 _13012_ ( .A1(_05278_ ), .A2(_05285_ ), .ZN(_05286_ ) );
INV_X1 _13013_ ( .A(_05286_ ), .ZN(_05287_ ) );
OAI21_X1 _13014_ ( .A(_05077_ ), .B1(_04672_ ), .B2(_04673_ ), .ZN(_05288_ ) );
NAND2_X1 _13015_ ( .A1(_03197_ ), .A2(fanout_net_8 ), .ZN(_05289_ ) );
NAND2_X1 _13016_ ( .A1(_05288_ ), .A2(_05289_ ), .ZN(_05290_ ) );
INV_X1 _13017_ ( .A(_03196_ ), .ZN(_05291_ ) );
NOR2_X1 _13018_ ( .A1(_05290_ ), .A2(_05291_ ), .ZN(_05292_ ) );
AOI21_X1 _13019_ ( .A(_03196_ ), .B1(_05288_ ), .B2(_05289_ ), .ZN(_05293_ ) );
NOR2_X1 _13020_ ( .A1(_05292_ ), .A2(_05293_ ), .ZN(_05294_ ) );
NAND3_X1 _13021_ ( .A1(_04632_ ), .A2(_05077_ ), .A3(_04651_ ), .ZN(_05295_ ) );
NAND2_X1 _13022_ ( .A1(_03016_ ), .A2(fanout_net_8 ), .ZN(_05296_ ) );
NAND2_X1 _13023_ ( .A1(_05295_ ), .A2(_05296_ ), .ZN(_05297_ ) );
NOR2_X1 _13024_ ( .A1(_05297_ ), .A2(_03040_ ), .ZN(_05298_ ) );
AOI21_X1 _13025_ ( .A(_03039_ ), .B1(_05295_ ), .B2(_05296_ ), .ZN(_05299_ ) );
NOR2_X1 _13026_ ( .A1(_05298_ ), .A2(_05299_ ), .ZN(_05300_ ) );
NOR4_X1 _13027_ ( .A1(_05274_ ), .A2(_05287_ ), .A3(_05294_ ), .A4(_05300_ ), .ZN(_05301_ ) );
OAI211_X1 _13028_ ( .A(_05290_ ), .B(_03196_ ), .C1(_05298_ ), .C2(_05299_ ), .ZN(_05302_ ) );
NAND2_X1 _13029_ ( .A1(_05297_ ), .A2(_03039_ ), .ZN(_05303_ ) );
AOI21_X1 _13030_ ( .A(_05287_ ), .B1(_05302_ ), .B2(_05303_ ), .ZN(_05304_ ) );
INV_X1 _13031_ ( .A(_05278_ ), .ZN(_05305_ ) );
AND3_X1 _13032_ ( .A1(_05305_ ), .A2(_03063_ ), .A3(_05281_ ), .ZN(_05306_ ) );
INV_X1 _13033_ ( .A(_02348_ ), .ZN(_05307_ ) );
AOI21_X1 _13034_ ( .A(_05307_ ), .B1(_05275_ ), .B2(_05276_ ), .ZN(_05308_ ) );
OR3_X1 _13035_ ( .A1(_05304_ ), .A2(_05306_ ), .A3(_05308_ ), .ZN(_05309_ ) );
OAI21_X1 _13036_ ( .A(_05103_ ), .B1(_05301_ ), .B2(_05309_ ), .ZN(_05310_ ) );
NOR2_X1 _13037_ ( .A1(_05080_ ), .A2(_02297_ ), .ZN(_05311_ ) );
AND2_X1 _13038_ ( .A1(_05088_ ), .A2(_05311_ ), .ZN(_05312_ ) );
INV_X1 _13039_ ( .A(_05084_ ), .ZN(_05313_ ) );
INV_X1 _13040_ ( .A(_05099_ ), .ZN(_05314_ ) );
NAND3_X1 _13041_ ( .A1(_05096_ ), .A2(_03095_ ), .A3(_05314_ ), .ZN(_05315_ ) );
OAI21_X1 _13042_ ( .A(_05315_ ), .B1(_05094_ ), .B2(_05093_ ), .ZN(_05316_ ) );
AOI221_X4 _13043_ ( .A(_05312_ ), .B1(_05085_ ), .B2(_05313_ ), .C1(_05316_ ), .C2(_05090_ ), .ZN(_05317_ ) );
AND2_X1 _13044_ ( .A1(_05310_ ), .A2(_05317_ ), .ZN(_05318_ ) );
INV_X1 _13045_ ( .A(\ID_EX_typ [1] ), .ZN(_05319_ ) );
NOR2_X1 _13046_ ( .A1(_05319_ ), .A2(fanout_net_7 ), .ZN(_05320_ ) );
INV_X1 _13047_ ( .A(\ID_EX_typ [2] ), .ZN(_05321_ ) );
AND2_X1 _13048_ ( .A1(_05320_ ), .A2(_05321_ ), .ZN(_05322_ ) );
BUF_X4 _13049_ ( .A(_05322_ ), .Z(_05323_ ) );
INV_X1 _13050_ ( .A(_05323_ ), .ZN(_05324_ ) );
OAI21_X2 _13051_ ( .A(_05074_ ), .B1(_05318_ ), .B2(_05324_ ), .ZN(_05325_ ) );
BUF_X4 _13052_ ( .A(_05321_ ), .Z(_05326_ ) );
NOR3_X1 _13053_ ( .A1(_05326_ ), .A2(\ID_EX_typ [1] ), .A3(fanout_net_7 ), .ZN(_05327_ ) );
NAND3_X1 _13054_ ( .A1(_05310_ ), .A2(_05317_ ), .A3(_05327_ ), .ZN(_05328_ ) );
AND2_X1 _13055_ ( .A1(\ID_EX_typ [1] ), .A2(fanout_net_7 ), .ZN(_05329_ ) );
AND2_X2 _13056_ ( .A1(_05329_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05330_ ) );
INV_X1 _13057_ ( .A(_05330_ ), .ZN(_05331_ ) );
AND2_X2 _13058_ ( .A1(_05071_ ), .A2(\ID_EX_typ [2] ), .ZN(_05332_ ) );
INV_X1 _13059_ ( .A(_05332_ ), .ZN(_05333_ ) );
NAND2_X1 _13060_ ( .A1(_04493_ ), .A2(_04677_ ), .ZN(_05334_ ) );
AND2_X1 _13061_ ( .A1(_04731_ ), .A2(_02838_ ), .ZN(_05335_ ) );
AND2_X1 _13062_ ( .A1(_04707_ ), .A2(_05335_ ), .ZN(_05336_ ) );
AND2_X1 _13063_ ( .A1(_04829_ ), .A2(_02571_ ), .ZN(_05337_ ) );
AND2_X1 _13064_ ( .A1(_04807_ ), .A2(_05337_ ), .ZN(_05338_ ) );
AOI21_X1 _13065_ ( .A(_05338_ ), .B1(_04783_ ), .B2(_04806_ ), .ZN(_05339_ ) );
AND2_X1 _13066_ ( .A1(_04877_ ), .A2(_02498_ ), .ZN(_05340_ ) );
AND2_X1 _13067_ ( .A1(_04855_ ), .A2(_05340_ ), .ZN(_05341_ ) );
AOI21_X1 _13068_ ( .A(_05341_ ), .B1(_04832_ ), .B2(_04854_ ), .ZN(_05342_ ) );
INV_X1 _13069_ ( .A(_04831_ ), .ZN(_05343_ ) );
OAI21_X1 _13070_ ( .A(_05339_ ), .B1(_05342_ ), .B2(_05343_ ), .ZN(_05344_ ) );
NAND2_X1 _13071_ ( .A1(_05344_ ), .A2(_04782_ ), .ZN(_05345_ ) );
NOR2_X1 _13072_ ( .A1(_04780_ ), .A2(_04758_ ), .ZN(_05346_ ) );
AND2_X1 _13073_ ( .A1(_04780_ ), .A2(_04758_ ), .ZN(_05347_ ) );
INV_X1 _13074_ ( .A(_05347_ ), .ZN(_05348_ ) );
NAND2_X1 _13075_ ( .A1(_04756_ ), .A2(_02886_ ), .ZN(_05349_ ) );
AOI21_X1 _13076_ ( .A(_05346_ ), .B1(_05348_ ), .B2(_05349_ ), .ZN(_05350_ ) );
NAND3_X1 _13077_ ( .A1(_05350_ ), .A2(_04707_ ), .A3(_04732_ ), .ZN(_05351_ ) );
NAND2_X1 _13078_ ( .A1(_05345_ ), .A2(_05351_ ), .ZN(_05352_ ) );
AOI211_X1 _13079_ ( .A(_05336_ ), .B(_05352_ ), .C1(_02815_ ), .C2(_04706_ ), .ZN(_05353_ ) );
AND2_X1 _13080_ ( .A1(_05067_ ), .A2(_04998_ ), .ZN(_05354_ ) );
AND2_X1 _13081_ ( .A1(_02704_ ), .A2(_04997_ ), .ZN(_05355_ ) );
OAI21_X1 _13082_ ( .A(_05021_ ), .B1(_05354_ ), .B2(_05355_ ), .ZN(_05356_ ) );
AND2_X1 _13083_ ( .A1(_05020_ ), .A2(_02774_ ), .ZN(_05357_ ) );
INV_X1 _13084_ ( .A(_05357_ ), .ZN(_05358_ ) );
OAI211_X1 _13085_ ( .A(_05356_ ), .B(_05358_ ), .C1(_02781_ ), .C2(_05041_ ), .ZN(_05359_ ) );
NAND3_X1 _13086_ ( .A1(_05041_ ), .A2(_02731_ ), .A3(_02751_ ), .ZN(_05360_ ) );
NAND3_X1 _13087_ ( .A1(_05359_ ), .A2(_05360_ ), .A3(_04975_ ), .ZN(_05361_ ) );
AND3_X1 _13088_ ( .A1(_04929_ ), .A2(_02670_ ), .A3(_04904_ ), .ZN(_05362_ ) );
AND2_X1 _13089_ ( .A1(_02622_ ), .A2(_04951_ ), .ZN(_05363_ ) );
NAND2_X1 _13090_ ( .A1(_04974_ ), .A2(_05363_ ), .ZN(_05364_ ) );
OAI21_X1 _13091_ ( .A(_05364_ ), .B1(_05172_ ), .B2(_04973_ ), .ZN(_05365_ ) );
AOI221_X4 _13092_ ( .A(_05362_ ), .B1(_04906_ ), .B2(_04928_ ), .C1(_05365_ ), .C2(_04930_ ), .ZN(_05366_ ) );
AND2_X1 _13093_ ( .A1(_05361_ ), .A2(_05366_ ), .ZN(_05367_ ) );
INV_X1 _13094_ ( .A(_05367_ ), .ZN(_05368_ ) );
NAND2_X1 _13095_ ( .A1(_05368_ ), .A2(_04881_ ), .ZN(_05369_ ) );
AOI21_X1 _13096_ ( .A(_05334_ ), .B1(_05353_ ), .B2(_05369_ ), .ZN(_05370_ ) );
NOR2_X1 _13097_ ( .A1(_05100_ ), .A2(_04514_ ), .ZN(_05371_ ) );
AND3_X1 _13098_ ( .A1(_03118_ ), .A2(_04516_ ), .A3(_04535_ ), .ZN(_05372_ ) );
NOR2_X1 _13099_ ( .A1(_05371_ ), .A2(_05372_ ), .ZN(_05373_ ) );
AOI21_X1 _13100_ ( .A(_03118_ ), .B1(_04516_ ), .B2(_04535_ ), .ZN(_05374_ ) );
NOR2_X1 _13101_ ( .A1(_05373_ ), .A2(_05374_ ), .ZN(_05375_ ) );
AND3_X1 _13102_ ( .A1(_04583_ ), .A2(_05375_ ), .A3(_04560_ ), .ZN(_05376_ ) );
AND3_X1 _13103_ ( .A1(_04394_ ), .A2(_02472_ ), .A3(_04370_ ), .ZN(_05377_ ) );
AND2_X1 _13104_ ( .A1(_04393_ ), .A2(_02965_ ), .ZN(_05378_ ) );
OAI21_X1 _13105_ ( .A(_04341_ ), .B1(_05377_ ), .B2(_05378_ ), .ZN(_05379_ ) );
AND2_X1 _13106_ ( .A1(_02940_ ), .A2(_04312_ ), .ZN(_05380_ ) );
INV_X1 _13107_ ( .A(_05380_ ), .ZN(_05381_ ) );
NAND3_X1 _13108_ ( .A1(_04313_ ), .A2(_02917_ ), .A3(_04338_ ), .ZN(_05382_ ) );
AND3_X2 _13109_ ( .A1(_05379_ ), .A2(_05381_ ), .A3(_05382_ ), .ZN(_05383_ ) );
INV_X1 _13110_ ( .A(_04492_ ), .ZN(_05384_ ) );
NOR2_X1 _13111_ ( .A1(_05383_ ), .A2(_05384_ ), .ZN(_05385_ ) );
NAND3_X1 _13112_ ( .A1(_04442_ ), .A2(_02373_ ), .A3(_04418_ ), .ZN(_05386_ ) );
INV_X1 _13113_ ( .A(_04441_ ), .ZN(_05387_ ) );
OAI21_X1 _13114_ ( .A(_05386_ ), .B1(_04420_ ), .B2(_05387_ ), .ZN(_05388_ ) );
AND2_X1 _13115_ ( .A1(_04490_ ), .A2(_04468_ ), .ZN(_05389_ ) );
NOR2_X1 _13116_ ( .A1(_04490_ ), .A2(_04468_ ), .ZN(_05390_ ) );
NAND2_X1 _13117_ ( .A1(_04466_ ), .A2(_02422_ ), .ZN(_05391_ ) );
NOR3_X1 _13118_ ( .A1(_05389_ ), .A2(_05390_ ), .A3(_05391_ ), .ZN(_05392_ ) );
OR2_X1 _13119_ ( .A1(_05392_ ), .A2(_05389_ ), .ZN(_05393_ ) );
AND2_X1 _13120_ ( .A1(_05393_ ), .A2(_04443_ ), .ZN(_05394_ ) );
NOR3_X4 _13121_ ( .A1(_05385_ ), .A2(_05388_ ), .A3(_05394_ ), .ZN(_05395_ ) );
INV_X1 _13122_ ( .A(_04677_ ), .ZN(_05396_ ) );
NOR2_X1 _13123_ ( .A1(_05395_ ), .A2(_05396_ ), .ZN(_05397_ ) );
INV_X1 _13124_ ( .A(_04584_ ), .ZN(_05398_ ) );
NOR2_X1 _13125_ ( .A1(_05282_ ), .A2(_04605_ ), .ZN(_05399_ ) );
NAND2_X1 _13126_ ( .A1(_04629_ ), .A2(_05399_ ), .ZN(_05400_ ) );
OAI21_X1 _13127_ ( .A(_05400_ ), .B1(_05307_ ), .B2(_04628_ ), .ZN(_05401_ ) );
AND3_X1 _13128_ ( .A1(_03039_ ), .A2(_04632_ ), .A3(_04651_ ), .ZN(_05402_ ) );
NOR2_X1 _13129_ ( .A1(_04674_ ), .A2(_05291_ ), .ZN(_05403_ ) );
AOI21_X1 _13130_ ( .A(_05402_ ), .B1(_04653_ ), .B2(_05403_ ), .ZN(_05404_ ) );
INV_X1 _13131_ ( .A(_05404_ ), .ZN(_05405_ ) );
AOI21_X1 _13132_ ( .A(_05401_ ), .B1(_04630_ ), .B2(_05405_ ), .ZN(_05406_ ) );
NOR2_X1 _13133_ ( .A1(_05398_ ), .A2(_05406_ ), .ZN(_05407_ ) );
NOR2_X1 _13134_ ( .A1(_02297_ ), .A2(_04581_ ), .ZN(_05408_ ) );
NAND2_X1 _13135_ ( .A1(_05408_ ), .A2(_04560_ ), .ZN(_05409_ ) );
OAI21_X1 _13136_ ( .A(_05409_ ), .B1(_05085_ ), .B2(_04559_ ), .ZN(_05410_ ) );
OR3_X1 _13137_ ( .A1(_05397_ ), .A2(_05407_ ), .A3(_05410_ ), .ZN(_05411_ ) );
NOR3_X1 _13138_ ( .A1(_05370_ ), .A2(_05376_ ), .A3(_05411_ ), .ZN(_05412_ ) );
MUX2_X1 _13139_ ( .A(_05331_ ), .B(_05333_ ), .S(_05412_ ), .Z(_05413_ ) );
NAND2_X1 _13140_ ( .A1(_05328_ ), .A2(_05413_ ), .ZN(_05414_ ) );
OAI221_X2 _13141_ ( .A(_04255_ ), .B1(_05070_ ), .B2(_05074_ ), .C1(_05325_ ), .C2(_05414_ ), .ZN(_05415_ ) );
NAND4_X1 _13142_ ( .A1(_05069_ ), .A2(_04975_ ), .A3(_04782_ ), .A4(_04880_ ), .ZN(_05416_ ) );
OAI21_X1 _13143_ ( .A(_04254_ ), .B1(_05334_ ), .B2(_05416_ ), .ZN(_05417_ ) );
AND2_X4 _13144_ ( .A1(_05415_ ), .A2(_05417_ ), .ZN(_05418_ ) );
BUF_X4 _13145_ ( .A(_05418_ ), .Z(_05419_ ) );
MUX2_X1 _13146_ ( .A(_04130_ ), .B(_04252_ ), .S(_05419_ ), .Z(_05420_ ) );
INV_X1 _13147_ ( .A(\ID_EX_typ [3] ), .ZN(_05421_ ) );
BUF_X4 _13148_ ( .A(_05421_ ), .Z(_05422_ ) );
MUX2_X1 _13149_ ( .A(_04110_ ), .B(_05420_ ), .S(_05422_ ), .Z(_05423_ ) );
INV_X2 _13150_ ( .A(_04018_ ), .ZN(_05424_ ) );
BUF_X4 _13151_ ( .A(_05424_ ), .Z(_05425_ ) );
BUF_X4 _13152_ ( .A(_05425_ ), .Z(_05426_ ) );
NAND2_X1 _13153_ ( .A1(_05423_ ), .A2(_05426_ ), .ZN(_05427_ ) );
BUF_X2 _13154_ ( .A(_04019_ ), .Z(_05428_ ) );
OR2_X1 _13155_ ( .A1(_03156_ ), .A2(_05428_ ), .ZN(_05429_ ) );
BUF_X2 _13156_ ( .A(_04018_ ), .Z(_05430_ ) );
BUF_X4 _13157_ ( .A(_05430_ ), .Z(_05431_ ) );
OAI211_X1 _13158_ ( .A(_05429_ ), .B(_05431_ ), .C1(fanout_net_7 ), .C2(_04252_ ), .ZN(_05432_ ) );
AOI21_X1 _13159_ ( .A(_04032_ ), .B1(_05427_ ), .B2(_05432_ ), .ZN(_00158_ ) );
CLKBUF_X2 _13160_ ( .A(_04018_ ), .Z(_05433_ ) );
INV_X4 _13161_ ( .A(_05418_ ), .ZN(_05434_ ) );
BUF_X4 _13162_ ( .A(_05434_ ), .Z(_05435_ ) );
AND4_X1 _13163_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [15] ), .A4(\ID_EX_pc [14] ), .ZN(_05436_ ) );
AND4_X1 _13164_ ( .A1(\ID_EX_pc [13] ), .A2(_05436_ ), .A3(\ID_EX_pc [12] ), .A4(_04118_ ), .ZN(_05437_ ) );
AND2_X1 _13165_ ( .A1(_04117_ ), .A2(_05437_ ), .ZN(_05438_ ) );
AND4_X1 _13166_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [23] ), .A4(\ID_EX_pc [22] ), .ZN(_05439_ ) );
AND2_X1 _13167_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_05440_ ) );
AND4_X1 _13168_ ( .A1(\ID_EX_pc [21] ), .A2(_05439_ ), .A3(\ID_EX_pc [20] ), .A4(_05440_ ), .ZN(_05441_ ) );
AND2_X1 _13169_ ( .A1(_05438_ ), .A2(_05441_ ), .ZN(_05442_ ) );
NAND3_X1 _13170_ ( .A1(_05442_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_pc [26] ), .ZN(_05443_ ) );
INV_X1 _13171_ ( .A(\ID_EX_pc [28] ), .ZN(_05444_ ) );
NOR2_X1 _13172_ ( .A1(_05443_ ), .A2(_05444_ ), .ZN(_05445_ ) );
XNOR2_X1 _13173_ ( .A(_05445_ ), .B(_04247_ ), .ZN(_05446_ ) );
AOI21_X1 _13174_ ( .A(\ID_EX_typ [3] ), .B1(_05435_ ), .B2(_05446_ ), .ZN(_05447_ ) );
NAND3_X1 _13175_ ( .A1(_04076_ ), .A2(\mepc [29] ), .A3(_04081_ ), .ZN(_05448_ ) );
NAND3_X1 _13176_ ( .A1(_04076_ ), .A2(\mycsreg.CSReg[3][29] ), .A3(_04085_ ), .ZN(_05449_ ) );
NAND3_X1 _13177_ ( .A1(_04091_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_04104_ ), .ZN(_05450_ ) );
NAND3_X1 _13178_ ( .A1(_04092_ ), .A2(\mtvec [29] ), .A3(_04095_ ), .ZN(_05451_ ) );
NAND4_X1 _13179_ ( .A1(_05448_ ), .A2(_05449_ ), .A3(_05450_ ), .A4(_05451_ ), .ZN(_05452_ ) );
AOI211_X1 _13180_ ( .A(_04102_ ), .B(_05452_ ), .C1(_04054_ ), .C2(_04066_ ), .ZN(_05453_ ) );
INV_X1 _13181_ ( .A(\EX_LS_result_csreg_mem [29] ), .ZN(_05454_ ) );
AND3_X1 _13182_ ( .A1(_04054_ ), .A2(_05454_ ), .A3(_04066_ ), .ZN(_05455_ ) );
OR2_X1 _13183_ ( .A1(_05453_ ), .A2(_05455_ ), .ZN(_05456_ ) );
AOI211_X1 _13184_ ( .A(_05433_ ), .B(_05447_ ), .C1(\ID_EX_typ [3] ), .C2(_05456_ ), .ZN(_05457_ ) );
NAND2_X1 _13185_ ( .A1(_04245_ ), .A2(_04246_ ), .ZN(_05458_ ) );
XOR2_X1 _13186_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .Z(_05459_ ) );
XNOR2_X1 _13187_ ( .A(_05458_ ), .B(_05459_ ), .ZN(_05460_ ) );
BUF_X4 _13188_ ( .A(_05418_ ), .Z(_05461_ ) );
BUF_X4 _13189_ ( .A(_05461_ ), .Z(_05462_ ) );
NOR4_X1 _13190_ ( .A1(_04063_ ), .A2(_02056_ ), .A3(_02148_ ), .A4(\EX_LS_flag [0] ), .ZN(_05463_ ) );
NAND2_X1 _13191_ ( .A1(_04055_ ), .A2(\ID_EX_csr [9] ), .ZN(_05464_ ) );
AND4_X1 _13192_ ( .A1(_04033_ ), .A2(_05463_ ), .A3(_04051_ ), .A4(_05464_ ), .ZN(_05465_ ) );
XNOR2_X1 _13193_ ( .A(fanout_net_5 ), .B(\ID_EX_csr [0] ), .ZN(_05466_ ) );
AND3_X1 _13194_ ( .A1(_05466_ ), .A2(_04037_ ), .A3(_04048_ ), .ZN(_05467_ ) );
XNOR2_X1 _13195_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_05468_ ) );
AND4_X1 _13196_ ( .A1(_04035_ ), .A2(_05467_ ), .A3(_04039_ ), .A4(_05468_ ), .ZN(_05469_ ) );
XOR2_X1 _13197_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .Z(_05470_ ) );
NOR2_X1 _13198_ ( .A1(_04064_ ), .A2(_05470_ ), .ZN(_05471_ ) );
NAND2_X1 _13199_ ( .A1(_05471_ ), .A2(_04058_ ), .ZN(_05472_ ) );
NAND2_X1 _13200_ ( .A1(_04053_ ), .A2(_04041_ ), .ZN(_05473_ ) );
NOR3_X2 _13201_ ( .A1(_05472_ ), .A2(_04065_ ), .A3(_05473_ ), .ZN(_05474_ ) );
AND4_X1 _13202_ ( .A1(_05454_ ), .A2(_05465_ ), .A3(_05469_ ), .A4(_05474_ ), .ZN(_05475_ ) );
NAND2_X1 _13203_ ( .A1(_05448_ ), .A2(_05450_ ), .ZN(_05476_ ) );
AND2_X2 _13204_ ( .A1(_05465_ ), .A2(_05469_ ), .ZN(_05477_ ) );
BUF_X4 _13205_ ( .A(_05477_ ), .Z(_05478_ ) );
BUF_X2 _13206_ ( .A(_05474_ ), .Z(_05479_ ) );
AOI21_X1 _13207_ ( .A(_05476_ ), .B1(_05478_ ), .B2(_05479_ ), .ZN(_05480_ ) );
AND3_X1 _13208_ ( .A1(_05449_ ), .A2(_04103_ ), .A3(_05451_ ), .ZN(_05481_ ) );
AOI21_X1 _13209_ ( .A(_05475_ ), .B1(_05480_ ), .B2(_05481_ ), .ZN(_05482_ ) );
OAI211_X1 _13210_ ( .A(_05462_ ), .B(_05424_ ), .C1(_05422_ ), .C2(_05482_ ), .ZN(_05483_ ) );
INV_X1 _13211_ ( .A(_04020_ ), .ZN(_05484_ ) );
AOI21_X1 _13212_ ( .A(_05460_ ), .B1(_05483_ ), .B2(_05484_ ), .ZN(_05485_ ) );
NOR2_X1 _13213_ ( .A1(_05457_ ), .A2(_05485_ ), .ZN(_05486_ ) );
BUF_X4 _13214_ ( .A(_04019_ ), .Z(_05487_ ) );
BUF_X2 _13215_ ( .A(_05487_ ), .Z(_05488_ ) );
OR3_X1 _13216_ ( .A1(_03188_ ), .A2(_05488_ ), .A3(_05425_ ), .ZN(_05489_ ) );
AOI21_X1 _13217_ ( .A(_04032_ ), .B1(_05486_ ), .B2(_05489_ ), .ZN(_00159_ ) );
BUF_X2 _13218_ ( .A(_04054_ ), .Z(_05490_ ) );
INV_X1 _13219_ ( .A(\EX_LS_result_csreg_mem [20] ), .ZN(_05491_ ) );
BUF_X2 _13220_ ( .A(_04066_ ), .Z(_05492_ ) );
AND3_X1 _13221_ ( .A1(_05490_ ), .A2(_05491_ ), .A3(_05492_ ), .ZN(_05493_ ) );
NOR2_X1 _13222_ ( .A1(_04068_ ), .A2(_04102_ ), .ZN(_05494_ ) );
AND2_X1 _13223_ ( .A1(_04101_ ), .A2(_04085_ ), .ZN(_05495_ ) );
INV_X1 _13224_ ( .A(_05495_ ), .ZN(_05496_ ) );
AND2_X1 _13225_ ( .A1(_05494_ ), .A2(_05496_ ), .ZN(_05497_ ) );
BUF_X4 _13226_ ( .A(_04076_ ), .Z(_05498_ ) );
BUF_X2 _13227_ ( .A(_05498_ ), .Z(_05499_ ) );
BUF_X2 _13228_ ( .A(_04085_ ), .Z(_05500_ ) );
NAND3_X1 _13229_ ( .A1(_05499_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_05500_ ), .ZN(_05501_ ) );
BUF_X2 _13230_ ( .A(_04076_ ), .Z(_05502_ ) );
NAND3_X1 _13231_ ( .A1(_05502_ ), .A2(\mepc [20] ), .A3(_04082_ ), .ZN(_05503_ ) );
BUF_X2 _13232_ ( .A(_04092_ ), .Z(_05504_ ) );
BUF_X2 _13233_ ( .A(_04104_ ), .Z(_05505_ ) );
NAND3_X1 _13234_ ( .A1(_05504_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_05505_ ), .ZN(_05506_ ) );
BUF_X2 _13235_ ( .A(_04095_ ), .Z(_05507_ ) );
NAND3_X1 _13236_ ( .A1(_05504_ ), .A2(\mtvec [20] ), .A3(_05507_ ), .ZN(_05508_ ) );
AND4_X1 _13237_ ( .A1(_05501_ ), .A2(_05503_ ), .A3(_05506_ ), .A4(_05508_ ), .ZN(_05509_ ) );
AOI21_X1 _13238_ ( .A(_05493_ ), .B1(_05497_ ), .B2(_05509_ ), .ZN(_05510_ ) );
NAND3_X1 _13239_ ( .A1(_04117_ ), .A2(_05437_ ), .A3(_05440_ ), .ZN(_05511_ ) );
XNOR2_X1 _13240_ ( .A(_05511_ ), .B(\ID_EX_pc [20] ), .ZN(_05512_ ) );
OAI21_X1 _13241_ ( .A(_04143_ ), .B1(_04189_ ), .B2(_04208_ ), .ZN(_05513_ ) );
NAND2_X1 _13242_ ( .A1(_05513_ ), .A2(_04219_ ), .ZN(_05514_ ) );
XOR2_X1 _13243_ ( .A(_05514_ ), .B(_04134_ ), .Z(_05515_ ) );
MUX2_X1 _13244_ ( .A(_05512_ ), .B(_05515_ ), .S(_05419_ ), .Z(_05516_ ) );
MUX2_X1 _13245_ ( .A(_05510_ ), .B(_05516_ ), .S(_05422_ ), .Z(_05517_ ) );
NAND2_X1 _13246_ ( .A1(_05517_ ), .A2(_05426_ ), .ZN(_05518_ ) );
AND2_X2 _13247_ ( .A1(_04018_ ), .A2(fanout_net_7 ), .ZN(_05519_ ) );
AND3_X1 _13248_ ( .A1(_03163_ ), .A2(_03160_ ), .A3(_05519_ ), .ZN(_05520_ ) );
BUF_X4 _13249_ ( .A(_04020_ ), .Z(_05521_ ) );
AOI21_X1 _13250_ ( .A(_05520_ ), .B1(_05521_ ), .B2(_05515_ ), .ZN(_05522_ ) );
AOI21_X1 _13251_ ( .A(_04032_ ), .B1(_05518_ ), .B2(_05522_ ), .ZN(_00160_ ) );
NOR2_X1 _13252_ ( .A1(_04189_ ), .A2(_04208_ ), .ZN(_05523_ ) );
NOR2_X1 _13253_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_05524_ ) );
NOR3_X1 _13254_ ( .A1(_05523_ ), .A2(_04215_ ), .A3(_05524_ ), .ZN(_05525_ ) );
AND2_X1 _13255_ ( .A1(_05525_ ), .A2(_04141_ ), .ZN(_05526_ ) );
OAI21_X1 _13256_ ( .A(_04139_ ), .B1(_05526_ ), .B2(_04218_ ), .ZN(_05527_ ) );
NAND2_X1 _13257_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_05528_ ) );
AND2_X1 _13258_ ( .A1(_05527_ ), .A2(_05528_ ), .ZN(_05529_ ) );
XNOR2_X1 _13259_ ( .A(_05529_ ), .B(_04138_ ), .ZN(_05530_ ) );
AOI21_X1 _13260_ ( .A(\ID_EX_typ [3] ), .B1(_05461_ ), .B2(_05530_ ), .ZN(_05531_ ) );
NAND3_X1 _13261_ ( .A1(_04117_ ), .A2(\ID_EX_pc [18] ), .A3(_05437_ ), .ZN(_05532_ ) );
XNOR2_X1 _13262_ ( .A(_05532_ ), .B(_04213_ ), .ZN(_05533_ ) );
OAI21_X1 _13263_ ( .A(_05531_ ), .B1(_05462_ ), .B2(_05533_ ), .ZN(_05534_ ) );
BUF_X4 _13264_ ( .A(_05425_ ), .Z(_05535_ ) );
BUF_X4 _13265_ ( .A(_05421_ ), .Z(_05536_ ) );
BUF_X4 _13266_ ( .A(_05536_ ), .Z(_05537_ ) );
NAND3_X1 _13267_ ( .A1(_04077_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_04086_ ), .ZN(_05538_ ) );
BUF_X2 _13268_ ( .A(_04092_ ), .Z(_05539_ ) );
NAND3_X1 _13269_ ( .A1(_05539_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_04105_ ), .ZN(_05540_ ) );
AND2_X1 _13270_ ( .A1(_05538_ ), .A2(_05540_ ), .ZN(_05541_ ) );
NAND3_X1 _13271_ ( .A1(_05504_ ), .A2(\mtvec [19] ), .A3(_05507_ ), .ZN(_05542_ ) );
BUF_X4 _13272_ ( .A(_04081_ ), .Z(_05543_ ) );
BUF_X4 _13273_ ( .A(_05543_ ), .Z(_05544_ ) );
NAND3_X1 _13274_ ( .A1(_05502_ ), .A2(\mepc [19] ), .A3(_05544_ ), .ZN(_05545_ ) );
NAND4_X1 _13275_ ( .A1(_05541_ ), .A2(_05496_ ), .A3(_05542_ ), .A4(_05545_ ), .ZN(_05546_ ) );
NAND2_X1 _13276_ ( .A1(_04069_ ), .A2(_05546_ ), .ZN(_05547_ ) );
BUF_X2 _13277_ ( .A(_04054_ ), .Z(_05548_ ) );
BUF_X2 _13278_ ( .A(_04066_ ), .Z(_05549_ ) );
NAND3_X1 _13279_ ( .A1(_05548_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_05549_ ), .ZN(_05550_ ) );
AND2_X1 _13280_ ( .A1(_05547_ ), .A2(_05550_ ), .ZN(_05551_ ) );
INV_X1 _13281_ ( .A(_05551_ ), .ZN(_05552_ ) );
OAI211_X1 _13282_ ( .A(_05534_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05552_ ), .ZN(_05553_ ) );
NOR3_X1 _13283_ ( .A1(_03169_ ), .A2(_05488_ ), .A3(_05425_ ), .ZN(_05554_ ) );
AOI21_X1 _13284_ ( .A(_05554_ ), .B1(_05521_ ), .B2(_05530_ ), .ZN(_05555_ ) );
AOI21_X1 _13285_ ( .A(_04032_ ), .B1(_05553_ ), .B2(_05555_ ), .ZN(_00161_ ) );
INV_X1 _13286_ ( .A(\ID_EX_pc [18] ), .ZN(_05556_ ) );
XNOR2_X1 _13287_ ( .A(_05438_ ), .B(_05556_ ), .ZN(_05557_ ) );
OR3_X1 _13288_ ( .A1(_05526_ ), .A2(_04139_ ), .A3(_04218_ ), .ZN(_05558_ ) );
AND2_X1 _13289_ ( .A1(_05558_ ), .A2(_05527_ ), .ZN(_05559_ ) );
MUX2_X1 _13290_ ( .A(_05557_ ), .B(_05559_ ), .S(_05419_ ), .Z(_05560_ ) );
OR2_X1 _13291_ ( .A1(_05560_ ), .A2(\ID_EX_typ [3] ), .ZN(_05561_ ) );
BUF_X2 _13292_ ( .A(_05490_ ), .Z(_05562_ ) );
BUF_X2 _13293_ ( .A(_05492_ ), .Z(_05563_ ) );
NAND3_X1 _13294_ ( .A1(_05562_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_05563_ ), .ZN(_05564_ ) );
BUF_X2 _13295_ ( .A(_04068_ ), .Z(_05565_ ) );
BUF_X4 _13296_ ( .A(_04077_ ), .Z(_05566_ ) );
NAND3_X1 _13297_ ( .A1(_05566_ ), .A2(\mepc [18] ), .A3(_05544_ ), .ZN(_05567_ ) );
BUF_X2 _13298_ ( .A(_05539_ ), .Z(_05568_ ) );
NAND3_X1 _13299_ ( .A1(_05568_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_04106_ ), .ZN(_05569_ ) );
NAND3_X1 _13300_ ( .A1(_04094_ ), .A2(\mtvec [18] ), .A3(_04097_ ), .ZN(_05570_ ) );
NAND3_X1 _13301_ ( .A1(_05567_ ), .A2(_05569_ ), .A3(_05570_ ), .ZN(_05571_ ) );
BUF_X2 _13302_ ( .A(_04086_ ), .Z(_05572_ ) );
NAND3_X1 _13303_ ( .A1(_05566_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_05572_ ), .ZN(_05573_ ) );
BUF_X2 _13304_ ( .A(_05496_ ), .Z(_05574_ ) );
NAND2_X1 _13305_ ( .A1(_05573_ ), .A2(_05574_ ), .ZN(_05575_ ) );
NOR2_X1 _13306_ ( .A1(_05571_ ), .A2(_05575_ ), .ZN(_05576_ ) );
OAI21_X1 _13307_ ( .A(_05564_ ), .B1(_05565_ ), .B2(_05576_ ), .ZN(_05577_ ) );
OAI211_X1 _13308_ ( .A(_05561_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05577_ ), .ZN(_05578_ ) );
BUF_X4 _13309_ ( .A(_05519_ ), .Z(_05579_ ) );
BUF_X4 _13310_ ( .A(_04020_ ), .Z(_05580_ ) );
AOI22_X1 _13311_ ( .A1(_03170_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05559_ ), .ZN(_05581_ ) );
AOI21_X1 _13312_ ( .A(_04032_ ), .B1(_05578_ ), .B2(_05581_ ), .ZN(_00162_ ) );
BUF_X4 _13313_ ( .A(_05425_ ), .Z(_05582_ ) );
BUF_X4 _13314_ ( .A(_05422_ ), .Z(_05583_ ) );
AND3_X1 _13315_ ( .A1(_04092_ ), .A2(\mtvec [17] ), .A3(_04095_ ), .ZN(_05584_ ) );
AOI21_X1 _13316_ ( .A(_05584_ ), .B1(_05477_ ), .B2(_05474_ ), .ZN(_05585_ ) );
NOR2_X1 _13317_ ( .A1(_04102_ ), .A2(_05495_ ), .ZN(_05586_ ) );
NAND3_X1 _13318_ ( .A1(_05502_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_05500_ ), .ZN(_05587_ ) );
NAND3_X1 _13319_ ( .A1(_05498_ ), .A2(\mepc [17] ), .A3(_05543_ ), .ZN(_05588_ ) );
NAND3_X1 _13320_ ( .A1(_04093_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_04105_ ), .ZN(_05589_ ) );
AND2_X1 _13321_ ( .A1(_05588_ ), .A2(_05589_ ), .ZN(_05590_ ) );
NAND4_X1 _13322_ ( .A1(_05585_ ), .A2(_05586_ ), .A3(_05587_ ), .A4(_05590_ ), .ZN(_05591_ ) );
INV_X1 _13323_ ( .A(\EX_LS_result_csreg_mem [17] ), .ZN(_05592_ ) );
NAND4_X1 _13324_ ( .A1(_05465_ ), .A2(_05474_ ), .A3(_05592_ ), .A4(_05469_ ), .ZN(_05593_ ) );
AND2_X1 _13325_ ( .A1(_05591_ ), .A2(_05593_ ), .ZN(_05594_ ) );
OR2_X1 _13326_ ( .A1(_05525_ ), .A2(_04215_ ), .ZN(_05595_ ) );
XNOR2_X1 _13327_ ( .A(_05595_ ), .B(_04141_ ), .ZN(_05596_ ) );
OAI21_X1 _13328_ ( .A(_05536_ ), .B1(_05435_ ), .B2(_05596_ ), .ZN(_05597_ ) );
NAND3_X1 _13329_ ( .A1(_04121_ ), .A2(\ID_EX_pc [15] ), .A3(\ID_EX_pc [14] ), .ZN(_05598_ ) );
INV_X1 _13330_ ( .A(\ID_EX_pc [16] ), .ZN(_05599_ ) );
NOR2_X1 _13331_ ( .A1(_05598_ ), .A2(_05599_ ), .ZN(_05600_ ) );
XNOR2_X1 _13332_ ( .A(_05600_ ), .B(\ID_EX_pc [17] ), .ZN(_05601_ ) );
AOI21_X1 _13333_ ( .A(_05601_ ), .B1(_05415_ ), .B2(_05417_ ), .ZN(_05602_ ) );
OAI221_X1 _13334_ ( .A(_05582_ ), .B1(_05583_ ), .B2(_05594_ ), .C1(_05597_ ), .C2(_05602_ ), .ZN(_05603_ ) );
BUF_X2 _13335_ ( .A(_05487_ ), .Z(_05604_ ) );
BUF_X4 _13336_ ( .A(_05424_ ), .Z(_05605_ ) );
NOR3_X1 _13337_ ( .A1(_03172_ ), .A2(_05604_ ), .A3(_05605_ ), .ZN(_05606_ ) );
NOR2_X1 _13338_ ( .A1(_05596_ ), .A2(_05484_ ), .ZN(_05607_ ) );
NOR2_X1 _13339_ ( .A1(_05606_ ), .A2(_05607_ ), .ZN(_05608_ ) );
AOI21_X1 _13340_ ( .A(_04032_ ), .B1(_05603_ ), .B2(_05608_ ), .ZN(_00163_ ) );
XNOR2_X1 _13341_ ( .A(_05598_ ), .B(\ID_EX_pc [16] ), .ZN(_05609_ ) );
XNOR2_X1 _13342_ ( .A(_05523_ ), .B(_04142_ ), .ZN(_05610_ ) );
MUX2_X1 _13343_ ( .A(_05609_ ), .B(_05610_ ), .S(_05419_ ), .Z(_05611_ ) );
OR2_X1 _13344_ ( .A1(_05611_ ), .A2(\ID_EX_typ [3] ), .ZN(_05612_ ) );
INV_X1 _13345_ ( .A(\EX_LS_result_csreg_mem [16] ), .ZN(_05613_ ) );
AND3_X1 _13346_ ( .A1(_05548_ ), .A2(_05613_ ), .A3(_05549_ ), .ZN(_05614_ ) );
NAND3_X1 _13347_ ( .A1(_05566_ ), .A2(\mepc [16] ), .A3(_05544_ ), .ZN(_05615_ ) );
NAND3_X1 _13348_ ( .A1(_05566_ ), .A2(\mycsreg.CSReg[3][16] ), .A3(_05572_ ), .ZN(_05616_ ) );
NAND3_X1 _13349_ ( .A1(_05568_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_04106_ ), .ZN(_05617_ ) );
NAND3_X1 _13350_ ( .A1(_05568_ ), .A2(\mtvec [16] ), .A3(_04097_ ), .ZN(_05618_ ) );
AND4_X1 _13351_ ( .A1(_05615_ ), .A2(_05616_ ), .A3(_05617_ ), .A4(_05618_ ), .ZN(_05619_ ) );
AOI21_X1 _13352_ ( .A(_05614_ ), .B1(_05497_ ), .B2(_05619_ ), .ZN(_05620_ ) );
OAI211_X1 _13353_ ( .A(_05612_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05620_ ), .ZN(_05621_ ) );
NOR4_X1 _13354_ ( .A1(_03173_ ), .A2(_02896_ ), .A3(_05487_ ), .A4(_05424_ ), .ZN(_05622_ ) );
AOI21_X1 _13355_ ( .A(_05622_ ), .B1(_05610_ ), .B2(_05521_ ), .ZN(_05623_ ) );
AOI21_X1 _13356_ ( .A(_04032_ ), .B1(_05621_ ), .B2(_05623_ ), .ZN(_00164_ ) );
NAND3_X1 _13357_ ( .A1(_05548_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_05549_ ), .ZN(_05624_ ) );
AND3_X1 _13358_ ( .A1(_05539_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_04105_ ), .ZN(_05625_ ) );
INV_X1 _13359_ ( .A(_05625_ ), .ZN(_05626_ ) );
NAND3_X1 _13360_ ( .A1(_05499_ ), .A2(\mepc [15] ), .A3(_05544_ ), .ZN(_05627_ ) );
NAND3_X1 _13361_ ( .A1(_05499_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_05572_ ), .ZN(_05628_ ) );
NAND3_X1 _13362_ ( .A1(_05626_ ), .A2(_05627_ ), .A3(_05628_ ), .ZN(_05629_ ) );
NAND3_X1 _13363_ ( .A1(_04094_ ), .A2(\mtvec [15] ), .A3(_04097_ ), .ZN(_05630_ ) );
NAND2_X1 _13364_ ( .A1(_05574_ ), .A2(_05630_ ), .ZN(_05631_ ) );
NOR2_X1 _13365_ ( .A1(_05629_ ), .A2(_05631_ ), .ZN(_05632_ ) );
OAI21_X1 _13366_ ( .A(_05624_ ), .B1(_05565_ ), .B2(_05632_ ), .ZN(_05633_ ) );
AND2_X1 _13367_ ( .A1(_04121_ ), .A2(\ID_EX_pc [14] ), .ZN(_05634_ ) );
INV_X1 _13368_ ( .A(\ID_EX_pc [15] ), .ZN(_05635_ ) );
XNOR2_X1 _13369_ ( .A(_05634_ ), .B(_05635_ ), .ZN(_05636_ ) );
INV_X1 _13370_ ( .A(_04179_ ), .ZN(_05637_ ) );
AND2_X1 _13371_ ( .A1(_04173_ ), .A2(_04188_ ), .ZN(_05638_ ) );
OAI21_X1 _13372_ ( .A(_04177_ ), .B1(_05638_ ), .B2(_04197_ ), .ZN(_05639_ ) );
AOI21_X1 _13373_ ( .A(_05637_ ), .B1(_05639_ ), .B2(_04201_ ), .ZN(_05640_ ) );
NOR2_X1 _13374_ ( .A1(_05640_ ), .A2(_04204_ ), .ZN(_05641_ ) );
XNOR2_X1 _13375_ ( .A(_05641_ ), .B(_04178_ ), .ZN(_05642_ ) );
MUX2_X1 _13376_ ( .A(_05636_ ), .B(_05642_ ), .S(_05419_ ), .Z(_05643_ ) );
MUX2_X1 _13377_ ( .A(_05633_ ), .B(_05643_ ), .S(_05422_ ), .Z(_05644_ ) );
NAND2_X1 _13378_ ( .A1(_05644_ ), .A2(_05426_ ), .ZN(_05645_ ) );
NOR3_X1 _13379_ ( .A1(_03181_ ), .A2(_05488_ ), .A3(_05425_ ), .ZN(_05646_ ) );
AOI21_X1 _13380_ ( .A(_05646_ ), .B1(_05521_ ), .B2(_05642_ ), .ZN(_05647_ ) );
AOI21_X1 _13381_ ( .A(_04032_ ), .B1(_05645_ ), .B2(_05647_ ), .ZN(_00165_ ) );
BUF_X4 _13382_ ( .A(_05430_ ), .Z(_05648_ ) );
NAND3_X1 _13383_ ( .A1(_04076_ ), .A2(\mepc [14] ), .A3(_04081_ ), .ZN(_05649_ ) );
NAND3_X1 _13384_ ( .A1(_04091_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_04104_ ), .ZN(_05650_ ) );
AND2_X1 _13385_ ( .A1(_05649_ ), .A2(_05650_ ), .ZN(_05651_ ) );
INV_X1 _13386_ ( .A(_05651_ ), .ZN(_05652_ ) );
AOI21_X1 _13387_ ( .A(_05652_ ), .B1(_05477_ ), .B2(_05474_ ), .ZN(_05653_ ) );
BUF_X2 _13388_ ( .A(_04092_ ), .Z(_05654_ ) );
NAND3_X1 _13389_ ( .A1(_05654_ ), .A2(\mtvec [14] ), .A3(_05507_ ), .ZN(_05655_ ) );
BUF_X4 _13390_ ( .A(_04076_ ), .Z(_05656_ ) );
NAND3_X1 _13391_ ( .A1(_05656_ ), .A2(\mycsreg.CSReg[3][14] ), .A3(_05500_ ), .ZN(_05657_ ) );
AND4_X1 _13392_ ( .A1(_05586_ ), .A2(_05653_ ), .A3(_05655_ ), .A4(_05657_ ), .ZN(_05658_ ) );
INV_X1 _13393_ ( .A(\EX_LS_result_csreg_mem [14] ), .ZN(_05659_ ) );
AND4_X1 _13394_ ( .A1(_05659_ ), .A2(_05465_ ), .A3(_05469_ ), .A4(_05474_ ), .ZN(_05660_ ) );
NOR2_X1 _13395_ ( .A1(_05658_ ), .A2(_05660_ ), .ZN(_05661_ ) );
INV_X1 _13396_ ( .A(_05661_ ), .ZN(_05662_ ) );
AOI21_X1 _13397_ ( .A(_05648_ ), .B1(_05662_ ), .B2(\ID_EX_typ [3] ), .ZN(_05663_ ) );
INV_X1 _13398_ ( .A(\ID_EX_pc [14] ), .ZN(_05664_ ) );
XNOR2_X1 _13399_ ( .A(_04121_ ), .B(_05664_ ), .ZN(_05665_ ) );
NAND2_X1 _13400_ ( .A1(_05639_ ), .A2(_04201_ ), .ZN(_05666_ ) );
XNOR2_X1 _13401_ ( .A(_05666_ ), .B(_05637_ ), .ZN(_05667_ ) );
MUX2_X1 _13402_ ( .A(_05665_ ), .B(_05667_ ), .S(_05461_ ), .Z(_05668_ ) );
OAI21_X1 _13403_ ( .A(_05663_ ), .B1(_05668_ ), .B2(\ID_EX_typ [3] ), .ZN(_05669_ ) );
AND3_X1 _13404_ ( .A1(_03182_ ), .A2(_03178_ ), .A3(_05519_ ), .ZN(_05670_ ) );
AOI21_X1 _13405_ ( .A(_05670_ ), .B1(_05521_ ), .B2(_05667_ ), .ZN(_05671_ ) );
AOI21_X1 _13406_ ( .A(_04032_ ), .B1(_05669_ ), .B2(_05671_ ), .ZN(_00166_ ) );
NAND3_X1 _13407_ ( .A1(_04077_ ), .A2(\mepc [13] ), .A3(_05543_ ), .ZN(_05672_ ) );
NAND3_X1 _13408_ ( .A1(_05539_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_05505_ ), .ZN(_05673_ ) );
AND2_X1 _13409_ ( .A1(_05672_ ), .A2(_05673_ ), .ZN(_05674_ ) );
NAND3_X1 _13410_ ( .A1(_04094_ ), .A2(\mtvec [13] ), .A3(_04097_ ), .ZN(_05675_ ) );
NAND3_X1 _13411_ ( .A1(_05499_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_05572_ ), .ZN(_05676_ ) );
AND4_X1 _13412_ ( .A1(_05494_ ), .A2(_05674_ ), .A3(_05675_ ), .A4(_05676_ ), .ZN(_05677_ ) );
INV_X1 _13413_ ( .A(\EX_LS_result_csreg_mem [13] ), .ZN(_05678_ ) );
AND3_X1 _13414_ ( .A1(_05490_ ), .A2(_05678_ ), .A3(_05492_ ), .ZN(_05679_ ) );
NOR2_X1 _13415_ ( .A1(_05677_ ), .A2(_05679_ ), .ZN(_05680_ ) );
XNOR2_X1 _13416_ ( .A(_04120_ ), .B(\ID_EX_pc [13] ), .ZN(_05681_ ) );
OAI21_X1 _13417_ ( .A(_05536_ ), .B1(_05462_ ), .B2(_05681_ ), .ZN(_05682_ ) );
OAI21_X1 _13418_ ( .A(_04174_ ), .B1(_05638_ ), .B2(_04197_ ), .ZN(_05683_ ) );
NAND2_X1 _13419_ ( .A1(_05683_ ), .A2(_04199_ ), .ZN(_05684_ ) );
XNOR2_X1 _13420_ ( .A(_05684_ ), .B(_04176_ ), .ZN(_05685_ ) );
AND3_X1 _13421_ ( .A1(_05415_ ), .A2(_05417_ ), .A3(_05685_ ), .ZN(_05686_ ) );
OAI221_X1 _13422_ ( .A(_05582_ ), .B1(_05583_ ), .B2(_05680_ ), .C1(_05682_ ), .C2(_05686_ ), .ZN(_05687_ ) );
AOI22_X1 _13423_ ( .A1(_05685_ ), .A2(_05521_ ), .B1(_03185_ ), .B2(_05519_ ), .ZN(_05688_ ) );
AOI21_X1 _13424_ ( .A(_04032_ ), .B1(_05687_ ), .B2(_05688_ ), .ZN(_00167_ ) );
BUF_X4 _13425_ ( .A(_04031_ ), .Z(_05689_ ) );
INV_X1 _13426_ ( .A(\ID_EX_pc [12] ), .ZN(_05690_ ) );
XNOR2_X1 _13427_ ( .A(_04119_ ), .B(_05690_ ), .ZN(_05691_ ) );
OR3_X1 _13428_ ( .A1(_05638_ ), .A2(_04174_ ), .A3(_04197_ ), .ZN(_05692_ ) );
AND2_X1 _13429_ ( .A1(_05683_ ), .A2(_05692_ ), .ZN(_05693_ ) );
MUX2_X1 _13430_ ( .A(_05691_ ), .B(_05693_ ), .S(_05461_ ), .Z(_05694_ ) );
AND2_X1 _13431_ ( .A1(_05694_ ), .A2(_05536_ ), .ZN(_05695_ ) );
NAND3_X1 _13432_ ( .A1(_05502_ ), .A2(\mepc [12] ), .A3(_04082_ ), .ZN(_05696_ ) );
NAND3_X1 _13433_ ( .A1(_05654_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_05505_ ), .ZN(_05697_ ) );
NAND2_X1 _13434_ ( .A1(_05696_ ), .A2(_05697_ ), .ZN(_05698_ ) );
BUF_X2 _13435_ ( .A(_05474_ ), .Z(_05699_ ) );
AOI21_X1 _13436_ ( .A(_05698_ ), .B1(_05478_ ), .B2(_05699_ ), .ZN(_05700_ ) );
NAND3_X1 _13437_ ( .A1(_05654_ ), .A2(\mtvec [12] ), .A3(_05507_ ), .ZN(_05701_ ) );
NAND3_X1 _13438_ ( .A1(_05656_ ), .A2(\mycsreg.CSReg[3][12] ), .A3(_05500_ ), .ZN(_05702_ ) );
NAND4_X1 _13439_ ( .A1(_05700_ ), .A2(_05586_ ), .A3(_05701_ ), .A4(_05702_ ), .ZN(_05703_ ) );
BUF_X2 _13440_ ( .A(_05465_ ), .Z(_05704_ ) );
INV_X1 _13441_ ( .A(\EX_LS_result_csreg_mem [12] ), .ZN(_05705_ ) );
BUF_X2 _13442_ ( .A(_05469_ ), .Z(_05706_ ) );
NAND4_X1 _13443_ ( .A1(_05704_ ), .A2(_05699_ ), .A3(_05705_ ), .A4(_05706_ ), .ZN(_05707_ ) );
NAND3_X1 _13444_ ( .A1(_05703_ ), .A2(\ID_EX_typ [3] ), .A3(_05707_ ), .ZN(_05708_ ) );
INV_X1 _13445_ ( .A(_05708_ ), .ZN(_05709_ ) );
OAI21_X1 _13446_ ( .A(_05426_ ), .B1(_05695_ ), .B2(_05709_ ), .ZN(_05710_ ) );
AOI22_X1 _13447_ ( .A1(_05693_ ), .A2(_05521_ ), .B1(_03186_ ), .B2(_05519_ ), .ZN(_05711_ ) );
AOI21_X1 _13448_ ( .A(_05689_ ), .B1(_05710_ ), .B2(_05711_ ), .ZN(_00168_ ) );
AND2_X1 _13449_ ( .A1(_04117_ ), .A2(\ID_EX_pc [10] ), .ZN(_05712_ ) );
INV_X1 _13450_ ( .A(\ID_EX_pc [11] ), .ZN(_05713_ ) );
XNOR2_X1 _13451_ ( .A(_05712_ ), .B(_05713_ ), .ZN(_05714_ ) );
AOI21_X1 _13452_ ( .A(\ID_EX_typ [3] ), .B1(_05435_ ), .B2(_05714_ ), .ZN(_05715_ ) );
INV_X1 _13453_ ( .A(_04183_ ), .ZN(_05716_ ) );
OAI21_X1 _13454_ ( .A(_04187_ ), .B1(_04170_ ), .B2(_04171_ ), .ZN(_05717_ ) );
AOI21_X1 _13455_ ( .A(_05716_ ), .B1(_05717_ ), .B2(_04195_ ), .ZN(_05718_ ) );
OR2_X1 _13456_ ( .A1(_05718_ ), .A2(_04190_ ), .ZN(_05719_ ) );
XNOR2_X1 _13457_ ( .A(_05719_ ), .B(_04182_ ), .ZN(_05720_ ) );
OAI21_X1 _13458_ ( .A(_05715_ ), .B1(_05435_ ), .B2(_05720_ ), .ZN(_05721_ ) );
BUF_X4 _13459_ ( .A(_04103_ ), .Z(_05722_ ) );
NAND3_X1 _13460_ ( .A1(_04077_ ), .A2(\mepc [11] ), .A3(_05543_ ), .ZN(_05723_ ) );
NAND3_X1 _13461_ ( .A1(_04077_ ), .A2(\mycsreg.CSReg[3][11] ), .A3(_04086_ ), .ZN(_05724_ ) );
NAND3_X1 _13462_ ( .A1(_04093_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_04105_ ), .ZN(_05725_ ) );
NAND3_X1 _13463_ ( .A1(_04093_ ), .A2(\mtvec [11] ), .A3(_04096_ ), .ZN(_05726_ ) );
AND4_X1 _13464_ ( .A1(_05723_ ), .A2(_05724_ ), .A3(_05725_ ), .A4(_05726_ ), .ZN(_05727_ ) );
NAND4_X1 _13465_ ( .A1(_04069_ ), .A2(_05722_ ), .A3(_05574_ ), .A4(_05727_ ), .ZN(_05728_ ) );
INV_X1 _13466_ ( .A(\EX_LS_result_csreg_mem [11] ), .ZN(_05729_ ) );
NAND3_X1 _13467_ ( .A1(_05548_ ), .A2(_05729_ ), .A3(_05549_ ), .ZN(_05730_ ) );
AND2_X1 _13468_ ( .A1(_05728_ ), .A2(_05730_ ), .ZN(_05731_ ) );
OAI211_X1 _13469_ ( .A(_05721_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05731_ ), .ZN(_05732_ ) );
NOR2_X1 _13470_ ( .A1(_05720_ ), .A2(_05484_ ), .ZN(_05733_ ) );
AND2_X1 _13471_ ( .A1(_02677_ ), .A2(_02783_ ), .ZN(_05734_ ) );
INV_X1 _13472_ ( .A(_05734_ ), .ZN(_05735_ ) );
AOI21_X1 _13473_ ( .A(_02787_ ), .B1(_05735_ ), .B2(_02525_ ), .ZN(_05736_ ) );
AOI21_X1 _13474_ ( .A(\ID_EX_imm [10] ), .B1(_02569_ ), .B2(_02570_ ), .ZN(_05737_ ) );
NOR3_X1 _13475_ ( .A1(_05736_ ), .A2(_02789_ ), .A3(_05737_ ), .ZN(_05738_ ) );
NOR2_X1 _13476_ ( .A1(_05738_ ), .A2(_02789_ ), .ZN(_05739_ ) );
XNOR2_X1 _13477_ ( .A(_05739_ ), .B(_02549_ ), .ZN(_05740_ ) );
AOI21_X1 _13478_ ( .A(_05733_ ), .B1(_05740_ ), .B2(_05579_ ), .ZN(_05741_ ) );
AOI21_X1 _13479_ ( .A(_05689_ ), .B1(_05732_ ), .B2(_05741_ ), .ZN(_00169_ ) );
XNOR2_X1 _13480_ ( .A(_05443_ ), .B(\ID_EX_pc [28] ), .ZN(_05742_ ) );
XOR2_X1 _13481_ ( .A(_04243_ ), .B(_04244_ ), .Z(_05743_ ) );
MUX2_X1 _13482_ ( .A(_05742_ ), .B(_05743_ ), .S(_05419_ ), .Z(_05744_ ) );
OR2_X1 _13483_ ( .A1(_05744_ ), .A2(\ID_EX_typ [3] ), .ZN(_05745_ ) );
INV_X1 _13484_ ( .A(\EX_LS_result_csreg_mem [28] ), .ZN(_05746_ ) );
AND3_X1 _13485_ ( .A1(_05562_ ), .A2(_05746_ ), .A3(_05563_ ), .ZN(_05747_ ) );
NAND3_X1 _13486_ ( .A1(_05566_ ), .A2(\mycsreg.CSReg[3][28] ), .A3(_05572_ ), .ZN(_05748_ ) );
NAND3_X1 _13487_ ( .A1(_05499_ ), .A2(\mepc [28] ), .A3(_05544_ ), .ZN(_05749_ ) );
NAND2_X1 _13488_ ( .A1(_05748_ ), .A2(_05749_ ), .ZN(_05750_ ) );
AND3_X1 _13489_ ( .A1(_05568_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_04106_ ), .ZN(_05751_ ) );
AND3_X1 _13490_ ( .A1(_05504_ ), .A2(\mtvec [28] ), .A3(_05507_ ), .ZN(_05752_ ) );
NOR3_X1 _13491_ ( .A1(_05750_ ), .A2(_05751_ ), .A3(_05752_ ), .ZN(_05753_ ) );
AOI21_X1 _13492_ ( .A(_05747_ ), .B1(_05494_ ), .B2(_05753_ ), .ZN(_05754_ ) );
OAI211_X1 _13493_ ( .A(_05745_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05754_ ), .ZN(_05755_ ) );
NAND2_X1 _13494_ ( .A1(_03189_ ), .A2(fanout_net_7 ), .ZN(_05756_ ) );
OAI211_X1 _13495_ ( .A(_05756_ ), .B(_05431_ ), .C1(fanout_net_7 ), .C2(_05743_ ), .ZN(_05757_ ) );
AOI21_X1 _13496_ ( .A(_05689_ ), .B1(_05755_ ), .B2(_05757_ ), .ZN(_00170_ ) );
INV_X1 _13497_ ( .A(\ID_EX_pc [10] ), .ZN(_05758_ ) );
XNOR2_X1 _13498_ ( .A(_04117_ ), .B(_05758_ ), .ZN(_05759_ ) );
AOI21_X1 _13499_ ( .A(\ID_EX_typ [3] ), .B1(_05435_ ), .B2(_05759_ ), .ZN(_05760_ ) );
NAND2_X1 _13500_ ( .A1(_05717_ ), .A2(_04195_ ), .ZN(_05761_ ) );
XNOR2_X1 _13501_ ( .A(_05761_ ), .B(_05716_ ), .ZN(_05762_ ) );
INV_X1 _13502_ ( .A(_05762_ ), .ZN(_05763_ ) );
OAI21_X1 _13503_ ( .A(_05760_ ), .B1(_05435_ ), .B2(_05763_ ), .ZN(_05764_ ) );
NAND3_X1 _13504_ ( .A1(_05562_ ), .A2(\EX_LS_result_csreg_mem [10] ), .A3(_05563_ ), .ZN(_05765_ ) );
NAND3_X1 _13505_ ( .A1(_05499_ ), .A2(\mepc [10] ), .A3(_05544_ ), .ZN(_05766_ ) );
NAND3_X1 _13506_ ( .A1(_04094_ ), .A2(\mycsreg.CSReg[0][10] ), .A3(_04106_ ), .ZN(_05767_ ) );
NAND2_X1 _13507_ ( .A1(_05766_ ), .A2(_05767_ ), .ZN(_05768_ ) );
AND3_X1 _13508_ ( .A1(_05502_ ), .A2(\mycsreg.CSReg[3][10] ), .A3(_05500_ ), .ZN(_05769_ ) );
AND3_X1 _13509_ ( .A1(_05654_ ), .A2(\mtvec [10] ), .A3(_04096_ ), .ZN(_05770_ ) );
NOR4_X1 _13510_ ( .A1(_05768_ ), .A2(_05769_ ), .A3(_05495_ ), .A4(_05770_ ), .ZN(_05771_ ) );
OAI21_X1 _13511_ ( .A(_05765_ ), .B1(_05565_ ), .B2(_05771_ ), .ZN(_05772_ ) );
OAI211_X1 _13512_ ( .A(_05764_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05772_ ), .ZN(_05773_ ) );
XNOR2_X1 _13513_ ( .A(_05736_ ), .B(_02573_ ), .ZN(_05774_ ) );
AOI22_X1 _13514_ ( .A1(_05774_ ), .A2(_05579_ ), .B1(_05762_ ), .B2(_04020_ ), .ZN(_05775_ ) );
AOI21_X1 _13515_ ( .A(_05689_ ), .B1(_05773_ ), .B2(_05775_ ), .ZN(_00171_ ) );
NAND3_X1 _13516_ ( .A1(_05548_ ), .A2(\EX_LS_result_csreg_mem [9] ), .A3(_05549_ ), .ZN(_05776_ ) );
NAND3_X1 _13517_ ( .A1(_05656_ ), .A2(\mepc [9] ), .A3(_04082_ ), .ZN(_05777_ ) );
NAND3_X1 _13518_ ( .A1(_05654_ ), .A2(\mycsreg.CSReg[0][9] ), .A3(_05505_ ), .ZN(_05778_ ) );
NAND2_X1 _13519_ ( .A1(_05777_ ), .A2(_05778_ ), .ZN(_05779_ ) );
AND3_X1 _13520_ ( .A1(_04077_ ), .A2(\mycsreg.CSReg[3][9] ), .A3(_04086_ ), .ZN(_05780_ ) );
AND3_X1 _13521_ ( .A1(_05539_ ), .A2(\mtvec [9] ), .A3(_04096_ ), .ZN(_05781_ ) );
NOR4_X1 _13522_ ( .A1(_05779_ ), .A2(_05780_ ), .A3(_05495_ ), .A4(_05781_ ), .ZN(_05782_ ) );
OAI21_X1 _13523_ ( .A(_05776_ ), .B1(_05565_ ), .B2(_05782_ ), .ZN(_05783_ ) );
INV_X1 _13524_ ( .A(\ID_EX_pc [9] ), .ZN(_05784_ ) );
XNOR2_X1 _13525_ ( .A(_04116_ ), .B(_05784_ ), .ZN(_05785_ ) );
AND2_X1 _13526_ ( .A1(_04173_ ), .A2(_04185_ ), .ZN(_05786_ ) );
NOR2_X1 _13527_ ( .A1(_05786_ ), .A2(_04193_ ), .ZN(_05787_ ) );
XNOR2_X1 _13528_ ( .A(_05787_ ), .B(_04186_ ), .ZN(_05788_ ) );
MUX2_X1 _13529_ ( .A(_05785_ ), .B(_05788_ ), .S(_05419_ ), .Z(_05789_ ) );
MUX2_X1 _13530_ ( .A(_05783_ ), .B(_05789_ ), .S(_05422_ ), .Z(_05790_ ) );
NAND2_X1 _13531_ ( .A1(_05790_ ), .A2(_05426_ ), .ZN(_05791_ ) );
AOI21_X1 _13532_ ( .A(\ID_EX_imm [8] ), .B1(_02496_ ), .B2(_02497_ ), .ZN(_05792_ ) );
NOR3_X1 _13533_ ( .A1(_05734_ ), .A2(_02785_ ), .A3(_05792_ ), .ZN(_05793_ ) );
OR2_X1 _13534_ ( .A1(_05793_ ), .A2(_02785_ ), .ZN(_05794_ ) );
XNOR2_X1 _13535_ ( .A(_05794_ ), .B(_02524_ ), .ZN(_05795_ ) );
NOR3_X1 _13536_ ( .A1(_05795_ ), .A2(_05488_ ), .A3(_05425_ ), .ZN(_05796_ ) );
AOI21_X1 _13537_ ( .A(_05796_ ), .B1(_05521_ ), .B2(_05788_ ), .ZN(_05797_ ) );
AOI21_X1 _13538_ ( .A(_05689_ ), .B1(_05791_ ), .B2(_05797_ ), .ZN(_00172_ ) );
NAND3_X1 _13539_ ( .A1(_05498_ ), .A2(\mepc [8] ), .A3(_05543_ ), .ZN(_05798_ ) );
NAND3_X1 _13540_ ( .A1(_05498_ ), .A2(\mycsreg.CSReg[3][8] ), .A3(_04086_ ), .ZN(_05799_ ) );
NAND3_X1 _13541_ ( .A1(_04093_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_04105_ ), .ZN(_05800_ ) );
NAND3_X1 _13542_ ( .A1(_04093_ ), .A2(\mtvec [8] ), .A3(_04096_ ), .ZN(_05801_ ) );
AND4_X1 _13543_ ( .A1(_05798_ ), .A2(_05799_ ), .A3(_05800_ ), .A4(_05801_ ), .ZN(_05802_ ) );
NAND4_X1 _13544_ ( .A1(_04069_ ), .A2(_05722_ ), .A3(_05574_ ), .A4(_05802_ ), .ZN(_05803_ ) );
INV_X1 _13545_ ( .A(\EX_LS_result_csreg_mem [8] ), .ZN(_05804_ ) );
NAND3_X1 _13546_ ( .A1(_05490_ ), .A2(_05804_ ), .A3(_05492_ ), .ZN(_05805_ ) );
NAND2_X1 _13547_ ( .A1(_05803_ ), .A2(_05805_ ), .ZN(_05806_ ) );
AOI21_X1 _13548_ ( .A(_05648_ ), .B1(_05806_ ), .B2(\ID_EX_typ [3] ), .ZN(_05807_ ) );
INV_X1 _13549_ ( .A(\ID_EX_pc [8] ), .ZN(_05808_ ) );
XNOR2_X1 _13550_ ( .A(_04115_ ), .B(_05808_ ), .ZN(_05809_ ) );
XNOR2_X1 _13551_ ( .A(_04172_ ), .B(_04185_ ), .ZN(_05810_ ) );
MUX2_X1 _13552_ ( .A(_05809_ ), .B(_05810_ ), .S(_05461_ ), .Z(_05811_ ) );
OAI21_X1 _13553_ ( .A(_05807_ ), .B1(_05811_ ), .B2(\ID_EX_typ [3] ), .ZN(_05812_ ) );
XNOR2_X1 _13554_ ( .A(_05734_ ), .B(_02500_ ), .ZN(_05813_ ) );
AOI22_X1 _13555_ ( .A1(_05813_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05810_ ), .ZN(_05814_ ) );
AOI21_X1 _13556_ ( .A(_05689_ ), .B1(_05812_ ), .B2(_05814_ ), .ZN(_00173_ ) );
NOR2_X1 _13557_ ( .A1(_04171_ ), .A2(_04169_ ), .ZN(_05815_ ) );
XNOR2_X1 _13558_ ( .A(_04168_ ), .B(_05815_ ), .ZN(_05816_ ) );
AOI21_X1 _13559_ ( .A(\ID_EX_typ [3] ), .B1(_05461_ ), .B2(_05816_ ), .ZN(_05817_ ) );
XNOR2_X1 _13560_ ( .A(_04114_ ), .B(\ID_EX_pc [7] ), .ZN(_05818_ ) );
OAI21_X1 _13561_ ( .A(_05817_ ), .B1(_05462_ ), .B2(_05818_ ), .ZN(_05819_ ) );
NAND3_X1 _13562_ ( .A1(_05490_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_05492_ ), .ZN(_05820_ ) );
NAND3_X1 _13563_ ( .A1(_04077_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_04086_ ), .ZN(_05821_ ) );
NAND3_X1 _13564_ ( .A1(_04077_ ), .A2(\mepc [7] ), .A3(_05543_ ), .ZN(_05822_ ) );
NAND3_X1 _13565_ ( .A1(_05539_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_04105_ ), .ZN(_05823_ ) );
NAND3_X1 _13566_ ( .A1(_05539_ ), .A2(\mtvec [7] ), .A3(_04096_ ), .ZN(_05824_ ) );
AND4_X1 _13567_ ( .A1(_05821_ ), .A2(_05822_ ), .A3(_05823_ ), .A4(_05824_ ), .ZN(_05825_ ) );
OAI21_X1 _13568_ ( .A(_05820_ ), .B1(_05565_ ), .B2(_05825_ ), .ZN(_05826_ ) );
OAI211_X1 _13569_ ( .A(_05819_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05826_ ), .ZN(_05827_ ) );
OAI21_X1 _13570_ ( .A(_02680_ ), .B1(_02778_ ), .B2(_02782_ ), .ZN(_05828_ ) );
NAND2_X1 _13571_ ( .A1(_05828_ ), .A2(_02626_ ), .ZN(_05829_ ) );
NAND2_X1 _13572_ ( .A1(_05829_ ), .A2(_02672_ ), .ZN(_05830_ ) );
AND2_X1 _13573_ ( .A1(_05830_ ), .A2(_02675_ ), .ZN(_05831_ ) );
XNOR2_X1 _13574_ ( .A(_05831_ ), .B(_02681_ ), .ZN(_05832_ ) );
AOI22_X1 _13575_ ( .A1(_05832_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05816_ ), .ZN(_05833_ ) );
AOI21_X1 _13576_ ( .A(_05689_ ), .B1(_05827_ ), .B2(_05833_ ), .ZN(_00174_ ) );
INV_X1 _13577_ ( .A(\ID_EX_pc [6] ), .ZN(_05834_ ) );
XNOR2_X1 _13578_ ( .A(_04113_ ), .B(_05834_ ), .ZN(_05835_ ) );
XOR2_X1 _13579_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_05836_ ) );
XNOR2_X1 _13580_ ( .A(_04164_ ), .B(_05836_ ), .ZN(_05837_ ) );
MUX2_X1 _13581_ ( .A(_05835_ ), .B(_05837_ ), .S(_05419_ ), .Z(_05838_ ) );
OR2_X1 _13582_ ( .A1(_05838_ ), .A2(\ID_EX_typ [3] ), .ZN(_05839_ ) );
INV_X1 _13583_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_05840_ ) );
AND3_X1 _13584_ ( .A1(_05548_ ), .A2(_05840_ ), .A3(_05549_ ), .ZN(_05841_ ) );
NAND3_X1 _13585_ ( .A1(_05566_ ), .A2(\mycsreg.CSReg[3][6] ), .A3(_05572_ ), .ZN(_05842_ ) );
NAND3_X1 _13586_ ( .A1(_05566_ ), .A2(\mepc [6] ), .A3(_05544_ ), .ZN(_05843_ ) );
NAND3_X1 _13587_ ( .A1(_05568_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_04106_ ), .ZN(_05844_ ) );
NAND3_X1 _13588_ ( .A1(_05568_ ), .A2(\mtvec [6] ), .A3(_04097_ ), .ZN(_05845_ ) );
AND4_X1 _13589_ ( .A1(_05842_ ), .A2(_05843_ ), .A3(_05844_ ), .A4(_05845_ ), .ZN(_05846_ ) );
AOI21_X1 _13590_ ( .A(_05841_ ), .B1(_05494_ ), .B2(_05846_ ), .ZN(_05847_ ) );
OAI211_X1 _13591_ ( .A(_05839_ ), .B(_05535_ ), .C1(_05537_ ), .C2(_05847_ ), .ZN(_05848_ ) );
XNOR2_X1 _13592_ ( .A(_05829_ ), .B(_02673_ ), .ZN(_05849_ ) );
AOI22_X1 _13593_ ( .A1(_05849_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05837_ ), .ZN(_05850_ ) );
AOI21_X1 _13594_ ( .A(_05689_ ), .B1(_05848_ ), .B2(_05850_ ), .ZN(_00175_ ) );
NAND3_X1 _13595_ ( .A1(_05502_ ), .A2(\mycsreg.CSReg[3][5] ), .A3(_05500_ ), .ZN(_05851_ ) );
NAND3_X1 _13596_ ( .A1(_05502_ ), .A2(\mepc [5] ), .A3(_04082_ ), .ZN(_05852_ ) );
NAND2_X1 _13597_ ( .A1(_05851_ ), .A2(_05852_ ), .ZN(_05853_ ) );
AND3_X1 _13598_ ( .A1(_05654_ ), .A2(\mtvec [5] ), .A3(_04096_ ), .ZN(_05854_ ) );
AND3_X1 _13599_ ( .A1(_05539_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_05505_ ), .ZN(_05855_ ) );
NOR3_X1 _13600_ ( .A1(_05853_ ), .A2(_05854_ ), .A3(_05855_ ), .ZN(_05856_ ) );
NAND3_X1 _13601_ ( .A1(_04069_ ), .A2(_05722_ ), .A3(_05856_ ), .ZN(_05857_ ) );
INV_X1 _13602_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_05858_ ) );
NAND3_X1 _13603_ ( .A1(_05562_ ), .A2(_05858_ ), .A3(_05563_ ), .ZN(_05859_ ) );
AND2_X1 _13604_ ( .A1(_05857_ ), .A2(_05859_ ), .ZN(_05860_ ) );
XNOR2_X1 _13605_ ( .A(_04112_ ), .B(\ID_EX_pc [5] ), .ZN(_05861_ ) );
OAI21_X1 _13606_ ( .A(_05536_ ), .B1(_05462_ ), .B2(_05861_ ), .ZN(_05862_ ) );
NOR2_X1 _13607_ ( .A1(_04163_ ), .A2(_04161_ ), .ZN(_05863_ ) );
XNOR2_X1 _13608_ ( .A(_04160_ ), .B(_05863_ ), .ZN(_05864_ ) );
AND3_X1 _13609_ ( .A1(_05415_ ), .A2(_05417_ ), .A3(_05864_ ), .ZN(_05865_ ) );
OAI221_X1 _13610_ ( .A(_05582_ ), .B1(_05583_ ), .B2(_05860_ ), .C1(_05862_ ), .C2(_05865_ ), .ZN(_05866_ ) );
NOR2_X1 _13611_ ( .A1(_02778_ ), .A2(_02782_ ), .ZN(_05867_ ) );
NOR2_X1 _13612_ ( .A1(_05867_ ), .A2(_02679_ ), .ZN(_05868_ ) );
AND3_X1 _13613_ ( .A1(_02620_ ), .A2(\ID_EX_imm [4] ), .A3(_02621_ ), .ZN(_05869_ ) );
OR2_X1 _13614_ ( .A1(_05868_ ), .A2(_05869_ ), .ZN(_05870_ ) );
XNOR2_X1 _13615_ ( .A(_05870_ ), .B(_02599_ ), .ZN(_05871_ ) );
AOI22_X1 _13616_ ( .A1(_05871_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05864_ ), .ZN(_05872_ ) );
AOI21_X1 _13617_ ( .A(_05689_ ), .B1(_05866_ ), .B2(_05872_ ), .ZN(_00176_ ) );
XNOR2_X1 _13618_ ( .A(_04111_ ), .B(\ID_EX_pc [4] ), .ZN(_05873_ ) );
XOR2_X1 _13619_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_05874_ ) );
XNOR2_X1 _13620_ ( .A(_04156_ ), .B(_05874_ ), .ZN(_05875_ ) );
INV_X1 _13621_ ( .A(_05875_ ), .ZN(_05876_ ) );
MUX2_X1 _13622_ ( .A(_05873_ ), .B(_05876_ ), .S(_05461_ ), .Z(_05877_ ) );
NAND2_X1 _13623_ ( .A1(_05877_ ), .A2(_05583_ ), .ZN(_05878_ ) );
AND3_X1 _13624_ ( .A1(_04092_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_04104_ ), .ZN(_05879_ ) );
NAND3_X1 _13625_ ( .A1(_05498_ ), .A2(\mycsreg.CSReg[3][4] ), .A3(_04085_ ), .ZN(_05880_ ) );
NAND3_X1 _13626_ ( .A1(_04076_ ), .A2(\mepc [4] ), .A3(_05543_ ), .ZN(_05881_ ) );
NAND3_X1 _13627_ ( .A1(_04092_ ), .A2(\mtvec [4] ), .A3(_04095_ ), .ZN(_05882_ ) );
NAND4_X1 _13628_ ( .A1(_05880_ ), .A2(_05881_ ), .A3(_05882_ ), .A4(_05722_ ), .ZN(_05883_ ) );
AOI211_X1 _13629_ ( .A(_05879_ ), .B(_05883_ ), .C1(_05478_ ), .C2(_05699_ ), .ZN(_05884_ ) );
INV_X1 _13630_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_05885_ ) );
AND4_X1 _13631_ ( .A1(_05885_ ), .A2(_05704_ ), .A3(_05706_ ), .A4(_05699_ ), .ZN(_05886_ ) );
NOR2_X1 _13632_ ( .A1(_05884_ ), .A2(_05886_ ), .ZN(_05887_ ) );
OAI211_X1 _13633_ ( .A(_05878_ ), .B(_05582_ ), .C1(_05537_ ), .C2(_05887_ ), .ZN(_05888_ ) );
XNOR2_X1 _13634_ ( .A(_05867_ ), .B(_02678_ ), .ZN(_05889_ ) );
AOI22_X1 _13635_ ( .A1(_05889_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05875_ ), .ZN(_05890_ ) );
AOI21_X1 _13636_ ( .A(_05689_ ), .B1(_05888_ ), .B2(_05890_ ), .ZN(_00177_ ) );
BUF_X4 _13637_ ( .A(_04031_ ), .Z(_05891_ ) );
NAND3_X1 _13638_ ( .A1(_05498_ ), .A2(\mepc [3] ), .A3(_05543_ ), .ZN(_05892_ ) );
NAND3_X1 _13639_ ( .A1(_04093_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_04105_ ), .ZN(_05893_ ) );
AND2_X1 _13640_ ( .A1(_05892_ ), .A2(_05893_ ), .ZN(_05894_ ) );
NAND3_X1 _13641_ ( .A1(_05654_ ), .A2(\mtvec [3] ), .A3(_05507_ ), .ZN(_05895_ ) );
NAND3_X1 _13642_ ( .A1(_05656_ ), .A2(\mycsreg.CSReg[3][3] ), .A3(_04086_ ), .ZN(_05896_ ) );
AND4_X1 _13643_ ( .A1(_05494_ ), .A2(_05894_ ), .A3(_05895_ ), .A4(_05896_ ), .ZN(_05897_ ) );
INV_X1 _13644_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_05898_ ) );
AND3_X1 _13645_ ( .A1(_05490_ ), .A2(_05898_ ), .A3(_05492_ ), .ZN(_05899_ ) );
NOR2_X1 _13646_ ( .A1(_05897_ ), .A2(_05899_ ), .ZN(_05900_ ) );
XNOR2_X1 _13647_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .ZN(_05901_ ) );
OAI21_X1 _13648_ ( .A(_05536_ ), .B1(_05462_ ), .B2(_05901_ ), .ZN(_05902_ ) );
NOR2_X1 _13649_ ( .A1(_04155_ ), .A2(_04153_ ), .ZN(_05903_ ) );
XNOR2_X1 _13650_ ( .A(_04152_ ), .B(_05903_ ), .ZN(_05904_ ) );
AND3_X1 _13651_ ( .A1(_05415_ ), .A2(_05417_ ), .A3(_05904_ ), .ZN(_05905_ ) );
OAI221_X1 _13652_ ( .A(_05582_ ), .B1(_05583_ ), .B2(_05900_ ), .C1(_05902_ ), .C2(_05905_ ), .ZN(_05906_ ) );
OAI21_X1 _13653_ ( .A(_02780_ ), .B1(_02730_ ), .B2(_02777_ ), .ZN(_05907_ ) );
XNOR2_X1 _13654_ ( .A(_05907_ ), .B(_02753_ ), .ZN(_05908_ ) );
AOI22_X1 _13655_ ( .A1(_05908_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05904_ ), .ZN(_05909_ ) );
AOI21_X1 _13656_ ( .A(_05891_ ), .B1(_05906_ ), .B2(_05909_ ), .ZN(_00178_ ) );
NAND3_X1 _13657_ ( .A1(_05562_ ), .A2(\EX_LS_result_csreg_mem [2] ), .A3(_05563_ ), .ZN(_05910_ ) );
AND3_X1 _13658_ ( .A1(_05539_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_04105_ ), .ZN(_05911_ ) );
INV_X1 _13659_ ( .A(_05911_ ), .ZN(_05912_ ) );
NAND3_X1 _13660_ ( .A1(_05499_ ), .A2(\mepc [2] ), .A3(_05544_ ), .ZN(_05913_ ) );
NAND3_X1 _13661_ ( .A1(_05499_ ), .A2(\mycsreg.CSReg[3][2] ), .A3(_05572_ ), .ZN(_05914_ ) );
NAND3_X1 _13662_ ( .A1(_05912_ ), .A2(_05913_ ), .A3(_05914_ ), .ZN(_05915_ ) );
NAND3_X1 _13663_ ( .A1(_04094_ ), .A2(\mtvec [2] ), .A3(_04097_ ), .ZN(_05916_ ) );
NAND2_X1 _13664_ ( .A1(_05574_ ), .A2(_05916_ ), .ZN(_05917_ ) );
NOR2_X1 _13665_ ( .A1(_05915_ ), .A2(_05917_ ), .ZN(_05918_ ) );
OAI21_X1 _13666_ ( .A(_05910_ ), .B1(_05565_ ), .B2(_05918_ ), .ZN(_05919_ ) );
AOI211_X1 _13667_ ( .A(_04148_ ), .B(_04144_ ), .C1(_04146_ ), .C2(_04145_ ), .ZN(_05920_ ) );
NOR2_X1 _13668_ ( .A1(_04150_ ), .A2(_05920_ ), .ZN(_05921_ ) );
MUX2_X1 _13669_ ( .A(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .B(_05921_ ), .S(_05419_ ), .Z(_05922_ ) );
MUX2_X1 _13670_ ( .A(_05919_ ), .B(_05922_ ), .S(_05422_ ), .Z(_05923_ ) );
NAND2_X1 _13671_ ( .A1(_05923_ ), .A2(_05426_ ), .ZN(_05924_ ) );
XNOR2_X1 _13672_ ( .A(_02730_ ), .B(_02776_ ), .ZN(_05925_ ) );
AOI22_X1 _13673_ ( .A1(_05925_ ), .A2(_05579_ ), .B1(_05580_ ), .B2(_05921_ ), .ZN(_05926_ ) );
AOI21_X1 _13674_ ( .A(_05891_ ), .B1(_05924_ ), .B2(_05926_ ), .ZN(_00179_ ) );
XOR2_X1 _13675_ ( .A(_04145_ ), .B(_04146_ ), .Z(_05927_ ) );
AOI21_X1 _13676_ ( .A(\ID_EX_typ [3] ), .B1(_05461_ ), .B2(_05927_ ), .ZN(_05928_ ) );
INV_X1 _13677_ ( .A(\ID_EX_pc [1] ), .ZN(_05929_ ) );
OAI21_X1 _13678_ ( .A(_05928_ ), .B1(_05929_ ), .B2(_05462_ ), .ZN(_05930_ ) );
NAND3_X1 _13679_ ( .A1(_05498_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_04086_ ), .ZN(_05931_ ) );
NAND3_X1 _13680_ ( .A1(_05498_ ), .A2(\mepc [1] ), .A3(_05543_ ), .ZN(_05932_ ) );
NAND3_X1 _13681_ ( .A1(_04093_ ), .A2(\mtvec [1] ), .A3(_04096_ ), .ZN(_05933_ ) );
NAND3_X1 _13682_ ( .A1(_04092_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_04104_ ), .ZN(_05934_ ) );
AND4_X1 _13683_ ( .A1(_05931_ ), .A2(_05932_ ), .A3(_05933_ ), .A4(_05934_ ), .ZN(_05935_ ) );
OR2_X1 _13684_ ( .A1(_05565_ ), .A2(_05935_ ), .ZN(_05936_ ) );
NAND3_X1 _13685_ ( .A1(_05548_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_05549_ ), .ZN(_05937_ ) );
AND2_X1 _13686_ ( .A1(_05936_ ), .A2(_05937_ ), .ZN(_05938_ ) );
INV_X1 _13687_ ( .A(_05938_ ), .ZN(_05939_ ) );
OAI211_X1 _13688_ ( .A(_05930_ ), .B(_05582_ ), .C1(_05537_ ), .C2(_05939_ ), .ZN(_05940_ ) );
XOR2_X1 _13689_ ( .A(_02706_ ), .B(_02728_ ), .Z(_05941_ ) );
AOI22_X1 _13690_ ( .A1(_05941_ ), .A2(_05519_ ), .B1(_05580_ ), .B2(_05927_ ), .ZN(_05942_ ) );
AOI21_X1 _13691_ ( .A(_05891_ ), .B1(_05940_ ), .B2(_05942_ ), .ZN(_00180_ ) );
NAND3_X1 _13692_ ( .A1(_05438_ ), .A2(\ID_EX_pc [26] ), .A3(_05441_ ), .ZN(_05943_ ) );
XNOR2_X1 _13693_ ( .A(_05943_ ), .B(\ID_EX_pc [27] ), .ZN(_05944_ ) );
NAND2_X1 _13694_ ( .A1(_05435_ ), .A2(_05944_ ), .ZN(_05945_ ) );
AND2_X1 _13695_ ( .A1(_04227_ ), .A2(_04235_ ), .ZN(_05946_ ) );
OAI21_X1 _13696_ ( .A(_04229_ ), .B1(_05946_ ), .B2(_04241_ ), .ZN(_05947_ ) );
NAND2_X1 _13697_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_05948_ ) );
NAND2_X1 _13698_ ( .A1(_05947_ ), .A2(_05948_ ), .ZN(_05949_ ) );
XNOR2_X1 _13699_ ( .A(_05949_ ), .B(_04228_ ), .ZN(_05950_ ) );
OAI211_X1 _13700_ ( .A(_05945_ ), .B(_05536_ ), .C1(_05435_ ), .C2(_05950_ ), .ZN(_05951_ ) );
INV_X1 _13701_ ( .A(\EX_LS_result_csreg_mem [27] ), .ZN(_05952_ ) );
AND3_X1 _13702_ ( .A1(_05562_ ), .A2(_05952_ ), .A3(_05563_ ), .ZN(_05953_ ) );
NAND3_X1 _13703_ ( .A1(_05566_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_05572_ ), .ZN(_05954_ ) );
NAND3_X1 _13704_ ( .A1(_05499_ ), .A2(\mepc [27] ), .A3(_05544_ ), .ZN(_05955_ ) );
NAND2_X1 _13705_ ( .A1(_05954_ ), .A2(_05955_ ), .ZN(_05956_ ) );
AND3_X1 _13706_ ( .A1(_05568_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_04106_ ), .ZN(_05957_ ) );
AND3_X1 _13707_ ( .A1(_05504_ ), .A2(\mtvec [27] ), .A3(_05507_ ), .ZN(_05958_ ) );
NOR3_X1 _13708_ ( .A1(_05956_ ), .A2(_05957_ ), .A3(_05958_ ), .ZN(_05959_ ) );
AOI21_X1 _13709_ ( .A(_05953_ ), .B1(_05494_ ), .B2(_05959_ ), .ZN(_05960_ ) );
OAI211_X1 _13710_ ( .A(_05951_ ), .B(_05582_ ), .C1(_05583_ ), .C2(_05960_ ), .ZN(_05961_ ) );
MUX2_X1 _13711_ ( .A(_05950_ ), .B(_03192_ ), .S(fanout_net_7 ), .Z(_05962_ ) );
BUF_X2 _13712_ ( .A(_05424_ ), .Z(_05963_ ) );
OR2_X1 _13713_ ( .A1(_05962_ ), .A2(_05963_ ), .ZN(_05964_ ) );
AOI21_X1 _13714_ ( .A(_05891_ ), .B1(_05961_ ), .B2(_05964_ ), .ZN(_00181_ ) );
XOR2_X1 _13715_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05965_ ) );
OAI21_X1 _13716_ ( .A(_05422_ ), .B1(_05435_ ), .B2(_05965_ ), .ZN(_05966_ ) );
INV_X1 _13717_ ( .A(\ID_EX_pc [0] ), .ZN(_05967_ ) );
AOI21_X1 _13718_ ( .A(_05966_ ), .B1(_05967_ ), .B2(_05435_ ), .ZN(_05968_ ) );
AND3_X1 _13719_ ( .A1(_04091_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_04104_ ), .ZN(_05969_ ) );
INV_X1 _13720_ ( .A(_05969_ ), .ZN(_05970_ ) );
NAND3_X1 _13721_ ( .A1(_04076_ ), .A2(\mepc [0] ), .A3(_04081_ ), .ZN(_05971_ ) );
NAND3_X1 _13722_ ( .A1(_04076_ ), .A2(\mycsreg.CSReg[3][0] ), .A3(_04085_ ), .ZN(_05972_ ) );
NAND3_X1 _13723_ ( .A1(_05970_ ), .A2(_05971_ ), .A3(_05972_ ), .ZN(_05973_ ) );
NAND3_X1 _13724_ ( .A1(_04092_ ), .A2(\mtvec [0] ), .A3(_04095_ ), .ZN(_05974_ ) );
NAND2_X1 _13725_ ( .A1(_05496_ ), .A2(_05974_ ), .ZN(_05975_ ) );
NOR2_X1 _13726_ ( .A1(_05973_ ), .A2(_05975_ ), .ZN(_05976_ ) );
OR2_X1 _13727_ ( .A1(_05565_ ), .A2(_05976_ ), .ZN(_05977_ ) );
NAND3_X1 _13728_ ( .A1(_05490_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_05492_ ), .ZN(_05978_ ) );
AOI21_X1 _13729_ ( .A(_05536_ ), .B1(_05977_ ), .B2(_05978_ ), .ZN(_05979_ ) );
OAI21_X1 _13730_ ( .A(_05426_ ), .B1(_05968_ ), .B2(_05979_ ), .ZN(_05980_ ) );
BUF_X4 _13731_ ( .A(_05487_ ), .Z(_05981_ ) );
NAND3_X1 _13732_ ( .A1(_05965_ ), .A2(_05981_ ), .A3(_05431_ ), .ZN(_05982_ ) );
AOI21_X1 _13733_ ( .A(_05891_ ), .B1(_05980_ ), .B2(_05982_ ), .ZN(_00182_ ) );
AND2_X2 _13734_ ( .A1(_05477_ ), .A2(_05474_ ), .ZN(_05983_ ) );
INV_X1 _13735_ ( .A(_05983_ ), .ZN(_05984_ ) );
NOR2_X1 _13736_ ( .A1(_05984_ ), .A2(\EX_LS_result_csreg_mem [26] ), .ZN(_05985_ ) );
NAND3_X1 _13737_ ( .A1(_05656_ ), .A2(\mycsreg.CSReg[3][26] ), .A3(_05500_ ), .ZN(_05986_ ) );
NAND3_X1 _13738_ ( .A1(_05656_ ), .A2(\mepc [26] ), .A3(_04082_ ), .ZN(_05987_ ) );
NAND3_X1 _13739_ ( .A1(_05654_ ), .A2(\mtvec [26] ), .A3(_05507_ ), .ZN(_05988_ ) );
NAND3_X1 _13740_ ( .A1(_05654_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_05505_ ), .ZN(_05989_ ) );
NAND4_X1 _13741_ ( .A1(_05986_ ), .A2(_05987_ ), .A3(_05988_ ), .A4(_05989_ ), .ZN(_05990_ ) );
AOI21_X1 _13742_ ( .A(_05990_ ), .B1(_05478_ ), .B2(_05479_ ), .ZN(_05991_ ) );
NOR2_X1 _13743_ ( .A1(_05985_ ), .A2(_05991_ ), .ZN(_05992_ ) );
INV_X1 _13744_ ( .A(\ID_EX_pc [26] ), .ZN(_05993_ ) );
XNOR2_X1 _13745_ ( .A(_05442_ ), .B(_05993_ ), .ZN(_05994_ ) );
OR3_X1 _13746_ ( .A1(_05946_ ), .A2(_04229_ ), .A3(_04241_ ), .ZN(_05995_ ) );
AND2_X1 _13747_ ( .A1(_05995_ ), .A2(_05947_ ), .ZN(_05996_ ) );
MUX2_X1 _13748_ ( .A(_05994_ ), .B(_05996_ ), .S(_05418_ ), .Z(_05997_ ) );
MUX2_X1 _13749_ ( .A(_05992_ ), .B(_05997_ ), .S(_05422_ ), .Z(_05998_ ) );
NAND2_X1 _13750_ ( .A1(_05998_ ), .A2(_05426_ ), .ZN(_05999_ ) );
OAI21_X1 _13751_ ( .A(fanout_net_7 ), .B1(_03190_ ), .B2(_03193_ ), .ZN(_06000_ ) );
OAI211_X1 _13752_ ( .A(_06000_ ), .B(_05431_ ), .C1(fanout_net_7 ), .C2(_05996_ ), .ZN(_06001_ ) );
AOI21_X1 _13753_ ( .A(_05891_ ), .B1(_05999_ ), .B2(_06001_ ), .ZN(_00183_ ) );
AND3_X1 _13754_ ( .A1(_05440_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_06002_ ) );
AND2_X1 _13755_ ( .A1(_05438_ ), .A2(_06002_ ), .ZN(_06003_ ) );
NAND3_X1 _13756_ ( .A1(_06003_ ), .A2(\ID_EX_pc [23] ), .A3(\ID_EX_pc [22] ), .ZN(_06004_ ) );
INV_X1 _13757_ ( .A(\ID_EX_pc [24] ), .ZN(_06005_ ) );
NOR2_X1 _13758_ ( .A1(_06004_ ), .A2(_06005_ ), .ZN(_06006_ ) );
XNOR2_X1 _13759_ ( .A(_06006_ ), .B(_04240_ ), .ZN(_06007_ ) );
NAND2_X1 _13760_ ( .A1(_04227_ ), .A2(_04231_ ), .ZN(_06008_ ) );
AND2_X1 _13761_ ( .A1(_06008_ ), .A2(_04238_ ), .ZN(_06009_ ) );
XNOR2_X1 _13762_ ( .A(_06009_ ), .B(_04234_ ), .ZN(_06010_ ) );
MUX2_X1 _13763_ ( .A(_06007_ ), .B(_06010_ ), .S(_05419_ ), .Z(_06011_ ) );
OR2_X1 _13764_ ( .A1(_06011_ ), .A2(\ID_EX_typ [3] ), .ZN(_06012_ ) );
NAND3_X1 _13765_ ( .A1(_05562_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_05563_ ), .ZN(_06013_ ) );
NAND3_X1 _13766_ ( .A1(_05502_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_05500_ ), .ZN(_06014_ ) );
NAND3_X1 _13767_ ( .A1(_05502_ ), .A2(\mepc [25] ), .A3(_04082_ ), .ZN(_06015_ ) );
NAND3_X1 _13768_ ( .A1(_05504_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_05505_ ), .ZN(_06016_ ) );
NAND3_X1 _13769_ ( .A1(_05504_ ), .A2(\mtvec [25] ), .A3(_05507_ ), .ZN(_06017_ ) );
AND4_X1 _13770_ ( .A1(_06014_ ), .A2(_06015_ ), .A3(_06016_ ), .A4(_06017_ ), .ZN(_06018_ ) );
OAI21_X1 _13771_ ( .A(_06013_ ), .B1(_05565_ ), .B2(_06018_ ), .ZN(_06019_ ) );
OAI211_X1 _13772_ ( .A(_06012_ ), .B(_05582_ ), .C1(_05583_ ), .C2(_06019_ ), .ZN(_06020_ ) );
NOR3_X1 _13773_ ( .A1(_03195_ ), .A2(_05488_ ), .A3(_05425_ ), .ZN(_06021_ ) );
AOI21_X1 _13774_ ( .A(_06021_ ), .B1(_05521_ ), .B2(_06010_ ), .ZN(_06022_ ) );
AOI21_X1 _13775_ ( .A(_05891_ ), .B1(_06020_ ), .B2(_06022_ ), .ZN(_00184_ ) );
XOR2_X1 _13776_ ( .A(_04227_ ), .B(_04231_ ), .Z(_06023_ ) );
AOI21_X1 _13777_ ( .A(\ID_EX_typ [3] ), .B1(_05461_ ), .B2(_06023_ ), .ZN(_06024_ ) );
XNOR2_X1 _13778_ ( .A(_06004_ ), .B(_06005_ ), .ZN(_06025_ ) );
OAI21_X1 _13779_ ( .A(_06024_ ), .B1(_05462_ ), .B2(_06025_ ), .ZN(_06026_ ) );
OR2_X1 _13780_ ( .A1(_04069_ ), .A2(\EX_LS_result_csreg_mem [24] ), .ZN(_06027_ ) );
NAND3_X1 _13781_ ( .A1(_05656_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_05500_ ), .ZN(_06028_ ) );
NAND3_X1 _13782_ ( .A1(_05656_ ), .A2(\mepc [24] ), .A3(_04082_ ), .ZN(_06029_ ) );
NAND3_X1 _13783_ ( .A1(_05654_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_05505_ ), .ZN(_06030_ ) );
NAND3_X1 _13784_ ( .A1(_05539_ ), .A2(\mtvec [24] ), .A3(_04096_ ), .ZN(_06031_ ) );
AND4_X1 _13785_ ( .A1(_06028_ ), .A2(_06029_ ), .A3(_06030_ ), .A4(_06031_ ), .ZN(_06032_ ) );
NAND4_X1 _13786_ ( .A1(_04069_ ), .A2(_05722_ ), .A3(_05574_ ), .A4(_06032_ ), .ZN(_06033_ ) );
AND2_X1 _13787_ ( .A1(_06027_ ), .A2(_06033_ ), .ZN(_06034_ ) );
OAI211_X1 _13788_ ( .A(_06026_ ), .B(_05582_ ), .C1(_05583_ ), .C2(_06034_ ), .ZN(_06035_ ) );
AOI22_X1 _13789_ ( .A1(_03199_ ), .A2(_05519_ ), .B1(_06023_ ), .B2(_04020_ ), .ZN(_06036_ ) );
AOI21_X1 _13790_ ( .A(_05891_ ), .B1(_06035_ ), .B2(_06036_ ), .ZN(_00185_ ) );
NAND2_X1 _13791_ ( .A1(_05514_ ), .A2(_04136_ ), .ZN(_06037_ ) );
NAND2_X1 _13792_ ( .A1(_06037_ ), .A2(_04224_ ), .ZN(_06038_ ) );
NAND2_X1 _13793_ ( .A1(_06038_ ), .A2(_04132_ ), .ZN(_06039_ ) );
NAND2_X1 _13794_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_06040_ ) );
AND2_X1 _13795_ ( .A1(_06039_ ), .A2(_06040_ ), .ZN(_06041_ ) );
XNOR2_X1 _13796_ ( .A(_06041_ ), .B(_04131_ ), .ZN(_06042_ ) );
NAND3_X1 _13797_ ( .A1(_05415_ ), .A2(_05417_ ), .A3(_06042_ ), .ZN(_06043_ ) );
NAND3_X1 _13798_ ( .A1(_05438_ ), .A2(\ID_EX_pc [22] ), .A3(_06002_ ), .ZN(_06044_ ) );
XNOR2_X1 _13799_ ( .A(_06044_ ), .B(_04211_ ), .ZN(_06045_ ) );
OAI211_X1 _13800_ ( .A(_05536_ ), .B(_06043_ ), .C1(_05462_ ), .C2(_06045_ ), .ZN(_06046_ ) );
NAND3_X1 _13801_ ( .A1(_05566_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_05572_ ), .ZN(_06047_ ) );
NAND3_X1 _13802_ ( .A1(_05566_ ), .A2(\mepc [23] ), .A3(_05544_ ), .ZN(_06048_ ) );
NAND3_X1 _13803_ ( .A1(_05568_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_04106_ ), .ZN(_06049_ ) );
NAND3_X1 _13804_ ( .A1(_05568_ ), .A2(\mtvec [23] ), .A3(_04097_ ), .ZN(_06050_ ) );
NAND4_X1 _13805_ ( .A1(_06047_ ), .A2(_06048_ ), .A3(_06049_ ), .A4(_06050_ ), .ZN(_06051_ ) );
MUX2_X1 _13806_ ( .A(_06051_ ), .B(\EX_LS_result_csreg_mem [23] ), .S(_05983_ ), .Z(_06052_ ) );
OAI211_X1 _13807_ ( .A(_06046_ ), .B(_05582_ ), .C1(_05583_ ), .C2(_06052_ ), .ZN(_06053_ ) );
NAND2_X1 _13808_ ( .A1(_03205_ ), .A2(fanout_net_7 ), .ZN(_06054_ ) );
OAI211_X1 _13809_ ( .A(_06054_ ), .B(_05431_ ), .C1(fanout_net_7 ), .C2(_06042_ ), .ZN(_06055_ ) );
AOI21_X1 _13810_ ( .A(_05891_ ), .B1(_06053_ ), .B2(_06055_ ), .ZN(_00186_ ) );
BUF_X4 _13811_ ( .A(_05425_ ), .Z(_06056_ ) );
INV_X1 _13812_ ( .A(\EX_LS_result_csreg_mem [22] ), .ZN(_06057_ ) );
AND3_X1 _13813_ ( .A1(_05548_ ), .A2(_06057_ ), .A3(_05549_ ), .ZN(_06058_ ) );
NAND3_X1 _13814_ ( .A1(_05656_ ), .A2(\mepc [22] ), .A3(_04082_ ), .ZN(_06059_ ) );
NAND3_X1 _13815_ ( .A1(_05504_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_05505_ ), .ZN(_06060_ ) );
NAND2_X1 _13816_ ( .A1(_06059_ ), .A2(_06060_ ), .ZN(_06061_ ) );
AND3_X1 _13817_ ( .A1(_05499_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_05572_ ), .ZN(_06062_ ) );
AND3_X1 _13818_ ( .A1(_04094_ ), .A2(\mtvec [22] ), .A3(_04097_ ), .ZN(_06063_ ) );
NOR3_X1 _13819_ ( .A1(_06061_ ), .A2(_06062_ ), .A3(_06063_ ), .ZN(_06064_ ) );
AOI21_X1 _13820_ ( .A(_06058_ ), .B1(_05497_ ), .B2(_06064_ ), .ZN(_06065_ ) );
XNOR2_X1 _13821_ ( .A(_06003_ ), .B(\ID_EX_pc [22] ), .ZN(_06066_ ) );
OAI21_X1 _13822_ ( .A(_05536_ ), .B1(_05462_ ), .B2(_06066_ ), .ZN(_06067_ ) );
XOR2_X1 _13823_ ( .A(_06038_ ), .B(_04132_ ), .Z(_06068_ ) );
AND3_X1 _13824_ ( .A1(_05415_ ), .A2(_05417_ ), .A3(_06068_ ), .ZN(_06069_ ) );
OAI221_X1 _13825_ ( .A(_06056_ ), .B1(_05583_ ), .B2(_06065_ ), .C1(_06067_ ), .C2(_06069_ ), .ZN(_06070_ ) );
AOI22_X1 _13826_ ( .A1(_03206_ ), .A2(_05519_ ), .B1(_05580_ ), .B2(_06068_ ), .ZN(_06071_ ) );
AOI21_X1 _13827_ ( .A(_05891_ ), .B1(_06070_ ), .B2(_06071_ ), .ZN(_00187_ ) );
INV_X1 _13828_ ( .A(\EX_LS_result_csreg_mem [21] ), .ZN(_06072_ ) );
AND3_X1 _13829_ ( .A1(_05490_ ), .A2(_06072_ ), .A3(_05492_ ), .ZN(_06073_ ) );
NAND3_X1 _13830_ ( .A1(_05504_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_05505_ ), .ZN(_06074_ ) );
NAND3_X1 _13831_ ( .A1(_05502_ ), .A2(\mepc [21] ), .A3(_04082_ ), .ZN(_06075_ ) );
NAND3_X1 _13832_ ( .A1(_05656_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_05500_ ), .ZN(_06076_ ) );
NAND3_X1 _13833_ ( .A1(_05504_ ), .A2(\mtvec [21] ), .A3(_05507_ ), .ZN(_06077_ ) );
AND4_X1 _13834_ ( .A1(_06074_ ), .A2(_06075_ ), .A3(_06076_ ), .A4(_06077_ ), .ZN(_06078_ ) );
AOI21_X1 _13835_ ( .A(_06073_ ), .B1(_05494_ ), .B2(_06078_ ), .ZN(_06079_ ) );
INV_X1 _13836_ ( .A(\ID_EX_pc [20] ), .ZN(_06080_ ) );
NOR2_X1 _13837_ ( .A1(_05511_ ), .A2(_06080_ ), .ZN(_06081_ ) );
INV_X1 _13838_ ( .A(\ID_EX_pc [21] ), .ZN(_06082_ ) );
XNOR2_X1 _13839_ ( .A(_06081_ ), .B(_06082_ ), .ZN(_06083_ ) );
AND2_X1 _13840_ ( .A1(_05514_ ), .A2(_04134_ ), .ZN(_06084_ ) );
NOR2_X1 _13841_ ( .A1(_06084_ ), .A2(_04223_ ), .ZN(_06085_ ) );
XNOR2_X1 _13842_ ( .A(_06085_ ), .B(_04135_ ), .ZN(_06086_ ) );
MUX2_X1 _13843_ ( .A(_06083_ ), .B(_06086_ ), .S(_05418_ ), .Z(_06087_ ) );
MUX2_X1 _13844_ ( .A(_06079_ ), .B(_06087_ ), .S(_05422_ ), .Z(_06088_ ) );
NAND2_X1 _13845_ ( .A1(_06088_ ), .A2(_05426_ ), .ZN(_06089_ ) );
NOR3_X1 _13846_ ( .A1(_03162_ ), .A2(_05488_ ), .A3(_05424_ ), .ZN(_06090_ ) );
AOI21_X1 _13847_ ( .A(_06090_ ), .B1(_05521_ ), .B2(_06086_ ), .ZN(_06091_ ) );
AOI21_X1 _13848_ ( .A(_04031_ ), .B1(_06089_ ), .B2(_06091_ ), .ZN(_00188_ ) );
NOR3_X1 _13849_ ( .A1(_03152_ ), .A2(_05428_ ), .A3(_05424_ ), .ZN(_06092_ ) );
OAI21_X1 _13850_ ( .A(_04251_ ), .B1(_04248_ ), .B2(_04249_ ), .ZN(_06093_ ) );
NAND2_X1 _13851_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_06094_ ) );
NAND2_X1 _13852_ ( .A1(_06093_ ), .A2(_06094_ ), .ZN(_06095_ ) );
XNOR2_X1 _13853_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_06096_ ) );
XOR2_X1 _13854_ ( .A(_06095_ ), .B(_06096_ ), .Z(_06097_ ) );
NAND3_X1 _13855_ ( .A1(_05490_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_05492_ ), .ZN(_06098_ ) );
NAND3_X1 _13856_ ( .A1(_05498_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_04086_ ), .ZN(_06099_ ) );
NAND3_X1 _13857_ ( .A1(_05498_ ), .A2(\mepc [31] ), .A3(_05543_ ), .ZN(_06100_ ) );
NAND3_X1 _13858_ ( .A1(_04093_ ), .A2(\mtvec [31] ), .A3(_04096_ ), .ZN(_06101_ ) );
NAND3_X1 _13859_ ( .A1(_04093_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04105_ ), .ZN(_06102_ ) );
AND4_X1 _13860_ ( .A1(_06099_ ), .A2(_06100_ ), .A3(_06101_ ), .A4(_06102_ ), .ZN(_06103_ ) );
OAI21_X1 _13861_ ( .A(_06098_ ), .B1(_05565_ ), .B2(_06103_ ), .ZN(_06104_ ) );
OAI211_X1 _13862_ ( .A(_05461_ ), .B(_05424_ ), .C1(_05421_ ), .C2(_06104_ ), .ZN(_06105_ ) );
AOI21_X1 _13863_ ( .A(_06097_ ), .B1(_06105_ ), .B2(_05484_ ), .ZN(_06106_ ) );
AND3_X1 _13864_ ( .A1(_04128_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_06107_ ) );
NAND2_X1 _13865_ ( .A1(_06107_ ), .A2(\ID_EX_pc [30] ), .ZN(_06108_ ) );
XNOR2_X1 _13866_ ( .A(_06108_ ), .B(\ID_EX_pc [31] ), .ZN(_06109_ ) );
AOI21_X1 _13867_ ( .A(\ID_EX_typ [3] ), .B1(_05434_ ), .B2(_06109_ ), .ZN(_06110_ ) );
NAND4_X1 _13868_ ( .A1(_06099_ ), .A2(_06100_ ), .A3(_06101_ ), .A4(_06102_ ), .ZN(_06111_ ) );
OR2_X1 _13869_ ( .A1(_05983_ ), .A2(_06111_ ), .ZN(_06112_ ) );
OAI21_X1 _13870_ ( .A(_06112_ ), .B1(\EX_LS_result_csreg_mem [31] ), .B2(_05984_ ), .ZN(_06113_ ) );
AOI211_X1 _13871_ ( .A(_04018_ ), .B(_06110_ ), .C1(\ID_EX_typ [3] ), .C2(_06113_ ), .ZN(_06114_ ) );
OR4_X1 _13872_ ( .A1(_04031_ ), .A2(_06092_ ), .A3(_06106_ ), .A4(_06114_ ), .ZN(_00189_ ) );
AND3_X1 _13873_ ( .A1(_04030_ ), .A2(\ID_EX_pc [31] ), .A3(_03239_ ), .ZN(_00190_ ) );
AND3_X1 _13874_ ( .A1(_04030_ ), .A2(\ID_EX_pc [30] ), .A3(_03239_ ), .ZN(_00191_ ) );
CLKBUF_X2 _13875_ ( .A(_03221_ ), .Z(_06115_ ) );
AND3_X1 _13876_ ( .A1(_04030_ ), .A2(\ID_EX_pc [21] ), .A3(_06115_ ), .ZN(_00192_ ) );
AND3_X1 _13877_ ( .A1(_04030_ ), .A2(\ID_EX_pc [20] ), .A3(_06115_ ), .ZN(_00193_ ) );
AND3_X1 _13878_ ( .A1(_04030_ ), .A2(\ID_EX_pc [19] ), .A3(_06115_ ), .ZN(_00194_ ) );
CLKBUF_X2 _13879_ ( .A(_04029_ ), .Z(_06116_ ) );
AND3_X1 _13880_ ( .A1(_06116_ ), .A2(\ID_EX_pc [18] ), .A3(_06115_ ), .ZN(_00195_ ) );
AND3_X1 _13881_ ( .A1(_06116_ ), .A2(\ID_EX_pc [17] ), .A3(_06115_ ), .ZN(_00196_ ) );
AND3_X1 _13882_ ( .A1(_06116_ ), .A2(\ID_EX_pc [16] ), .A3(_06115_ ), .ZN(_00197_ ) );
AND3_X1 _13883_ ( .A1(_06116_ ), .A2(\ID_EX_pc [15] ), .A3(_06115_ ), .ZN(_00198_ ) );
AND3_X1 _13884_ ( .A1(_06116_ ), .A2(\ID_EX_pc [14] ), .A3(_06115_ ), .ZN(_00199_ ) );
AND3_X1 _13885_ ( .A1(_06116_ ), .A2(\ID_EX_pc [13] ), .A3(_06115_ ), .ZN(_00200_ ) );
AND3_X1 _13886_ ( .A1(_06116_ ), .A2(\ID_EX_pc [12] ), .A3(_06115_ ), .ZN(_00201_ ) );
CLKBUF_X2 _13887_ ( .A(_03221_ ), .Z(_06117_ ) );
AND3_X1 _13888_ ( .A1(_06116_ ), .A2(\ID_EX_pc [29] ), .A3(_06117_ ), .ZN(_00202_ ) );
AND3_X1 _13889_ ( .A1(_06116_ ), .A2(\ID_EX_pc [11] ), .A3(_06117_ ), .ZN(_00203_ ) );
AND3_X1 _13890_ ( .A1(_06116_ ), .A2(\ID_EX_pc [10] ), .A3(_06117_ ), .ZN(_00204_ ) );
CLKBUF_X2 _13891_ ( .A(_04024_ ), .Z(_06118_ ) );
AND3_X1 _13892_ ( .A1(_06118_ ), .A2(\ID_EX_pc [9] ), .A3(_06117_ ), .ZN(_00205_ ) );
AND3_X1 _13893_ ( .A1(_06118_ ), .A2(\ID_EX_pc [8] ), .A3(_06117_ ), .ZN(_00206_ ) );
AND3_X1 _13894_ ( .A1(_06118_ ), .A2(\ID_EX_pc [7] ), .A3(_06117_ ), .ZN(_00207_ ) );
AND3_X1 _13895_ ( .A1(_06118_ ), .A2(\ID_EX_pc [6] ), .A3(_06117_ ), .ZN(_00208_ ) );
AND3_X1 _13896_ ( .A1(_06118_ ), .A2(\ID_EX_pc [5] ), .A3(_06117_ ), .ZN(_00209_ ) );
AND3_X1 _13897_ ( .A1(_06118_ ), .A2(\ID_EX_pc [4] ), .A3(_06117_ ), .ZN(_00210_ ) );
AND3_X1 _13898_ ( .A1(_06118_ ), .A2(\ID_EX_pc [3] ), .A3(_06117_ ), .ZN(_00211_ ) );
CLKBUF_X2 _13899_ ( .A(_03221_ ), .Z(_06119_ ) );
AND3_X1 _13900_ ( .A1(_06118_ ), .A2(\ID_EX_pc [2] ), .A3(_06119_ ), .ZN(_00212_ ) );
AND3_X1 _13901_ ( .A1(_06118_ ), .A2(\ID_EX_pc [28] ), .A3(_06119_ ), .ZN(_00213_ ) );
AND3_X1 _13902_ ( .A1(_06118_ ), .A2(\ID_EX_pc [1] ), .A3(_06119_ ), .ZN(_00214_ ) );
CLKBUF_X2 _13903_ ( .A(_04024_ ), .Z(_06120_ ) );
AND3_X1 _13904_ ( .A1(_06120_ ), .A2(\ID_EX_pc [0] ), .A3(_06119_ ), .ZN(_00215_ ) );
AND3_X1 _13905_ ( .A1(_06120_ ), .A2(\ID_EX_pc [27] ), .A3(_06119_ ), .ZN(_00216_ ) );
AND3_X1 _13906_ ( .A1(_06120_ ), .A2(\ID_EX_pc [26] ), .A3(_06119_ ), .ZN(_00217_ ) );
AND3_X1 _13907_ ( .A1(_06120_ ), .A2(\ID_EX_pc [25] ), .A3(_06119_ ), .ZN(_00218_ ) );
AND3_X1 _13908_ ( .A1(_06120_ ), .A2(\ID_EX_pc [24] ), .A3(_06119_ ), .ZN(_00219_ ) );
AND3_X1 _13909_ ( .A1(_06120_ ), .A2(\ID_EX_pc [23] ), .A3(_06119_ ), .ZN(_00220_ ) );
AND3_X1 _13910_ ( .A1(_06120_ ), .A2(\ID_EX_pc [22] ), .A3(_06119_ ), .ZN(_00221_ ) );
CLKBUF_X2 _13911_ ( .A(_03221_ ), .Z(_06121_ ) );
AND3_X1 _13912_ ( .A1(_06120_ ), .A2(\ID_EX_typ [7] ), .A3(_06121_ ), .ZN(_00222_ ) );
INV_X1 _13913_ ( .A(io_master_awready ), .ZN(_06122_ ) );
NAND3_X1 _13914_ ( .A1(_03988_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A3(_06122_ ), .ZN(_06123_ ) );
OAI21_X1 _13915_ ( .A(_06123_ ), .B1(\mylsu.state [4] ), .B2(\mylsu.state [0] ), .ZN(_06124_ ) );
AND3_X1 _13916_ ( .A1(_02170_ ), .A2(\myclint.rvalid ), .A3(_02173_ ), .ZN(_06125_ ) );
INV_X1 _13917_ ( .A(_06125_ ), .ZN(_06126_ ) );
OAI21_X1 _13918_ ( .A(_06126_ ), .B1(_02174_ ), .B2(io_master_arready ), .ZN(_06127_ ) );
INV_X1 _13919_ ( .A(_02076_ ), .ZN(_06128_ ) );
BUF_X4 _13920_ ( .A(_06128_ ), .Z(_06129_ ) );
BUF_X4 _13921_ ( .A(_06129_ ), .Z(_06130_ ) );
BUF_X2 _13922_ ( .A(_06130_ ), .Z(_06131_ ) );
OR2_X1 _13923_ ( .A1(_06127_ ), .A2(_06131_ ), .ZN(_06132_ ) );
AOI21_X1 _13924_ ( .A(_06124_ ), .B1(_06132_ ), .B2(_02134_ ), .ZN(_06133_ ) );
INV_X1 _13925_ ( .A(EXU_valid_LSU ), .ZN(_06134_ ) );
OR2_X1 _13926_ ( .A1(_06133_ ), .A2(_06134_ ), .ZN(_06135_ ) );
AOI21_X1 _13927_ ( .A(_04031_ ), .B1(_06135_ ), .B2(_04027_ ), .ZN(_00223_ ) );
AND3_X1 _13928_ ( .A1(_06120_ ), .A2(\ID_EX_typ [6] ), .A3(_06121_ ), .ZN(_00224_ ) );
AND3_X1 _13929_ ( .A1(_06120_ ), .A2(\ID_EX_typ [5] ), .A3(_06121_ ), .ZN(_00225_ ) );
AND3_X1 _13930_ ( .A1(_04029_ ), .A2(fanout_net_8 ), .A3(_06121_ ), .ZN(_00226_ ) );
AND3_X1 _13931_ ( .A1(_04029_ ), .A2(\ID_EX_typ [3] ), .A3(_06121_ ), .ZN(_00227_ ) );
AND3_X1 _13932_ ( .A1(_04029_ ), .A2(\ID_EX_typ [2] ), .A3(_06121_ ), .ZN(_00228_ ) );
AND3_X1 _13933_ ( .A1(_04029_ ), .A2(\ID_EX_typ [1] ), .A3(_06121_ ), .ZN(_00229_ ) );
AND3_X1 _13934_ ( .A1(_04029_ ), .A2(fanout_net_7 ), .A3(_06121_ ), .ZN(_00230_ ) );
AND2_X1 _13935_ ( .A1(_02162_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_06136_ ) );
CLKBUF_X2 _13936_ ( .A(_06136_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _13937_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .ZN(_06137_ ) );
BUF_X2 _13938_ ( .A(_06137_ ), .Z(_06138_ ) );
AND3_X1 _13939_ ( .A1(_02162_ ), .A2(_06138_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00278_ ) );
BUF_X4 _13940_ ( .A(_03426_ ), .Z(_06139_ ) );
CLKBUF_X2 _13941_ ( .A(_06139_ ), .Z(_06140_ ) );
BUF_X2 _13942_ ( .A(_06140_ ), .Z(_06141_ ) );
AND3_X1 _13943_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06141_ ), .A3(fanout_net_9 ), .ZN(_00279_ ) );
INV_X1 _13944_ ( .A(fanout_net_9 ), .ZN(_06142_ ) );
BUF_X8 _13945_ ( .A(_06142_ ), .Z(_06143_ ) );
BUF_X2 _13946_ ( .A(_06143_ ), .Z(_06144_ ) );
AND3_X1 _13947_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_13 ), .A3(_06144_ ), .ZN(_00280_ ) );
AND3_X1 _13948_ ( .A1(_04029_ ), .A2(\EX_LS_pc [2] ), .A3(_06121_ ), .ZN(_00318_ ) );
AND3_X1 _13949_ ( .A1(_04024_ ), .A2(fanout_net_45 ), .A3(_03221_ ), .ZN(_00319_ ) );
NOR2_X1 _13950_ ( .A1(_04031_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_06145_ ) );
NOR2_X1 _13951_ ( .A1(fanout_net_45 ), .A2(\mylsu.state [1] ), .ZN(_06146_ ) );
NAND2_X1 _13952_ ( .A1(_06145_ ), .A2(_06146_ ), .ZN(_06147_ ) );
BUF_X2 _13953_ ( .A(_02150_ ), .Z(_06148_ ) );
AOI21_X1 _13954_ ( .A(_02218_ ), .B1(_06148_ ), .B2(_02220_ ), .ZN(_06149_ ) );
OAI21_X1 _13955_ ( .A(_02148_ ), .B1(_02224_ ), .B2(_02225_ ), .ZN(_06150_ ) );
OR2_X1 _13956_ ( .A1(_06150_ ), .A2(_02228_ ), .ZN(_06151_ ) );
AOI21_X1 _13957_ ( .A(_03982_ ), .B1(_06151_ ), .B2(\EX_LS_flag [2] ), .ZN(_06152_ ) );
AOI21_X1 _13958_ ( .A(_06147_ ), .B1(_06149_ ), .B2(_06152_ ), .ZN(_00332_ ) );
NOR2_X1 _13959_ ( .A1(_03988_ ), .A2(_03978_ ), .ZN(_06153_ ) );
AOI21_X1 _13960_ ( .A(_02218_ ), .B1(_06151_ ), .B2(_06153_ ), .ZN(_06154_ ) );
AOI21_X1 _13961_ ( .A(_06147_ ), .B1(_06154_ ), .B2(_03986_ ), .ZN(_00333_ ) );
NOR2_X1 _13962_ ( .A1(_02226_ ), .A2(_02228_ ), .ZN(_06155_ ) );
NAND3_X1 _13963_ ( .A1(_06155_ ), .A2(\EX_LS_flag [2] ), .A3(_02130_ ), .ZN(_06156_ ) );
NOR2_X1 _13964_ ( .A1(_06156_ ), .A2(_06147_ ), .ZN(_00334_ ) );
AOI21_X1 _13965_ ( .A(_06147_ ), .B1(_03975_ ), .B2(_02147_ ), .ZN(_00335_ ) );
AOI21_X1 _13966_ ( .A(_06147_ ), .B1(_03986_ ), .B2(_06156_ ), .ZN(_00336_ ) );
NAND3_X1 _13967_ ( .A1(_04026_ ), .A2(EXU_valid_LSU ), .A3(_06146_ ), .ZN(_06157_ ) );
OR3_X1 _13968_ ( .A1(_02158_ ), .A2(_03982_ ), .A3(_06157_ ), .ZN(_06158_ ) );
INV_X1 _13969_ ( .A(_02133_ ), .ZN(_06159_ ) );
OR3_X1 _13970_ ( .A1(_06159_ ), .A2(_02158_ ), .A3(_02146_ ), .ZN(_06160_ ) );
AND3_X1 _13971_ ( .A1(_06150_ ), .A2(_02227_ ), .A3(_06153_ ), .ZN(_06161_ ) );
NOR2_X1 _13972_ ( .A1(_02152_ ), .A2(_06161_ ), .ZN(_06162_ ) );
AOI21_X1 _13973_ ( .A(_06158_ ), .B1(_06160_ ), .B2(_06162_ ), .ZN(_00337_ ) );
INV_X1 _13974_ ( .A(_00319_ ), .ZN(_06163_ ) );
OAI211_X1 _13975_ ( .A(EXU_valid_LSU ), .B(_06146_ ), .C1(_02129_ ), .C2(_02151_ ), .ZN(_06164_ ) );
BUF_X4 _13976_ ( .A(_03976_ ), .Z(_06165_ ) );
OAI21_X1 _13977_ ( .A(_04026_ ), .B1(_06165_ ), .B2(_02230_ ), .ZN(_06166_ ) );
OAI21_X1 _13978_ ( .A(_06163_ ), .B1(_06164_ ), .B2(_06166_ ), .ZN(_00338_ ) );
CLKBUF_X2 _13979_ ( .A(_02176_ ), .Z(\io_master_arburst [0] ) );
BUF_X2 _13980_ ( .A(_02077_ ), .Z(_06167_ ) );
NOR3_X1 _13981_ ( .A1(_06167_ ), .A2(fanout_net_6 ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06168_ ) );
BUF_X4 _13982_ ( .A(_06130_ ), .Z(_06169_ ) );
INV_X1 _13983_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_06170_ ) );
INV_X1 _13984_ ( .A(_02079_ ), .ZN(_06171_ ) );
BUF_X4 _13985_ ( .A(_06171_ ), .Z(_06172_ ) );
AOI211_X1 _13986_ ( .A(_06168_ ), .B(_06169_ ), .C1(_06170_ ), .C2(_06172_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _13987_ ( .A1(_06167_ ), .A2(fanout_net_5 ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06173_ ) );
INV_X1 _13988_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_06174_ ) );
AOI211_X1 _13989_ ( .A(_06173_ ), .B(_06169_ ), .C1(_06174_ ), .C2(_06172_ ), .ZN(\io_master_araddr [0] ) );
BUF_X4 _13990_ ( .A(_06169_ ), .Z(_06175_ ) );
AND2_X1 _13991_ ( .A1(_02177_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .ZN(_06176_ ) );
AOI21_X1 _13992_ ( .A(_06176_ ), .B1(\mylsu.araddr_tmp [15] ), .B2(_06172_ ), .ZN(_06177_ ) );
BUF_X4 _13993_ ( .A(_02087_ ), .Z(_06178_ ) );
BUF_X4 _13994_ ( .A(_06178_ ), .Z(_06179_ ) );
OAI22_X1 _13995_ ( .A1(_06175_ ), .A2(_06177_ ), .B1(_03660_ ), .B2(_06179_ ), .ZN(\io_master_araddr [15] ) );
OR3_X1 _13996_ ( .A1(_06167_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06180_ ) );
OAI21_X1 _13997_ ( .A(_06180_ ), .B1(\mylsu.araddr_tmp [14] ), .B2(_02177_ ), .ZN(_06181_ ) );
OAI22_X1 _13998_ ( .A1(_06175_ ), .A2(_06181_ ), .B1(_03670_ ), .B2(_06179_ ), .ZN(\io_master_araddr [14] ) );
OR3_X1 _13999_ ( .A1(_06167_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06182_ ) );
OAI21_X1 _14000_ ( .A(_06182_ ), .B1(\mylsu.araddr_tmp [5] ), .B2(_02177_ ), .ZN(_06183_ ) );
OAI22_X1 _14001_ ( .A1(_06175_ ), .A2(_06183_ ), .B1(_03610_ ), .B2(_06179_ ), .ZN(\io_master_araddr [5] ) );
NOR3_X1 _14002_ ( .A1(_06167_ ), .A2(_04038_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06184_ ) );
AOI21_X1 _14003_ ( .A(_06184_ ), .B1(_06172_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_06185_ ) );
OAI22_X1 _14004_ ( .A1(_06175_ ), .A2(_06185_ ), .B1(_06141_ ), .B2(_06179_ ), .ZN(\io_master_araddr [4] ) );
NOR3_X1 _14005_ ( .A1(_06167_ ), .A2(_04052_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06186_ ) );
AOI21_X1 _14006_ ( .A(_06186_ ), .B1(_06172_ ), .B2(\mylsu.araddr_tmp [3] ), .ZN(_06187_ ) );
OAI22_X1 _14007_ ( .A1(_06175_ ), .A2(_06187_ ), .B1(_06144_ ), .B2(_06179_ ), .ZN(\io_master_araddr [3] ) );
AND2_X1 _14008_ ( .A1(_02177_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .ZN(_06188_ ) );
AOI21_X1 _14009_ ( .A(_06188_ ), .B1(\mylsu.araddr_tmp [13] ), .B2(_06172_ ), .ZN(_06189_ ) );
OAI22_X1 _14010_ ( .A1(_06175_ ), .A2(_06189_ ), .B1(_01886_ ), .B2(_06179_ ), .ZN(\io_master_araddr [13] ) );
AND2_X1 _14011_ ( .A1(_02177_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .ZN(_06190_ ) );
AOI21_X1 _14012_ ( .A(_06190_ ), .B1(\mylsu.araddr_tmp [12] ), .B2(_06172_ ), .ZN(_06191_ ) );
BUF_X4 _14013_ ( .A(_02087_ ), .Z(_06192_ ) );
OAI22_X1 _14014_ ( .A1(_06175_ ), .A2(_06191_ ), .B1(_02004_ ), .B2(_06192_ ), .ZN(\io_master_araddr [12] ) );
AND2_X1 _14015_ ( .A1(_02177_ ), .A2(\EX_LS_dest_csreg_mem [11] ), .ZN(_06193_ ) );
AOI21_X1 _14016_ ( .A(_06193_ ), .B1(\mylsu.araddr_tmp [11] ), .B2(_06172_ ), .ZN(_06194_ ) );
OAI22_X1 _14017_ ( .A1(_06175_ ), .A2(_06194_ ), .B1(_03708_ ), .B2(_06192_ ), .ZN(\io_master_araddr [11] ) );
OR3_X1 _14018_ ( .A1(_06167_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06195_ ) );
OAI21_X1 _14019_ ( .A(_06195_ ), .B1(\mylsu.araddr_tmp [10] ), .B2(_02177_ ), .ZN(_06196_ ) );
OAI22_X1 _14020_ ( .A1(_06175_ ), .A2(_06196_ ), .B1(_03701_ ), .B2(_06192_ ), .ZN(\io_master_araddr [10] ) );
NOR3_X1 _14021_ ( .A1(_06167_ ), .A2(_04055_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06197_ ) );
AOI21_X1 _14022_ ( .A(_06197_ ), .B1(_06172_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_06198_ ) );
OAI22_X1 _14023_ ( .A1(_06175_ ), .A2(_06198_ ), .B1(_03693_ ), .B2(_06192_ ), .ZN(\io_master_araddr [9] ) );
AND2_X1 _14024_ ( .A1(_02177_ ), .A2(\EX_LS_dest_csreg_mem [8] ), .ZN(_06199_ ) );
AOI21_X1 _14025_ ( .A(_06199_ ), .B1(\mylsu.araddr_tmp [8] ), .B2(_06171_ ), .ZN(_06200_ ) );
OAI22_X1 _14026_ ( .A1(_06169_ ), .A2(_06200_ ), .B1(_03654_ ), .B2(_06192_ ), .ZN(\io_master_araddr [8] ) );
NOR3_X1 _14027_ ( .A1(_06167_ ), .A2(_04056_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06201_ ) );
AOI21_X1 _14028_ ( .A(_06201_ ), .B1(_06172_ ), .B2(\mylsu.araddr_tmp [7] ), .ZN(_06202_ ) );
OAI22_X1 _14029_ ( .A1(_06169_ ), .A2(_06202_ ), .B1(_02021_ ), .B2(_06192_ ), .ZN(\io_master_araddr [7] ) );
AND2_X1 _14030_ ( .A1(_02177_ ), .A2(\EX_LS_dest_csreg_mem [6] ), .ZN(_06203_ ) );
AOI21_X1 _14031_ ( .A(_06203_ ), .B1(\mylsu.araddr_tmp [6] ), .B2(_06171_ ), .ZN(_06204_ ) );
OAI22_X1 _14032_ ( .A1(_06169_ ), .A2(_06204_ ), .B1(_01875_ ), .B2(_06192_ ), .ZN(\io_master_araddr [6] ) );
INV_X1 _14033_ ( .A(_02060_ ), .ZN(_06205_ ) );
OR3_X1 _14034_ ( .A1(_06167_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .ZN(_06206_ ) );
OAI211_X1 _14035_ ( .A(_06205_ ), .B(_06206_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_02079_ ), .ZN(_06207_ ) );
NOR2_X1 _14036_ ( .A1(_02055_ ), .A2(_06207_ ), .ZN(_06208_ ) );
BUF_X4 _14037_ ( .A(_06208_ ), .Z(_06209_ ) );
BUF_X4 _14038_ ( .A(_06209_ ), .Z(_06210_ ) );
BUF_X2 _14039_ ( .A(_06210_ ), .Z(\io_master_araddr [2] ) );
BUF_X2 _14040_ ( .A(_02076_ ), .Z(_06211_ ) );
CLKBUF_X2 _14041_ ( .A(_06211_ ), .Z(\io_master_arid [1] ) );
NOR3_X1 _14042_ ( .A1(\io_master_arburst [0] ), .A2(_02138_ ), .A3(_02060_ ), .ZN(\io_master_arsize [2] ) );
NOR3_X1 _14043_ ( .A1(\io_master_arburst [0] ), .A2(_02137_ ), .A3(_02060_ ), .ZN(\io_master_arsize [0] ) );
INV_X1 _14044_ ( .A(\EX_LS_typ [2] ), .ZN(_06212_ ) );
OAI22_X1 _14045_ ( .A1(_02053_ ), .A2(_02054_ ), .B1(_06212_ ), .B2(_02060_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _14046_ ( .A(_02178_ ), .B(_02179_ ), .C1(_02170_ ), .C2(_02173_ ), .ZN(io_master_arvalid ) );
AND2_X1 _14047_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ) );
AND2_X1 _14048_ ( .A1(_06148_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .ZN(_06213_ ) );
BUF_X4 _14049_ ( .A(_06213_ ), .Z(_06214_ ) );
BUF_X4 _14050_ ( .A(_06214_ ), .Z(_06215_ ) );
MUX2_X1 _14051_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_06215_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _14052_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_06215_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _14053_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_06215_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _14054_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_06215_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _14055_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_06215_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _14056_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_06215_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _14057_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_06215_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _14058_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_06215_ ), .Z(\io_master_awaddr [16] ) );
MUX2_X1 _14059_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_06215_ ), .Z(\io_master_awaddr [15] ) );
BUF_X4 _14060_ ( .A(_06214_ ), .Z(_06216_ ) );
MUX2_X1 _14061_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_06216_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _14062_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_06216_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _14063_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_06216_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _14064_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_06216_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _14065_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_06216_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _14066_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_06216_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _14067_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_06216_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _14068_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_06216_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _14069_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_06216_ ), .Z(\io_master_awaddr [7] ) );
MUX2_X1 _14070_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_06216_ ), .Z(\io_master_awaddr [6] ) );
BUF_X4 _14071_ ( .A(_06214_ ), .Z(_06217_ ) );
MUX2_X1 _14072_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_06217_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _14073_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_06217_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _14074_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_06217_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _14075_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_06217_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _14076_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_06217_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _14077_ ( .A(\mylsu.awaddr_tmp [1] ), .B(fanout_net_6 ), .S(_06217_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _14078_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_5 ), .S(_06217_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _14079_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_06217_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _14080_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_06217_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _14081_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_06217_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _14082_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_06214_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _14083_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_06214_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _14084_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_06214_ ), .Z(\io_master_awaddr [22] ) );
AND3_X1 _14085_ ( .A1(_02157_ ), .A2(\EX_LS_typ [1] ), .A3(_02141_ ), .ZN(\io_master_awsize [0] ) );
NAND2_X1 _14086_ ( .A1(_02157_ ), .A2(_02141_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _14087_ ( .A1(_02147_ ), .A2(_02159_ ), .A3(_06215_ ), .ZN(_06218_ ) );
INV_X1 _14088_ ( .A(\mylsu.state [4] ), .ZN(_06219_ ) );
NAND2_X1 _14089_ ( .A1(_06218_ ), .A2(_06219_ ), .ZN(io_master_awvalid ) );
INV_X1 _14090_ ( .A(\mylsu.state [2] ), .ZN(_06220_ ) );
INV_X1 _14091_ ( .A(\mylsu.state [1] ), .ZN(_06221_ ) );
NAND4_X1 _14092_ ( .A1(_06218_ ), .A2(_06220_ ), .A3(_06219_ ), .A4(_06221_ ), .ZN(io_master_bready ) );
NOR3_X1 _14093_ ( .A1(_02059_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_06222_ ) );
NOR2_X1 _14094_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_06223_ ) );
AND2_X1 _14095_ ( .A1(_06223_ ), .A2(io_master_bvalid ), .ZN(_06224_ ) );
NAND2_X1 _14096_ ( .A1(\io_master_bid [1] ), .A2(\io_master_bid [0] ), .ZN(_06225_ ) );
NOR3_X1 _14097_ ( .A1(_06225_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bid [2] ), .ZN(_06226_ ) );
AND2_X1 _14098_ ( .A1(_06224_ ), .A2(_06226_ ), .ZN(_06227_ ) );
INV_X1 _14099_ ( .A(_06227_ ), .ZN(_06228_ ) );
NAND4_X1 _14100_ ( .A1(_02173_ ), .A2(_06211_ ), .A3(_02168_ ), .A4(_02169_ ), .ZN(_06229_ ) );
NOR2_X1 _14101_ ( .A1(_03963_ ), .A2(\io_master_rid [0] ), .ZN(_06230_ ) );
NAND4_X1 _14102_ ( .A1(_06230_ ), .A2(_03961_ ), .A3(_03962_ ), .A4(io_master_rlast ), .ZN(_06231_ ) );
OAI21_X1 _14103_ ( .A(_06229_ ), .B1(_06130_ ), .B2(_06231_ ), .ZN(_06232_ ) );
AND2_X1 _14104_ ( .A1(_03960_ ), .A2(_06232_ ), .ZN(_06233_ ) );
INV_X1 _14105_ ( .A(_06233_ ), .ZN(_06234_ ) );
AOI221_X4 _14106_ ( .A(_06222_ ), .B1(\mylsu.state [1] ), .B2(_06228_ ), .C1(_06234_ ), .C2(fanout_net_45 ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _14107_ ( .A(_02161_ ), .B(_02164_ ), .C1(_02170_ ), .C2(_02173_ ), .ZN(io_master_rready ) );
MUX2_X1 _14108_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_5 ), .Z(_06235_ ) );
CLKBUF_X2 _14109_ ( .A(_04036_ ), .Z(_06236_ ) );
AND2_X1 _14110_ ( .A1(_06235_ ), .A2(_06236_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _14111_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_5 ), .Z(_06237_ ) );
AND2_X1 _14112_ ( .A1(_06237_ ), .A2(_06236_ ), .ZN(\io_master_wdata [14] ) );
NOR3_X1 _14113_ ( .A1(_05858_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [5] ) );
NOR3_X1 _14114_ ( .A1(_05885_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [4] ) );
NOR3_X1 _14115_ ( .A1(_05898_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [3] ) );
INV_X1 _14116_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_06238_ ) );
NOR3_X1 _14117_ ( .A1(_06238_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [2] ) );
INV_X1 _14118_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_06239_ ) );
NOR3_X1 _14119_ ( .A1(_06239_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [1] ) );
INV_X1 _14120_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_06240_ ) );
NOR3_X1 _14121_ ( .A1(_06240_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _14122_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_5 ), .Z(_06241_ ) );
AND2_X1 _14123_ ( .A1(_06241_ ), .A2(_06236_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _14124_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_5 ), .Z(_06242_ ) );
AND2_X1 _14125_ ( .A1(_06242_ ), .A2(_06236_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _14126_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_5 ), .Z(_06243_ ) );
AND2_X1 _14127_ ( .A1(_06243_ ), .A2(_06236_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _14128_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_5 ), .Z(_06244_ ) );
AND2_X1 _14129_ ( .A1(_06244_ ), .A2(_06236_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _14130_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_5 ), .Z(_06245_ ) );
AND2_X1 _14131_ ( .A1(_06245_ ), .A2(_06236_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _14132_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_5 ), .Z(_06246_ ) );
AND2_X1 _14133_ ( .A1(_06246_ ), .A2(_06236_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _14134_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_06247_ ) );
NOR3_X1 _14135_ ( .A1(_06247_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [7] ) );
NOR3_X1 _14136_ ( .A1(_05840_ ), .A2(fanout_net_5 ), .A3(fanout_net_6 ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _14137_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_5 ), .Z(_06248_ ) );
MUX2_X1 _14138_ ( .A(_06248_ ), .B(_06235_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _14139_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_5 ), .Z(_06249_ ) );
MUX2_X1 _14140_ ( .A(_06249_ ), .B(_06237_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [30] ) );
MUX2_X1 _14141_ ( .A(_06072_ ), .B(_05678_ ), .S(fanout_net_5 ), .Z(_06250_ ) );
NOR2_X1 _14142_ ( .A1(_04036_ ), .A2(fanout_net_5 ), .ZN(_06251_ ) );
INV_X1 _14143_ ( .A(_06251_ ), .ZN(_06252_ ) );
OAI22_X1 _14144_ ( .A1(_06250_ ), .A2(fanout_net_6 ), .B1(_06252_ ), .B2(_05858_ ), .ZN(\io_master_wdata [21] ) );
MUX2_X1 _14145_ ( .A(_05491_ ), .B(_05705_ ), .S(fanout_net_5 ), .Z(_06253_ ) );
OAI22_X1 _14146_ ( .A1(_06253_ ), .A2(fanout_net_6 ), .B1(_06252_ ), .B2(_05885_ ), .ZN(\io_master_wdata [20] ) );
INV_X1 _14147_ ( .A(\EX_LS_result_csreg_mem [19] ), .ZN(_06254_ ) );
MUX2_X1 _14148_ ( .A(_06254_ ), .B(_05729_ ), .S(fanout_net_5 ), .Z(_06255_ ) );
OAI22_X1 _14149_ ( .A1(_06255_ ), .A2(fanout_net_6 ), .B1(_06252_ ), .B2(_05898_ ), .ZN(\io_master_wdata [19] ) );
OAI21_X1 _14150_ ( .A(_04036_ ), .B1(_04043_ ), .B2(\EX_LS_result_csreg_mem [10] ), .ZN(_06256_ ) );
NOR2_X1 _14151_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [18] ), .ZN(_06257_ ) );
OAI22_X1 _14152_ ( .A1(_06252_ ), .A2(_06238_ ), .B1(_06256_ ), .B2(_06257_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _14153_ ( .A(_04036_ ), .B1(_04043_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_06258_ ) );
NOR2_X1 _14154_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_06259_ ) );
OAI22_X1 _14155_ ( .A1(_06252_ ), .A2(_06239_ ), .B1(_06258_ ), .B2(_06259_ ), .ZN(\io_master_wdata [17] ) );
MUX2_X1 _14156_ ( .A(_05613_ ), .B(_05804_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06260_ ) );
OAI22_X1 _14157_ ( .A1(_06260_ ), .A2(fanout_net_6 ), .B1(_06252_ ), .B2(_06240_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _14158_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06261_ ) );
MUX2_X1 _14159_ ( .A(_06261_ ), .B(_06241_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _14160_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06262_ ) );
MUX2_X1 _14161_ ( .A(_06262_ ), .B(_06242_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _14162_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06263_ ) );
MUX2_X1 _14163_ ( .A(_06263_ ), .B(_06243_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _14164_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06264_ ) );
MUX2_X1 _14165_ ( .A(_06264_ ), .B(_06244_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _14166_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06265_ ) );
MUX2_X1 _14167_ ( .A(_06265_ ), .B(_06245_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _14168_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06266_ ) );
MUX2_X1 _14169_ ( .A(_06266_ ), .B(_06246_ ), .S(fanout_net_6 ), .Z(\io_master_wdata [24] ) );
INV_X1 _14170_ ( .A(\EX_LS_result_csreg_mem [23] ), .ZN(_06267_ ) );
INV_X1 _14171_ ( .A(\EX_LS_result_csreg_mem [15] ), .ZN(_06268_ ) );
MUX2_X1 _14172_ ( .A(_06267_ ), .B(_06268_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06269_ ) );
OAI22_X1 _14173_ ( .A1(_06269_ ), .A2(fanout_net_6 ), .B1(_06252_ ), .B2(_06247_ ), .ZN(\io_master_wdata [23] ) );
MUX2_X1 _14174_ ( .A(_06057_ ), .B(_05659_ ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06270_ ) );
OAI22_X1 _14175_ ( .A1(_06270_ ), .A2(fanout_net_6 ), .B1(_06252_ ), .B2(_05840_ ), .ZN(\io_master_wdata [22] ) );
MUX2_X1 _14176_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06271_ ) );
AND2_X1 _14177_ ( .A1(_06271_ ), .A2(_06236_ ), .ZN(\io_master_wstrb [1] ) );
AND3_X1 _14178_ ( .A1(_04043_ ), .A2(_06236_ ), .A3(\EX_LS_typ [0] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _14179_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_06272_ ) );
MUX2_X1 _14180_ ( .A(_06272_ ), .B(_06271_ ), .S(fanout_net_6 ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _14181_ ( .A1(_04036_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_06273_ ) );
NAND3_X1 _14182_ ( .A1(_04043_ ), .A2(fanout_net_6 ), .A3(\EX_LS_typ [0] ), .ZN(_06274_ ) );
OAI211_X1 _14183_ ( .A(_06273_ ), .B(_06274_ ), .C1(_02136_ ), .C2(_06212_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _14184_ ( .A1(_06218_ ), .A2(_06220_ ), .ZN(io_master_wvalid ) );
AND2_X1 _14185_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_06275_ ) );
NOR2_X1 _14186_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_06276_ ) );
AND2_X1 _14187_ ( .A1(_06275_ ), .A2(_06276_ ), .ZN(_06277_ ) );
NOR4_X1 _14188_ ( .A1(\LS_WB_waddr_csreg [7] ), .A2(\LS_WB_waddr_csreg [6] ), .A3(\LS_WB_waddr_csreg [5] ), .A4(\LS_WB_waddr_csreg [4] ), .ZN(_06278_ ) );
NAND2_X1 _14189_ ( .A1(_06277_ ), .A2(_06278_ ), .ZN(_06279_ ) );
INV_X1 _14190_ ( .A(\LS_WB_wen_csreg [7] ), .ZN(_06280_ ) );
NOR2_X1 _14191_ ( .A1(_06280_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_06281_ ) );
INV_X1 _14192_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_06282_ ) );
INV_X1 _14193_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_06283_ ) );
INV_X1 _14194_ ( .A(\LS_WB_waddr_csreg [2] ), .ZN(_06284_ ) );
NAND4_X1 _14195_ ( .A1(_06281_ ), .A2(_06282_ ), .A3(_06283_ ), .A4(_06284_ ), .ZN(_06285_ ) );
NOR2_X1 _14196_ ( .A1(_06279_ ), .A2(_06285_ ), .ZN(\mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ) );
NAND4_X1 _14197_ ( .A1(_06281_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(_06283_ ), .A4(\LS_WB_waddr_csreg [2] ), .ZN(_06286_ ) );
NOR2_X1 _14198_ ( .A1(_06279_ ), .A2(_06286_ ), .ZN(\mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _14199_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_06287_ ) );
NAND2_X1 _14200_ ( .A1(_06287_ ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_06288_ ) );
NOR2_X1 _14201_ ( .A1(_06288_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_06289_ ) );
AND4_X1 _14202_ ( .A1(\LS_WB_waddr_csreg [0] ), .A2(_06289_ ), .A3(_06283_ ), .A4(_06281_ ), .ZN(_06290_ ) );
AND3_X1 _14203_ ( .A1(_06290_ ), .A2(_06284_ ), .A3(_06277_ ), .ZN(\mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14204_ ( .A(_06289_ ), .ZN(_06291_ ) );
NOR4_X1 _14205_ ( .A1(_06291_ ), .A2(\LS_WB_waddr_csreg [0] ), .A3(_06283_ ), .A4(\LS_WB_waddr_csreg [3] ), .ZN(_06292_ ) );
NAND3_X1 _14206_ ( .A1(_06292_ ), .A2(_06284_ ), .A3(_06277_ ), .ZN(_06293_ ) );
AOI21_X1 _14207_ ( .A(_06280_ ), .B1(_06293_ ), .B2(_02213_ ), .ZN(\mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ) );
INV_X1 _14208_ ( .A(_02160_ ), .ZN(_06294_ ) );
NOR2_X1 _14209_ ( .A1(_06155_ ), .A2(exception_quest_IDU ), .ZN(_06295_ ) );
OR2_X2 _14210_ ( .A1(_06294_ ), .A2(_06295_ ), .ZN(_06296_ ) );
BUF_X4 _14211_ ( .A(_06296_ ), .Z(_06297_ ) );
MUX2_X1 _14212_ ( .A(\ID_EX_pc [21] ), .B(\EX_LS_pc [21] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _14213_ ( .A(\ID_EX_pc [20] ), .B(\EX_LS_pc [20] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _14214_ ( .A(\ID_EX_pc [19] ), .B(\EX_LS_pc [19] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _14215_ ( .A(\ID_EX_pc [18] ), .B(\EX_LS_pc [18] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _14216_ ( .A(\ID_EX_pc [17] ), .B(\EX_LS_pc [17] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _14217_ ( .A(\ID_EX_pc [16] ), .B(\EX_LS_pc [16] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _14218_ ( .A(\ID_EX_pc [15] ), .B(\EX_LS_pc [15] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _14219_ ( .A(\ID_EX_pc [14] ), .B(\EX_LS_pc [14] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _14220_ ( .A(\ID_EX_pc [13] ), .B(\EX_LS_pc [13] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _14221_ ( .A(\ID_EX_pc [12] ), .B(\EX_LS_pc [12] ), .S(_06297_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _14222_ ( .A(_06296_ ), .Z(_06298_ ) );
MUX2_X1 _14223_ ( .A(\ID_EX_pc [30] ), .B(\EX_LS_pc [30] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _14224_ ( .A(\ID_EX_pc [11] ), .B(\EX_LS_pc [11] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _14225_ ( .A(\ID_EX_pc [10] ), .B(\EX_LS_pc [10] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _14226_ ( .A(\ID_EX_pc [9] ), .B(\EX_LS_pc [9] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _14227_ ( .A(\ID_EX_pc [8] ), .B(\EX_LS_pc [8] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _14228_ ( .A(\ID_EX_pc [7] ), .B(\EX_LS_pc [7] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _14229_ ( .A(\ID_EX_pc [6] ), .B(\EX_LS_pc [6] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _14230_ ( .A(\ID_EX_pc [5] ), .B(\EX_LS_pc [5] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _14231_ ( .A(\ID_EX_pc [4] ), .B(\EX_LS_pc [4] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _14232_ ( .A(\ID_EX_pc [3] ), .B(\EX_LS_pc [3] ), .S(_06298_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _14233_ ( .A(_06296_ ), .Z(_06299_ ) );
MUX2_X1 _14234_ ( .A(\ID_EX_pc [2] ), .B(\EX_LS_pc [2] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _14235_ ( .A(\ID_EX_pc [29] ), .B(\EX_LS_pc [29] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _14236_ ( .A(\ID_EX_pc [1] ), .B(\EX_LS_pc [1] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _14237_ ( .A(\ID_EX_pc [0] ), .B(\EX_LS_pc [0] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _14238_ ( .A(\ID_EX_pc [28] ), .B(\EX_LS_pc [28] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _14239_ ( .A(\ID_EX_pc [27] ), .B(\EX_LS_pc [27] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _14240_ ( .A(\ID_EX_pc [26] ), .B(\EX_LS_pc [26] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _14241_ ( .A(\ID_EX_pc [25] ), .B(\EX_LS_pc [25] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _14242_ ( .A(\ID_EX_pc [24] ), .B(\EX_LS_pc [24] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _14243_ ( .A(\ID_EX_pc [23] ), .B(\EX_LS_pc [23] ), .S(_06299_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _14244_ ( .A(\ID_EX_pc [22] ), .B(\EX_LS_pc [22] ), .S(_06296_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _14245_ ( .A(\ID_EX_pc [31] ), .B(\EX_LS_pc [31] ), .S(_06296_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
INV_X1 _14246_ ( .A(_02221_ ), .ZN(_06300_ ) );
NOR4_X1 _14247_ ( .A1(_06294_ ), .A2(exception_quest_IDU ), .A3(_06300_ ), .A4(_06295_ ), .ZN(_06301_ ) );
XNOR2_X1 _14248_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_06302_ ) );
XNOR2_X1 _14249_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_06303_ ) );
XNOR2_X1 _14250_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_06304_ ) );
XNOR2_X1 _14251_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_06305_ ) );
AND4_X1 _14252_ ( .A1(_06302_ ), .A2(_06303_ ), .A3(_06304_ ), .A4(_06305_ ), .ZN(_06306_ ) );
XNOR2_X1 _14253_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_06307_ ) );
XNOR2_X1 _14254_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_06308_ ) );
XNOR2_X1 _14255_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_06309_ ) );
XNOR2_X1 _14256_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_06310_ ) );
AND4_X1 _14257_ ( .A1(_06307_ ), .A2(_06308_ ), .A3(_06309_ ), .A4(_06310_ ), .ZN(_06311_ ) );
XNOR2_X1 _14258_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_06312_ ) );
XNOR2_X1 _14259_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_06313_ ) );
XNOR2_X1 _14260_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_06314_ ) );
XNOR2_X1 _14261_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_06315_ ) );
AND4_X1 _14262_ ( .A1(_06312_ ), .A2(_06313_ ), .A3(_06314_ ), .A4(_06315_ ), .ZN(_06316_ ) );
XNOR2_X1 _14263_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_06317_ ) );
XNOR2_X1 _14264_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_06318_ ) );
XNOR2_X1 _14265_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_06319_ ) );
XNOR2_X1 _14266_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_06320_ ) );
AND4_X1 _14267_ ( .A1(_06317_ ), .A2(_06318_ ), .A3(_06319_ ), .A4(_06320_ ), .ZN(_06321_ ) );
AND4_X1 _14268_ ( .A1(_06306_ ), .A2(_06311_ ), .A3(_06316_ ), .A4(_06321_ ), .ZN(_06322_ ) );
XNOR2_X1 _14269_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_06323_ ) );
XNOR2_X1 _14270_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_06324_ ) );
XNOR2_X1 _14271_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_06325_ ) );
XNOR2_X1 _14272_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_06326_ ) );
XNOR2_X1 _14273_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_06327_ ) );
AND4_X1 _14274_ ( .A1(_06324_ ), .A2(_06325_ ), .A3(_06326_ ), .A4(_06327_ ), .ZN(_06328_ ) );
XNOR2_X1 _14275_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_06329_ ) );
XOR2_X1 _14276_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .Z(_06330_ ) );
XOR2_X1 _14277_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .Z(_06331_ ) );
NOR2_X1 _14278_ ( .A1(_06330_ ), .A2(_06331_ ), .ZN(_06332_ ) );
AND4_X1 _14279_ ( .A1(_06323_ ), .A2(_06328_ ), .A3(_06329_ ), .A4(_06332_ ), .ZN(_06333_ ) );
XNOR2_X1 _14280_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_06334_ ) );
XNOR2_X1 _14281_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_06335_ ) );
XNOR2_X1 _14282_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_06336_ ) );
XNOR2_X1 _14283_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_06337_ ) );
NAND4_X1 _14284_ ( .A1(_06334_ ), .A2(_06335_ ), .A3(_06336_ ), .A4(_06337_ ), .ZN(_06338_ ) );
XNOR2_X1 _14285_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_06339_ ) );
XNOR2_X1 _14286_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_06340_ ) );
XNOR2_X1 _14287_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_06341_ ) );
XNOR2_X1 _14288_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_06342_ ) );
NAND4_X1 _14289_ ( .A1(_06339_ ), .A2(_06340_ ), .A3(_06341_ ), .A4(_06342_ ), .ZN(_06343_ ) );
NOR2_X1 _14290_ ( .A1(_06338_ ), .A2(_06343_ ), .ZN(_06344_ ) );
NAND4_X1 _14291_ ( .A1(_06322_ ), .A2(_06333_ ), .A3(excp_written ), .A4(_06344_ ), .ZN(_06345_ ) );
AOI21_X1 _14292_ ( .A(_06301_ ), .B1(_06300_ ), .B2(_06345_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
AND4_X1 _14293_ ( .A1(\ID_EX_typ [7] ), .A2(_04015_ ), .A3(_06134_ ), .A4(IDU_valid_EXU ), .ZN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NAND2_X1 _14294_ ( .A1(_05941_ ), .A2(_03157_ ), .ZN(_06346_ ) );
AND2_X1 _14295_ ( .A1(_03153_ ), .A2(_04017_ ), .ZN(_06347_ ) );
INV_X1 _14296_ ( .A(_06347_ ), .ZN(_06348_ ) );
BUF_X2 _14297_ ( .A(_06348_ ), .Z(_06349_ ) );
BUF_X4 _14298_ ( .A(_06349_ ), .Z(_06350_ ) );
OAI21_X1 _14299_ ( .A(_06346_ ), .B1(_04047_ ), .B2(_06350_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
XNOR2_X1 _14300_ ( .A(_05044_ ), .B(\ID_EX_imm [0] ), .ZN(_06351_ ) );
BUF_X4 _14301_ ( .A(_06347_ ), .Z(_06352_ ) );
BUF_X4 _14302_ ( .A(_06352_ ), .Z(_06353_ ) );
BUF_X4 _14303_ ( .A(_06353_ ), .Z(_06354_ ) );
AOI22_X1 _14304_ ( .A1(_06351_ ), .A2(_03158_ ), .B1(_04059_ ), .B2(_06354_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AND2_X2 _14305_ ( .A1(_03494_ ), .A2(\ID_EX_typ [7] ), .ZN(_06355_ ) );
INV_X1 _14306_ ( .A(_06355_ ), .ZN(_06356_ ) );
BUF_X4 _14307_ ( .A(_06356_ ), .Z(_06357_ ) );
AND2_X1 _14308_ ( .A1(_05774_ ), .A2(_06357_ ), .ZN(_06358_ ) );
BUF_X4 _14309_ ( .A(_06348_ ), .Z(_06359_ ) );
BUF_X4 _14310_ ( .A(_06359_ ), .Z(_06360_ ) );
MUX2_X1 _14311_ ( .A(\ID_EX_csr [10] ), .B(_06358_ ), .S(_06360_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
AOI22_X1 _14312_ ( .A1(_05795_ ), .A2(_03158_ ), .B1(_04050_ ), .B2(_06354_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR2_X1 _14313_ ( .A1(_05813_ ), .A2(_06355_ ), .ZN(_06361_ ) );
MUX2_X1 _14314_ ( .A(\ID_EX_csr [8] ), .B(_06361_ ), .S(_06360_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _14315_ ( .A1(_05832_ ), .A2(_03157_ ), .ZN(_06362_ ) );
OAI21_X1 _14316_ ( .A(_06362_ ), .B1(_04060_ ), .B2(_06350_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
NOR2_X1 _14317_ ( .A1(_05849_ ), .A2(_03153_ ), .ZN(_06363_ ) );
BUF_X4 _14318_ ( .A(_06352_ ), .Z(_06364_ ) );
BUF_X4 _14319_ ( .A(_06364_ ), .Z(_06365_ ) );
AOI21_X1 _14320_ ( .A(_06363_ ), .B1(_04073_ ), .B2(_06365_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _14321_ ( .A1(_05871_ ), .A2(_03157_ ), .ZN(_06366_ ) );
OAI21_X1 _14322_ ( .A(_06366_ ), .B1(_04044_ ), .B2(_06350_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _14323_ ( .A1(_05889_ ), .A2(_03157_ ), .ZN(_06367_ ) );
OAI21_X1 _14324_ ( .A(_06367_ ), .B1(_04034_ ), .B2(_06350_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _14325_ ( .A1(_05908_ ), .A2(_03157_ ), .ZN(_06368_ ) );
OAI21_X1 _14326_ ( .A(_06368_ ), .B1(_04040_ ), .B2(_06350_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _14327_ ( .A1(_05925_ ), .A2(_03157_ ), .ZN(_06369_ ) );
OAI21_X1 _14328_ ( .A(_06369_ ), .B1(_04078_ ), .B2(_06350_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
NAND2_X1 _14329_ ( .A1(_05740_ ), .A2(_03157_ ), .ZN(_06370_ ) );
OAI21_X1 _14330_ ( .A(_06370_ ), .B1(_04070_ ), .B2(_06350_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
BUF_X4 _14331_ ( .A(_06352_ ), .Z(_06371_ ) );
AND3_X1 _14332_ ( .A1(_02443_ ), .A2(_05487_ ), .A3(_02444_ ), .ZN(_06372_ ) );
AND2_X1 _14333_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [21] ), .ZN(_06373_ ) );
BUF_X4 _14334_ ( .A(_05326_ ), .Z(_06374_ ) );
OAI221_X1 _14335_ ( .A(_06371_ ), .B1(_06372_ ), .B2(_06373_ ), .C1(_06079_ ), .C2(_06374_ ), .ZN(_06375_ ) );
NAND2_X1 _14336_ ( .A1(_06075_ ), .A2(_06074_ ), .ZN(_06376_ ) );
AOI21_X1 _14337_ ( .A(_06376_ ), .B1(_05478_ ), .B2(_05699_ ), .ZN(_06377_ ) );
NAND4_X1 _14338_ ( .A1(_06377_ ), .A2(_05722_ ), .A3(_06077_ ), .A4(_06076_ ), .ZN(_06378_ ) );
NOR2_X1 _14339_ ( .A1(_05319_ ), .A2(\ID_EX_typ [2] ), .ZN(_06379_ ) );
BUF_X4 _14340_ ( .A(_06379_ ), .Z(_06380_ ) );
NAND4_X1 _14341_ ( .A1(_05704_ ), .A2(_05699_ ), .A3(_06072_ ), .A4(_05706_ ), .ZN(_06381_ ) );
NAND4_X1 _14342_ ( .A1(_06378_ ), .A2(_06380_ ), .A3(_06381_ ), .A4(_06371_ ), .ZN(_06382_ ) );
MUX2_X1 _14343_ ( .A(_06082_ ), .B(_04490_ ), .S(_06357_ ), .Z(_06383_ ) );
BUF_X4 _14344_ ( .A(_06353_ ), .Z(_06384_ ) );
OAI211_X1 _14345_ ( .A(_06375_ ), .B(_06382_ ), .C1(_06383_ ), .C2(_06384_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
BUF_X4 _14346_ ( .A(_06352_ ), .Z(_06385_ ) );
NAND3_X1 _14347_ ( .A1(_05510_ ), .A2(_06380_ ), .A3(_06385_ ), .ZN(_06386_ ) );
BUF_X4 _14348_ ( .A(_06356_ ), .Z(_06387_ ) );
MUX2_X1 _14349_ ( .A(_06080_ ), .B(_04466_ ), .S(_06387_ ), .Z(_06388_ ) );
OAI221_X1 _14350_ ( .A(_06364_ ), .B1(_05981_ ), .B2(\ID_EX_imm [20] ), .C1(_05510_ ), .C2(_06374_ ), .ZN(_06389_ ) );
AOI21_X1 _14351_ ( .A(fanout_net_7 ), .B1(_02420_ ), .B2(_02421_ ), .ZN(_06390_ ) );
OAI221_X1 _14352_ ( .A(_06386_ ), .B1(_06354_ ), .B2(_06388_ ), .C1(_06389_ ), .C2(_06390_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
INV_X1 _14353_ ( .A(_06379_ ), .ZN(_06391_ ) );
AOI21_X1 _14354_ ( .A(_06391_ ), .B1(_05547_ ), .B2(_05550_ ), .ZN(_06392_ ) );
AOI22_X1 _14355_ ( .A1(_05551_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02941_ ), .ZN(_06393_ ) );
OR2_X1 _14356_ ( .A1(_02940_ ), .A2(fanout_net_7 ), .ZN(_06394_ ) );
AOI211_X1 _14357_ ( .A(_06349_ ), .B(_06392_ ), .C1(_06393_ ), .C2(_06394_ ), .ZN(_06395_ ) );
MUX2_X1 _14358_ ( .A(_04213_ ), .B(_04312_ ), .S(_06357_ ), .Z(_06396_ ) );
AOI21_X1 _14359_ ( .A(_06395_ ), .B1(_06350_ ), .B2(_06396_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _14360_ ( .A1(_05577_ ), .A2(_06380_ ), .A3(_06385_ ), .ZN(_06397_ ) );
AND3_X1 _14361_ ( .A1(_02897_ ), .A2(_05488_ ), .A3(_02916_ ), .ZN(_06398_ ) );
OAI221_X1 _14362_ ( .A(_06353_ ), .B1(_05488_ ), .B2(\ID_EX_imm [18] ), .C1(_05577_ ), .C2(_06374_ ), .ZN(_06399_ ) );
MUX2_X1 _14363_ ( .A(_05556_ ), .B(_04338_ ), .S(_06357_ ), .Z(_06400_ ) );
OAI221_X1 _14364_ ( .A(_06397_ ), .B1(_06398_ ), .B2(_06399_ ), .C1(_06400_ ), .C2(_06354_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
BUF_X4 _14365_ ( .A(_06352_ ), .Z(_06401_ ) );
OAI22_X1 _14366_ ( .A1(_05594_ ), .A2(_05326_ ), .B1(_05487_ ), .B2(\ID_EX_imm [17] ), .ZN(_06402_ ) );
AOI21_X1 _14367_ ( .A(_06402_ ), .B1(_05604_ ), .B2(_04372_ ), .ZN(_06403_ ) );
BUF_X4 _14368_ ( .A(_06379_ ), .Z(_06404_ ) );
NAND3_X1 _14369_ ( .A1(_05591_ ), .A2(_06404_ ), .A3(_05593_ ), .ZN(_06405_ ) );
INV_X1 _14370_ ( .A(_06405_ ), .ZN(_06406_ ) );
OAI21_X1 _14371_ ( .A(_06401_ ), .B1(_06403_ ), .B2(_06406_ ), .ZN(_06407_ ) );
AND4_X1 _14372_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06408_ ) );
INV_X1 _14373_ ( .A(_04393_ ), .ZN(_06409_ ) );
BUF_X4 _14374_ ( .A(_06387_ ), .Z(_06410_ ) );
AOI21_X1 _14375_ ( .A(_06408_ ), .B1(_06409_ ), .B2(_06410_ ), .ZN(_06411_ ) );
OAI21_X1 _14376_ ( .A(_06407_ ), .B1(_06365_ ), .B2(_06411_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
NAND3_X1 _14377_ ( .A1(_05620_ ), .A2(_06380_ ), .A3(_06385_ ), .ZN(_06412_ ) );
MUX2_X1 _14378_ ( .A(_05599_ ), .B(_04370_ ), .S(_06387_ ), .Z(_06413_ ) );
OAI221_X1 _14379_ ( .A(_06364_ ), .B1(_05981_ ), .B2(\ID_EX_imm [16] ), .C1(_05620_ ), .C2(_06374_ ), .ZN(_06414_ ) );
AOI21_X1 _14380_ ( .A(fanout_net_7 ), .B1(_02470_ ), .B2(_02471_ ), .ZN(_06415_ ) );
OAI221_X1 _14381_ ( .A(_06412_ ), .B1(_06354_ ), .B2(_06413_ ), .C1(_06414_ ), .C2(_06415_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
AND3_X1 _14382_ ( .A1(_02813_ ), .A2(_05428_ ), .A3(_02814_ ), .ZN(_06416_ ) );
AND2_X1 _14383_ ( .A1(fanout_net_7 ), .A2(\ID_EX_imm [15] ), .ZN(_06417_ ) );
OAI221_X1 _14384_ ( .A(_06371_ ), .B1(_05633_ ), .B2(_06374_ ), .C1(_06416_ ), .C2(_06417_ ), .ZN(_06418_ ) );
AOI21_X1 _14385_ ( .A(_05625_ ), .B1(_05478_ ), .B2(_05699_ ), .ZN(_06419_ ) );
AND2_X1 _14386_ ( .A1(_05628_ ), .A2(_05574_ ), .ZN(_06420_ ) );
NAND4_X1 _14387_ ( .A1(_06419_ ), .A2(_05630_ ), .A3(_05627_ ), .A4(_06420_ ), .ZN(_06421_ ) );
NAND4_X1 _14388_ ( .A1(_05704_ ), .A2(_05699_ ), .A3(_06268_ ), .A4(_05706_ ), .ZN(_06422_ ) );
NAND4_X1 _14389_ ( .A1(_06421_ ), .A2(_06404_ ), .A3(_06422_ ), .A4(_06371_ ), .ZN(_06423_ ) );
MUX2_X1 _14390_ ( .A(_05635_ ), .B(_04706_ ), .S(_06357_ ), .Z(_06424_ ) );
OAI211_X1 _14391_ ( .A(_06418_ ), .B(_06423_ ), .C1(_06424_ ), .C2(_06354_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
OAI22_X1 _14392_ ( .A1(_05661_ ), .A2(_05326_ ), .B1(_05487_ ), .B2(\ID_EX_imm [14] ), .ZN(_06425_ ) );
AOI21_X1 _14393_ ( .A(_06425_ ), .B1(_05604_ ), .B2(_04708_ ), .ZN(_06426_ ) );
OR3_X1 _14394_ ( .A1(_05658_ ), .A2(_06391_ ), .A3(_05660_ ), .ZN(_06427_ ) );
INV_X1 _14395_ ( .A(_06427_ ), .ZN(_06428_ ) );
OAI21_X1 _14396_ ( .A(_06401_ ), .B1(_06426_ ), .B2(_06428_ ), .ZN(_06429_ ) );
MUX2_X1 _14397_ ( .A(_05664_ ), .B(_04731_ ), .S(_06357_ ), .Z(_06430_ ) );
OAI21_X1 _14398_ ( .A(_06429_ ), .B1(_06365_ ), .B2(_06430_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OR3_X1 _14399_ ( .A1(_05677_ ), .A2(_06391_ ), .A3(_05679_ ), .ZN(_06431_ ) );
OAI22_X1 _14400_ ( .A1(_05680_ ), .A2(_05326_ ), .B1(_05428_ ), .B2(\ID_EX_imm [13] ), .ZN(_06432_ ) );
AOI21_X1 _14401_ ( .A(fanout_net_7 ), .B1(_02860_ ), .B2(_02861_ ), .ZN(_06433_ ) );
OAI211_X1 _14402_ ( .A(_06353_ ), .B(_06431_ ), .C1(_06432_ ), .C2(_06433_ ), .ZN(_06434_ ) );
NAND4_X1 _14403_ ( .A1(\ID_EX_pc [13] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06435_ ) );
OAI211_X1 _14404_ ( .A(_06349_ ), .B(_06435_ ), .C1(_04780_ ), .C2(_06355_ ), .ZN(_06436_ ) );
AND2_X1 _14405_ ( .A1(_06434_ ), .A2(_06436_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AND4_X1 _14406_ ( .A1(_05696_ ), .A2(_05702_ ), .A3(_05697_ ), .A4(_05701_ ), .ZN(_06437_ ) );
NAND4_X1 _14407_ ( .A1(_04069_ ), .A2(_05722_ ), .A3(_05574_ ), .A4(_06437_ ), .ZN(_06438_ ) );
NAND3_X1 _14408_ ( .A1(_05562_ ), .A2(_05705_ ), .A3(_05563_ ), .ZN(_06439_ ) );
NAND4_X1 _14409_ ( .A1(_06438_ ), .A2(_06404_ ), .A3(_06439_ ), .A4(_06353_ ), .ZN(_06440_ ) );
BUF_X4 _14410_ ( .A(_06352_ ), .Z(_06441_ ) );
MUX2_X1 _14411_ ( .A(_05690_ ), .B(_04756_ ), .S(_06387_ ), .Z(_06442_ ) );
AND2_X1 _14412_ ( .A1(_06438_ ), .A2(_06439_ ), .ZN(_06443_ ) );
OAI221_X1 _14413_ ( .A(_06371_ ), .B1(_05981_ ), .B2(\ID_EX_imm [12] ), .C1(_06443_ ), .C2(_06374_ ), .ZN(_06444_ ) );
AOI21_X1 _14414_ ( .A(fanout_net_7 ), .B1(_02884_ ), .B2(_02885_ ), .ZN(_06445_ ) );
OAI221_X1 _14415_ ( .A(_06440_ ), .B1(_06441_ ), .B2(_06442_ ), .C1(_06444_ ), .C2(_06445_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
NAND3_X1 _14416_ ( .A1(_04110_ ), .A2(_06380_ ), .A3(_06385_ ), .ZN(_06446_ ) );
AND4_X1 _14417_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06447_ ) );
AOI21_X1 _14418_ ( .A(_06447_ ), .B1(_04581_ ), .B2(_06410_ ), .ZN(_06448_ ) );
OAI221_X1 _14419_ ( .A(_06371_ ), .B1(_05604_ ), .B2(\ID_EX_imm [30] ), .C1(_04110_ ), .C2(_06374_ ), .ZN(_06449_ ) );
AND3_X1 _14420_ ( .A1(_02295_ ), .A2(_05604_ ), .A3(_02296_ ), .ZN(_06450_ ) );
OAI221_X1 _14421_ ( .A(_06446_ ), .B1(_06441_ ), .B2(_06448_ ), .C1(_06449_ ), .C2(_06450_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
NOR2_X1 _14422_ ( .A1(_05487_ ), .A2(\ID_EX_imm [11] ), .ZN(_06451_ ) );
NAND2_X1 _14423_ ( .A1(_05728_ ), .A2(_05730_ ), .ZN(_06452_ ) );
AOI21_X1 _14424_ ( .A(_06451_ ), .B1(_06452_ ), .B2(\ID_EX_typ [2] ), .ZN(_06453_ ) );
OR2_X1 _14425_ ( .A1(_04783_ ), .A2(fanout_net_7 ), .ZN(_06454_ ) );
AND2_X1 _14426_ ( .A1(_06453_ ), .A2(_06454_ ), .ZN(_06455_ ) );
AND3_X1 _14427_ ( .A1(_05728_ ), .A2(_06379_ ), .A3(_05730_ ), .ZN(_06456_ ) );
OAI21_X1 _14428_ ( .A(_06401_ ), .B1(_06455_ ), .B2(_06456_ ), .ZN(_06457_ ) );
MUX2_X1 _14429_ ( .A(_05713_ ), .B(_04806_ ), .S(_06357_ ), .Z(_06458_ ) );
OAI21_X1 _14430_ ( .A(_06457_ ), .B1(_06365_ ), .B2(_06458_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
NAND3_X1 _14431_ ( .A1(_05772_ ), .A2(_06380_ ), .A3(_06385_ ), .ZN(_06459_ ) );
AOI21_X1 _14432_ ( .A(fanout_net_7 ), .B1(_02569_ ), .B2(_02570_ ), .ZN(_06460_ ) );
OAI221_X1 _14433_ ( .A(_06353_ ), .B1(_05488_ ), .B2(\ID_EX_imm [10] ), .C1(_05772_ ), .C2(_06374_ ), .ZN(_06461_ ) );
MUX2_X1 _14434_ ( .A(_05758_ ), .B(_04829_ ), .S(_06387_ ), .Z(_06462_ ) );
OAI221_X1 _14435_ ( .A(_06459_ ), .B1(_06460_ ), .B2(_06461_ ), .C1(_06462_ ), .C2(_06354_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
NAND3_X1 _14436_ ( .A1(_05783_ ), .A2(_06380_ ), .A3(_06385_ ), .ZN(_06463_ ) );
AOI21_X1 _14437_ ( .A(fanout_net_7 ), .B1(_02520_ ), .B2(_02521_ ), .ZN(_06464_ ) );
OAI221_X1 _14438_ ( .A(_06352_ ), .B1(_05488_ ), .B2(\ID_EX_imm [9] ), .C1(_05783_ ), .C2(_05326_ ), .ZN(_06465_ ) );
MUX2_X1 _14439_ ( .A(_05784_ ), .B(_04854_ ), .S(_06387_ ), .Z(_06466_ ) );
OAI221_X1 _14440_ ( .A(_06463_ ), .B1(_06464_ ), .B2(_06465_ ), .C1(_06466_ ), .C2(_06354_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
BUF_X4 _14441_ ( .A(_06352_ ), .Z(_06467_ ) );
AOI22_X1 _14442_ ( .A1(_05806_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02499_ ), .ZN(_06468_ ) );
OR2_X1 _14443_ ( .A1(_02498_ ), .A2(fanout_net_7 ), .ZN(_06469_ ) );
AND2_X1 _14444_ ( .A1(_06468_ ), .A2(_06469_ ), .ZN(_06470_ ) );
AND3_X1 _14445_ ( .A1(_05803_ ), .A2(_06379_ ), .A3(_05805_ ), .ZN(_06471_ ) );
OAI21_X1 _14446_ ( .A(_06467_ ), .B1(_06470_ ), .B2(_06471_ ), .ZN(_06472_ ) );
MUX2_X1 _14447_ ( .A(_05808_ ), .B(_04877_ ), .S(_06357_ ), .Z(_06473_ ) );
OAI21_X1 _14448_ ( .A(_06472_ ), .B1(_06365_ ), .B2(_06473_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
OAI22_X1 _14449_ ( .A1(_05826_ ), .A2(_05326_ ), .B1(_05487_ ), .B2(\ID_EX_imm [7] ), .ZN(_06474_ ) );
AOI211_X1 _14450_ ( .A(_06359_ ), .B(_06474_ ), .C1(_05604_ ), .C2(_04907_ ), .ZN(_06475_ ) );
NAND2_X1 _14451_ ( .A1(_04928_ ), .A2(_06356_ ), .ZN(_06476_ ) );
OR4_X1 _14452_ ( .A1(\ID_EX_pc [7] ), .A2(_03495_ ), .A3(_04015_ ), .A4(_04017_ ), .ZN(_06477_ ) );
AND3_X1 _14453_ ( .A1(_06476_ ), .A2(_06359_ ), .A3(_06477_ ), .ZN(_06478_ ) );
NAND4_X1 _14454_ ( .A1(_05821_ ), .A2(_05822_ ), .A3(_05823_ ), .A4(_05824_ ), .ZN(_06479_ ) );
AOI21_X1 _14455_ ( .A(_06479_ ), .B1(_05478_ ), .B2(_05699_ ), .ZN(_06480_ ) );
AND4_X1 _14456_ ( .A1(_06247_ ), .A2(_05465_ ), .A3(_05469_ ), .A4(_05479_ ), .ZN(_06481_ ) );
NOR4_X1 _14457_ ( .A1(_06480_ ), .A2(_06481_ ), .A3(_06391_ ), .A4(_06348_ ), .ZN(_06482_ ) );
OR3_X1 _14458_ ( .A1(_06475_ ), .A2(_06478_ ), .A3(_06482_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
NAND3_X1 _14459_ ( .A1(_05847_ ), .A2(_06380_ ), .A3(_06385_ ), .ZN(_06483_ ) );
MUX2_X1 _14460_ ( .A(_05834_ ), .B(_04904_ ), .S(_06387_ ), .Z(_06484_ ) );
AND3_X1 _14461_ ( .A1(_02650_ ), .A2(_05604_ ), .A3(_02669_ ), .ZN(_06485_ ) );
OAI221_X1 _14462_ ( .A(_06353_ ), .B1(_05604_ ), .B2(\ID_EX_imm [6] ), .C1(_05847_ ), .C2(_06374_ ), .ZN(_06486_ ) );
OAI221_X1 _14463_ ( .A(_06483_ ), .B1(_06484_ ), .B2(_06401_ ), .C1(_06485_ ), .C2(_06486_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
AND4_X1 _14464_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06487_ ) );
AOI211_X1 _14465_ ( .A(_06352_ ), .B(_06487_ ), .C1(_04973_ ), .C2(_06410_ ), .ZN(_06488_ ) );
NAND3_X1 _14466_ ( .A1(_05857_ ), .A2(_06404_ ), .A3(_05859_ ), .ZN(_06489_ ) );
INV_X1 _14467_ ( .A(_06489_ ), .ZN(_06490_ ) );
NOR2_X1 _14468_ ( .A1(_05428_ ), .A2(\ID_EX_imm [5] ), .ZN(_06491_ ) );
NAND2_X1 _14469_ ( .A1(_05857_ ), .A2(_05859_ ), .ZN(_06492_ ) );
AOI21_X1 _14470_ ( .A(_06491_ ), .B1(_06492_ ), .B2(\ID_EX_typ [2] ), .ZN(_06493_ ) );
OR2_X1 _14471_ ( .A1(_02598_ ), .A2(fanout_net_7 ), .ZN(_06494_ ) );
AOI21_X1 _14472_ ( .A(_06490_ ), .B1(_06493_ ), .B2(_06494_ ), .ZN(_06495_ ) );
AOI21_X1 _14473_ ( .A(_06488_ ), .B1(_06495_ ), .B2(_06365_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
INV_X1 _14474_ ( .A(_05879_ ), .ZN(_06496_ ) );
NAND4_X1 _14475_ ( .A1(_06496_ ), .A2(_05880_ ), .A3(_05881_ ), .A4(_05882_ ), .ZN(_06497_ ) );
AOI211_X1 _14476_ ( .A(_04102_ ), .B(_06497_ ), .C1(_05490_ ), .C2(_05492_ ), .ZN(_06498_ ) );
AND3_X1 _14477_ ( .A1(_04054_ ), .A2(_05885_ ), .A3(_04066_ ), .ZN(_06499_ ) );
OR3_X1 _14478_ ( .A1(_06498_ ), .A2(_06391_ ), .A3(_06499_ ), .ZN(_06500_ ) );
INV_X1 _14479_ ( .A(_06500_ ), .ZN(_06501_ ) );
OR2_X1 _14480_ ( .A1(_06498_ ), .A2(_06499_ ), .ZN(_06502_ ) );
AOI22_X1 _14481_ ( .A1(_06502_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_7 ), .B2(_02600_ ), .ZN(_06503_ ) );
OR2_X1 _14482_ ( .A1(_02622_ ), .A2(\ID_EX_typ [0] ), .ZN(_06504_ ) );
AOI21_X1 _14483_ ( .A(_06501_ ), .B1(_06503_ ), .B2(_06504_ ), .ZN(_06505_ ) );
NAND2_X1 _14484_ ( .A1(_06505_ ), .A2(_06385_ ), .ZN(_06506_ ) );
NAND4_X1 _14485_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06507_ ) );
OAI211_X1 _14486_ ( .A(_06349_ ), .B(_06507_ ), .C1(_04951_ ), .C2(_06355_ ), .ZN(_06508_ ) );
AND2_X1 _14487_ ( .A1(_06506_ ), .A2(_06508_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
OAI22_X1 _14488_ ( .A1(_05900_ ), .A2(_05326_ ), .B1(_05487_ ), .B2(\ID_EX_imm [3] ), .ZN(_06509_ ) );
AOI21_X1 _14489_ ( .A(_06509_ ), .B1(_05604_ ), .B2(_02781_ ), .ZN(_06510_ ) );
NOR3_X1 _14490_ ( .A1(_05897_ ), .A2(_06391_ ), .A3(_05899_ ), .ZN(_06511_ ) );
OAI21_X1 _14491_ ( .A(_06467_ ), .B1(_06510_ ), .B2(_06511_ ), .ZN(_06512_ ) );
AND4_X1 _14492_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06513_ ) );
AOI21_X1 _14493_ ( .A(_06513_ ), .B1(_05041_ ), .B2(_06410_ ), .ZN(_06514_ ) );
OAI21_X1 _14494_ ( .A(_06512_ ), .B1(_06365_ ), .B2(_06514_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
AOI21_X1 _14495_ ( .A(_05911_ ), .B1(_05478_ ), .B2(_05479_ ), .ZN(_06515_ ) );
AND2_X1 _14496_ ( .A1(_05914_ ), .A2(_05574_ ), .ZN(_06516_ ) );
NAND4_X1 _14497_ ( .A1(_06515_ ), .A2(_05916_ ), .A3(_05913_ ), .A4(_06516_ ), .ZN(_06517_ ) );
NAND4_X1 _14498_ ( .A1(_05704_ ), .A2(_05699_ ), .A3(_06238_ ), .A4(_05706_ ), .ZN(_06518_ ) );
NAND2_X1 _14499_ ( .A1(_06517_ ), .A2(_06518_ ), .ZN(_06519_ ) );
AOI22_X1 _14500_ ( .A1(_06519_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02775_ ), .ZN(_06520_ ) );
OAI211_X1 _14501_ ( .A(_06520_ ), .B(_06467_ ), .C1(\ID_EX_typ [0] ), .C2(_02774_ ), .ZN(_06521_ ) );
BUF_X4 _14502_ ( .A(_06359_ ), .Z(_06522_ ) );
AND3_X1 _14503_ ( .A1(_05000_ ), .A2(_05019_ ), .A3(_06387_ ), .ZN(_06523_ ) );
AND3_X1 _14504_ ( .A1(_03494_ ), .A2(\ID_EX_pc [2] ), .A3(\ID_EX_typ [7] ), .ZN(_06524_ ) );
OAI21_X1 _14505_ ( .A(_06522_ ), .B1(_06523_ ), .B2(_06524_ ), .ZN(_06525_ ) );
NAND4_X1 _14506_ ( .A1(_06517_ ), .A2(_06380_ ), .A3(_06518_ ), .A4(_06385_ ), .ZN(_06526_ ) );
NAND3_X1 _14507_ ( .A1(_06521_ ), .A2(_06525_ ), .A3(_06526_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
AOI221_X4 _14508_ ( .A(_06348_ ), .B1(\ID_EX_typ [0] ), .B2(_03119_ ), .C1(_05456_ ), .C2(\ID_EX_typ [2] ), .ZN(_06527_ ) );
OAI21_X1 _14509_ ( .A(_06527_ ), .B1(\ID_EX_typ [0] ), .B2(_03118_ ), .ZN(_06528_ ) );
NOR3_X1 _14510_ ( .A1(_05453_ ), .A2(_05455_ ), .A3(_06359_ ), .ZN(_06529_ ) );
NAND2_X1 _14511_ ( .A1(_06529_ ), .A2(_06380_ ), .ZN(_06530_ ) );
AND4_X1 _14512_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06531_ ) );
AOI21_X1 _14513_ ( .A(_06531_ ), .B1(_04536_ ), .B2(_06410_ ), .ZN(_06532_ ) );
OAI211_X1 _14514_ ( .A(_06528_ ), .B(_06530_ ), .C1(_06365_ ), .C2(_06532_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
NAND4_X1 _14515_ ( .A1(_05704_ ), .A2(_05479_ ), .A3(_06239_ ), .A4(_05706_ ), .ZN(_06533_ ) );
NAND4_X1 _14516_ ( .A1(_05931_ ), .A2(_05932_ ), .A3(_05933_ ), .A4(_05934_ ), .ZN(_06534_ ) );
OAI211_X1 _14517_ ( .A(_06379_ ), .B(_06533_ ), .C1(_05983_ ), .C2(_06534_ ), .ZN(_06535_ ) );
INV_X1 _14518_ ( .A(_06535_ ), .ZN(_06536_ ) );
AOI22_X1 _14519_ ( .A1(_05938_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02705_ ), .ZN(_06537_ ) );
OR2_X1 _14520_ ( .A1(_02704_ ), .A2(\ID_EX_typ [0] ), .ZN(_06538_ ) );
AOI211_X1 _14521_ ( .A(_06349_ ), .B(_06536_ ), .C1(_06537_ ), .C2(_06538_ ), .ZN(_06539_ ) );
MUX2_X1 _14522_ ( .A(_05929_ ), .B(_04997_ ), .S(_06357_ ), .Z(_06540_ ) );
AOI21_X1 _14523_ ( .A(_06539_ ), .B1(_06350_ ), .B2(_06540_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
AOI21_X1 _14524_ ( .A(_06391_ ), .B1(_05977_ ), .B2(_05978_ ), .ZN(_06541_ ) );
AOI21_X1 _14525_ ( .A(_06541_ ), .B1(\ID_EX_typ [0] ), .B2(\ID_EX_imm [0] ), .ZN(_06542_ ) );
OAI21_X1 _14526_ ( .A(_06542_ ), .B1(\ID_EX_typ [0] ), .B2(_05158_ ), .ZN(_06543_ ) );
AND2_X1 _14527_ ( .A1(_05977_ ), .A2(_05978_ ), .ZN(_06544_ ) );
AOI21_X1 _14528_ ( .A(_06359_ ), .B1(_06544_ ), .B2(\ID_EX_typ [2] ), .ZN(_06545_ ) );
AND2_X1 _14529_ ( .A1(_06543_ ), .A2(_06545_ ), .ZN(_06546_ ) );
AND4_X1 _14530_ ( .A1(_05967_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06547_ ) );
AOI211_X1 _14531_ ( .A(_06352_ ), .B(_06547_ ), .C1(_05065_ ), .C2(_06357_ ), .ZN(_06548_ ) );
OR2_X1 _14532_ ( .A1(_06546_ ), .A2(_06548_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
AOI21_X1 _14533_ ( .A(_05752_ ), .B1(_05478_ ), .B2(_05479_ ), .ZN(_06549_ ) );
NAND3_X1 _14534_ ( .A1(_04094_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_04106_ ), .ZN(_06550_ ) );
AND2_X1 _14535_ ( .A1(_05749_ ), .A2(_06550_ ), .ZN(_06551_ ) );
NAND4_X1 _14536_ ( .A1(_06549_ ), .A2(_05722_ ), .A3(_05748_ ), .A4(_06551_ ), .ZN(_06552_ ) );
NAND4_X1 _14537_ ( .A1(_05704_ ), .A2(_05479_ ), .A3(_05746_ ), .A4(_05706_ ), .ZN(_06553_ ) );
NAND2_X1 _14538_ ( .A1(_06552_ ), .A2(_06553_ ), .ZN(_06554_ ) );
AOI22_X1 _14539_ ( .A1(_06554_ ), .A2(\ID_EX_typ [2] ), .B1(_05100_ ), .B2(_05428_ ), .ZN(_06555_ ) );
OAI211_X1 _14540_ ( .A(_06555_ ), .B(_06364_ ), .C1(_05981_ ), .C2(\ID_EX_imm [28] ), .ZN(_06556_ ) );
NAND4_X1 _14541_ ( .A1(_06552_ ), .A2(_06404_ ), .A3(_06553_ ), .A4(_06371_ ), .ZN(_06557_ ) );
AND3_X1 _14542_ ( .A1(_03494_ ), .A2(\ID_EX_pc [28] ), .A3(\ID_EX_typ [7] ), .ZN(_06558_ ) );
AOI21_X1 _14543_ ( .A(_06558_ ), .B1(_04514_ ), .B2(_06410_ ), .ZN(_06559_ ) );
OAI211_X1 _14544_ ( .A(_06556_ ), .B(_06557_ ), .C1(_06365_ ), .C2(_06559_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _14545_ ( .A(_05958_ ), .B1(_05478_ ), .B2(_05474_ ), .ZN(_06560_ ) );
NAND3_X1 _14546_ ( .A1(_04094_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_04106_ ), .ZN(_06561_ ) );
AND2_X1 _14547_ ( .A1(_05955_ ), .A2(_06561_ ), .ZN(_06562_ ) );
NAND4_X1 _14548_ ( .A1(_06560_ ), .A2(_05722_ ), .A3(_05954_ ), .A4(_06562_ ), .ZN(_06563_ ) );
NAND4_X1 _14549_ ( .A1(_05704_ ), .A2(_05479_ ), .A3(_05952_ ), .A4(_05706_ ), .ZN(_06564_ ) );
NAND2_X1 _14550_ ( .A1(_06563_ ), .A2(_06564_ ), .ZN(_06565_ ) );
AOI22_X1 _14551_ ( .A1(_06565_ ), .A2(\ID_EX_typ [2] ), .B1(_05307_ ), .B2(_05428_ ), .ZN(_06566_ ) );
OAI211_X1 _14552_ ( .A(_06566_ ), .B(_06364_ ), .C1(_05981_ ), .C2(\ID_EX_imm [27] ), .ZN(_06567_ ) );
NAND4_X1 _14553_ ( .A1(_06563_ ), .A2(_06404_ ), .A3(_06564_ ), .A4(_06371_ ), .ZN(_06568_ ) );
AND3_X1 _14554_ ( .A1(_03494_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_06569_ ) );
AOI21_X1 _14555_ ( .A(_06569_ ), .B1(_04628_ ), .B2(_06410_ ), .ZN(_06570_ ) );
OAI211_X1 _14556_ ( .A(_06567_ ), .B(_06568_ ), .C1(_06365_ ), .C2(_06570_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
AND3_X1 _14557_ ( .A1(_05548_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_05549_ ), .ZN(_06571_ ) );
AND2_X1 _14558_ ( .A1(_05986_ ), .A2(_05988_ ), .ZN(_06572_ ) );
AND2_X1 _14559_ ( .A1(_05987_ ), .A2(_05989_ ), .ZN(_06573_ ) );
AOI22_X1 _14560_ ( .A1(_05548_ ), .A2(_05549_ ), .B1(_06572_ ), .B2(_06573_ ), .ZN(_06574_ ) );
NOR2_X1 _14561_ ( .A1(_06571_ ), .A2(_06574_ ), .ZN(_06575_ ) );
AOI22_X1 _14562_ ( .A1(_06575_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_03064_ ), .ZN(_06576_ ) );
OAI211_X1 _14563_ ( .A(_06576_ ), .B(_06364_ ), .C1(\ID_EX_typ [0] ), .C2(_03063_ ), .ZN(_06577_ ) );
OR2_X1 _14564_ ( .A1(_05984_ ), .A2(\EX_LS_result_csreg_mem [26] ), .ZN(_06578_ ) );
OR2_X1 _14565_ ( .A1(_05983_ ), .A2(_05990_ ), .ZN(_06579_ ) );
NAND4_X1 _14566_ ( .A1(_06578_ ), .A2(_06404_ ), .A3(_06579_ ), .A4(_06371_ ), .ZN(_06580_ ) );
AND3_X1 _14567_ ( .A1(_03494_ ), .A2(\ID_EX_pc [26] ), .A3(\ID_EX_typ [7] ), .ZN(_06581_ ) );
AOI21_X1 _14568_ ( .A(_06581_ ), .B1(_04605_ ), .B2(_06410_ ), .ZN(_06582_ ) );
OAI211_X1 _14569_ ( .A(_06577_ ), .B(_06580_ ), .C1(_06384_ ), .C2(_06582_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND4_X1 _14570_ ( .A1(_06014_ ), .A2(_06015_ ), .A3(_06016_ ), .A4(_06017_ ), .ZN(_06583_ ) );
OR2_X1 _14571_ ( .A1(_05983_ ), .A2(_06583_ ), .ZN(_06584_ ) );
OAI21_X1 _14572_ ( .A(_06584_ ), .B1(\EX_LS_result_csreg_mem [25] ), .B2(_05984_ ), .ZN(_06585_ ) );
AOI22_X1 _14573_ ( .A1(_06585_ ), .A2(\ID_EX_typ [2] ), .B1(_05428_ ), .B2(_03040_ ), .ZN(_06586_ ) );
OAI211_X1 _14574_ ( .A(_06586_ ), .B(_06364_ ), .C1(_05981_ ), .C2(\ID_EX_imm [25] ), .ZN(_06587_ ) );
OR2_X1 _14575_ ( .A1(_05984_ ), .A2(\EX_LS_result_csreg_mem [25] ), .ZN(_06588_ ) );
NAND4_X1 _14576_ ( .A1(_06588_ ), .A2(_06404_ ), .A3(_06584_ ), .A4(_06371_ ), .ZN(_06589_ ) );
AND3_X1 _14577_ ( .A1(_03494_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06590_ ) );
AOI21_X1 _14578_ ( .A(_06590_ ), .B1(_04652_ ), .B2(_06410_ ), .ZN(_06591_ ) );
OAI211_X1 _14579_ ( .A(_06587_ ), .B(_06589_ ), .C1(_06384_ ), .C2(_06591_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
NAND4_X1 _14580_ ( .A1(_06005_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06592_ ) );
OAI211_X1 _14581_ ( .A(_06360_ ), .B(_06592_ ), .C1(_04674_ ), .C2(_06355_ ), .ZN(_06593_ ) );
NAND3_X1 _14582_ ( .A1(_06027_ ), .A2(_06379_ ), .A3(_06033_ ), .ZN(_06594_ ) );
OAI21_X1 _14583_ ( .A(_06594_ ), .B1(_05604_ ), .B2(_03197_ ), .ZN(_06595_ ) );
AOI21_X1 _14584_ ( .A(_06595_ ), .B1(_05981_ ), .B2(_03196_ ), .ZN(_06596_ ) );
OAI21_X1 _14585_ ( .A(_06467_ ), .B1(_06034_ ), .B2(_06374_ ), .ZN(_06597_ ) );
OAI21_X1 _14586_ ( .A(_06593_ ), .B1(_06596_ ), .B2(_06597_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND4_X1 _14587_ ( .A1(_05704_ ), .A2(_05479_ ), .A3(_06267_ ), .A4(_05706_ ), .ZN(_06598_ ) );
OAI21_X1 _14588_ ( .A(_06598_ ), .B1(_05983_ ), .B2(_06051_ ), .ZN(_06599_ ) );
AOI22_X1 _14589_ ( .A1(_06599_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(_02397_ ), .ZN(_06600_ ) );
OAI211_X1 _14590_ ( .A(_06600_ ), .B(_06364_ ), .C1(\ID_EX_typ [0] ), .C2(_02396_ ), .ZN(_06601_ ) );
OR3_X1 _14591_ ( .A1(_06599_ ), .A2(_06391_ ), .A3(_06359_ ), .ZN(_06602_ ) );
MUX2_X1 _14592_ ( .A(_04211_ ), .B(_04441_ ), .S(_06387_ ), .Z(_06603_ ) );
OAI211_X1 _14593_ ( .A(_06601_ ), .B(_06602_ ), .C1(_06384_ ), .C2(_06603_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
AOI21_X1 _14594_ ( .A(_06061_ ), .B1(_05477_ ), .B2(_05474_ ), .ZN(_06604_ ) );
INV_X1 _14595_ ( .A(_06063_ ), .ZN(_06605_ ) );
INV_X1 _14596_ ( .A(_06062_ ), .ZN(_06606_ ) );
NAND4_X1 _14597_ ( .A1(_06604_ ), .A2(_05586_ ), .A3(_06605_ ), .A4(_06606_ ), .ZN(_06607_ ) );
NAND4_X1 _14598_ ( .A1(_05704_ ), .A2(_05479_ ), .A3(_06057_ ), .A4(_05706_ ), .ZN(_06608_ ) );
NAND2_X1 _14599_ ( .A1(_06607_ ), .A2(_06608_ ), .ZN(_06609_ ) );
AOI22_X1 _14600_ ( .A1(_06609_ ), .A2(\ID_EX_typ [2] ), .B1(_04396_ ), .B2(_05428_ ), .ZN(_06610_ ) );
OAI211_X1 _14601_ ( .A(_06610_ ), .B(_06364_ ), .C1(_05981_ ), .C2(\ID_EX_imm [22] ), .ZN(_06611_ ) );
NAND4_X1 _14602_ ( .A1(_06607_ ), .A2(_06404_ ), .A3(_06608_ ), .A4(_06353_ ), .ZN(_06612_ ) );
AND3_X1 _14603_ ( .A1(_04397_ ), .A2(_04417_ ), .A3(_06387_ ), .ZN(_06613_ ) );
AOI21_X1 _14604_ ( .A(_06613_ ), .B1(\ID_EX_pc [22] ), .B2(_06355_ ), .ZN(_06614_ ) );
OAI211_X1 _14605_ ( .A(_06611_ ), .B(_06612_ ), .C1(_06384_ ), .C2(_06614_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
AOI22_X1 _14606_ ( .A1(_06113_ ), .A2(\ID_EX_typ [2] ), .B1(_05428_ ), .B2(_05085_ ), .ZN(_06615_ ) );
OAI211_X1 _14607_ ( .A(_06615_ ), .B(_06364_ ), .C1(_05981_ ), .C2(\ID_EX_imm [31] ), .ZN(_06616_ ) );
OR2_X1 _14608_ ( .A1(_05984_ ), .A2(\EX_LS_result_csreg_mem [31] ), .ZN(_06617_ ) );
NAND4_X1 _14609_ ( .A1(_06617_ ), .A2(_06404_ ), .A3(_06112_ ), .A4(_06353_ ), .ZN(_06618_ ) );
AND3_X1 _14610_ ( .A1(_03494_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06619_ ) );
AOI21_X1 _14611_ ( .A(_06619_ ), .B1(_04559_ ), .B2(_06410_ ), .ZN(_06620_ ) );
OAI211_X1 _14612_ ( .A(_06616_ ), .B(_06618_ ), .C1(_06384_ ), .C2(_06620_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
NAND2_X1 _14613_ ( .A1(_06079_ ), .A2(_06441_ ), .ZN(_06621_ ) );
AND2_X1 _14614_ ( .A1(_05353_ ), .A2(_05369_ ), .ZN(_06622_ ) );
INV_X1 _14615_ ( .A(_06622_ ), .ZN(_06623_ ) );
NAND2_X1 _14616_ ( .A1(_06623_ ), .A2(_04395_ ), .ZN(_06624_ ) );
AND2_X1 _14617_ ( .A1(_06624_ ), .A2(_05383_ ), .ZN(_06625_ ) );
INV_X1 _14618_ ( .A(_04467_ ), .ZN(_06626_ ) );
OR2_X1 _14619_ ( .A1(_06625_ ), .A2(_06626_ ), .ZN(_06627_ ) );
AND2_X1 _14620_ ( .A1(_06627_ ), .A2(_05391_ ), .ZN(_06628_ ) );
XNOR2_X1 _14621_ ( .A(_06628_ ), .B(_04491_ ), .ZN(_06629_ ) );
AND3_X1 _14622_ ( .A1(_04253_ ), .A2(\ID_EX_typ [3] ), .A3(_05326_ ), .ZN(_06630_ ) );
AND2_X1 _14623_ ( .A1(_06630_ ), .A2(_05077_ ), .ZN(_06631_ ) );
BUF_X4 _14624_ ( .A(_06631_ ), .Z(_06632_ ) );
NAND2_X1 _14625_ ( .A1(_06629_ ), .A2(_06632_ ), .ZN(_06633_ ) );
NOR3_X1 _14626_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06634_ ) );
AND2_X2 _14627_ ( .A1(\ID_EX_typ [3] ), .A2(\ID_EX_typ [2] ), .ZN(_06635_ ) );
AND2_X2 _14628_ ( .A1(_06634_ ), .A2(_06635_ ), .ZN(_06636_ ) );
BUF_X4 _14629_ ( .A(_06636_ ), .Z(_06637_ ) );
NOR3_X1 _14630_ ( .A1(_05319_ ), .A2(\ID_EX_typ [0] ), .A3(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_06638_ ) );
AND2_X2 _14631_ ( .A1(_06638_ ), .A2(_06635_ ), .ZN(_06639_ ) );
BUF_X4 _14632_ ( .A(_06639_ ), .Z(_06640_ ) );
AOI22_X1 _14633_ ( .A1(_06086_ ), .A2(_06637_ ), .B1(\ID_EX_imm [21] ), .B2(_06640_ ), .ZN(_06641_ ) );
AND2_X1 _14634_ ( .A1(_06633_ ), .A2(_06641_ ), .ZN(_06642_ ) );
NOR2_X1 _14635_ ( .A1(_04017_ ), .A2(\ID_EX_typ [6] ), .ZN(_06643_ ) );
AND2_X1 _14636_ ( .A1(_06643_ ), .A2(_03495_ ), .ZN(_06644_ ) );
BUF_X4 _14637_ ( .A(_06644_ ), .Z(_06645_ ) );
INV_X2 _14638_ ( .A(_06645_ ), .ZN(_06646_ ) );
BUF_X4 _14639_ ( .A(_06646_ ), .Z(_06647_ ) );
OAI21_X1 _14640_ ( .A(_05605_ ), .B1(_06642_ ), .B2(_06647_ ), .ZN(_06648_ ) );
INV_X1 _14641_ ( .A(_05239_ ), .ZN(_06649_ ) );
AND2_X1 _14642_ ( .A1(_05137_ ), .A2(_05142_ ), .ZN(_06650_ ) );
INV_X1 _14643_ ( .A(_06650_ ), .ZN(_06651_ ) );
NOR2_X1 _14644_ ( .A1(_05151_ ), .A2(_04999_ ), .ZN(_06652_ ) );
INV_X1 _14645_ ( .A(_06652_ ), .ZN(_06653_ ) );
INV_X1 _14646_ ( .A(_05147_ ), .ZN(_06654_ ) );
NAND2_X4 _14647_ ( .A1(_05159_ ), .A2(_05160_ ), .ZN(_06655_ ) );
NOR2_X4 _14648_ ( .A1(_06655_ ), .A2(_05158_ ), .ZN(_06656_ ) );
AND3_X1 _14649_ ( .A1(_05153_ ), .A2(_02704_ ), .A3(_05154_ ), .ZN(_06657_ ) );
INV_X1 _14650_ ( .A(_06657_ ), .ZN(_06658_ ) );
NAND2_X1 _14651_ ( .A1(_05155_ ), .A2(_04976_ ), .ZN(_06659_ ) );
AND3_X1 _14652_ ( .A1(_06656_ ), .A2(_06658_ ), .A3(_06659_ ), .ZN(_06660_ ) );
NOR2_X2 _14653_ ( .A1(_06660_ ), .A2(_06657_ ), .ZN(_06661_ ) );
INV_X1 _14654_ ( .A(_05152_ ), .ZN(_06662_ ) );
OAI221_X2 _14655_ ( .A(_06653_ ), .B1(_02781_ ), .B2(_06654_ ), .C1(_06661_ ), .C2(_06662_ ), .ZN(_06663_ ) );
NOR2_X1 _14656_ ( .A1(_05147_ ), .A2(_02752_ ), .ZN(_06664_ ) );
INV_X1 _14657_ ( .A(_06664_ ), .ZN(_06665_ ) );
AND2_X1 _14658_ ( .A1(_05177_ ), .A2(_05182_ ), .ZN(_06666_ ) );
AND2_X1 _14659_ ( .A1(_05173_ ), .A2(_05187_ ), .ZN(_06667_ ) );
NAND4_X4 _14660_ ( .A1(_06663_ ), .A2(_06665_ ), .A3(_06666_ ), .A4(_06667_ ), .ZN(_06668_ ) );
NOR2_X1 _14661_ ( .A1(_05181_ ), .A2(_04883_ ), .ZN(_06669_ ) );
AND2_X1 _14662_ ( .A1(_05177_ ), .A2(_06669_ ), .ZN(_06670_ ) );
INV_X1 _14663_ ( .A(_05176_ ), .ZN(_06671_ ) );
AND3_X1 _14664_ ( .A1(_05172_ ), .A2(_05169_ ), .A3(_05170_ ), .ZN(_06672_ ) );
AND2_X1 _14665_ ( .A1(_05171_ ), .A2(_02598_ ), .ZN(_06673_ ) );
INV_X1 _14666_ ( .A(_06673_ ), .ZN(_06674_ ) );
NOR2_X1 _14667_ ( .A1(_05185_ ), .A2(_02623_ ), .ZN(_06675_ ) );
INV_X1 _14668_ ( .A(_06675_ ), .ZN(_06676_ ) );
AOI21_X1 _14669_ ( .A(_06672_ ), .B1(_06674_ ), .B2(_06676_ ), .ZN(_06677_ ) );
AOI221_X4 _14670_ ( .A(_06670_ ), .B1(_04906_ ), .B2(_06671_ ), .C1(_06666_ ), .C2(_06677_ ), .ZN(_06678_ ) );
AOI21_X2 _14671_ ( .A(_06651_ ), .B1(_06668_ ), .B2(_06678_ ), .ZN(_06679_ ) );
AND2_X1 _14672_ ( .A1(_05122_ ), .A2(_05117_ ), .ZN(_06680_ ) );
AND2_X1 _14673_ ( .A1(_05112_ ), .A2(_05108_ ), .ZN(_06681_ ) );
AND2_X1 _14674_ ( .A1(_06680_ ), .A2(_06681_ ), .ZN(_06682_ ) );
AND2_X1 _14675_ ( .A1(_05132_ ), .A2(_05128_ ), .ZN(_06683_ ) );
NAND3_X2 _14676_ ( .A1(_06679_ ), .A2(_06682_ ), .A3(_06683_ ), .ZN(_06684_ ) );
NOR2_X1 _14677_ ( .A1(_05136_ ), .A2(_04833_ ), .ZN(_06685_ ) );
AND2_X1 _14678_ ( .A1(_05136_ ), .A2(_04833_ ), .ZN(_06686_ ) );
INV_X1 _14679_ ( .A(_06686_ ), .ZN(_06687_ ) );
NOR2_X1 _14680_ ( .A1(_05141_ ), .A2(_04856_ ), .ZN(_06688_ ) );
AOI21_X1 _14681_ ( .A(_06685_ ), .B1(_06687_ ), .B2(_06688_ ), .ZN(_06689_ ) );
INV_X1 _14682_ ( .A(_06689_ ), .ZN(_06690_ ) );
NAND2_X1 _14683_ ( .A1(_06690_ ), .A2(_06683_ ), .ZN(_06691_ ) );
NOR2_X1 _14684_ ( .A1(_05131_ ), .A2(_04784_ ), .ZN(_06692_ ) );
INV_X1 _14685_ ( .A(_06692_ ), .ZN(_06693_ ) );
NAND3_X1 _14686_ ( .A1(_05132_ ), .A2(_02571_ ), .A3(_05208_ ), .ZN(_06694_ ) );
AND3_X1 _14687_ ( .A1(_06691_ ), .A2(_06693_ ), .A3(_06694_ ), .ZN(_06695_ ) );
INV_X1 _14688_ ( .A(_06682_ ), .ZN(_06696_ ) );
NOR2_X1 _14689_ ( .A1(_06695_ ), .A2(_06696_ ), .ZN(_06697_ ) );
NOR2_X1 _14690_ ( .A1(_05111_ ), .A2(_04678_ ), .ZN(_06698_ ) );
NOR2_X1 _14691_ ( .A1(_05116_ ), .A2(_04759_ ), .ZN(_06699_ ) );
NOR2_X1 _14692_ ( .A1(_05121_ ), .A2(_04734_ ), .ZN(_06700_ ) );
AOI21_X1 _14693_ ( .A(_06699_ ), .B1(_05117_ ), .B2(_06700_ ), .ZN(_06701_ ) );
INV_X1 _14694_ ( .A(_05112_ ), .ZN(_06702_ ) );
INV_X1 _14695_ ( .A(_05108_ ), .ZN(_06703_ ) );
NOR3_X1 _14696_ ( .A1(_06701_ ), .A2(_06702_ ), .A3(_06703_ ), .ZN(_06704_ ) );
NOR2_X1 _14697_ ( .A1(_05107_ ), .A2(_04708_ ), .ZN(_06705_ ) );
AND2_X1 _14698_ ( .A1(_05112_ ), .A2(_06705_ ), .ZN(_06706_ ) );
NOR4_X1 _14699_ ( .A1(_06697_ ), .A2(_06698_ ), .A3(_06704_ ), .A4(_06706_ ), .ZN(_06707_ ) );
AND2_X1 _14700_ ( .A1(_06684_ ), .A2(_06707_ ), .ZN(_06708_ ) );
INV_X1 _14701_ ( .A(_06708_ ), .ZN(_06709_ ) );
AND2_X1 _14702_ ( .A1(_05248_ ), .A2(_05253_ ), .ZN(_06710_ ) );
AND2_X1 _14703_ ( .A1(_05225_ ), .A2(_05220_ ), .ZN(_06711_ ) );
NAND3_X1 _14704_ ( .A1(_06709_ ), .A2(_06710_ ), .A3(_06711_ ), .ZN(_06712_ ) );
NOR2_X1 _14705_ ( .A1(_05224_ ), .A2(_04342_ ), .ZN(_06713_ ) );
AOI21_X1 _14706_ ( .A(_05259_ ), .B1(_05220_ ), .B2(_06713_ ), .ZN(_06714_ ) );
NOR3_X1 _14707_ ( .A1(_06714_ ), .A2(_05249_ ), .A3(_05254_ ), .ZN(_06715_ ) );
NOR2_X1 _14708_ ( .A1(_05252_ ), .A2(_04256_ ), .ZN(_06716_ ) );
INV_X1 _14709_ ( .A(_02917_ ), .ZN(_06717_ ) );
NOR2_X1 _14710_ ( .A1(_05247_ ), .A2(_06717_ ), .ZN(_06718_ ) );
AND2_X1 _14711_ ( .A1(_05253_ ), .A2(_06718_ ), .ZN(_06719_ ) );
NOR3_X1 _14712_ ( .A1(_06715_ ), .A2(_06716_ ), .A3(_06719_ ), .ZN(_06720_ ) );
AOI21_X1 _14713_ ( .A(_06649_ ), .B1(_06712_ ), .B2(_06720_ ), .ZN(_06721_ ) );
NOR2_X1 _14714_ ( .A1(_05238_ ), .A2(_04444_ ), .ZN(_06722_ ) );
NOR3_X1 _14715_ ( .A1(_06721_ ), .A2(_05243_ ), .A3(_06722_ ), .ZN(_06723_ ) );
NOR2_X1 _14716_ ( .A1(\ID_EX_typ [2] ), .A2(\ID_EX_typ [1] ), .ZN(_06724_ ) );
INV_X1 _14717_ ( .A(_06724_ ), .ZN(_06725_ ) );
NOR2_X1 _14718_ ( .A1(_05073_ ), .A2(_06725_ ), .ZN(_06726_ ) );
INV_X1 _14719_ ( .A(_06726_ ), .ZN(_06727_ ) );
NOR2_X1 _14720_ ( .A1(_06723_ ), .A2(_06727_ ), .ZN(_06728_ ) );
OAI21_X1 _14721_ ( .A(_05243_ ), .B1(_06721_ ), .B2(_06722_ ), .ZN(_06729_ ) );
NAND2_X1 _14722_ ( .A1(_06728_ ), .A2(_06729_ ), .ZN(_06730_ ) );
AND2_X1 _14723_ ( .A1(_05329_ ), .A2(\ID_EX_typ [2] ), .ZN(_06731_ ) );
BUF_X4 _14724_ ( .A(_06731_ ), .Z(_06732_ ) );
OR2_X1 _14725_ ( .A1(_05238_ ), .A2(_05252_ ), .ZN(_06733_ ) );
NOR3_X1 _14726_ ( .A1(_06733_ ), .A2(_05242_ ), .A3(_05247_ ), .ZN(_06734_ ) );
AOI22_X1 _14727_ ( .A1(_05223_ ), .A2(_05222_ ), .B1(_05109_ ), .B2(_05110_ ), .ZN(_06735_ ) );
NAND4_X1 _14728_ ( .A1(_06734_ ), .A2(_05200_ ), .A3(_05261_ ), .A4(_06735_ ), .ZN(_06736_ ) );
NAND2_X1 _14729_ ( .A1(_05202_ ), .A2(_06671_ ), .ZN(_06737_ ) );
OR3_X1 _14730_ ( .A1(_06737_ ), .A2(_05136_ ), .A3(_05181_ ), .ZN(_06738_ ) );
NOR4_X1 _14731_ ( .A1(_06736_ ), .A2(_06738_ ), .A3(_05116_ ), .A4(_05127_ ), .ZN(_06739_ ) );
NAND4_X1 _14732_ ( .A1(_06739_ ), .A2(_05119_ ), .A3(_05120_ ), .A4(_05206_ ), .ZN(_06740_ ) );
INV_X1 _14733_ ( .A(_05171_ ), .ZN(_06741_ ) );
AND2_X1 _14734_ ( .A1(_06655_ ), .A2(_05156_ ), .ZN(_06742_ ) );
AND2_X1 _14735_ ( .A1(_06742_ ), .A2(_05151_ ), .ZN(_06743_ ) );
BUF_X2 _14736_ ( .A(_06654_ ), .Z(_06744_ ) );
AND2_X1 _14737_ ( .A1(_06743_ ), .A2(_06744_ ), .ZN(_06745_ ) );
AND2_X2 _14738_ ( .A1(_06745_ ), .A2(_05186_ ), .ZN(_06746_ ) );
NOR3_X1 _14739_ ( .A1(_06740_ ), .A2(_06741_ ), .A3(_06746_ ), .ZN(_06747_ ) );
AND2_X1 _14740_ ( .A1(_05136_ ), .A2(_05141_ ), .ZN(_06748_ ) );
AND3_X1 _14741_ ( .A1(_06748_ ), .A2(_05131_ ), .A3(_05127_ ), .ZN(_06749_ ) );
AND2_X1 _14742_ ( .A1(_05121_ ), .A2(_05116_ ), .ZN(_06750_ ) );
AND4_X1 _14743_ ( .A1(_05111_ ), .A2(_06749_ ), .A3(_05107_ ), .A4(_06750_ ), .ZN(_06751_ ) );
AND4_X1 _14744_ ( .A1(_05176_ ), .A2(_05171_ ), .A3(_05181_ ), .A4(_05186_ ), .ZN(_06752_ ) );
BUF_X2 _14745_ ( .A(_05151_ ), .Z(_06753_ ) );
NAND4_X1 _14746_ ( .A1(_06752_ ), .A2(_06744_ ), .A3(_06753_ ), .A4(_06742_ ), .ZN(_06754_ ) );
NAND4_X1 _14747_ ( .A1(_05169_ ), .A2(_05176_ ), .A3(_05181_ ), .A4(_05170_ ), .ZN(_06755_ ) );
NAND2_X1 _14748_ ( .A1(_06754_ ), .A2(_06755_ ), .ZN(_06756_ ) );
AND2_X1 _14749_ ( .A1(_05224_ ), .A2(_05219_ ), .ZN(_06757_ ) );
AND2_X1 _14750_ ( .A1(_05247_ ), .A2(_05252_ ), .ZN(_06758_ ) );
AND2_X1 _14751_ ( .A1(_05242_ ), .A2(_05238_ ), .ZN(_06759_ ) );
AND3_X1 _14752_ ( .A1(_06757_ ), .A2(_06758_ ), .A3(_06759_ ), .ZN(_06760_ ) );
AND3_X1 _14753_ ( .A1(_06751_ ), .A2(_06756_ ), .A3(_06760_ ), .ZN(_06761_ ) );
OAI21_X1 _14754_ ( .A(_03150_ ), .B1(_06747_ ), .B2(_06761_ ), .ZN(_06762_ ) );
INV_X1 _14755_ ( .A(_06761_ ), .ZN(_06763_ ) );
OR3_X1 _14756_ ( .A1(_06763_ ), .A2(_05272_ ), .A3(_05233_ ), .ZN(_06764_ ) );
NAND3_X1 _14757_ ( .A1(_06763_ ), .A2(_05272_ ), .A3(_05233_ ), .ZN(_06765_ ) );
AOI21_X1 _14758_ ( .A(_06762_ ), .B1(_06764_ ), .B2(_06765_ ), .ZN(_06766_ ) );
AND4_X1 _14759_ ( .A1(_05111_ ), .A2(_05107_ ), .A3(_05131_ ), .A4(_05127_ ), .ZN(_06767_ ) );
NAND4_X1 _14760_ ( .A1(_06767_ ), .A2(_05176_ ), .A3(_05181_ ), .A4(_06748_ ), .ZN(_06768_ ) );
NAND4_X1 _14761_ ( .A1(_06750_ ), .A2(_06757_ ), .A3(_06758_ ), .A4(_06759_ ), .ZN(_06769_ ) );
NOR2_X1 _14762_ ( .A1(_06768_ ), .A2(_06769_ ), .ZN(_06770_ ) );
OAI21_X1 _14763_ ( .A(_06770_ ), .B1(_06746_ ), .B2(_06741_ ), .ZN(_06771_ ) );
NOR3_X1 _14764_ ( .A1(_06771_ ), .A2(_05272_ ), .A3(_05233_ ), .ZN(_06772_ ) );
NOR4_X1 _14765_ ( .A1(_05093_ ), .A2(_05313_ ), .A3(_05099_ ), .A4(_05080_ ), .ZN(_06773_ ) );
INV_X1 _14766_ ( .A(_05297_ ), .ZN(_06774_ ) );
AOI21_X1 _14767_ ( .A(_06774_ ), .B1(_05288_ ), .B2(_05289_ ), .ZN(_06775_ ) );
AND4_X1 _14768_ ( .A1(_05277_ ), .A2(_06773_ ), .A3(_05281_ ), .A4(_06775_ ), .ZN(_06776_ ) );
NAND2_X1 _14769_ ( .A1(_06772_ ), .A2(_06776_ ), .ZN(_06777_ ) );
NOR4_X1 _14770_ ( .A1(_05290_ ), .A2(_05277_ ), .A3(_05281_ ), .A4(_05297_ ), .ZN(_06778_ ) );
AND4_X1 _14771_ ( .A1(_05093_ ), .A2(_05313_ ), .A3(_05099_ ), .A4(_05080_ ), .ZN(_06779_ ) );
NAND2_X1 _14772_ ( .A1(_06778_ ), .A2(_06779_ ), .ZN(_06780_ ) );
OAI21_X1 _14773_ ( .A(_06777_ ), .B1(_06772_ ), .B2(_06780_ ), .ZN(_06781_ ) );
AND2_X2 _14774_ ( .A1(_06766_ ), .A2(_06781_ ), .ZN(_06782_ ) );
XNOR2_X1 _14775_ ( .A(_06746_ ), .B(_05171_ ), .ZN(_06783_ ) );
NAND2_X1 _14776_ ( .A1(_06782_ ), .A2(_06783_ ), .ZN(_06784_ ) );
XNOR2_X1 _14777_ ( .A(_06745_ ), .B(_05186_ ), .ZN(_06785_ ) );
NOR2_X1 _14778_ ( .A1(_06785_ ), .A2(_05171_ ), .ZN(_06786_ ) );
INV_X1 _14779_ ( .A(_06786_ ), .ZN(_06787_ ) );
INV_X1 _14780_ ( .A(_06785_ ), .ZN(_06788_ ) );
BUF_X2 _14781_ ( .A(_06781_ ), .Z(_06789_ ) );
NAND4_X1 _14782_ ( .A1(_05200_ ), .A2(_05208_ ), .A3(_05214_ ), .A4(_05206_ ), .ZN(_06790_ ) );
NOR4_X1 _14783_ ( .A1(_06790_ ), .A2(_06737_ ), .A3(_05136_ ), .A4(_05181_ ), .ZN(_06791_ ) );
NOR4_X1 _14784_ ( .A1(_05121_ ), .A2(_05224_ ), .A3(_05116_ ), .A4(_05219_ ), .ZN(_06792_ ) );
AND3_X1 _14785_ ( .A1(_06791_ ), .A2(_06734_ ), .A3(_06792_ ), .ZN(_06793_ ) );
INV_X1 _14786_ ( .A(_06745_ ), .ZN(_06794_ ) );
OAI211_X1 _14787_ ( .A(_05171_ ), .B(_06793_ ), .C1(_06794_ ), .C2(_05192_ ), .ZN(_06795_ ) );
NAND2_X1 _14788_ ( .A1(_06771_ ), .A2(_06795_ ), .ZN(_06796_ ) );
NAND2_X1 _14789_ ( .A1(_06796_ ), .A2(_03150_ ), .ZN(_06797_ ) );
AOI21_X1 _14790_ ( .A(_06797_ ), .B1(_06764_ ), .B2(_06765_ ), .ZN(_06798_ ) );
BUF_X4 _14791_ ( .A(_06655_ ), .Z(_06799_ ) );
BUF_X2 _14792_ ( .A(_05156_ ), .Z(_06800_ ) );
BUF_X2 _14793_ ( .A(_06800_ ), .Z(_06801_ ) );
XNOR2_X1 _14794_ ( .A(_06799_ ), .B(_06801_ ), .ZN(_06802_ ) );
BUF_X2 _14795_ ( .A(_05166_ ), .Z(_06803_ ) );
BUF_X2 _14796_ ( .A(_06803_ ), .Z(_06804_ ) );
BUF_X2 _14797_ ( .A(_06804_ ), .Z(_06805_ ) );
OR2_X1 _14798_ ( .A1(_06802_ ), .A2(_06805_ ), .ZN(_06806_ ) );
XNOR2_X1 _14799_ ( .A(_06743_ ), .B(_05147_ ), .ZN(_06807_ ) );
INV_X1 _14800_ ( .A(_06807_ ), .ZN(_06808_ ) );
NAND4_X1 _14801_ ( .A1(_06789_ ), .A2(_06798_ ), .A3(_06806_ ), .A4(_06808_ ), .ZN(_06809_ ) );
AOI22_X1 _14802_ ( .A1(_06784_ ), .A2(_06787_ ), .B1(_06788_ ), .B2(_06809_ ), .ZN(_06810_ ) );
BUF_X4 _14803_ ( .A(_06803_ ), .Z(_06811_ ) );
BUF_X2 _14804_ ( .A(_05159_ ), .Z(_06812_ ) );
BUF_X2 _14805_ ( .A(_06812_ ), .Z(_06813_ ) );
BUF_X2 _14806_ ( .A(_05160_ ), .Z(_06814_ ) );
BUF_X2 _14807_ ( .A(_06814_ ), .Z(_06815_ ) );
AND3_X1 _14808_ ( .A1(_06813_ ), .A2(_05282_ ), .A3(_06815_ ), .ZN(_06816_ ) );
AOI21_X1 _14809_ ( .A(_03039_ ), .B1(_06813_ ), .B2(_06815_ ), .ZN(_06817_ ) );
INV_X1 _14810_ ( .A(_05156_ ), .ZN(_06818_ ) );
BUF_X2 _14811_ ( .A(_06818_ ), .Z(_06819_ ) );
BUF_X4 _14812_ ( .A(_06819_ ), .Z(_06820_ ) );
NOR3_X1 _14813_ ( .A1(_06816_ ), .A2(_06817_ ), .A3(_06820_ ), .ZN(_06821_ ) );
BUF_X2 _14814_ ( .A(_05159_ ), .Z(_06822_ ) );
BUF_X2 _14815_ ( .A(_05160_ ), .Z(_06823_ ) );
AND3_X1 _14816_ ( .A1(_06822_ ), .A2(_05100_ ), .A3(_06823_ ), .ZN(_06824_ ) );
AOI21_X1 _14817_ ( .A(_02348_ ), .B1(_06822_ ), .B2(_06823_ ), .ZN(_06825_ ) );
BUF_X2 _14818_ ( .A(_05156_ ), .Z(_06826_ ) );
BUF_X2 _14819_ ( .A(_06826_ ), .Z(_06827_ ) );
NOR3_X1 _14820_ ( .A1(_06824_ ), .A2(_06825_ ), .A3(_06827_ ), .ZN(_06828_ ) );
OAI21_X1 _14821_ ( .A(_06811_ ), .B1(_06821_ ), .B2(_06828_ ), .ZN(_06829_ ) );
BUF_X4 _14822_ ( .A(_06818_ ), .Z(_06830_ ) );
BUF_X4 _14823_ ( .A(_06830_ ), .Z(_06831_ ) );
AND3_X1 _14824_ ( .A1(_05291_ ), .A2(_06813_ ), .A3(_06815_ ), .ZN(_06832_ ) );
AOI21_X1 _14825_ ( .A(_02396_ ), .B1(_06813_ ), .B2(_06815_ ), .ZN(_06833_ ) );
OAI21_X1 _14826_ ( .A(_06831_ ), .B1(_06832_ ), .B2(_06833_ ), .ZN(_06834_ ) );
CLKBUF_X2 _14827_ ( .A(_05159_ ), .Z(_06835_ ) );
CLKBUF_X2 _14828_ ( .A(_05160_ ), .Z(_06836_ ) );
AND3_X1 _14829_ ( .A1(_06835_ ), .A2(_04396_ ), .A3(_06836_ ), .ZN(_06837_ ) );
AOI21_X1 _14830_ ( .A(_04468_ ), .B1(_06813_ ), .B2(_06815_ ), .ZN(_06838_ ) );
OAI21_X1 _14831_ ( .A(_06801_ ), .B1(_06837_ ), .B2(_06838_ ), .ZN(_06839_ ) );
BUF_X2 _14832_ ( .A(_06753_ ), .Z(_06840_ ) );
BUF_X2 _14833_ ( .A(_06840_ ), .Z(_06841_ ) );
NAND3_X1 _14834_ ( .A1(_06834_ ), .A2(_06839_ ), .A3(_06841_ ), .ZN(_06842_ ) );
NAND2_X1 _14835_ ( .A1(_06829_ ), .A2(_06842_ ), .ZN(_06843_ ) );
NAND2_X1 _14836_ ( .A1(_06655_ ), .A2(_05094_ ), .ZN(_06844_ ) );
NAND3_X1 _14837_ ( .A1(_06835_ ), .A2(_02297_ ), .A3(_06836_ ), .ZN(_06845_ ) );
AND3_X1 _14838_ ( .A1(_06844_ ), .A2(_06800_ ), .A3(_06845_ ), .ZN(_06846_ ) );
AND2_X1 _14839_ ( .A1(_06799_ ), .A2(_03150_ ), .ZN(_06847_ ) );
AOI21_X1 _14840_ ( .A(_06846_ ), .B1(_06831_ ), .B2(_06847_ ), .ZN(_06848_ ) );
NOR2_X1 _14841_ ( .A1(_06848_ ), .A2(_06805_ ), .ZN(_06849_ ) );
BUF_X4 _14842_ ( .A(_05147_ ), .Z(_06850_ ) );
BUF_X4 _14843_ ( .A(_06850_ ), .Z(_06851_ ) );
MUX2_X1 _14844_ ( .A(_06843_ ), .B(_06849_ ), .S(_06851_ ), .Z(_06852_ ) );
BUF_X2 _14845_ ( .A(_05186_ ), .Z(_06853_ ) );
BUF_X2 _14846_ ( .A(_06853_ ), .Z(_06854_ ) );
AND2_X1 _14847_ ( .A1(_06852_ ), .A2(_06854_ ), .ZN(_06855_ ) );
OAI21_X1 _14848_ ( .A(_06732_ ), .B1(_06810_ ), .B2(_06855_ ), .ZN(_06856_ ) );
BUF_X2 _14849_ ( .A(_05186_ ), .Z(_06857_ ) );
BUF_X2 _14850_ ( .A(_06857_ ), .Z(_06858_ ) );
CLKBUF_X2 _14851_ ( .A(_06822_ ), .Z(_06859_ ) );
BUF_X2 _14852_ ( .A(_06836_ ), .Z(_06860_ ) );
AND3_X1 _14853_ ( .A1(_04856_ ), .A2(_06859_ ), .A3(_06860_ ), .ZN(_06861_ ) );
BUF_X2 _14854_ ( .A(_06835_ ), .Z(_06862_ ) );
AOI21_X1 _14855_ ( .A(_04832_ ), .B1(_06862_ ), .B2(_06860_ ), .ZN(_06863_ ) );
BUF_X2 _14856_ ( .A(_06820_ ), .Z(_06864_ ) );
NOR3_X1 _14857_ ( .A1(_06861_ ), .A2(_06863_ ), .A3(_06864_ ), .ZN(_06865_ ) );
AND3_X1 _14858_ ( .A1(_06813_ ), .A2(_04883_ ), .A3(_06815_ ), .ZN(_06866_ ) );
BUF_X2 _14859_ ( .A(_06823_ ), .Z(_06867_ ) );
AOI21_X1 _14860_ ( .A(_04906_ ), .B1(_06859_ ), .B2(_06867_ ), .ZN(_06868_ ) );
BUF_X2 _14861_ ( .A(_06827_ ), .Z(_06869_ ) );
NOR3_X1 _14862_ ( .A1(_06866_ ), .A2(_06868_ ), .A3(_06869_ ), .ZN(_06870_ ) );
NOR2_X1 _14863_ ( .A1(_06865_ ), .A2(_06870_ ), .ZN(_06871_ ) );
BUF_X2 _14864_ ( .A(_06841_ ), .Z(_06872_ ) );
NOR2_X1 _14865_ ( .A1(_06871_ ), .A2(_06872_ ), .ZN(_06873_ ) );
BUF_X4 _14866_ ( .A(_06744_ ), .Z(_06874_ ) );
BUF_X2 _14867_ ( .A(_06874_ ), .Z(_06875_ ) );
BUF_X4 _14868_ ( .A(_06811_ ), .Z(_06876_ ) );
AND3_X1 _14869_ ( .A1(_04734_ ), .A2(_06859_ ), .A3(_06867_ ), .ZN(_06877_ ) );
AOI21_X1 _14870_ ( .A(_04758_ ), .B1(_06862_ ), .B2(_06860_ ), .ZN(_06878_ ) );
OR3_X1 _14871_ ( .A1(_06877_ ), .A2(_06878_ ), .A3(_06864_ ), .ZN(_06879_ ) );
AOI21_X1 _14872_ ( .A(_04783_ ), .B1(_06862_ ), .B2(_06860_ ), .ZN(_06880_ ) );
INV_X1 _14873_ ( .A(_06880_ ), .ZN(_06881_ ) );
BUF_X4 _14874_ ( .A(_06831_ ), .Z(_06882_ ) );
OAI211_X1 _14875_ ( .A(_06881_ ), .B(_06882_ ), .C1(_02571_ ), .C2(_06799_ ), .ZN(_06883_ ) );
AOI21_X1 _14876_ ( .A(_06876_ ), .B1(_06879_ ), .B2(_06883_ ), .ZN(_06884_ ) );
NOR3_X1 _14877_ ( .A1(_06873_ ), .A2(_06875_ ), .A3(_06884_ ), .ZN(_06885_ ) );
BUF_X4 _14878_ ( .A(_06753_ ), .Z(_06886_ ) );
BUF_X4 _14879_ ( .A(_06886_ ), .Z(_06887_ ) );
AND3_X1 _14880_ ( .A1(_04342_ ), .A2(_06862_ ), .A3(_06860_ ), .ZN(_06888_ ) );
AOI21_X1 _14881_ ( .A(_02965_ ), .B1(_06862_ ), .B2(_06860_ ), .ZN(_06889_ ) );
OR3_X1 _14882_ ( .A1(_06888_ ), .A2(_06864_ ), .A3(_06889_ ), .ZN(_06890_ ) );
AND3_X1 _14883_ ( .A1(_04708_ ), .A2(_06859_ ), .A3(_06867_ ), .ZN(_06891_ ) );
AOI21_X1 _14884_ ( .A(_02815_ ), .B1(_06862_ ), .B2(_06860_ ), .ZN(_06892_ ) );
OR3_X1 _14885_ ( .A1(_06891_ ), .A2(_06892_ ), .A3(_06869_ ), .ZN(_06893_ ) );
AOI21_X1 _14886_ ( .A(_06887_ ), .B1(_06890_ ), .B2(_06893_ ), .ZN(_06894_ ) );
BUF_X2 _14887_ ( .A(_06801_ ), .Z(_06895_ ) );
AND3_X1 _14888_ ( .A1(_04444_ ), .A2(_06835_ ), .A3(_06836_ ), .ZN(_06896_ ) );
OAI21_X1 _14889_ ( .A(_06895_ ), .B1(_06896_ ), .B2(_06838_ ), .ZN(_06897_ ) );
AND3_X1 _14890_ ( .A1(_06859_ ), .A2(_06717_ ), .A3(_06867_ ), .ZN(_06898_ ) );
AOI21_X1 _14891_ ( .A(_02940_ ), .B1(_06813_ ), .B2(_06815_ ), .ZN(_06899_ ) );
OAI21_X1 _14892_ ( .A(_06864_ ), .B1(_06898_ ), .B2(_06899_ ), .ZN(_06900_ ) );
AND3_X1 _14893_ ( .A1(_06897_ ), .A2(_06900_ ), .A3(_06887_ ), .ZN(_06901_ ) );
BUF_X4 _14894_ ( .A(_06851_ ), .Z(_06902_ ) );
NOR3_X1 _14895_ ( .A1(_06894_ ), .A2(_06901_ ), .A3(_06902_ ), .ZN(_06903_ ) );
OAI21_X1 _14896_ ( .A(_06858_ ), .B1(_06885_ ), .B2(_06903_ ), .ZN(_06904_ ) );
BUF_X2 _14897_ ( .A(_05192_ ), .Z(_06905_ ) );
BUF_X2 _14898_ ( .A(_06905_ ), .Z(_06906_ ) );
AND3_X1 _14899_ ( .A1(_02623_ ), .A2(_06859_ ), .A3(_06867_ ), .ZN(_06907_ ) );
AOI21_X1 _14900_ ( .A(_02598_ ), .B1(_06859_ ), .B2(_06867_ ), .ZN(_06908_ ) );
OR3_X1 _14901_ ( .A1(_06907_ ), .A2(_06830_ ), .A3(_06908_ ), .ZN(_06909_ ) );
AND3_X1 _14902_ ( .A1(_06859_ ), .A2(_04999_ ), .A3(_06867_ ), .ZN(_06910_ ) );
AOI21_X1 _14903_ ( .A(_02752_ ), .B1(_06862_ ), .B2(_06867_ ), .ZN(_06911_ ) );
OR3_X1 _14904_ ( .A1(_06910_ ), .A2(_06911_ ), .A3(_06827_ ), .ZN(_06912_ ) );
NAND3_X1 _14905_ ( .A1(_06909_ ), .A2(_06912_ ), .A3(_06841_ ), .ZN(_06913_ ) );
BUF_X2 _14906_ ( .A(_06886_ ), .Z(_06914_ ) );
AOI21_X1 _14907_ ( .A(_02704_ ), .B1(_06859_ ), .B2(_06867_ ), .ZN(_06915_ ) );
NOR3_X1 _14908_ ( .A1(_05161_ ), .A2(_06915_ ), .A3(_06831_ ), .ZN(_06916_ ) );
OAI21_X1 _14909_ ( .A(_06913_ ), .B1(_06914_ ), .B2(_06916_ ), .ZN(_06917_ ) );
BUF_X4 _14910_ ( .A(_06850_ ), .Z(_06918_ ) );
BUF_X4 _14911_ ( .A(_06918_ ), .Z(_06919_ ) );
OAI21_X1 _14912_ ( .A(_06906_ ), .B1(_06917_ ), .B2(_06919_ ), .ZN(_06920_ ) );
NAND3_X1 _14913_ ( .A1(_06904_ ), .A2(_05332_ ), .A3(_06920_ ), .ZN(_06921_ ) );
BUF_X2 _14914_ ( .A(_05330_ ), .Z(_06922_ ) );
NOR2_X1 _14915_ ( .A1(_05242_ ), .A2(_04469_ ), .ZN(_06923_ ) );
AOI22_X1 _14916_ ( .A1(_05243_ ), .A2(_06922_ ), .B1(_05073_ ), .B2(_06923_ ), .ZN(_06924_ ) );
NAND4_X1 _14917_ ( .A1(_06730_ ), .A2(_06856_ ), .A3(_06921_ ), .A4(_06924_ ), .ZN(_06925_ ) );
BUF_X2 _14918_ ( .A(_06854_ ), .Z(_06926_ ) );
AND2_X1 _14919_ ( .A1(_05320_ ), .A2(\ID_EX_typ [2] ), .ZN(_06927_ ) );
BUF_X2 _14920_ ( .A(_06927_ ), .Z(_06928_ ) );
AND3_X1 _14921_ ( .A1(_06852_ ), .A2(_06926_ ), .A3(_06928_ ), .ZN(_06929_ ) );
BUF_X4 _14922_ ( .A(_05324_ ), .Z(_06930_ ) );
AOI21_X1 _14923_ ( .A(_06930_ ), .B1(_05242_ ), .B2(_04469_ ), .ZN(_06931_ ) );
OR3_X1 _14924_ ( .A1(_06925_ ), .A2(_06929_ ), .A3(_06931_ ), .ZN(_06932_ ) );
INV_X1 _14925_ ( .A(_06631_ ), .ZN(_06933_ ) );
OAI21_X1 _14926_ ( .A(_06635_ ), .B1(_06638_ ), .B2(_06634_ ), .ZN(_06934_ ) );
NAND2_X1 _14927_ ( .A1(_06933_ ), .A2(_06934_ ), .ZN(_06935_ ) );
AND4_X1 _14928_ ( .A1(\ID_EX_typ [3] ), .A2(_05326_ ), .A3(_05319_ ), .A4(\ID_EX_typ [0] ), .ZN(_06936_ ) );
MUX2_X1 _14929_ ( .A(_06936_ ), .B(_06630_ ), .S(\ID_EX_typ [4] ), .Z(_06937_ ) );
NOR2_X1 _14930_ ( .A1(_06935_ ), .A2(_06937_ ), .ZN(_06938_ ) );
NOR2_X2 _14931_ ( .A1(_06938_ ), .A2(_06646_ ), .ZN(_06939_ ) );
INV_X1 _14932_ ( .A(_06939_ ), .ZN(_06940_ ) );
BUF_X4 _14933_ ( .A(_06940_ ), .Z(_06941_ ) );
BUF_X4 _14934_ ( .A(_06941_ ), .Z(_06942_ ) );
AOI21_X1 _14935_ ( .A(_06648_ ), .B1(_06932_ ), .B2(_06942_ ), .ZN(_06943_ ) );
OAI21_X1 _14936_ ( .A(_06522_ ), .B1(_06083_ ), .B2(_06056_ ), .ZN(_06944_ ) );
OAI21_X1 _14937_ ( .A(_06621_ ), .B1(_06943_ ), .B2(_06944_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
NAND2_X1 _14938_ ( .A1(_05510_ ), .A2(_06441_ ), .ZN(_06945_ ) );
BUF_X4 _14939_ ( .A(_06646_ ), .Z(_06946_ ) );
NAND3_X1 _14940_ ( .A1(_06624_ ), .A2(_06626_ ), .A3(_05383_ ), .ZN(_06947_ ) );
NAND3_X1 _14941_ ( .A1(_06627_ ), .A2(_06632_ ), .A3(_06947_ ), .ZN(_06948_ ) );
BUF_X2 _14942_ ( .A(_06636_ ), .Z(_06949_ ) );
BUF_X4 _14943_ ( .A(_06639_ ), .Z(_06950_ ) );
AOI22_X1 _14944_ ( .A1(_05515_ ), .A2(_06949_ ), .B1(\ID_EX_imm [20] ), .B2(_06950_ ), .ZN(_06951_ ) );
AOI21_X1 _14945_ ( .A(_06946_ ), .B1(_06948_ ), .B2(_06951_ ), .ZN(_06952_ ) );
OR2_X1 _14946_ ( .A1(_06952_ ), .A2(_05433_ ), .ZN(_06953_ ) );
BUF_X4 _14947_ ( .A(_06727_ ), .Z(_06954_ ) );
NOR2_X1 _14948_ ( .A1(_06721_ ), .A2(_06954_ ), .ZN(_06955_ ) );
AND2_X1 _14949_ ( .A1(_06712_ ), .A2(_06720_ ), .ZN(_06956_ ) );
INV_X2 _14950_ ( .A(_06956_ ), .ZN(_06957_ ) );
OAI21_X1 _14951_ ( .A(_06955_ ), .B1(_05239_ ), .B2(_06957_ ), .ZN(_06958_ ) );
BUF_X4 _14952_ ( .A(_06732_ ), .Z(_06959_ ) );
AND2_X1 _14953_ ( .A1(_06781_ ), .A2(_06798_ ), .ZN(_06960_ ) );
BUF_X2 _14954_ ( .A(_06960_ ), .Z(_06961_ ) );
BUF_X2 _14955_ ( .A(_06808_ ), .Z(_06962_ ) );
INV_X1 _14956_ ( .A(_06655_ ), .ZN(_06963_ ) );
OAI21_X1 _14957_ ( .A(_06887_ ), .B1(_06963_ ), .B2(_06882_ ), .ZN(_06964_ ) );
NAND3_X1 _14958_ ( .A1(_06961_ ), .A2(_06962_ ), .A3(_06964_ ), .ZN(_06965_ ) );
AOI22_X1 _14959_ ( .A1(_06784_ ), .A2(_06787_ ), .B1(_06965_ ), .B2(_06788_ ), .ZN(_06966_ ) );
AOI21_X1 _14960_ ( .A(_03063_ ), .B1(_05159_ ), .B2(_05160_ ), .ZN(_06967_ ) );
INV_X1 _14961_ ( .A(_06967_ ), .ZN(_06968_ ) );
NAND3_X1 _14962_ ( .A1(_06822_ ), .A2(_05307_ ), .A3(_06823_ ), .ZN(_06969_ ) );
AND3_X1 _14963_ ( .A1(_06968_ ), .A2(_06819_ ), .A3(_06969_ ), .ZN(_06970_ ) );
AND3_X1 _14964_ ( .A1(_03040_ ), .A2(_06812_ ), .A3(_06814_ ), .ZN(_06971_ ) );
AOI21_X1 _14965_ ( .A(_03196_ ), .B1(_06822_ ), .B2(_06823_ ), .ZN(_06972_ ) );
NOR3_X1 _14966_ ( .A1(_06971_ ), .A2(_06972_ ), .A3(_06819_ ), .ZN(_06973_ ) );
NOR3_X1 _14967_ ( .A1(_06970_ ), .A2(_06973_ ), .A3(_06753_ ), .ZN(_06974_ ) );
AND3_X1 _14968_ ( .A1(_04469_ ), .A2(_06835_ ), .A3(_06836_ ), .ZN(_06975_ ) );
AOI21_X1 _14969_ ( .A(_02422_ ), .B1(_06813_ ), .B2(_06815_ ), .ZN(_06976_ ) );
OAI21_X1 _14970_ ( .A(_06800_ ), .B1(_06975_ ), .B2(_06976_ ), .ZN(_06977_ ) );
AND3_X1 _14971_ ( .A1(_04420_ ), .A2(_06822_ ), .A3(_06823_ ), .ZN(_06978_ ) );
AOI21_X1 _14972_ ( .A(_02373_ ), .B1(_06822_ ), .B2(_06823_ ), .ZN(_06979_ ) );
OAI21_X1 _14973_ ( .A(_06830_ ), .B1(_06978_ ), .B2(_06979_ ), .ZN(_06980_ ) );
AOI21_X1 _14974_ ( .A(_06803_ ), .B1(_06977_ ), .B2(_06980_ ), .ZN(_06981_ ) );
NOR2_X1 _14975_ ( .A1(_06974_ ), .A2(_06981_ ), .ZN(_06982_ ) );
INV_X1 _14976_ ( .A(_02297_ ), .ZN(_06983_ ) );
AOI21_X1 _14977_ ( .A(_06983_ ), .B1(_06835_ ), .B2(_06836_ ), .ZN(_06984_ ) );
AOI21_X1 _14978_ ( .A(_06984_ ), .B1(_05085_ ), .B2(_06963_ ), .ZN(_06985_ ) );
NAND2_X1 _14979_ ( .A1(_06985_ ), .A2(_06819_ ), .ZN(_06986_ ) );
NAND2_X1 _14980_ ( .A1(_06655_ ), .A2(_05100_ ), .ZN(_06987_ ) );
NAND3_X1 _14981_ ( .A1(_06812_ ), .A2(_05094_ ), .A3(_06814_ ), .ZN(_06988_ ) );
NAND2_X1 _14982_ ( .A1(_06987_ ), .A2(_06988_ ), .ZN(_06989_ ) );
OAI21_X1 _14983_ ( .A(_06986_ ), .B1(_06830_ ), .B2(_06989_ ), .ZN(_06990_ ) );
AND2_X1 _14984_ ( .A1(_06990_ ), .A2(_06840_ ), .ZN(_06991_ ) );
MUX2_X1 _14985_ ( .A(_06982_ ), .B(_06991_ ), .S(_06850_ ), .Z(_06992_ ) );
AND2_X1 _14986_ ( .A1(_06992_ ), .A2(_06926_ ), .ZN(_06993_ ) );
OAI21_X1 _14987_ ( .A(_06959_ ), .B1(_06966_ ), .B2(_06993_ ), .ZN(_06994_ ) );
AND3_X1 _14988_ ( .A1(_06992_ ), .A2(_06858_ ), .A3(_06928_ ), .ZN(_06995_ ) );
AND3_X1 _14989_ ( .A1(_04759_ ), .A2(_06812_ ), .A3(_06814_ ), .ZN(_06996_ ) );
AOI21_X1 _14990_ ( .A(_02838_ ), .B1(_06812_ ), .B2(_06814_ ), .ZN(_06997_ ) );
OR3_X1 _14991_ ( .A1(_06996_ ), .A2(_06997_ ), .A3(_06800_ ), .ZN(_06998_ ) );
AND3_X1 _14992_ ( .A1(_04678_ ), .A2(_06812_ ), .A3(_06814_ ), .ZN(_06999_ ) );
AOI21_X1 _14993_ ( .A(_02472_ ), .B1(_06822_ ), .B2(_06823_ ), .ZN(_07000_ ) );
OR3_X1 _14994_ ( .A1(_06999_ ), .A2(_07000_ ), .A3(_06819_ ), .ZN(_07001_ ) );
AOI21_X1 _14995_ ( .A(_06887_ ), .B1(_06998_ ), .B2(_07001_ ), .ZN(_07002_ ) );
AND3_X1 _14996_ ( .A1(_04256_ ), .A2(_06835_ ), .A3(_06836_ ), .ZN(_07003_ ) );
OAI21_X1 _14997_ ( .A(_06869_ ), .B1(_07003_ ), .B2(_06976_ ), .ZN(_07004_ ) );
AND3_X1 _14998_ ( .A1(_04372_ ), .A2(_05159_ ), .A3(_05160_ ), .ZN(_07005_ ) );
AOI21_X1 _14999_ ( .A(_02917_ ), .B1(_06812_ ), .B2(_06814_ ), .ZN(_07006_ ) );
OAI21_X1 _15000_ ( .A(_06864_ ), .B1(_07005_ ), .B2(_07006_ ), .ZN(_07007_ ) );
AND3_X1 _15001_ ( .A1(_07004_ ), .A2(_07007_ ), .A3(_06914_ ), .ZN(_07008_ ) );
OR3_X1 _15002_ ( .A1(_07002_ ), .A2(_07008_ ), .A3(_06902_ ), .ZN(_07009_ ) );
AND3_X1 _15003_ ( .A1(_04833_ ), .A2(_06835_ ), .A3(_06836_ ), .ZN(_07010_ ) );
AOI21_X1 _15004_ ( .A(_02571_ ), .B1(_06813_ ), .B2(_06815_ ), .ZN(_07011_ ) );
OR3_X1 _15005_ ( .A1(_07010_ ), .A2(_06826_ ), .A3(_07011_ ), .ZN(_07012_ ) );
AOI21_X1 _15006_ ( .A(_02886_ ), .B1(_06822_ ), .B2(_06823_ ), .ZN(_07013_ ) );
INV_X1 _15007_ ( .A(_07013_ ), .ZN(_07014_ ) );
OAI211_X1 _15008_ ( .A(_07014_ ), .B(_06827_ ), .C1(_04783_ ), .C2(_06799_ ), .ZN(_07015_ ) );
AND3_X1 _15009_ ( .A1(_07012_ ), .A2(_07015_ ), .A3(_06914_ ), .ZN(_07016_ ) );
AND3_X1 _15010_ ( .A1(_04907_ ), .A2(_06835_ ), .A3(_06836_ ), .ZN(_07017_ ) );
AOI21_X1 _15011_ ( .A(_02498_ ), .B1(_06835_ ), .B2(_06836_ ), .ZN(_07018_ ) );
NOR3_X1 _15012_ ( .A1(_07017_ ), .A2(_07018_ ), .A3(_06830_ ), .ZN(_07019_ ) );
AND3_X1 _15013_ ( .A1(_05172_ ), .A2(_06812_ ), .A3(_06814_ ), .ZN(_07020_ ) );
AOI21_X1 _15014_ ( .A(_02670_ ), .B1(_06822_ ), .B2(_06823_ ), .ZN(_07021_ ) );
NOR3_X1 _15015_ ( .A1(_07020_ ), .A2(_07021_ ), .A3(_06800_ ), .ZN(_07022_ ) );
NOR3_X1 _15016_ ( .A1(_07019_ ), .A2(_07022_ ), .A3(_06914_ ), .ZN(_07023_ ) );
OAI21_X1 _15017_ ( .A(_06919_ ), .B1(_07016_ ), .B2(_07023_ ), .ZN(_07024_ ) );
NAND3_X1 _15018_ ( .A1(_07009_ ), .A2(_06858_ ), .A3(_07024_ ), .ZN(_07025_ ) );
AOI21_X1 _15019_ ( .A(_05158_ ), .B1(_06862_ ), .B2(_06860_ ), .ZN(_07026_ ) );
AND2_X1 _15020_ ( .A1(_07026_ ), .A2(_06801_ ), .ZN(_07027_ ) );
INV_X1 _15021_ ( .A(_07027_ ), .ZN(_07028_ ) );
AND3_X1 _15022_ ( .A1(_04976_ ), .A2(_06813_ ), .A3(_06815_ ), .ZN(_07029_ ) );
AOI21_X1 _15023_ ( .A(_02774_ ), .B1(_06859_ ), .B2(_06867_ ), .ZN(_07030_ ) );
OAI21_X1 _15024_ ( .A(_06820_ ), .B1(_07029_ ), .B2(_07030_ ), .ZN(_07031_ ) );
BUF_X4 _15025_ ( .A(_06826_ ), .Z(_07032_ ) );
AND3_X1 _15026_ ( .A1(_06812_ ), .A2(_02781_ ), .A3(_06814_ ), .ZN(_07033_ ) );
AOI21_X1 _15027_ ( .A(_02622_ ), .B1(_06812_ ), .B2(_06814_ ), .ZN(_07034_ ) );
OAI21_X1 _15028_ ( .A(_07032_ ), .B1(_07033_ ), .B2(_07034_ ), .ZN(_07035_ ) );
NAND2_X1 _15029_ ( .A1(_07031_ ), .A2(_07035_ ), .ZN(_07036_ ) );
MUX2_X1 _15030_ ( .A(_07028_ ), .B(_07036_ ), .S(_06841_ ), .Z(_07037_ ) );
BUF_X2 _15031_ ( .A(_06853_ ), .Z(_07038_ ) );
OR3_X1 _15032_ ( .A1(_07037_ ), .A2(_07038_ ), .A3(_06902_ ), .ZN(_07039_ ) );
AOI21_X1 _15033_ ( .A(_05333_ ), .B1(_07025_ ), .B2(_07039_ ), .ZN(_07040_ ) );
AOI21_X1 _15034_ ( .A(_06930_ ), .B1(_05238_ ), .B2(_04444_ ), .ZN(_07041_ ) );
OR3_X1 _15035_ ( .A1(_05238_ ), .A2(_04444_ ), .A3(_05074_ ), .ZN(_07042_ ) );
OAI21_X1 _15036_ ( .A(_07042_ ), .B1(_06649_ ), .B2(_05331_ ), .ZN(_07043_ ) );
NOR4_X1 _15037_ ( .A1(_06995_ ), .A2(_07040_ ), .A3(_07041_ ), .A4(_07043_ ), .ZN(_07044_ ) );
NAND3_X1 _15038_ ( .A1(_06958_ ), .A2(_06994_ ), .A3(_07044_ ), .ZN(_07045_ ) );
AOI21_X1 _15039_ ( .A(_06953_ ), .B1(_07045_ ), .B2(_06942_ ), .ZN(_07046_ ) );
OAI21_X1 _15040_ ( .A(_06522_ ), .B1(_05512_ ), .B2(_06056_ ), .ZN(_07047_ ) );
OAI21_X1 _15041_ ( .A(_06945_ ), .B1(_07046_ ), .B2(_07047_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
OR2_X1 _15042_ ( .A1(_05551_ ), .A2(_06349_ ), .ZN(_07048_ ) );
NAND2_X1 _15043_ ( .A1(_05533_ ), .A2(_05648_ ), .ZN(_07049_ ) );
AOI22_X1 _15044_ ( .A1(_05530_ ), .A2(_06637_ ), .B1(\ID_EX_imm [19] ), .B2(_06640_ ), .ZN(_07050_ ) );
BUF_X2 _15045_ ( .A(_06933_ ), .Z(_07051_ ) );
INV_X1 _15046_ ( .A(_04371_ ), .ZN(_07052_ ) );
INV_X1 _15047_ ( .A(_04394_ ), .ZN(_07053_ ) );
AOI211_X1 _15048_ ( .A(_07052_ ), .B(_07053_ ), .C1(_05353_ ), .C2(_05369_ ), .ZN(_07054_ ) );
NOR3_X1 _15049_ ( .A1(_07054_ ), .A2(_05378_ ), .A3(_05377_ ), .ZN(_07055_ ) );
XNOR2_X1 _15050_ ( .A(_04338_ ), .B(_02917_ ), .ZN(_07056_ ) );
OAI21_X1 _15051_ ( .A(_04339_ ), .B1(_07055_ ), .B2(_07056_ ), .ZN(_07057_ ) );
AOI21_X1 _15052_ ( .A(_07051_ ), .B1(_07057_ ), .B2(_04313_ ), .ZN(_07058_ ) );
OAI21_X1 _15053_ ( .A(_07058_ ), .B1(_04313_ ), .B2(_07057_ ), .ZN(_07059_ ) );
AOI21_X1 _15054_ ( .A(_06647_ ), .B1(_07050_ ), .B2(_07059_ ), .ZN(_07060_ ) );
OR2_X1 _15055_ ( .A1(_07060_ ), .A2(_05433_ ), .ZN(_07061_ ) );
INV_X1 _15056_ ( .A(_06731_ ), .ZN(_07062_ ) );
BUF_X4 _15057_ ( .A(_07062_ ), .Z(_07063_ ) );
AND2_X1 _15058_ ( .A1(_06783_ ), .A2(_06785_ ), .ZN(_07064_ ) );
AND2_X1 _15059_ ( .A1(_06782_ ), .A2(_07064_ ), .ZN(_07065_ ) );
OAI21_X1 _15060_ ( .A(_06800_ ), .B1(_06832_ ), .B2(_06833_ ), .ZN(_07066_ ) );
OAI21_X1 _15061_ ( .A(_06830_ ), .B1(_06816_ ), .B2(_06817_ ), .ZN(_07067_ ) );
NAND3_X1 _15062_ ( .A1(_07066_ ), .A2(_07067_ ), .A3(_06803_ ), .ZN(_07068_ ) );
OAI21_X1 _15063_ ( .A(_06800_ ), .B1(_06896_ ), .B2(_06899_ ), .ZN(_07069_ ) );
OAI21_X1 _15064_ ( .A(_06819_ ), .B1(_06837_ ), .B2(_06838_ ), .ZN(_07070_ ) );
NAND3_X1 _15065_ ( .A1(_07069_ ), .A2(_07070_ ), .A3(_06753_ ), .ZN(_07071_ ) );
NAND2_X1 _15066_ ( .A1(_07068_ ), .A2(_07071_ ), .ZN(_07072_ ) );
INV_X1 _15067_ ( .A(_06824_ ), .ZN(_07073_ ) );
INV_X1 _15068_ ( .A(_06825_ ), .ZN(_07074_ ) );
NAND3_X1 _15069_ ( .A1(_07073_ ), .A2(_07074_ ), .A3(_06826_ ), .ZN(_07075_ ) );
NAND3_X1 _15070_ ( .A1(_06844_ ), .A2(_06819_ ), .A3(_06845_ ), .ZN(_07076_ ) );
AOI21_X1 _15071_ ( .A(_05166_ ), .B1(_07075_ ), .B2(_07076_ ), .ZN(_07077_ ) );
AND4_X1 _15072_ ( .A1(_03150_ ), .A2(_06655_ ), .A3(_05166_ ), .A4(_06826_ ), .ZN(_07078_ ) );
OR2_X1 _15073_ ( .A1(_07077_ ), .A2(_07078_ ), .ZN(_07079_ ) );
MUX2_X1 _15074_ ( .A(_07072_ ), .B(_07079_ ), .S(_06850_ ), .Z(_07080_ ) );
AOI21_X1 _15075_ ( .A(_07065_ ), .B1(_06858_ ), .B2(_07080_ ), .ZN(_07081_ ) );
XNOR2_X1 _15076_ ( .A(_06742_ ), .B(_06840_ ), .ZN(_07082_ ) );
NAND4_X1 _15077_ ( .A1(_06961_ ), .A2(_06962_ ), .A3(_07082_ ), .A4(_06783_ ), .ZN(_07083_ ) );
AOI21_X1 _15078_ ( .A(_07063_ ), .B1(_07081_ ), .B2(_07083_ ), .ZN(_07084_ ) );
INV_X1 _15079_ ( .A(_06718_ ), .ZN(_07085_ ) );
AOI211_X1 _15080_ ( .A(_05221_ ), .B(_05226_ ), .C1(_06684_ ), .C2(_06707_ ), .ZN(_07086_ ) );
INV_X1 _15081_ ( .A(_07086_ ), .ZN(_07087_ ) );
AND2_X1 _15082_ ( .A1(_07087_ ), .A2(_06714_ ), .ZN(_07088_ ) );
OAI211_X1 _15083_ ( .A(_05253_ ), .B(_07085_ ), .C1(_07088_ ), .C2(_05249_ ), .ZN(_07089_ ) );
AOI21_X1 _15084_ ( .A(_05249_ ), .B1(_07087_ ), .B2(_06714_ ), .ZN(_07090_ ) );
OAI21_X1 _15085_ ( .A(_05254_ ), .B1(_07090_ ), .B2(_06718_ ), .ZN(_07091_ ) );
AOI21_X1 _15086_ ( .A(_06727_ ), .B1(_07089_ ), .B2(_07091_ ), .ZN(_07092_ ) );
OAI21_X1 _15087_ ( .A(_06830_ ), .B1(_05161_ ), .B2(_06915_ ), .ZN(_07093_ ) );
OAI21_X1 _15088_ ( .A(_06827_ ), .B1(_06910_ ), .B2(_06911_ ), .ZN(_07094_ ) );
AND3_X1 _15089_ ( .A1(_07093_ ), .A2(_07094_ ), .A3(_06841_ ), .ZN(_07095_ ) );
BUF_X4 _15090_ ( .A(_06874_ ), .Z(_07096_ ) );
AND2_X1 _15091_ ( .A1(_07095_ ), .A2(_07096_ ), .ZN(_07097_ ) );
OAI21_X1 _15092_ ( .A(_05332_ ), .B1(_07097_ ), .B2(_06854_ ), .ZN(_07098_ ) );
NOR3_X1 _15093_ ( .A1(_06907_ ), .A2(_06908_ ), .A3(_06800_ ), .ZN(_07099_ ) );
NOR3_X1 _15094_ ( .A1(_06866_ ), .A2(_06868_ ), .A3(_06830_ ), .ZN(_07100_ ) );
NOR2_X1 _15095_ ( .A1(_07099_ ), .A2(_07100_ ), .ZN(_07101_ ) );
NAND2_X1 _15096_ ( .A1(_07101_ ), .A2(_06876_ ), .ZN(_07102_ ) );
AND3_X1 _15097_ ( .A1(_04808_ ), .A2(_06862_ ), .A3(_06860_ ), .ZN(_07103_ ) );
OAI21_X1 _15098_ ( .A(_06801_ ), .B1(_07103_ ), .B2(_06880_ ), .ZN(_07104_ ) );
OAI21_X1 _15099_ ( .A(_06831_ ), .B1(_06861_ ), .B2(_06863_ ), .ZN(_07105_ ) );
NAND2_X1 _15100_ ( .A1(_07104_ ), .A2(_07105_ ), .ZN(_07106_ ) );
NAND2_X1 _15101_ ( .A1(_07106_ ), .A2(_06872_ ), .ZN(_07107_ ) );
NAND2_X1 _15102_ ( .A1(_07102_ ), .A2(_07107_ ), .ZN(_07108_ ) );
NOR3_X1 _15103_ ( .A1(_06898_ ), .A2(_06899_ ), .A3(_06820_ ), .ZN(_07109_ ) );
NOR3_X1 _15104_ ( .A1(_06888_ ), .A2(_06889_ ), .A3(_07032_ ), .ZN(_07110_ ) );
NOR2_X1 _15105_ ( .A1(_07109_ ), .A2(_07110_ ), .ZN(_07111_ ) );
NOR3_X1 _15106_ ( .A1(_06891_ ), .A2(_06892_ ), .A3(_06820_ ), .ZN(_07112_ ) );
NOR3_X1 _15107_ ( .A1(_06877_ ), .A2(_06878_ ), .A3(_07032_ ), .ZN(_07113_ ) );
NOR2_X1 _15108_ ( .A1(_07112_ ), .A2(_07113_ ), .ZN(_07114_ ) );
MUX2_X1 _15109_ ( .A(_07111_ ), .B(_07114_ ), .S(_06805_ ), .Z(_07115_ ) );
MUX2_X1 _15110_ ( .A(_07108_ ), .B(_07115_ ), .S(_07096_ ), .Z(_07116_ ) );
AOI21_X1 _15111_ ( .A(_07098_ ), .B1(_07116_ ), .B2(_06858_ ), .ZN(_07117_ ) );
OR3_X1 _15112_ ( .A1(_05252_ ), .A2(_04256_ ), .A3(_05074_ ), .ZN(_07118_ ) );
OAI21_X1 _15113_ ( .A(_07118_ ), .B1(_05254_ ), .B2(_05331_ ), .ZN(_07119_ ) );
NOR4_X1 _15114_ ( .A1(_07084_ ), .A2(_07092_ ), .A3(_07117_ ), .A4(_07119_ ), .ZN(_07120_ ) );
BUF_X2 _15115_ ( .A(_06928_ ), .Z(_07121_ ) );
AND3_X1 _15116_ ( .A1(_07080_ ), .A2(_06926_ ), .A3(_07121_ ), .ZN(_07122_ ) );
AOI21_X1 _15117_ ( .A(_06930_ ), .B1(_05252_ ), .B2(_04256_ ), .ZN(_07123_ ) );
NOR2_X1 _15118_ ( .A1(_07122_ ), .A2(_07123_ ), .ZN(_07124_ ) );
AOI21_X1 _15119_ ( .A(_06939_ ), .B1(_07120_ ), .B2(_07124_ ), .ZN(_07125_ ) );
OAI21_X1 _15120_ ( .A(_07049_ ), .B1(_07061_ ), .B2(_07125_ ), .ZN(_07126_ ) );
OAI21_X1 _15121_ ( .A(_07048_ ), .B1(_07126_ ), .B2(_06384_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
AND2_X1 _15122_ ( .A1(_06960_ ), .A2(_06783_ ), .ZN(_07127_ ) );
NOR2_X1 _15123_ ( .A1(_07127_ ), .A2(_06786_ ), .ZN(_07128_ ) );
NAND3_X1 _15124_ ( .A1(_06782_ ), .A2(_06808_ ), .A3(_07082_ ), .ZN(_07129_ ) );
NOR2_X1 _15125_ ( .A1(_06799_ ), .A2(_06882_ ), .ZN(_07130_ ) );
OR2_X1 _15126_ ( .A1(_07129_ ), .A2(_07130_ ), .ZN(_07131_ ) );
AOI21_X1 _15127_ ( .A(_07128_ ), .B1(_07131_ ), .B2(_06788_ ), .ZN(_07132_ ) );
OAI21_X1 _15128_ ( .A(_05156_ ), .B1(_06978_ ), .B2(_06979_ ), .ZN(_07133_ ) );
OAI21_X1 _15129_ ( .A(_06818_ ), .B1(_06971_ ), .B2(_06972_ ), .ZN(_07134_ ) );
NAND3_X1 _15130_ ( .A1(_07133_ ), .A2(_07134_ ), .A3(_06811_ ), .ZN(_07135_ ) );
OAI21_X1 _15131_ ( .A(_07032_ ), .B1(_07003_ ), .B2(_07006_ ), .ZN(_07136_ ) );
OAI21_X1 _15132_ ( .A(_06820_ ), .B1(_06975_ ), .B2(_06976_ ), .ZN(_07137_ ) );
NAND3_X1 _15133_ ( .A1(_07136_ ), .A2(_07137_ ), .A3(_06914_ ), .ZN(_07138_ ) );
NAND2_X1 _15134_ ( .A1(_07135_ ), .A2(_07138_ ), .ZN(_07139_ ) );
BUF_X2 _15135_ ( .A(_06744_ ), .Z(_07140_ ) );
BUF_X2 _15136_ ( .A(_07140_ ), .Z(_07141_ ) );
NAND2_X1 _15137_ ( .A1(_07139_ ), .A2(_07141_ ), .ZN(_07142_ ) );
AND3_X1 _15138_ ( .A1(_06985_ ), .A2(_06804_ ), .A3(_06801_ ), .ZN(_07143_ ) );
AOI21_X1 _15139_ ( .A(_06818_ ), .B1(_06968_ ), .B2(_06969_ ), .ZN(_07144_ ) );
AOI21_X1 _15140_ ( .A(_05156_ ), .B1(_06987_ ), .B2(_06988_ ), .ZN(_07145_ ) );
NOR3_X1 _15141_ ( .A1(_07144_ ), .A2(_07145_ ), .A3(_06804_ ), .ZN(_07146_ ) );
NOR2_X1 _15142_ ( .A1(_07143_ ), .A2(_07146_ ), .ZN(_07147_ ) );
OAI21_X1 _15143_ ( .A(_07142_ ), .B1(_07147_ ), .B2(_07096_ ), .ZN(_07148_ ) );
AND2_X1 _15144_ ( .A1(_07148_ ), .A2(_06854_ ), .ZN(_07149_ ) );
OAI21_X1 _15145_ ( .A(_06959_ ), .B1(_07132_ ), .B2(_07149_ ), .ZN(_07150_ ) );
NAND3_X1 _15146_ ( .A1(_07148_ ), .A2(_06926_ ), .A3(_07121_ ), .ZN(_07151_ ) );
NAND3_X1 _15147_ ( .A1(_05245_ ), .A2(_06717_ ), .A3(_05246_ ), .ZN(_07152_ ) );
BUF_X4 _15148_ ( .A(_05323_ ), .Z(_07153_ ) );
NAND2_X1 _15149_ ( .A1(_07152_ ), .A2(_07153_ ), .ZN(_07154_ ) );
OAI21_X1 _15150_ ( .A(_06827_ ), .B1(_07029_ ), .B2(_07030_ ), .ZN(_07155_ ) );
OAI21_X1 _15151_ ( .A(_07155_ ), .B1(_07032_ ), .B2(_07026_ ), .ZN(_07156_ ) );
NOR3_X1 _15152_ ( .A1(_07156_ ), .A2(_06850_ ), .A3(_06804_ ), .ZN(_07157_ ) );
OAI21_X1 _15153_ ( .A(_05332_ ), .B1(_07157_ ), .B2(_06853_ ), .ZN(_07158_ ) );
OR3_X1 _15154_ ( .A1(_07020_ ), .A2(_07021_ ), .A3(_06818_ ), .ZN(_07159_ ) );
OR3_X1 _15155_ ( .A1(_07033_ ), .A2(_07034_ ), .A3(_05156_ ), .ZN(_07160_ ) );
AND3_X1 _15156_ ( .A1(_07159_ ), .A2(_07160_ ), .A3(_05166_ ), .ZN(_07161_ ) );
OAI21_X1 _15157_ ( .A(_06826_ ), .B1(_07010_ ), .B2(_07011_ ), .ZN(_07162_ ) );
OAI21_X1 _15158_ ( .A(_06819_ ), .B1(_07017_ ), .B2(_07018_ ), .ZN(_07163_ ) );
AOI21_X1 _15159_ ( .A(_05166_ ), .B1(_07162_ ), .B2(_07163_ ), .ZN(_07164_ ) );
OR2_X1 _15160_ ( .A1(_07161_ ), .A2(_07164_ ), .ZN(_07165_ ) );
OR3_X1 _15161_ ( .A1(_06999_ ), .A2(_07000_ ), .A3(_05156_ ), .ZN(_07166_ ) );
OR3_X1 _15162_ ( .A1(_07005_ ), .A2(_07006_ ), .A3(_06818_ ), .ZN(_07167_ ) );
AND3_X1 _15163_ ( .A1(_07166_ ), .A2(_07167_ ), .A3(_06753_ ), .ZN(_07168_ ) );
OR3_X1 _15164_ ( .A1(_06996_ ), .A2(_06997_ ), .A3(_06818_ ), .ZN(_07169_ ) );
OAI211_X1 _15165_ ( .A(_07014_ ), .B(_06818_ ), .C1(_04783_ ), .C2(_06655_ ), .ZN(_07170_ ) );
AND3_X1 _15166_ ( .A1(_07169_ ), .A2(_05166_ ), .A3(_07170_ ), .ZN(_07171_ ) );
OR2_X1 _15167_ ( .A1(_07168_ ), .A2(_07171_ ), .ZN(_07172_ ) );
MUX2_X1 _15168_ ( .A(_07165_ ), .B(_07172_ ), .S(_06744_ ), .Z(_07173_ ) );
AOI21_X1 _15169_ ( .A(_07158_ ), .B1(_07173_ ), .B2(_06853_ ), .ZN(_07174_ ) );
AOI221_X4 _15170_ ( .A(_07174_ ), .B1(_05073_ ), .B2(_06718_ ), .C1(_05248_ ), .C2(_05330_ ), .ZN(_07175_ ) );
NAND4_X1 _15171_ ( .A1(_07150_ ), .A2(_07151_ ), .A3(_07154_ ), .A4(_07175_ ), .ZN(_07176_ ) );
OAI21_X1 _15172_ ( .A(_06726_ ), .B1(_07088_ ), .B2(_05249_ ), .ZN(_07177_ ) );
AOI21_X1 _15173_ ( .A(_07177_ ), .B1(_05249_ ), .B2(_07088_ ), .ZN(_07178_ ) );
OAI21_X1 _15174_ ( .A(_06940_ ), .B1(_07176_ ), .B2(_07178_ ), .ZN(_07179_ ) );
AOI22_X1 _15175_ ( .A1(_05559_ ), .A2(_06637_ ), .B1(\ID_EX_imm [18] ), .B2(_06640_ ), .ZN(_07180_ ) );
AND2_X1 _15176_ ( .A1(_07055_ ), .A2(_07056_ ), .ZN(_07181_ ) );
BUF_X2 _15177_ ( .A(_06631_ ), .Z(_07182_ ) );
OAI21_X1 _15178_ ( .A(_07182_ ), .B1(_07055_ ), .B2(_07056_ ), .ZN(_07183_ ) );
OAI21_X1 _15179_ ( .A(_07180_ ), .B1(_07181_ ), .B2(_07183_ ), .ZN(_07184_ ) );
NAND2_X1 _15180_ ( .A1(_07184_ ), .A2(_06645_ ), .ZN(_07185_ ) );
AOI21_X1 _15181_ ( .A(_05648_ ), .B1(_07179_ ), .B2(_07185_ ), .ZN(_07186_ ) );
AND2_X1 _15182_ ( .A1(_05557_ ), .A2(_05648_ ), .ZN(_07187_ ) );
OAI21_X1 _15183_ ( .A(_06522_ ), .B1(_07186_ ), .B2(_07187_ ), .ZN(_07188_ ) );
NAND2_X1 _15184_ ( .A1(_05577_ ), .A2(_06354_ ), .ZN(_07189_ ) );
NAND2_X1 _15185_ ( .A1(_07188_ ), .A2(_07189_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _15186_ ( .A1(_05568_ ), .A2(\mtvec [17] ), .A3(_04097_ ), .ZN(_07190_ ) );
AND4_X1 _15187_ ( .A1(_05587_ ), .A2(_05588_ ), .A3(_05589_ ), .A4(_07190_ ), .ZN(_07191_ ) );
NAND4_X1 _15188_ ( .A1(_04069_ ), .A2(_05722_ ), .A3(_05574_ ), .A4(_07191_ ), .ZN(_07192_ ) );
NAND3_X1 _15189_ ( .A1(_05562_ ), .A2(_05592_ ), .A3(_05563_ ), .ZN(_07193_ ) );
NAND3_X1 _15190_ ( .A1(_07192_ ), .A2(_07193_ ), .A3(_06467_ ), .ZN(_07194_ ) );
INV_X1 _15191_ ( .A(_06636_ ), .ZN(_07195_ ) );
INV_X1 _15192_ ( .A(_06639_ ), .ZN(_07196_ ) );
OAI22_X1 _15193_ ( .A1(_05596_ ), .A2(_07195_ ), .B1(_02966_ ), .B2(_07196_ ), .ZN(_07197_ ) );
OR2_X1 _15194_ ( .A1(_06622_ ), .A2(_07052_ ), .ZN(_07198_ ) );
NAND2_X1 _15195_ ( .A1(_04370_ ), .A2(_02472_ ), .ZN(_07199_ ) );
AND3_X1 _15196_ ( .A1(_07198_ ), .A2(_07199_ ), .A3(_07053_ ), .ZN(_07200_ ) );
AOI21_X1 _15197_ ( .A(_07053_ ), .B1(_07198_ ), .B2(_07199_ ), .ZN(_07201_ ) );
NOR3_X1 _15198_ ( .A1(_07200_ ), .A2(_07201_ ), .A3(_07051_ ), .ZN(_07202_ ) );
OAI21_X1 _15199_ ( .A(_06645_ ), .B1(_07197_ ), .B2(_07202_ ), .ZN(_07203_ ) );
NAND2_X1 _15200_ ( .A1(_07203_ ), .A2(_05605_ ), .ZN(_07204_ ) );
NAND4_X1 _15201_ ( .A1(_06961_ ), .A2(_06802_ ), .A3(_06962_ ), .A4(_07082_ ), .ZN(_07205_ ) );
AOI22_X1 _15202_ ( .A1(_06787_ ), .A2(_06784_ ), .B1(_07205_ ), .B2(_06788_ ), .ZN(_07206_ ) );
NOR2_X1 _15203_ ( .A1(_06821_ ), .A2(_06828_ ), .ZN(_07207_ ) );
MUX2_X1 _15204_ ( .A(_07207_ ), .B(_06848_ ), .S(_06804_ ), .Z(_07208_ ) );
NAND2_X1 _15205_ ( .A1(_07208_ ), .A2(_06918_ ), .ZN(_07209_ ) );
OAI21_X1 _15206_ ( .A(_06864_ ), .B1(_06896_ ), .B2(_06899_ ), .ZN(_07210_ ) );
OAI21_X1 _15207_ ( .A(_06869_ ), .B1(_06898_ ), .B2(_06889_ ), .ZN(_07211_ ) );
AOI21_X1 _15208_ ( .A(_06811_ ), .B1(_07210_ ), .B2(_07211_ ), .ZN(_07212_ ) );
AOI21_X1 _15209_ ( .A(_06914_ ), .B1(_06834_ ), .B2(_06839_ ), .ZN(_07213_ ) );
OAI21_X1 _15210_ ( .A(_07141_ ), .B1(_07212_ ), .B2(_07213_ ), .ZN(_07214_ ) );
AND3_X1 _15211_ ( .A1(_07209_ ), .A2(_06854_ ), .A3(_07214_ ), .ZN(_07215_ ) );
OAI21_X1 _15212_ ( .A(_06959_ ), .B1(_07206_ ), .B2(_07215_ ), .ZN(_07216_ ) );
AOI21_X1 _15213_ ( .A(_05226_ ), .B1(_06684_ ), .B2(_06707_ ), .ZN(_07217_ ) );
OR3_X1 _15214_ ( .A1(_07217_ ), .A2(_05220_ ), .A3(_06713_ ), .ZN(_07218_ ) );
BUF_X4 _15215_ ( .A(_06726_ ), .Z(_07219_ ) );
OAI21_X1 _15216_ ( .A(_05220_ ), .B1(_07217_ ), .B2(_06713_ ), .ZN(_07220_ ) );
NAND3_X1 _15217_ ( .A1(_07218_ ), .A2(_07219_ ), .A3(_07220_ ), .ZN(_07221_ ) );
AND2_X1 _15218_ ( .A1(_07215_ ), .A2(_07121_ ), .ZN(_07222_ ) );
AND2_X1 _15219_ ( .A1(_06916_ ), .A2(_06887_ ), .ZN(_07223_ ) );
AND2_X1 _15220_ ( .A1(_07223_ ), .A2(_07096_ ), .ZN(_07224_ ) );
OAI21_X1 _15221_ ( .A(_05332_ ), .B1(_07224_ ), .B2(_06858_ ), .ZN(_07225_ ) );
NAND2_X1 _15222_ ( .A1(_06871_ ), .A2(_06872_ ), .ZN(_07226_ ) );
NAND3_X1 _15223_ ( .A1(_06909_ ), .A2(_06912_ ), .A3(_06876_ ), .ZN(_07227_ ) );
NAND2_X1 _15224_ ( .A1(_07226_ ), .A2(_07227_ ), .ZN(_07228_ ) );
AOI21_X1 _15225_ ( .A(_06887_ ), .B1(_06879_ ), .B2(_06883_ ), .ZN(_07229_ ) );
AOI21_X1 _15226_ ( .A(_06876_ ), .B1(_06890_ ), .B2(_06893_ ), .ZN(_07230_ ) );
NOR2_X1 _15227_ ( .A1(_07229_ ), .A2(_07230_ ), .ZN(_07231_ ) );
MUX2_X1 _15228_ ( .A(_07228_ ), .B(_07231_ ), .S(_06875_ ), .Z(_07232_ ) );
AOI21_X1 _15229_ ( .A(_07225_ ), .B1(_07232_ ), .B2(_06926_ ), .ZN(_07233_ ) );
BUF_X2 _15230_ ( .A(_05074_ ), .Z(_07234_ ) );
NOR3_X1 _15231_ ( .A1(_05219_ ), .A2(_04372_ ), .A3(_07234_ ), .ZN(_07235_ ) );
OAI22_X1 _15232_ ( .A1(_05221_ ), .A2(_05331_ ), .B1(_05258_ ), .B2(_06930_ ), .ZN(_07236_ ) );
NOR4_X1 _15233_ ( .A1(_07222_ ), .A2(_07233_ ), .A3(_07235_ ), .A4(_07236_ ), .ZN(_07237_ ) );
NAND3_X1 _15234_ ( .A1(_07216_ ), .A2(_07221_ ), .A3(_07237_ ), .ZN(_07238_ ) );
AOI21_X1 _15235_ ( .A(_07204_ ), .B1(_07238_ ), .B2(_06942_ ), .ZN(_07239_ ) );
NAND2_X1 _15236_ ( .A1(_05601_ ), .A2(_05431_ ), .ZN(_07240_ ) );
NAND2_X1 _15237_ ( .A1(_07240_ ), .A2(_06522_ ), .ZN(_07241_ ) );
OAI21_X1 _15238_ ( .A(_07194_ ), .B1(_07239_ ), .B2(_07241_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
NAND2_X1 _15239_ ( .A1(_05620_ ), .A2(_06441_ ), .ZN(_07242_ ) );
OAI21_X1 _15240_ ( .A(_07182_ ), .B1(_06622_ ), .B2(_07052_ ), .ZN(_07243_ ) );
AOI21_X1 _15241_ ( .A(_07243_ ), .B1(_07052_ ), .B2(_06622_ ), .ZN(_07244_ ) );
AND2_X1 _15242_ ( .A1(_05610_ ), .A2(_06949_ ), .ZN(_07245_ ) );
AND3_X1 _15243_ ( .A1(_06638_ ), .A2(\ID_EX_imm [16] ), .A3(_06635_ ), .ZN(_07246_ ) );
NOR3_X1 _15244_ ( .A1(_07244_ ), .A2(_07245_ ), .A3(_07246_ ), .ZN(_07247_ ) );
OAI21_X1 _15245_ ( .A(_05605_ ), .B1(_07247_ ), .B2(_06647_ ), .ZN(_07248_ ) );
AOI21_X1 _15246_ ( .A(_06784_ ), .B1(_06926_ ), .B2(_06794_ ), .ZN(_07249_ ) );
OR3_X1 _15247_ ( .A1(_07003_ ), .A2(_07006_ ), .A3(_06826_ ), .ZN(_07250_ ) );
OR3_X1 _15248_ ( .A1(_07005_ ), .A2(_07000_ ), .A3(_06819_ ), .ZN(_07251_ ) );
AND3_X1 _15249_ ( .A1(_07250_ ), .A2(_07251_ ), .A3(_06840_ ), .ZN(_07252_ ) );
AOI21_X1 _15250_ ( .A(_06886_ ), .B1(_06977_ ), .B2(_06980_ ), .ZN(_07253_ ) );
OR3_X1 _15251_ ( .A1(_07252_ ), .A2(_06850_ ), .A3(_07253_ ), .ZN(_07254_ ) );
OAI211_X1 _15252_ ( .A(_06986_ ), .B(_06811_ ), .C1(_06882_ ), .C2(_06989_ ), .ZN(_07255_ ) );
OR3_X1 _15253_ ( .A1(_06970_ ), .A2(_06973_ ), .A3(_06803_ ), .ZN(_07256_ ) );
NAND3_X1 _15254_ ( .A1(_07255_ ), .A2(_07256_ ), .A3(_06851_ ), .ZN(_07257_ ) );
NAND2_X1 _15255_ ( .A1(_07254_ ), .A2(_07257_ ), .ZN(_07258_ ) );
AND2_X1 _15256_ ( .A1(_07258_ ), .A2(_06854_ ), .ZN(_07259_ ) );
OAI21_X1 _15257_ ( .A(_06959_ ), .B1(_07249_ ), .B2(_07259_ ), .ZN(_07260_ ) );
NOR2_X1 _15258_ ( .A1(_07217_ ), .A2(_06954_ ), .ZN(_07261_ ) );
OAI21_X1 _15259_ ( .A(_07261_ ), .B1(_05225_ ), .B2(_06709_ ), .ZN(_07262_ ) );
AOI21_X1 _15260_ ( .A(_06804_ ), .B1(_06998_ ), .B2(_07001_ ), .ZN(_07263_ ) );
AOI21_X1 _15261_ ( .A(_06840_ ), .B1(_07012_ ), .B2(_07015_ ), .ZN(_07264_ ) );
NOR3_X1 _15262_ ( .A1(_07263_ ), .A2(_07264_ ), .A3(_06850_ ), .ZN(_07265_ ) );
OR3_X1 _15263_ ( .A1(_07019_ ), .A2(_07022_ ), .A3(_06803_ ), .ZN(_07266_ ) );
NAND2_X1 _15264_ ( .A1(_07036_ ), .A2(_06811_ ), .ZN(_07267_ ) );
NAND2_X1 _15265_ ( .A1(_07266_ ), .A2(_07267_ ), .ZN(_07268_ ) );
AOI211_X1 _15266_ ( .A(_05192_ ), .B(_07265_ ), .C1(_06918_ ), .C2(_07268_ ), .ZN(_07269_ ) );
AND3_X1 _15267_ ( .A1(_07026_ ), .A2(_06886_ ), .A3(_06869_ ), .ZN(_07270_ ) );
AND3_X1 _15268_ ( .A1(_07270_ ), .A2(_05192_ ), .A3(_07140_ ), .ZN(_07271_ ) );
OAI21_X1 _15269_ ( .A(_05332_ ), .B1(_07269_ ), .B2(_07271_ ), .ZN(_07272_ ) );
INV_X1 _15270_ ( .A(_06713_ ), .ZN(_07273_ ) );
OAI221_X1 _15271_ ( .A(_07272_ ), .B1(_05074_ ), .B2(_07273_ ), .C1(_05226_ ), .C2(_05331_ ), .ZN(_07274_ ) );
NAND3_X1 _15272_ ( .A1(_05222_ ), .A2(_04342_ ), .A3(_05223_ ), .ZN(_07275_ ) );
AOI221_X4 _15273_ ( .A(_07274_ ), .B1(_07275_ ), .B2(_05323_ ), .C1(_06928_ ), .C2(_07259_ ), .ZN(_07276_ ) );
NAND3_X1 _15274_ ( .A1(_07260_ ), .A2(_07262_ ), .A3(_07276_ ), .ZN(_07277_ ) );
AOI21_X1 _15275_ ( .A(_07248_ ), .B1(_07277_ ), .B2(_06942_ ), .ZN(_07278_ ) );
BUF_X4 _15276_ ( .A(_06359_ ), .Z(_07279_ ) );
OAI21_X1 _15277_ ( .A(_07279_ ), .B1(_05609_ ), .B2(_06056_ ), .ZN(_07280_ ) );
OAI21_X1 _15278_ ( .A(_07242_ ), .B1(_07278_ ), .B2(_07280_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
NAND2_X1 _15279_ ( .A1(_05633_ ), .A2(_06441_ ), .ZN(_07281_ ) );
AND2_X1 _15280_ ( .A1(_06679_ ), .A2(_06683_ ), .ZN(_07282_ ) );
INV_X1 _15281_ ( .A(_07282_ ), .ZN(_07283_ ) );
AND2_X1 _15282_ ( .A1(_07283_ ), .A2(_06695_ ), .ZN(_07284_ ) );
AND2_X1 _15283_ ( .A1(_05116_ ), .A2(_04759_ ), .ZN(_07285_ ) );
OR4_X1 _15284_ ( .A1(_06699_ ), .A2(_07284_ ), .A3(_07285_ ), .A4(_05123_ ), .ZN(_07286_ ) );
AOI21_X1 _15285_ ( .A(_06703_ ), .B1(_07286_ ), .B2(_06701_ ), .ZN(_07287_ ) );
OR3_X1 _15286_ ( .A1(_07287_ ), .A2(_06702_ ), .A3(_06705_ ), .ZN(_07288_ ) );
OAI21_X1 _15287_ ( .A(_06702_ ), .B1(_07287_ ), .B2(_06705_ ), .ZN(_07289_ ) );
AOI21_X1 _15288_ ( .A(_06954_ ), .B1(_07288_ ), .B2(_07289_ ), .ZN(_07290_ ) );
BUF_X2 _15289_ ( .A(_07064_ ), .Z(_07291_ ) );
AOI21_X1 _15290_ ( .A(_06886_ ), .B1(_07075_ ), .B2(_07076_ ), .ZN(_07292_ ) );
AND3_X1 _15291_ ( .A1(_07066_ ), .A2(_07067_ ), .A3(_06840_ ), .ZN(_07293_ ) );
OAI21_X1 _15292_ ( .A(_06902_ ), .B1(_07292_ ), .B2(_07293_ ), .ZN(_07294_ ) );
OAI21_X1 _15293_ ( .A(_07032_ ), .B1(_06888_ ), .B2(_06892_ ), .ZN(_07295_ ) );
OAI21_X1 _15294_ ( .A(_06820_ ), .B1(_06898_ ), .B2(_06889_ ), .ZN(_07296_ ) );
NAND2_X1 _15295_ ( .A1(_07295_ ), .A2(_07296_ ), .ZN(_07297_ ) );
NAND2_X1 _15296_ ( .A1(_07297_ ), .A2(_06872_ ), .ZN(_07298_ ) );
NAND2_X1 _15297_ ( .A1(_07069_ ), .A2(_07070_ ), .ZN(_07299_ ) );
NAND2_X1 _15298_ ( .A1(_07299_ ), .A2(_06876_ ), .ZN(_07300_ ) );
NAND3_X1 _15299_ ( .A1(_07298_ ), .A2(_07300_ ), .A3(_07141_ ), .ZN(_07301_ ) );
NAND3_X1 _15300_ ( .A1(_07294_ ), .A2(_07301_ ), .A3(_07038_ ), .ZN(_07302_ ) );
NAND3_X1 _15301_ ( .A1(_06847_ ), .A2(_06841_ ), .A3(_06895_ ), .ZN(_07303_ ) );
OAI21_X1 _15302_ ( .A(_06906_ ), .B1(_07303_ ), .B2(_06902_ ), .ZN(_07304_ ) );
AOI22_X1 _15303_ ( .A1(_06782_ ), .A2(_07291_ ), .B1(_07302_ ), .B2(_07304_ ), .ZN(_07305_ ) );
NOR2_X1 _15304_ ( .A1(_07305_ ), .A2(_07063_ ), .ZN(_07306_ ) );
AND3_X1 _15305_ ( .A1(_07302_ ), .A2(_06928_ ), .A3(_07304_ ), .ZN(_07307_ ) );
AND2_X1 _15306_ ( .A1(_05186_ ), .A2(_05332_ ), .ZN(_07308_ ) );
BUF_X4 _15307_ ( .A(_07308_ ), .Z(_07309_ ) );
NAND2_X1 _15308_ ( .A1(_07093_ ), .A2(_07094_ ), .ZN(_07310_ ) );
MUX2_X1 _15309_ ( .A(_07310_ ), .B(_07101_ ), .S(_06886_ ), .Z(_07311_ ) );
NOR2_X1 _15310_ ( .A1(_07311_ ), .A2(_07096_ ), .ZN(_07312_ ) );
NAND2_X1 _15311_ ( .A1(_07114_ ), .A2(_06841_ ), .ZN(_07313_ ) );
NAND2_X1 _15312_ ( .A1(_07106_ ), .A2(_06811_ ), .ZN(_07314_ ) );
AND3_X1 _15313_ ( .A1(_07313_ ), .A2(_07314_ ), .A3(_07141_ ), .ZN(_07315_ ) );
OAI21_X1 _15314_ ( .A(_07309_ ), .B1(_07312_ ), .B2(_07315_ ), .ZN(_07316_ ) );
NAND3_X1 _15315_ ( .A1(_05214_ ), .A2(_02815_ ), .A3(_05073_ ), .ZN(_07317_ ) );
OAI211_X1 _15316_ ( .A(_07316_ ), .B(_07317_ ), .C1(_06702_ ), .C2(_05331_ ), .ZN(_07318_ ) );
NOR4_X1 _15317_ ( .A1(_07290_ ), .A2(_07306_ ), .A3(_07307_ ), .A4(_07318_ ), .ZN(_07319_ ) );
OAI21_X1 _15318_ ( .A(_07153_ ), .B1(_05214_ ), .B2(_02815_ ), .ZN(_07320_ ) );
AOI21_X1 _15319_ ( .A(_06939_ ), .B1(_07319_ ), .B2(_07320_ ), .ZN(_07321_ ) );
AOI21_X1 _15320_ ( .A(_05344_ ), .B1(_05368_ ), .B2(_04880_ ), .ZN(_07322_ ) );
INV_X1 _15321_ ( .A(_04757_ ), .ZN(_07323_ ) );
OR2_X1 _15322_ ( .A1(_07322_ ), .A2(_07323_ ), .ZN(_07324_ ) );
AND2_X1 _15323_ ( .A1(_07324_ ), .A2(_05349_ ), .ZN(_07325_ ) );
OAI21_X1 _15324_ ( .A(_05348_ ), .B1(_07325_ ), .B2(_05346_ ), .ZN(_07326_ ) );
AND2_X1 _15325_ ( .A1(_07326_ ), .A2(_04732_ ), .ZN(_07327_ ) );
OR3_X1 _15326_ ( .A1(_07327_ ), .A2(_04707_ ), .A3(_05335_ ), .ZN(_07328_ ) );
OAI21_X1 _15327_ ( .A(_04707_ ), .B1(_07327_ ), .B2(_05335_ ), .ZN(_07329_ ) );
NAND3_X1 _15328_ ( .A1(_07328_ ), .A2(_06632_ ), .A3(_07329_ ), .ZN(_07330_ ) );
AOI22_X1 _15329_ ( .A1(_05642_ ), .A2(_06949_ ), .B1(\ID_EX_imm [15] ), .B2(_06640_ ), .ZN(_07331_ ) );
AOI21_X1 _15330_ ( .A(_06946_ ), .B1(_07330_ ), .B2(_07331_ ), .ZN(_07332_ ) );
OR2_X1 _15331_ ( .A1(_07332_ ), .A2(_05433_ ), .ZN(_07333_ ) );
OAI22_X1 _15332_ ( .A1(_07321_ ), .A2(_07333_ ), .B1(_05963_ ), .B2(_05636_ ), .ZN(_07334_ ) );
OAI21_X1 _15333_ ( .A(_07281_ ), .B1(_07334_ ), .B2(_06384_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
NAND3_X1 _15334_ ( .A1(_05562_ ), .A2(_05659_ ), .A3(_05563_ ), .ZN(_07335_ ) );
INV_X1 _15335_ ( .A(_05497_ ), .ZN(_07336_ ) );
NAND4_X1 _15336_ ( .A1(_05649_ ), .A2(_05657_ ), .A3(_05650_ ), .A4(_05655_ ), .ZN(_07337_ ) );
OAI211_X1 _15337_ ( .A(_07335_ ), .B(_06385_ ), .C1(_07336_ ), .C2(_07337_ ), .ZN(_07338_ ) );
AOI21_X1 _15338_ ( .A(_07051_ ), .B1(_07326_ ), .B2(_04732_ ), .ZN(_07339_ ) );
OAI21_X1 _15339_ ( .A(_07339_ ), .B1(_04732_ ), .B2(_07326_ ), .ZN(_07340_ ) );
AOI22_X1 _15340_ ( .A1(_05667_ ), .A2(_06949_ ), .B1(\ID_EX_imm [14] ), .B2(_06950_ ), .ZN(_07341_ ) );
AOI21_X1 _15341_ ( .A(_06946_ ), .B1(_07340_ ), .B2(_07341_ ), .ZN(_07342_ ) );
OR2_X1 _15342_ ( .A1(_07342_ ), .A2(_05433_ ), .ZN(_07343_ ) );
AND3_X1 _15343_ ( .A1(_07286_ ), .A2(_06703_ ), .A3(_06701_ ), .ZN(_07344_ ) );
NOR3_X1 _15344_ ( .A1(_07344_ ), .A2(_07287_ ), .A3(_06954_ ), .ZN(_07345_ ) );
NAND3_X1 _15345_ ( .A1(_06963_ ), .A2(_06886_ ), .A3(_06801_ ), .ZN(_07346_ ) );
OAI211_X1 _15346_ ( .A(_06782_ ), .B(_07291_ ), .C1(_06962_ ), .C2(_07346_ ), .ZN(_07347_ ) );
OR3_X1 _15347_ ( .A1(_07005_ ), .A2(_07000_ ), .A3(_06826_ ), .ZN(_07348_ ) );
OR3_X1 _15348_ ( .A1(_06999_ ), .A2(_06997_ ), .A3(_06819_ ), .ZN(_07349_ ) );
AND3_X1 _15349_ ( .A1(_07348_ ), .A2(_07349_ ), .A3(_06840_ ), .ZN(_07350_ ) );
AOI21_X1 _15350_ ( .A(_06840_ ), .B1(_07136_ ), .B2(_07137_ ), .ZN(_07351_ ) );
OAI21_X1 _15351_ ( .A(_06744_ ), .B1(_07350_ ), .B2(_07351_ ), .ZN(_07352_ ) );
OR3_X1 _15352_ ( .A1(_07144_ ), .A2(_07145_ ), .A3(_06753_ ), .ZN(_07353_ ) );
NAND3_X1 _15353_ ( .A1(_07133_ ), .A2(_07134_ ), .A3(_06753_ ), .ZN(_07354_ ) );
NAND3_X1 _15354_ ( .A1(_07353_ ), .A2(_06850_ ), .A3(_07354_ ), .ZN(_07355_ ) );
AND4_X1 _15355_ ( .A1(_05184_ ), .A2(_07352_ ), .A3(_05183_ ), .A4(_07355_ ), .ZN(_07356_ ) );
AND3_X1 _15356_ ( .A1(_06985_ ), .A2(_06753_ ), .A3(_06827_ ), .ZN(_07357_ ) );
AND3_X1 _15357_ ( .A1(_07357_ ), .A2(_05192_ ), .A3(_07140_ ), .ZN(_07358_ ) );
NOR2_X1 _15358_ ( .A1(_07356_ ), .A2(_07358_ ), .ZN(_07359_ ) );
AOI21_X1 _15359_ ( .A(_07063_ ), .B1(_07347_ ), .B2(_07359_ ), .ZN(_07360_ ) );
INV_X1 _15360_ ( .A(_06927_ ), .ZN(_07361_ ) );
NOR2_X1 _15361_ ( .A1(_07359_ ), .A2(_07361_ ), .ZN(_07362_ ) );
AND2_X1 _15362_ ( .A1(_05108_ ), .A2(_05330_ ), .ZN(_07363_ ) );
INV_X1 _15363_ ( .A(_07308_ ), .ZN(_07364_ ) );
AND3_X1 _15364_ ( .A1(_07159_ ), .A2(_07160_ ), .A3(_06840_ ), .ZN(_07365_ ) );
AOI21_X1 _15365_ ( .A(_07365_ ), .B1(_06804_ ), .B2(_07156_ ), .ZN(_07366_ ) );
NAND2_X1 _15366_ ( .A1(_07366_ ), .A2(_06851_ ), .ZN(_07367_ ) );
AOI21_X1 _15367_ ( .A(_06804_ ), .B1(_07169_ ), .B2(_07170_ ), .ZN(_07368_ ) );
AND3_X1 _15368_ ( .A1(_07162_ ), .A2(_07163_ ), .A3(_06803_ ), .ZN(_07369_ ) );
OAI21_X1 _15369_ ( .A(_07140_ ), .B1(_07368_ ), .B2(_07369_ ), .ZN(_07370_ ) );
AOI21_X1 _15370_ ( .A(_07364_ ), .B1(_07367_ ), .B2(_07370_ ), .ZN(_07371_ ) );
NOR3_X1 _15371_ ( .A1(_05107_ ), .A2(_04708_ ), .A3(_05074_ ), .ZN(_07372_ ) );
OR2_X1 _15372_ ( .A1(_07371_ ), .A2(_07372_ ), .ZN(_07373_ ) );
AOI21_X1 _15373_ ( .A(_05324_ ), .B1(_05107_ ), .B2(_04708_ ), .ZN(_07374_ ) );
OR4_X1 _15374_ ( .A1(_07362_ ), .A2(_07363_ ), .A3(_07373_ ), .A4(_07374_ ), .ZN(_07375_ ) );
OR3_X1 _15375_ ( .A1(_07345_ ), .A2(_07360_ ), .A3(_07375_ ), .ZN(_07376_ ) );
AOI21_X1 _15376_ ( .A(_07343_ ), .B1(_07376_ ), .B2(_06942_ ), .ZN(_07377_ ) );
OAI21_X1 _15377_ ( .A(_07279_ ), .B1(_05665_ ), .B2(_06056_ ), .ZN(_07378_ ) );
OAI21_X1 _15378_ ( .A(_07338_ ), .B1(_07377_ ), .B2(_07378_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
OR3_X1 _15379_ ( .A1(_05677_ ), .A2(_05679_ ), .A3(_06359_ ), .ZN(_07379_ ) );
XNOR2_X1 _15380_ ( .A(_07325_ ), .B(_04781_ ), .ZN(_07380_ ) );
NAND2_X1 _15381_ ( .A1(_07380_ ), .A2(_06632_ ), .ZN(_07381_ ) );
AOI22_X1 _15382_ ( .A1(_05685_ ), .A2(_06949_ ), .B1(\ID_EX_imm [13] ), .B2(_06950_ ), .ZN(_07382_ ) );
AOI21_X1 _15383_ ( .A(_06946_ ), .B1(_07381_ ), .B2(_07382_ ), .ZN(_07383_ ) );
OR2_X1 _15384_ ( .A1(_07383_ ), .A2(_05433_ ), .ZN(_07384_ ) );
NAND2_X1 _15385_ ( .A1(_06843_ ), .A2(_06902_ ), .ZN(_07385_ ) );
OR3_X1 _15386_ ( .A1(_06888_ ), .A2(_06892_ ), .A3(_07032_ ), .ZN(_07386_ ) );
OR3_X1 _15387_ ( .A1(_06891_ ), .A2(_06878_ ), .A3(_06820_ ), .ZN(_07387_ ) );
NAND2_X1 _15388_ ( .A1(_07386_ ), .A2(_07387_ ), .ZN(_07388_ ) );
NAND2_X1 _15389_ ( .A1(_07388_ ), .A2(_06887_ ), .ZN(_07389_ ) );
NAND3_X1 _15390_ ( .A1(_07210_ ), .A2(_07211_ ), .A3(_06876_ ), .ZN(_07390_ ) );
NAND2_X1 _15391_ ( .A1(_07389_ ), .A2(_07390_ ), .ZN(_07391_ ) );
INV_X1 _15392_ ( .A(_07391_ ), .ZN(_07392_ ) );
OAI211_X1 _15393_ ( .A(_06854_ ), .B(_07385_ ), .C1(_07392_ ), .C2(_06919_ ), .ZN(_07393_ ) );
NOR3_X1 _15394_ ( .A1(_06848_ ), .A2(_06851_ ), .A3(_06805_ ), .ZN(_07394_ ) );
OR2_X1 _15395_ ( .A1(_07394_ ), .A2(_07038_ ), .ZN(_07395_ ) );
AND3_X1 _15396_ ( .A1(_07393_ ), .A2(_06928_ ), .A3(_07395_ ), .ZN(_07396_ ) );
OAI211_X1 _15397_ ( .A(_06961_ ), .B(_07291_ ), .C1(_06806_ ), .C2(_06962_ ), .ZN(_07397_ ) );
NAND2_X1 _15398_ ( .A1(_07393_ ), .A2(_07395_ ), .ZN(_07398_ ) );
AOI21_X1 _15399_ ( .A(_07063_ ), .B1(_07397_ ), .B2(_07398_ ), .ZN(_07399_ ) );
OAI21_X1 _15400_ ( .A(_06875_ ), .B1(_06873_ ), .B2(_06884_ ), .ZN(_07400_ ) );
BUF_X4 _15401_ ( .A(_07096_ ), .Z(_07401_ ) );
OAI21_X1 _15402_ ( .A(_07400_ ), .B1(_06917_ ), .B2(_07401_ ), .ZN(_07402_ ) );
AOI211_X1 _15403_ ( .A(_07396_ ), .B(_07399_ ), .C1(_07309_ ), .C2(_07402_ ), .ZN(_07403_ ) );
AOI21_X1 _15404_ ( .A(_05123_ ), .B1(_07283_ ), .B2(_06695_ ), .ZN(_07404_ ) );
OR3_X1 _15405_ ( .A1(_07404_ ), .A2(_05117_ ), .A3(_06700_ ), .ZN(_07405_ ) );
OAI21_X1 _15406_ ( .A(_05117_ ), .B1(_07404_ ), .B2(_06700_ ), .ZN(_07406_ ) );
NAND3_X1 _15407_ ( .A1(_07405_ ), .A2(_07219_ ), .A3(_07406_ ), .ZN(_07407_ ) );
OR3_X1 _15408_ ( .A1(_05116_ ), .A2(_04759_ ), .A3(_07234_ ), .ZN(_07408_ ) );
OAI21_X1 _15409_ ( .A(_07408_ ), .B1(_07285_ ), .B2(_06930_ ), .ZN(_07409_ ) );
BUF_X2 _15410_ ( .A(_06922_ ), .Z(_07410_ ) );
AOI21_X1 _15411_ ( .A(_07409_ ), .B1(_05117_ ), .B2(_07410_ ), .ZN(_07411_ ) );
NAND3_X1 _15412_ ( .A1(_07403_ ), .A2(_07407_ ), .A3(_07411_ ), .ZN(_07412_ ) );
AOI21_X1 _15413_ ( .A(_07384_ ), .B1(_07412_ ), .B2(_06942_ ), .ZN(_07413_ ) );
NAND2_X1 _15414_ ( .A1(_05681_ ), .A2(_05648_ ), .ZN(_07414_ ) );
NAND2_X1 _15415_ ( .A1(_07414_ ), .A2(_06522_ ), .ZN(_07415_ ) );
OAI21_X1 _15416_ ( .A(_07379_ ), .B1(_07413_ ), .B2(_07415_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
NAND2_X1 _15417_ ( .A1(_07322_ ), .A2(_07323_ ), .ZN(_07416_ ) );
NAND3_X1 _15418_ ( .A1(_07324_ ), .A2(_06632_ ), .A3(_07416_ ), .ZN(_07417_ ) );
NAND3_X1 _15419_ ( .A1(_05692_ ), .A2(_05683_ ), .A3(_06637_ ), .ZN(_07418_ ) );
NAND3_X1 _15420_ ( .A1(_06638_ ), .A2(\ID_EX_imm [12] ), .A3(_06635_ ), .ZN(_07419_ ) );
NAND3_X1 _15421_ ( .A1(_07417_ ), .A2(_07418_ ), .A3(_07419_ ), .ZN(_07420_ ) );
AOI21_X1 _15422_ ( .A(_05433_ ), .B1(_07420_ ), .B2(_06645_ ), .ZN(_07421_ ) );
OAI211_X1 _15423_ ( .A(_06961_ ), .B(_07291_ ), .C1(_06808_ ), .C2(_06964_ ), .ZN(_07422_ ) );
NAND3_X1 _15424_ ( .A1(_07250_ ), .A2(_07251_ ), .A3(_06803_ ), .ZN(_07423_ ) );
OR3_X1 _15425_ ( .A1(_06999_ ), .A2(_06997_ ), .A3(_06826_ ), .ZN(_07424_ ) );
OAI211_X1 _15426_ ( .A(_07014_ ), .B(_06800_ ), .C1(_04758_ ), .C2(_06799_ ), .ZN(_07425_ ) );
NAND3_X1 _15427_ ( .A1(_07424_ ), .A2(_06840_ ), .A3(_07425_ ), .ZN(_07426_ ) );
AND2_X1 _15428_ ( .A1(_07423_ ), .A2(_07426_ ), .ZN(_07427_ ) );
OR2_X1 _15429_ ( .A1(_07427_ ), .A2(_06850_ ), .ZN(_07428_ ) );
OAI211_X1 _15430_ ( .A(_07428_ ), .B(_06853_ ), .C1(_07141_ ), .C2(_06982_ ), .ZN(_07429_ ) );
NAND4_X1 _15431_ ( .A1(_06990_ ), .A2(_06905_ ), .A3(_06874_ ), .A4(_06872_ ), .ZN(_07430_ ) );
AND2_X1 _15432_ ( .A1(_07429_ ), .A2(_07430_ ), .ZN(_07431_ ) );
AOI21_X1 _15433_ ( .A(_07063_ ), .B1(_07422_ ), .B2(_07431_ ), .ZN(_07432_ ) );
AOI21_X1 _15434_ ( .A(_07361_ ), .B1(_07429_ ), .B2(_07430_ ), .ZN(_07433_ ) );
NOR2_X1 _15435_ ( .A1(_07037_ ), .A2(_07096_ ), .ZN(_07434_ ) );
NOR3_X1 _15436_ ( .A1(_07016_ ), .A2(_07023_ ), .A3(_06918_ ), .ZN(_07435_ ) );
NOR2_X1 _15437_ ( .A1(_07434_ ), .A2(_07435_ ), .ZN(_07436_ ) );
NOR2_X1 _15438_ ( .A1(_07436_ ), .A2(_07364_ ), .ZN(_07437_ ) );
OR3_X1 _15439_ ( .A1(_07432_ ), .A2(_07433_ ), .A3(_07437_ ), .ZN(_07438_ ) );
OAI21_X1 _15440_ ( .A(_06726_ ), .B1(_07284_ ), .B2(_05123_ ), .ZN(_07439_ ) );
AOI21_X1 _15441_ ( .A(_07439_ ), .B1(_05123_ ), .B2(_07284_ ), .ZN(_07440_ ) );
AND2_X1 _15442_ ( .A1(_05122_ ), .A2(_06922_ ), .ZN(_07441_ ) );
AOI21_X1 _15443_ ( .A(_05324_ ), .B1(_05121_ ), .B2(_04734_ ), .ZN(_07442_ ) );
NOR3_X1 _15444_ ( .A1(_05121_ ), .A2(_04734_ ), .A3(_07234_ ), .ZN(_07443_ ) );
OR3_X1 _15445_ ( .A1(_07441_ ), .A2(_07442_ ), .A3(_07443_ ), .ZN(_07444_ ) );
NOR3_X1 _15446_ ( .A1(_07438_ ), .A2(_07440_ ), .A3(_07444_ ), .ZN(_07445_ ) );
OAI21_X1 _15447_ ( .A(_07421_ ), .B1(_07445_ ), .B2(_06939_ ), .ZN(_07446_ ) );
OR2_X1 _15448_ ( .A1(_05691_ ), .A2(_05425_ ), .ZN(_07447_ ) );
NAND3_X1 _15449_ ( .A1(_07446_ ), .A2(_06350_ ), .A3(_07447_ ), .ZN(_07448_ ) );
NAND3_X1 _15450_ ( .A1(_06438_ ), .A2(_06439_ ), .A3(_06401_ ), .ZN(_07449_ ) );
NAND2_X1 _15451_ ( .A1(_07448_ ), .A2(_07449_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
OR2_X1 _15452_ ( .A1(_04109_ ), .A2(_06349_ ), .ZN(_07450_ ) );
INV_X1 _15453_ ( .A(_05285_ ), .ZN(_07451_ ) );
AND2_X1 _15454_ ( .A1(_05243_ ), .A2(_05239_ ), .ZN(_07452_ ) );
NAND4_X1 _15455_ ( .A1(_06957_ ), .A2(_05230_ ), .A3(_05234_ ), .A4(_07452_ ), .ZN(_07453_ ) );
AND2_X1 _15456_ ( .A1(_05243_ ), .A2(_06722_ ), .ZN(_07454_ ) );
OAI211_X1 _15457_ ( .A(_05230_ ), .B(_05234_ ), .C1(_07454_ ), .C2(_06923_ ), .ZN(_07455_ ) );
OR2_X1 _15458_ ( .A1(_05229_ ), .A2(_04420_ ), .ZN(_07456_ ) );
AND2_X1 _15459_ ( .A1(_05233_ ), .A2(_02373_ ), .ZN(_07457_ ) );
NAND2_X1 _15460_ ( .A1(_05230_ ), .A2(_07457_ ), .ZN(_07458_ ) );
AND3_X1 _15461_ ( .A1(_07455_ ), .A2(_07456_ ), .A3(_07458_ ), .ZN(_07459_ ) );
AND2_X1 _15462_ ( .A1(_07453_ ), .A2(_07459_ ), .ZN(_07460_ ) );
INV_X1 _15463_ ( .A(_07460_ ), .ZN(_07461_ ) );
NAND3_X2 _15464_ ( .A1(_07461_ ), .A2(_05294_ ), .A3(_05300_ ), .ZN(_07462_ ) );
INV_X1 _15465_ ( .A(_05299_ ), .ZN(_07463_ ) );
AOI21_X1 _15466_ ( .A(_05298_ ), .B1(_05292_ ), .B2(_07463_ ), .ZN(_07464_ ) );
AOI211_X2 _15467_ ( .A(_05305_ ), .B(_07451_ ), .C1(_07462_ ), .C2(_07464_ ), .ZN(_07465_ ) );
NOR2_X1 _15468_ ( .A1(_05277_ ), .A2(_05307_ ), .ZN(_07466_ ) );
AOI21_X1 _15469_ ( .A(_07466_ ), .B1(_05278_ ), .B2(_05283_ ), .ZN(_07467_ ) );
INV_X1 _15470_ ( .A(_07467_ ), .ZN(_07468_ ) );
OAI211_X1 _15471_ ( .A(_05095_ ), .B(_05101_ ), .C1(_07465_ ), .C2(_07468_ ), .ZN(_07469_ ) );
INV_X1 _15472_ ( .A(_05081_ ), .ZN(_07470_ ) );
AND2_X1 _15473_ ( .A1(_05099_ ), .A2(_03095_ ), .ZN(_07471_ ) );
AND2_X1 _15474_ ( .A1(_07471_ ), .A2(_05095_ ), .ZN(_07472_ ) );
AOI21_X1 _15475_ ( .A(_07472_ ), .B1(_03118_ ), .B2(_05093_ ), .ZN(_07473_ ) );
AND3_X1 _15476_ ( .A1(_07469_ ), .A2(_07470_ ), .A3(_07473_ ), .ZN(_07474_ ) );
AOI21_X1 _15477_ ( .A(_07470_ ), .B1(_07469_ ), .B2(_07473_ ), .ZN(_07475_ ) );
OR3_X2 _15478_ ( .A1(_07474_ ), .A2(_07475_ ), .A3(_06954_ ), .ZN(_07476_ ) );
NAND2_X1 _15479_ ( .A1(_05081_ ), .A2(_07410_ ), .ZN(_07477_ ) );
AND4_X1 _15480_ ( .A1(_06808_ ), .A2(_06766_ ), .A3(_06789_ ), .A4(_06786_ ), .ZN(_07478_ ) );
NOR2_X1 _15481_ ( .A1(_07065_ ), .A2(_07478_ ), .ZN(_07479_ ) );
INV_X1 _15482_ ( .A(_07479_ ), .ZN(_07480_ ) );
NAND3_X1 _15483_ ( .A1(_06766_ ), .A2(_06789_ ), .A3(_07346_ ), .ZN(_07481_ ) );
AOI21_X1 _15484_ ( .A(_07481_ ), .B1(_06784_ ), .B2(_06787_ ), .ZN(_07482_ ) );
AND2_X1 _15485_ ( .A1(_07357_ ), .A2(_06744_ ), .ZN(_07483_ ) );
AND2_X1 _15486_ ( .A1(_07483_ ), .A2(_05186_ ), .ZN(_07484_ ) );
OR2_X1 _15487_ ( .A1(_07482_ ), .A2(_07484_ ), .ZN(_07485_ ) );
OAI21_X1 _15488_ ( .A(_06732_ ), .B1(_07480_ ), .B2(_07485_ ), .ZN(_07486_ ) );
AOI21_X1 _15489_ ( .A(_06857_ ), .B1(_07367_ ), .B2(_07370_ ), .ZN(_07487_ ) );
OAI21_X1 _15490_ ( .A(_07032_ ), .B1(_06971_ ), .B2(_06967_ ), .ZN(_07488_ ) );
OAI21_X1 _15491_ ( .A(_06831_ ), .B1(_06978_ ), .B2(_06972_ ), .ZN(_07489_ ) );
AND3_X1 _15492_ ( .A1(_07488_ ), .A2(_07489_ ), .A3(_06804_ ), .ZN(_07490_ ) );
AND2_X1 _15493_ ( .A1(_06987_ ), .A2(_06969_ ), .ZN(_07491_ ) );
AOI21_X1 _15494_ ( .A(_06984_ ), .B1(_05094_ ), .B2(_06963_ ), .ZN(_07492_ ) );
MUX2_X1 _15495_ ( .A(_07491_ ), .B(_07492_ ), .S(_06869_ ), .Z(_07493_ ) );
AOI211_X1 _15496_ ( .A(_06850_ ), .B(_07490_ ), .C1(_07493_ ), .C2(_06887_ ), .ZN(_07494_ ) );
OAI21_X1 _15497_ ( .A(_06801_ ), .B1(_06975_ ), .B2(_06979_ ), .ZN(_07495_ ) );
OAI21_X1 _15498_ ( .A(_06831_ ), .B1(_07003_ ), .B2(_06976_ ), .ZN(_07496_ ) );
NAND2_X1 _15499_ ( .A1(_07495_ ), .A2(_07496_ ), .ZN(_07497_ ) );
NAND2_X1 _15500_ ( .A1(_07497_ ), .A2(_06914_ ), .ZN(_07498_ ) );
NAND3_X1 _15501_ ( .A1(_07166_ ), .A2(_07167_ ), .A3(_06811_ ), .ZN(_07499_ ) );
AOI21_X1 _15502_ ( .A(_07140_ ), .B1(_07498_ ), .B2(_07499_ ), .ZN(_07500_ ) );
NOR3_X1 _15503_ ( .A1(_07494_ ), .A2(_06905_ ), .A3(_07500_ ), .ZN(_07501_ ) );
OAI21_X1 _15504_ ( .A(_05332_ ), .B1(_07487_ ), .B2(_07501_ ), .ZN(_07502_ ) );
NAND3_X1 _15505_ ( .A1(_07483_ ), .A2(_06854_ ), .A3(_06928_ ), .ZN(_07503_ ) );
AND3_X1 _15506_ ( .A1(_07486_ ), .A2(_07502_ ), .A3(_07503_ ), .ZN(_07504_ ) );
BUF_X4 _15507_ ( .A(_05073_ ), .Z(_07505_ ) );
NAND3_X1 _15508_ ( .A1(_06983_ ), .A2(_07505_ ), .A3(_05080_ ), .ZN(_07506_ ) );
OAI21_X1 _15509_ ( .A(_05323_ ), .B1(_06983_ ), .B2(_05080_ ), .ZN(_07507_ ) );
AND4_X1 _15510_ ( .A1(_07477_ ), .A2(_07504_ ), .A3(_07506_ ), .A4(_07507_ ), .ZN(_07508_ ) );
AOI21_X1 _15511_ ( .A(_06939_ ), .B1(_07476_ ), .B2(_07508_ ), .ZN(_07509_ ) );
NAND2_X1 _15512_ ( .A1(_06623_ ), .A2(_04493_ ), .ZN(_07510_ ) );
AND2_X1 _15513_ ( .A1(_07510_ ), .A2(_05395_ ), .ZN(_07511_ ) );
INV_X1 _15514_ ( .A(_07511_ ), .ZN(_07512_ ) );
NAND2_X1 _15515_ ( .A1(_07512_ ), .A2(_04676_ ), .ZN(_07513_ ) );
AND2_X1 _15516_ ( .A1(_07513_ ), .A2(_05406_ ), .ZN(_07514_ ) );
INV_X1 _15517_ ( .A(_04515_ ), .ZN(_07515_ ) );
NOR2_X1 _15518_ ( .A1(_07514_ ), .A2(_07515_ ), .ZN(_07516_ ) );
INV_X1 _15519_ ( .A(_07516_ ), .ZN(_07517_ ) );
AOI21_X1 _15520_ ( .A(_05374_ ), .B1(_07517_ ), .B2(_05373_ ), .ZN(_07518_ ) );
AOI21_X1 _15521_ ( .A(_07051_ ), .B1(_07518_ ), .B2(_04583_ ), .ZN(_07519_ ) );
OAI21_X1 _15522_ ( .A(_07519_ ), .B1(_04583_ ), .B2(_07518_ ), .ZN(_07520_ ) );
AOI22_X1 _15523_ ( .A1(_04252_ ), .A2(_06949_ ), .B1(\ID_EX_imm [30] ), .B2(_06950_ ), .ZN(_07521_ ) );
AOI21_X1 _15524_ ( .A(_06946_ ), .B1(_07520_ ), .B2(_07521_ ), .ZN(_07522_ ) );
OR2_X1 _15525_ ( .A1(_07522_ ), .A2(_05433_ ), .ZN(_07523_ ) );
OAI22_X1 _15526_ ( .A1(_07509_ ), .A2(_07523_ ), .B1(_05963_ ), .B2(_04130_ ), .ZN(_07524_ ) );
OAI21_X1 _15527_ ( .A(_07450_ ), .B1(_07524_ ), .B2(_06384_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _15528_ ( .A1(_05728_ ), .A2(_05730_ ), .A3(_06467_ ), .ZN(_07525_ ) );
NAND2_X1 _15529_ ( .A1(_05368_ ), .A2(_04879_ ), .ZN(_07526_ ) );
NAND2_X1 _15530_ ( .A1(_07526_ ), .A2(_05342_ ), .ZN(_07527_ ) );
AND2_X1 _15531_ ( .A1(_07527_ ), .A2(_04830_ ), .ZN(_07528_ ) );
OR3_X1 _15532_ ( .A1(_07528_ ), .A2(_04807_ ), .A3(_05337_ ), .ZN(_07529_ ) );
OAI21_X1 _15533_ ( .A(_04807_ ), .B1(_07528_ ), .B2(_05337_ ), .ZN(_07530_ ) );
NAND3_X1 _15534_ ( .A1(_07529_ ), .A2(_06632_ ), .A3(_07530_ ), .ZN(_07531_ ) );
NOR2_X1 _15535_ ( .A1(_05720_ ), .A2(_07195_ ), .ZN(_07532_ ) );
AOI21_X1 _15536_ ( .A(_07532_ ), .B1(\ID_EX_imm [11] ), .B2(_06640_ ), .ZN(_07533_ ) );
AOI21_X1 _15537_ ( .A(_06946_ ), .B1(_07531_ ), .B2(_07533_ ), .ZN(_07534_ ) );
OR2_X1 _15538_ ( .A1(_07534_ ), .A2(_05433_ ), .ZN(_07535_ ) );
OAI211_X1 _15539_ ( .A(_06766_ ), .B(_06789_ ), .C1(_06962_ ), .C2(_07082_ ), .ZN(_07536_ ) );
INV_X1 _15540_ ( .A(_07064_ ), .ZN(_07537_ ) );
NOR2_X1 _15541_ ( .A1(_07536_ ), .A2(_07537_ ), .ZN(_07538_ ) );
NOR3_X1 _15542_ ( .A1(_06877_ ), .A2(_06880_ ), .A3(_06830_ ), .ZN(_07539_ ) );
NOR3_X1 _15543_ ( .A1(_06891_ ), .A2(_06878_ ), .A3(_06800_ ), .ZN(_07540_ ) );
OAI21_X1 _15544_ ( .A(_06886_ ), .B1(_07539_ ), .B2(_07540_ ), .ZN(_07541_ ) );
NAND3_X1 _15545_ ( .A1(_07295_ ), .A2(_07296_ ), .A3(_06803_ ), .ZN(_07542_ ) );
NAND2_X1 _15546_ ( .A1(_07541_ ), .A2(_07542_ ), .ZN(_07543_ ) );
MUX2_X1 _15547_ ( .A(_07072_ ), .B(_07543_ ), .S(_07140_ ), .Z(_07544_ ) );
AND2_X1 _15548_ ( .A1(_07544_ ), .A2(_06857_ ), .ZN(_07545_ ) );
AND3_X1 _15549_ ( .A1(_07079_ ), .A2(_06905_ ), .A3(_07141_ ), .ZN(_07546_ ) );
OR2_X1 _15550_ ( .A1(_07545_ ), .A2(_07546_ ), .ZN(_07547_ ) );
OAI21_X1 _15551_ ( .A(_06959_ ), .B1(_07538_ ), .B2(_07547_ ), .ZN(_07548_ ) );
OAI21_X1 _15552_ ( .A(_07121_ ), .B1(_07545_ ), .B2(_07546_ ), .ZN(_07549_ ) );
NAND3_X1 _15553_ ( .A1(_07102_ ), .A2(_07401_ ), .A3(_07107_ ), .ZN(_07550_ ) );
BUF_X4 _15554_ ( .A(_06887_ ), .Z(_07551_ ) );
NAND4_X1 _15555_ ( .A1(_07093_ ), .A2(_07094_ ), .A3(_06919_ ), .A4(_07551_ ), .ZN(_07552_ ) );
NAND2_X1 _15556_ ( .A1(_07550_ ), .A2(_07552_ ), .ZN(_07553_ ) );
NAND2_X1 _15557_ ( .A1(_07553_ ), .A2(_07309_ ), .ZN(_07554_ ) );
AOI22_X1 _15558_ ( .A1(_05132_ ), .A2(_07410_ ), .B1(_07505_ ), .B2(_06692_ ), .ZN(_07555_ ) );
AND4_X1 _15559_ ( .A1(_07548_ ), .A2(_07549_ ), .A3(_07554_ ), .A4(_07555_ ), .ZN(_07556_ ) );
OAI21_X1 _15560_ ( .A(_05128_ ), .B1(_06679_ ), .B2(_06690_ ), .ZN(_07557_ ) );
OR2_X1 _15561_ ( .A1(_05127_ ), .A2(_04808_ ), .ZN(_07558_ ) );
NAND2_X1 _15562_ ( .A1(_07557_ ), .A2(_07558_ ), .ZN(_07559_ ) );
AOI21_X1 _15563_ ( .A(_06954_ ), .B1(_07559_ ), .B2(_05132_ ), .ZN(_07560_ ) );
OAI21_X1 _15564_ ( .A(_07560_ ), .B1(_05132_ ), .B2(_07559_ ), .ZN(_07561_ ) );
OAI21_X1 _15565_ ( .A(_07153_ ), .B1(_05206_ ), .B2(_04783_ ), .ZN(_07562_ ) );
NAND3_X1 _15566_ ( .A1(_07556_ ), .A2(_07561_ ), .A3(_07562_ ), .ZN(_07563_ ) );
AOI21_X1 _15567_ ( .A(_07535_ ), .B1(_07563_ ), .B2(_06942_ ), .ZN(_07564_ ) );
OAI21_X1 _15568_ ( .A(_07279_ ), .B1(_05714_ ), .B2(_06056_ ), .ZN(_07565_ ) );
OAI21_X1 _15569_ ( .A(_07525_ ), .B1(_07564_ ), .B2(_07565_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
NAND2_X1 _15570_ ( .A1(_05772_ ), .A2(_06441_ ), .ZN(_07566_ ) );
AND2_X1 _15571_ ( .A1(_06960_ ), .A2(_07082_ ), .ZN(_07567_ ) );
OAI21_X1 _15572_ ( .A(_07567_ ), .B1(_06882_ ), .B2(_06799_ ), .ZN(_07568_ ) );
AND2_X1 _15573_ ( .A1(_06961_ ), .A2(_06962_ ), .ZN(_07569_ ) );
INV_X1 _15574_ ( .A(_07569_ ), .ZN(_07570_ ) );
AOI21_X1 _15575_ ( .A(_07537_ ), .B1(_07568_ ), .B2(_07570_ ), .ZN(_07571_ ) );
AND3_X1 _15576_ ( .A1(_07348_ ), .A2(_07349_ ), .A3(_06805_ ), .ZN(_07572_ ) );
NOR3_X1 _15577_ ( .A1(_06996_ ), .A2(_07013_ ), .A3(_06869_ ), .ZN(_07573_ ) );
AND3_X1 _15578_ ( .A1(_04784_ ), .A2(_06862_ ), .A3(_06860_ ), .ZN(_07574_ ) );
NOR3_X1 _15579_ ( .A1(_07574_ ), .A2(_07011_ ), .A3(_06864_ ), .ZN(_07575_ ) );
NOR3_X1 _15580_ ( .A1(_07573_ ), .A2(_07575_ ), .A3(_06805_ ), .ZN(_07576_ ) );
OAI21_X1 _15581_ ( .A(_07096_ ), .B1(_07572_ ), .B2(_07576_ ), .ZN(_07577_ ) );
OAI211_X1 _15582_ ( .A(_07577_ ), .B(_07038_ ), .C1(_06875_ ), .C2(_07139_ ), .ZN(_07578_ ) );
OAI211_X1 _15583_ ( .A(_06906_ ), .B(_06875_ ), .C1(_07146_ ), .C2(_07143_ ), .ZN(_07579_ ) );
NAND2_X1 _15584_ ( .A1(_07578_ ), .A2(_07579_ ), .ZN(_07580_ ) );
OAI21_X1 _15585_ ( .A(_06959_ ), .B1(_07571_ ), .B2(_07580_ ), .ZN(_07581_ ) );
OR3_X1 _15586_ ( .A1(_06679_ ), .A2(_05128_ ), .A3(_06690_ ), .ZN(_07582_ ) );
NAND3_X1 _15587_ ( .A1(_07582_ ), .A2(_06726_ ), .A3(_07557_ ), .ZN(_07583_ ) );
NAND2_X1 _15588_ ( .A1(_07580_ ), .A2(_07121_ ), .ZN(_07584_ ) );
OAI21_X1 _15589_ ( .A(_07153_ ), .B1(_05208_ ), .B2(_02571_ ), .ZN(_07585_ ) );
NOR3_X1 _15590_ ( .A1(_05127_ ), .A2(_04808_ ), .A3(_05074_ ), .ZN(_07586_ ) );
OR3_X1 _15591_ ( .A1(_07156_ ), .A2(_06744_ ), .A3(_06803_ ), .ZN(_07587_ ) );
OR3_X1 _15592_ ( .A1(_07161_ ), .A2(_05147_ ), .A3(_07164_ ), .ZN(_07588_ ) );
AND2_X1 _15593_ ( .A1(_07587_ ), .A2(_07588_ ), .ZN(_07589_ ) );
INV_X1 _15594_ ( .A(_07589_ ), .ZN(_07590_ ) );
AOI221_X4 _15595_ ( .A(_07586_ ), .B1(_05128_ ), .B2(_05330_ ), .C1(_07590_ ), .C2(_07308_ ), .ZN(_07591_ ) );
AND4_X1 _15596_ ( .A1(_07583_ ), .A2(_07584_ ), .A3(_07585_ ), .A4(_07591_ ), .ZN(_07592_ ) );
AOI21_X1 _15597_ ( .A(_06939_ ), .B1(_07581_ ), .B2(_07592_ ), .ZN(_07593_ ) );
NOR2_X1 _15598_ ( .A1(_07527_ ), .A2(_04830_ ), .ZN(_07594_ ) );
NOR3_X1 _15599_ ( .A1(_07528_ ), .A2(_07594_ ), .A3(_07051_ ), .ZN(_07595_ ) );
OAI22_X1 _15600_ ( .A1(_05763_ ), .A2(_07195_ ), .B1(_02572_ ), .B2(_07196_ ), .ZN(_07596_ ) );
OAI21_X1 _15601_ ( .A(_06645_ ), .B1(_07595_ ), .B2(_07596_ ), .ZN(_07597_ ) );
NAND2_X1 _15602_ ( .A1(_07597_ ), .A2(_05963_ ), .ZN(_07598_ ) );
OAI22_X1 _15603_ ( .A1(_07593_ ), .A2(_07598_ ), .B1(_05963_ ), .B2(_05759_ ), .ZN(_07599_ ) );
OAI21_X1 _15604_ ( .A(_07566_ ), .B1(_07599_ ), .B2(_06384_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
NAND2_X1 _15605_ ( .A1(_05783_ ), .A2(_06441_ ), .ZN(_07600_ ) );
AOI22_X1 _15606_ ( .A1(_05788_ ), .A2(_06637_ ), .B1(\ID_EX_imm [9] ), .B2(_06640_ ), .ZN(_07601_ ) );
INV_X1 _15607_ ( .A(_04878_ ), .ZN(_07602_ ) );
AOI21_X1 _15608_ ( .A(_07602_ ), .B1(_05361_ ), .B2(_05366_ ), .ZN(_07603_ ) );
OR3_X1 _15609_ ( .A1(_07603_ ), .A2(_04855_ ), .A3(_05340_ ), .ZN(_07604_ ) );
OAI21_X1 _15610_ ( .A(_04855_ ), .B1(_07603_ ), .B2(_05340_ ), .ZN(_07605_ ) );
NAND3_X1 _15611_ ( .A1(_07604_ ), .A2(_07182_ ), .A3(_07605_ ), .ZN(_07606_ ) );
AOI21_X1 _15612_ ( .A(_06946_ ), .B1(_07601_ ), .B2(_07606_ ), .ZN(_07607_ ) );
OR2_X1 _15613_ ( .A1(_07607_ ), .A2(_05433_ ), .ZN(_07608_ ) );
NAND3_X1 _15614_ ( .A1(_07567_ ), .A2(_06802_ ), .A3(_06807_ ), .ZN(_07609_ ) );
AOI21_X1 _15615_ ( .A(_07537_ ), .B1(_07609_ ), .B2(_07570_ ), .ZN(_07610_ ) );
OR3_X1 _15616_ ( .A1(_07208_ ), .A2(_06854_ ), .A3(_06919_ ), .ZN(_07611_ ) );
OAI21_X1 _15617_ ( .A(_06919_ ), .B1(_07212_ ), .B2(_07213_ ), .ZN(_07612_ ) );
NAND2_X1 _15618_ ( .A1(_07388_ ), .A2(_06805_ ), .ZN(_07613_ ) );
OAI21_X1 _15619_ ( .A(_06869_ ), .B1(_07103_ ), .B2(_06863_ ), .ZN(_07614_ ) );
OAI21_X1 _15620_ ( .A(_06864_ ), .B1(_06877_ ), .B2(_06880_ ), .ZN(_07615_ ) );
NAND3_X1 _15621_ ( .A1(_07614_ ), .A2(_07615_ ), .A3(_06914_ ), .ZN(_07616_ ) );
NAND2_X1 _15622_ ( .A1(_07613_ ), .A2(_07616_ ), .ZN(_07617_ ) );
BUF_X4 _15623_ ( .A(_06902_ ), .Z(_07618_ ) );
OAI211_X1 _15624_ ( .A(_06858_ ), .B(_07612_ ), .C1(_07617_ ), .C2(_07618_ ), .ZN(_07619_ ) );
NAND2_X1 _15625_ ( .A1(_07611_ ), .A2(_07619_ ), .ZN(_07620_ ) );
OAI21_X1 _15626_ ( .A(_06959_ ), .B1(_07610_ ), .B2(_07620_ ), .ZN(_07621_ ) );
AOI21_X1 _15627_ ( .A(_05143_ ), .B1(_06668_ ), .B2(_06678_ ), .ZN(_07622_ ) );
NOR2_X1 _15628_ ( .A1(_07622_ ), .A2(_06688_ ), .ZN(_07623_ ) );
AOI21_X1 _15629_ ( .A(_06954_ ), .B1(_07623_ ), .B2(_05138_ ), .ZN(_07624_ ) );
OAI21_X1 _15630_ ( .A(_07624_ ), .B1(_05138_ ), .B2(_07623_ ), .ZN(_07625_ ) );
AOI21_X1 _15631_ ( .A(_07361_ ), .B1(_07611_ ), .B2(_07619_ ), .ZN(_07626_ ) );
NAND3_X1 _15632_ ( .A1(_07226_ ), .A2(_07401_ ), .A3(_07227_ ), .ZN(_07627_ ) );
NAND3_X1 _15633_ ( .A1(_06916_ ), .A2(_07618_ ), .A3(_07551_ ), .ZN(_07628_ ) );
AOI21_X1 _15634_ ( .A(_07364_ ), .B1(_07627_ ), .B2(_07628_ ), .ZN(_07629_ ) );
NOR3_X1 _15635_ ( .A1(_05136_ ), .A2(_04833_ ), .A3(_07234_ ), .ZN(_07630_ ) );
OAI22_X1 _15636_ ( .A1(_05138_ ), .A2(_05331_ ), .B1(_06686_ ), .B2(_06930_ ), .ZN(_07631_ ) );
NOR4_X1 _15637_ ( .A1(_07626_ ), .A2(_07629_ ), .A3(_07630_ ), .A4(_07631_ ), .ZN(_07632_ ) );
NAND3_X1 _15638_ ( .A1(_07621_ ), .A2(_07625_ ), .A3(_07632_ ), .ZN(_07633_ ) );
AOI21_X1 _15639_ ( .A(_07608_ ), .B1(_07633_ ), .B2(_06942_ ), .ZN(_07634_ ) );
OAI21_X1 _15640_ ( .A(_07279_ ), .B1(_05785_ ), .B2(_06056_ ), .ZN(_07635_ ) );
OAI21_X1 _15641_ ( .A(_07600_ ), .B1(_07634_ ), .B2(_07635_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _15642_ ( .A1(_05803_ ), .A2(_05805_ ), .A3(_06467_ ), .ZN(_07636_ ) );
NOR2_X1 _15643_ ( .A1(_07603_ ), .A2(_07051_ ), .ZN(_07637_ ) );
OAI21_X1 _15644_ ( .A(_07637_ ), .B1(_04878_ ), .B2(_05368_ ), .ZN(_07638_ ) );
AOI22_X1 _15645_ ( .A1(_05810_ ), .A2(_06949_ ), .B1(\ID_EX_imm [8] ), .B2(_06950_ ), .ZN(_07639_ ) );
AOI21_X1 _15646_ ( .A(_06946_ ), .B1(_07638_ ), .B2(_07639_ ), .ZN(_07640_ ) );
OR2_X1 _15647_ ( .A1(_07640_ ), .A2(_05430_ ), .ZN(_07641_ ) );
NOR2_X1 _15648_ ( .A1(_06743_ ), .A2(_06902_ ), .ZN(_07642_ ) );
INV_X1 _15649_ ( .A(_07642_ ), .ZN(_07643_ ) );
NAND4_X1 _15650_ ( .A1(_06766_ ), .A2(_07643_ ), .A3(_06789_ ), .A4(_07291_ ), .ZN(_07644_ ) );
NOR3_X1 _15651_ ( .A1(_07252_ ), .A2(_07140_ ), .A3(_07253_ ), .ZN(_07645_ ) );
OAI21_X1 _15652_ ( .A(_07032_ ), .B1(_07010_ ), .B2(_07018_ ), .ZN(_07646_ ) );
OAI21_X1 _15653_ ( .A(_06820_ ), .B1(_07574_ ), .B2(_07011_ ), .ZN(_07647_ ) );
NAND2_X1 _15654_ ( .A1(_07646_ ), .A2(_07647_ ), .ZN(_07648_ ) );
NAND2_X1 _15655_ ( .A1(_07648_ ), .A2(_06841_ ), .ZN(_07649_ ) );
NAND3_X1 _15656_ ( .A1(_07424_ ), .A2(_06804_ ), .A3(_07425_ ), .ZN(_07650_ ) );
AND3_X1 _15657_ ( .A1(_07649_ ), .A2(_07650_ ), .A3(_06744_ ), .ZN(_07651_ ) );
OAI21_X1 _15658_ ( .A(_06857_ ), .B1(_07645_ ), .B2(_07651_ ), .ZN(_07652_ ) );
NAND4_X1 _15659_ ( .A1(_07255_ ), .A2(_07256_ ), .A3(_06905_ ), .A4(_06874_ ), .ZN(_07653_ ) );
AND2_X1 _15660_ ( .A1(_07652_ ), .A2(_07653_ ), .ZN(_07654_ ) );
AOI21_X1 _15661_ ( .A(_07063_ ), .B1(_07644_ ), .B2(_07654_ ), .ZN(_07655_ ) );
AND3_X1 _15662_ ( .A1(_06668_ ), .A2(_05143_ ), .A3(_06678_ ), .ZN(_07656_ ) );
NOR3_X1 _15663_ ( .A1(_07656_ ), .A2(_07622_ ), .A3(_06954_ ), .ZN(_07657_ ) );
OR2_X1 _15664_ ( .A1(_07654_ ), .A2(_07361_ ), .ZN(_07658_ ) );
NAND2_X1 _15665_ ( .A1(_07268_ ), .A2(_07401_ ), .ZN(_07659_ ) );
OR2_X1 _15666_ ( .A1(_07270_ ), .A2(_06875_ ), .ZN(_07660_ ) );
NAND3_X1 _15667_ ( .A1(_07659_ ), .A2(_07309_ ), .A3(_07660_ ), .ZN(_07661_ ) );
NAND3_X1 _15668_ ( .A1(_05202_ ), .A2(_02498_ ), .A3(_07505_ ), .ZN(_07662_ ) );
AOI21_X1 _15669_ ( .A(_05324_ ), .B1(_05141_ ), .B2(_04856_ ), .ZN(_07663_ ) );
AOI21_X1 _15670_ ( .A(_07663_ ), .B1(_05142_ ), .B2(_06922_ ), .ZN(_07664_ ) );
NAND4_X1 _15671_ ( .A1(_07658_ ), .A2(_07661_ ), .A3(_07662_ ), .A4(_07664_ ), .ZN(_07665_ ) );
OR3_X1 _15672_ ( .A1(_07655_ ), .A2(_07657_ ), .A3(_07665_ ), .ZN(_07666_ ) );
AOI21_X1 _15673_ ( .A(_07641_ ), .B1(_07666_ ), .B2(_06942_ ), .ZN(_07667_ ) );
OAI21_X1 _15674_ ( .A(_07279_ ), .B1(_05809_ ), .B2(_06056_ ), .ZN(_07668_ ) );
OAI21_X1 _15675_ ( .A(_07636_ ), .B1(_07667_ ), .B2(_07668_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
NAND2_X1 _15676_ ( .A1(_05826_ ), .A2(_06441_ ), .ZN(_07669_ ) );
AOI22_X1 _15677_ ( .A1(_05816_ ), .A2(_06637_ ), .B1(\ID_EX_imm [7] ), .B2(_06640_ ), .ZN(_07670_ ) );
AND4_X1 _15678_ ( .A1(_05360_ ), .A2(_05359_ ), .A3(_04952_ ), .A4(_04974_ ), .ZN(_07671_ ) );
OAI21_X1 _15679_ ( .A(_04905_ ), .B1(_07671_ ), .B2(_05365_ ), .ZN(_07672_ ) );
NAND2_X1 _15680_ ( .A1(_04904_ ), .A2(_02670_ ), .ZN(_07673_ ) );
AND2_X1 _15681_ ( .A1(_07672_ ), .A2(_07673_ ), .ZN(_07674_ ) );
XOR2_X1 _15682_ ( .A(_07674_ ), .B(_04929_ ), .Z(_07675_ ) );
OAI21_X1 _15683_ ( .A(_07670_ ), .B1(_07675_ ), .B2(_07051_ ), .ZN(_07676_ ) );
NAND2_X1 _15684_ ( .A1(_07676_ ), .A2(_06645_ ), .ZN(_07677_ ) );
NAND2_X1 _15685_ ( .A1(_07677_ ), .A2(_05605_ ), .ZN(_07678_ ) );
NAND4_X1 _15686_ ( .A1(_06766_ ), .A2(_06962_ ), .A3(_06789_ ), .A4(_07291_ ), .ZN(_07679_ ) );
NAND3_X1 _15687_ ( .A1(_07298_ ), .A2(_07300_ ), .A3(_06919_ ), .ZN(_07680_ ) );
NOR2_X1 _15688_ ( .A1(_07539_ ), .A2(_07540_ ), .ZN(_07681_ ) );
NOR3_X1 _15689_ ( .A1(_07103_ ), .A2(_06863_ ), .A3(_06827_ ), .ZN(_07682_ ) );
NOR3_X1 _15690_ ( .A1(_06861_ ), .A2(_06868_ ), .A3(_06830_ ), .ZN(_07683_ ) );
NOR2_X1 _15691_ ( .A1(_07682_ ), .A2(_07683_ ), .ZN(_07684_ ) );
MUX2_X1 _15692_ ( .A(_07681_ ), .B(_07684_ ), .S(_06872_ ), .Z(_07685_ ) );
OAI211_X1 _15693_ ( .A(_06858_ ), .B(_07680_ ), .C1(_07685_ ), .C2(_07618_ ), .ZN(_07686_ ) );
OAI21_X1 _15694_ ( .A(_07140_ ), .B1(_07292_ ), .B2(_07293_ ), .ZN(_07687_ ) );
OAI211_X1 _15695_ ( .A(_07687_ ), .B(_06906_ ), .C1(_07401_ ), .C2(_07303_ ), .ZN(_07688_ ) );
NAND2_X1 _15696_ ( .A1(_07686_ ), .A2(_07688_ ), .ZN(_07689_ ) );
AOI21_X1 _15697_ ( .A(_07063_ ), .B1(_07679_ ), .B2(_07689_ ), .ZN(_07690_ ) );
AND3_X1 _15698_ ( .A1(_07686_ ), .A2(_07121_ ), .A3(_07688_ ), .ZN(_07691_ ) );
NOR3_X1 _15699_ ( .A1(_07311_ ), .A2(_07618_ ), .A3(_07364_ ), .ZN(_07692_ ) );
NOR3_X1 _15700_ ( .A1(_07690_ ), .A2(_07691_ ), .A3(_07692_ ), .ZN(_07693_ ) );
NAND3_X1 _15701_ ( .A1(_06663_ ), .A2(_06665_ ), .A3(_06667_ ), .ZN(_07694_ ) );
INV_X1 _15702_ ( .A(_06677_ ), .ZN(_07695_ ) );
AOI21_X1 _15703_ ( .A(_05191_ ), .B1(_07694_ ), .B2(_07695_ ), .ZN(_07696_ ) );
OR3_X1 _15704_ ( .A1(_07696_ ), .A2(_05177_ ), .A3(_06669_ ), .ZN(_07697_ ) );
OAI21_X1 _15705_ ( .A(_05177_ ), .B1(_07696_ ), .B2(_06669_ ), .ZN(_07698_ ) );
NAND3_X1 _15706_ ( .A1(_07697_ ), .A2(_07219_ ), .A3(_07698_ ), .ZN(_07699_ ) );
NAND2_X1 _15707_ ( .A1(_05177_ ), .A2(_07410_ ), .ZN(_07700_ ) );
NAND3_X1 _15708_ ( .A1(_06671_ ), .A2(_04906_ ), .A3(_07505_ ), .ZN(_07701_ ) );
OAI21_X1 _15709_ ( .A(_07153_ ), .B1(_06671_ ), .B2(_04906_ ), .ZN(_07702_ ) );
AND3_X1 _15710_ ( .A1(_07700_ ), .A2(_07701_ ), .A3(_07702_ ), .ZN(_07703_ ) );
NAND3_X1 _15711_ ( .A1(_07693_ ), .A2(_07699_ ), .A3(_07703_ ), .ZN(_07704_ ) );
AOI21_X1 _15712_ ( .A(_07678_ ), .B1(_07704_ ), .B2(_06942_ ), .ZN(_07705_ ) );
NAND2_X1 _15713_ ( .A1(_05818_ ), .A2(_05648_ ), .ZN(_07706_ ) );
NAND2_X1 _15714_ ( .A1(_07706_ ), .A2(_06522_ ), .ZN(_07707_ ) );
OAI21_X1 _15715_ ( .A(_07669_ ), .B1(_07705_ ), .B2(_07707_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _15716_ ( .A1(_05847_ ), .A2(_06441_ ), .ZN(_07708_ ) );
OR3_X1 _15717_ ( .A1(_07671_ ), .A2(_04905_ ), .A3(_05365_ ), .ZN(_07709_ ) );
NAND3_X1 _15718_ ( .A1(_07709_ ), .A2(_07672_ ), .A3(_07182_ ), .ZN(_07710_ ) );
AOI22_X1 _15719_ ( .A1(_05837_ ), .A2(_06949_ ), .B1(\ID_EX_imm [6] ), .B2(_06950_ ), .ZN(_07711_ ) );
AOI21_X1 _15720_ ( .A(_06946_ ), .B1(_07710_ ), .B2(_07711_ ), .ZN(_07712_ ) );
OR2_X1 _15721_ ( .A1(_07712_ ), .A2(_05430_ ), .ZN(_07713_ ) );
NAND3_X1 _15722_ ( .A1(_06789_ ), .A2(_06798_ ), .A3(_07346_ ), .ZN(_07714_ ) );
NOR3_X1 _15723_ ( .A1(_07714_ ), .A2(_06807_ ), .A3(_07537_ ), .ZN(_07715_ ) );
AOI21_X1 _15724_ ( .A(_05147_ ), .B1(_07353_ ), .B2(_07354_ ), .ZN(_07716_ ) );
AND4_X1 _15725_ ( .A1(_05147_ ), .A2(_06985_ ), .A3(_06753_ ), .A4(_06826_ ), .ZN(_07717_ ) );
OAI21_X1 _15726_ ( .A(_06906_ ), .B1(_07716_ ), .B2(_07717_ ), .ZN(_07718_ ) );
OAI21_X1 _15727_ ( .A(_06918_ ), .B1(_07350_ ), .B2(_07351_ ), .ZN(_07719_ ) );
OR3_X1 _15728_ ( .A1(_07010_ ), .A2(_07018_ ), .A3(_06801_ ), .ZN(_07720_ ) );
OR3_X1 _15729_ ( .A1(_07017_ ), .A2(_07021_ ), .A3(_06831_ ), .ZN(_07721_ ) );
NAND2_X1 _15730_ ( .A1(_07720_ ), .A2(_07721_ ), .ZN(_07722_ ) );
NAND2_X1 _15731_ ( .A1(_07722_ ), .A2(_06872_ ), .ZN(_07723_ ) );
OAI21_X1 _15732_ ( .A(_06876_ ), .B1(_07573_ ), .B2(_07575_ ), .ZN(_07724_ ) );
NAND3_X1 _15733_ ( .A1(_07723_ ), .A2(_07141_ ), .A3(_07724_ ), .ZN(_07725_ ) );
NAND3_X1 _15734_ ( .A1(_07719_ ), .A2(_07038_ ), .A3(_07725_ ), .ZN(_07726_ ) );
NAND2_X1 _15735_ ( .A1(_07718_ ), .A2(_07726_ ), .ZN(_07727_ ) );
OAI21_X1 _15736_ ( .A(_06732_ ), .B1(_07715_ ), .B2(_07727_ ), .ZN(_07728_ ) );
NAND2_X1 _15737_ ( .A1(_07727_ ), .A2(_07121_ ), .ZN(_07729_ ) );
NAND2_X1 _15738_ ( .A1(_07366_ ), .A2(_07141_ ), .ZN(_07730_ ) );
OAI211_X1 _15739_ ( .A(_07728_ ), .B(_07729_ ), .C1(_07364_ ), .C2(_07730_ ), .ZN(_07731_ ) );
AND3_X1 _15740_ ( .A1(_07694_ ), .A2(_05191_ ), .A3(_07695_ ), .ZN(_07732_ ) );
NOR3_X1 _15741_ ( .A1(_07732_ ), .A2(_07696_ ), .A3(_06954_ ), .ZN(_07733_ ) );
AND2_X1 _15742_ ( .A1(_05182_ ), .A2(_06922_ ), .ZN(_07734_ ) );
NOR3_X1 _15743_ ( .A1(_05181_ ), .A2(_04883_ ), .A3(_07234_ ), .ZN(_07735_ ) );
AOI21_X1 _15744_ ( .A(_05324_ ), .B1(_05181_ ), .B2(_04883_ ), .ZN(_07736_ ) );
OR3_X1 _15745_ ( .A1(_07734_ ), .A2(_07735_ ), .A3(_07736_ ), .ZN(_07737_ ) );
OR3_X1 _15746_ ( .A1(_07731_ ), .A2(_07733_ ), .A3(_07737_ ), .ZN(_07738_ ) );
AOI21_X1 _15747_ ( .A(_07713_ ), .B1(_07738_ ), .B2(_06941_ ), .ZN(_07739_ ) );
OAI21_X1 _15748_ ( .A(_07279_ ), .B1(_05835_ ), .B2(_06056_ ), .ZN(_07740_ ) );
OAI21_X1 _15749_ ( .A(_07708_ ), .B1(_07739_ ), .B2(_07740_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
NAND3_X1 _15750_ ( .A1(_05857_ ), .A2(_05859_ ), .A3(_06467_ ), .ZN(_07741_ ) );
AND4_X1 _15751_ ( .A1(_06806_ ), .A2(_06961_ ), .A3(_06962_ ), .A4(_07291_ ), .ZN(_07742_ ) );
AND2_X1 _15752_ ( .A1(_06852_ ), .A2(_06906_ ), .ZN(_07743_ ) );
NAND3_X1 _15753_ ( .A1(_07614_ ), .A2(_07615_ ), .A3(_06805_ ), .ZN(_07744_ ) );
OAI21_X1 _15754_ ( .A(_06864_ ), .B1(_06861_ ), .B2(_06868_ ), .ZN(_07745_ ) );
OAI21_X1 _15755_ ( .A(_06869_ ), .B1(_06866_ ), .B2(_06908_ ), .ZN(_07746_ ) );
NAND3_X1 _15756_ ( .A1(_07745_ ), .A2(_07746_ ), .A3(_06914_ ), .ZN(_07747_ ) );
AND3_X1 _15757_ ( .A1(_07744_ ), .A2(_07747_ ), .A3(_06874_ ), .ZN(_07748_ ) );
AOI211_X1 _15758_ ( .A(_06905_ ), .B(_07748_ ), .C1(_07392_ ), .C2(_06919_ ), .ZN(_07749_ ) );
OR2_X1 _15759_ ( .A1(_07743_ ), .A2(_07749_ ), .ZN(_07750_ ) );
OAI21_X1 _15760_ ( .A(_06959_ ), .B1(_07742_ ), .B2(_07750_ ), .ZN(_07751_ ) );
NAND3_X1 _15761_ ( .A1(_06663_ ), .A2(_06665_ ), .A3(_05187_ ), .ZN(_07752_ ) );
AND3_X1 _15762_ ( .A1(_07752_ ), .A2(_05173_ ), .A3(_06676_ ), .ZN(_07753_ ) );
AOI21_X1 _15763_ ( .A(_05173_ ), .B1(_07752_ ), .B2(_06676_ ), .ZN(_07754_ ) );
OAI21_X1 _15764_ ( .A(_06726_ ), .B1(_07753_ ), .B2(_07754_ ), .ZN(_07755_ ) );
OAI21_X1 _15765_ ( .A(_06928_ ), .B1(_07743_ ), .B2(_07749_ ), .ZN(_07756_ ) );
OAI21_X1 _15766_ ( .A(_07153_ ), .B1(_05171_ ), .B2(_02598_ ), .ZN(_07757_ ) );
NOR3_X1 _15767_ ( .A1(_06917_ ), .A2(_06918_ ), .A3(_07364_ ), .ZN(_07758_ ) );
AOI221_X4 _15768_ ( .A(_07758_ ), .B1(_05073_ ), .B2(_06673_ ), .C1(_05173_ ), .C2(_05330_ ), .ZN(_07759_ ) );
AND4_X1 _15769_ ( .A1(_07755_ ), .A2(_07756_ ), .A3(_07757_ ), .A4(_07759_ ), .ZN(_07760_ ) );
AOI21_X1 _15770_ ( .A(_06939_ ), .B1(_07751_ ), .B2(_07760_ ), .ZN(_07761_ ) );
AND3_X1 _15771_ ( .A1(_05359_ ), .A2(_05360_ ), .A3(_04952_ ), .ZN(_07762_ ) );
OR3_X1 _15772_ ( .A1(_07762_ ), .A2(_05363_ ), .A3(_04974_ ), .ZN(_07763_ ) );
OAI21_X1 _15773_ ( .A(_04974_ ), .B1(_07762_ ), .B2(_05363_ ), .ZN(_07764_ ) );
NAND3_X1 _15774_ ( .A1(_07763_ ), .A2(_06632_ ), .A3(_07764_ ), .ZN(_07765_ ) );
AOI22_X1 _15775_ ( .A1(_05864_ ), .A2(_06637_ ), .B1(\ID_EX_imm [5] ), .B2(_06640_ ), .ZN(_07766_ ) );
AOI21_X1 _15776_ ( .A(_06647_ ), .B1(_07765_ ), .B2(_07766_ ), .ZN(_07767_ ) );
NOR3_X1 _15777_ ( .A1(_07761_ ), .A2(_05431_ ), .A3(_07767_ ), .ZN(_07768_ ) );
NAND2_X1 _15778_ ( .A1(_05861_ ), .A2(_05648_ ), .ZN(_07769_ ) );
NAND2_X1 _15779_ ( .A1(_07769_ ), .A2(_06522_ ), .ZN(_07770_ ) );
OAI21_X1 _15780_ ( .A(_07741_ ), .B1(_07768_ ), .B2(_07770_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
AND2_X1 _15781_ ( .A1(_05873_ ), .A2(_04018_ ), .ZN(_07771_ ) );
NAND4_X1 _15782_ ( .A1(_06961_ ), .A2(_06808_ ), .A3(_06964_ ), .A4(_07291_ ), .ZN(_07772_ ) );
AND2_X1 _15783_ ( .A1(_06992_ ), .A2(_06905_ ), .ZN(_07773_ ) );
AOI21_X1 _15784_ ( .A(_07140_ ), .B1(_07423_ ), .B2(_07426_ ), .ZN(_07774_ ) );
NOR3_X1 _15785_ ( .A1(_07017_ ), .A2(_07021_ ), .A3(_06827_ ), .ZN(_07775_ ) );
NOR3_X1 _15786_ ( .A1(_07020_ ), .A2(_07034_ ), .A3(_06820_ ), .ZN(_07776_ ) );
NOR2_X1 _15787_ ( .A1(_07775_ ), .A2(_07776_ ), .ZN(_07777_ ) );
MUX2_X1 _15788_ ( .A(_07648_ ), .B(_07777_ ), .S(_06886_ ), .Z(_07778_ ) );
AOI211_X1 _15789_ ( .A(_05192_ ), .B(_07774_ ), .C1(_07141_ ), .C2(_07778_ ), .ZN(_07779_ ) );
NOR2_X1 _15790_ ( .A1(_07773_ ), .A2(_07779_ ), .ZN(_07780_ ) );
AOI21_X1 _15791_ ( .A(_07062_ ), .B1(_07772_ ), .B2(_07780_ ), .ZN(_07781_ ) );
NOR3_X1 _15792_ ( .A1(_07037_ ), .A2(_06919_ ), .A3(_07364_ ), .ZN(_07782_ ) );
NAND2_X1 _15793_ ( .A1(_05187_ ), .A2(_06922_ ), .ZN(_07783_ ) );
NAND3_X1 _15794_ ( .A1(_06906_ ), .A2(_02622_ ), .A3(_05073_ ), .ZN(_07784_ ) );
NAND2_X1 _15795_ ( .A1(_07783_ ), .A2(_07784_ ), .ZN(_07785_ ) );
OR3_X1 _15796_ ( .A1(_07781_ ), .A2(_07782_ ), .A3(_07785_ ), .ZN(_07786_ ) );
AOI21_X1 _15797_ ( .A(_05187_ ), .B1(_06663_ ), .B2(_06665_ ), .ZN(_07787_ ) );
NOR2_X1 _15798_ ( .A1(_07787_ ), .A2(_06727_ ), .ZN(_07788_ ) );
NAND2_X1 _15799_ ( .A1(_07788_ ), .A2(_07752_ ), .ZN(_07789_ ) );
OAI21_X1 _15800_ ( .A(_05323_ ), .B1(_06906_ ), .B2(_02622_ ), .ZN(_07790_ ) );
OAI211_X1 _15801_ ( .A(_07789_ ), .B(_07790_ ), .C1(_07780_ ), .C2(_07361_ ), .ZN(_07791_ ) );
OAI21_X1 _15802_ ( .A(_06940_ ), .B1(_07786_ ), .B2(_07791_ ), .ZN(_07792_ ) );
AOI21_X1 _15803_ ( .A(_04952_ ), .B1(_05359_ ), .B2(_05360_ ), .ZN(_07793_ ) );
NOR3_X1 _15804_ ( .A1(_07762_ ), .A2(_07793_ ), .A3(_07051_ ), .ZN(_07794_ ) );
OAI22_X1 _15805_ ( .A1(_05876_ ), .A2(_07195_ ), .B1(_02600_ ), .B2(_07196_ ), .ZN(_07795_ ) );
OAI21_X1 _15806_ ( .A(_06645_ ), .B1(_07794_ ), .B2(_07795_ ), .ZN(_07796_ ) );
AND2_X1 _15807_ ( .A1(_07796_ ), .A2(_05424_ ), .ZN(_07797_ ) );
AOI21_X1 _15808_ ( .A(_07771_ ), .B1(_07792_ ), .B2(_07797_ ), .ZN(_07798_ ) );
MUX2_X1 _15809_ ( .A(_05887_ ), .B(_07798_ ), .S(_06360_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
AND2_X1 _15810_ ( .A1(_04018_ ), .A2(_05901_ ), .ZN(_07799_ ) );
NAND4_X1 _15811_ ( .A1(_06782_ ), .A2(_06962_ ), .A3(_07082_ ), .A4(_07291_ ), .ZN(_07800_ ) );
OR2_X1 _15812_ ( .A1(_07080_ ), .A2(_06853_ ), .ZN(_07801_ ) );
NAND2_X1 _15813_ ( .A1(_07543_ ), .A2(_06851_ ), .ZN(_07802_ ) );
NOR3_X1 _15814_ ( .A1(_06866_ ), .A2(_06908_ ), .A3(_06827_ ), .ZN(_07803_ ) );
NOR2_X1 _15815_ ( .A1(_06907_ ), .A2(_06911_ ), .ZN(_07804_ ) );
AOI21_X1 _15816_ ( .A(_07803_ ), .B1(_06801_ ), .B2(_07804_ ), .ZN(_07805_ ) );
MUX2_X1 _15817_ ( .A(_07684_ ), .B(_07805_ ), .S(_06886_ ), .Z(_07806_ ) );
OAI211_X1 _15818_ ( .A(_06853_ ), .B(_07802_ ), .C1(_07806_ ), .C2(_06918_ ), .ZN(_07807_ ) );
NAND2_X1 _15819_ ( .A1(_07801_ ), .A2(_07807_ ), .ZN(_07808_ ) );
AOI21_X1 _15820_ ( .A(_07063_ ), .B1(_07800_ ), .B2(_07808_ ), .ZN(_07809_ ) );
AND3_X1 _15821_ ( .A1(_07801_ ), .A2(_06927_ ), .A3(_07807_ ), .ZN(_07810_ ) );
INV_X1 _15822_ ( .A(_05148_ ), .ZN(_07811_ ) );
INV_X1 _15823_ ( .A(_06660_ ), .ZN(_07812_ ) );
AOI21_X1 _15824_ ( .A(_06662_ ), .B1(_07812_ ), .B2(_06658_ ), .ZN(_07813_ ) );
OAI21_X1 _15825_ ( .A(_07811_ ), .B1(_07813_ ), .B2(_06652_ ), .ZN(_07814_ ) );
OAI211_X1 _15826_ ( .A(_05148_ ), .B(_06653_ ), .C1(_06661_ ), .C2(_06662_ ), .ZN(_07815_ ) );
AOI21_X1 _15827_ ( .A(_06727_ ), .B1(_07814_ ), .B2(_07815_ ), .ZN(_07816_ ) );
AND3_X1 _15828_ ( .A1(_06902_ ), .A2(_02752_ ), .A3(_05073_ ), .ZN(_07817_ ) );
NAND3_X1 _15829_ ( .A1(_07095_ ), .A2(_06874_ ), .A3(_07308_ ), .ZN(_07818_ ) );
OAI221_X1 _15830_ ( .A(_07818_ ), .B1(_06664_ ), .B2(_05324_ ), .C1(_07811_ ), .C2(_05331_ ), .ZN(_07819_ ) );
OR4_X1 _15831_ ( .A1(_07810_ ), .A2(_07816_ ), .A3(_07817_ ), .A4(_07819_ ), .ZN(_07820_ ) );
OAI21_X1 _15832_ ( .A(_06940_ ), .B1(_07809_ ), .B2(_07820_ ), .ZN(_07821_ ) );
INV_X1 _15833_ ( .A(_05042_ ), .ZN(_07822_ ) );
AND3_X1 _15834_ ( .A1(_05356_ ), .A2(_07822_ ), .A3(_05358_ ), .ZN(_07823_ ) );
AOI21_X1 _15835_ ( .A(_07822_ ), .B1(_05356_ ), .B2(_05358_ ), .ZN(_07824_ ) );
OR3_X1 _15836_ ( .A1(_07823_ ), .A2(_07824_ ), .A3(_07051_ ), .ZN(_07825_ ) );
AOI22_X1 _15837_ ( .A1(_05904_ ), .A2(_06636_ ), .B1(\ID_EX_imm [3] ), .B2(_06950_ ), .ZN(_07826_ ) );
AOI21_X1 _15838_ ( .A(_06646_ ), .B1(_07825_ ), .B2(_07826_ ), .ZN(_07827_ ) );
NOR2_X1 _15839_ ( .A1(_07827_ ), .A2(_05430_ ), .ZN(_07828_ ) );
AOI21_X1 _15840_ ( .A(_07799_ ), .B1(_07821_ ), .B2(_07828_ ), .ZN(_07829_ ) );
MUX2_X1 _15841_ ( .A(_05900_ ), .B(_07829_ ), .S(_06360_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
NAND2_X1 _15842_ ( .A1(_05919_ ), .A2(_06401_ ), .ZN(_07830_ ) );
OR3_X1 _15843_ ( .A1(_05354_ ), .A2(_05355_ ), .A3(_05021_ ), .ZN(_07831_ ) );
NAND3_X1 _15844_ ( .A1(_07831_ ), .A2(_05356_ ), .A3(_07182_ ), .ZN(_07832_ ) );
AOI22_X1 _15845_ ( .A1(_05921_ ), .A2(_06949_ ), .B1(\ID_EX_imm [2] ), .B2(_06950_ ), .ZN(_07833_ ) );
AOI21_X1 _15846_ ( .A(_06946_ ), .B1(_07832_ ), .B2(_07833_ ), .ZN(_07834_ ) );
OR2_X1 _15847_ ( .A1(_07834_ ), .A2(_05430_ ), .ZN(_07835_ ) );
NOR3_X1 _15848_ ( .A1(_07129_ ), .A2(_07130_ ), .A3(_07537_ ), .ZN(_07836_ ) );
OAI21_X1 _15849_ ( .A(_07618_ ), .B1(_07572_ ), .B2(_07576_ ), .ZN(_07837_ ) );
NOR2_X1 _15850_ ( .A1(_07033_ ), .A2(_07030_ ), .ZN(_07838_ ) );
NOR2_X1 _15851_ ( .A1(_07020_ ), .A2(_07034_ ), .ZN(_07839_ ) );
MUX2_X1 _15852_ ( .A(_07838_ ), .B(_07839_ ), .S(_06882_ ), .Z(_07840_ ) );
MUX2_X1 _15853_ ( .A(_07722_ ), .B(_07840_ ), .S(_07551_ ), .Z(_07841_ ) );
OAI211_X1 _15854_ ( .A(_06858_ ), .B(_07837_ ), .C1(_07841_ ), .C2(_07618_ ), .ZN(_07842_ ) );
NAND2_X1 _15855_ ( .A1(_07148_ ), .A2(_06906_ ), .ZN(_07843_ ) );
NAND2_X1 _15856_ ( .A1(_07842_ ), .A2(_07843_ ), .ZN(_07844_ ) );
OAI21_X1 _15857_ ( .A(_06959_ ), .B1(_07836_ ), .B2(_07844_ ), .ZN(_07845_ ) );
NAND2_X1 _15858_ ( .A1(_07844_ ), .A2(_07121_ ), .ZN(_07846_ ) );
NAND2_X1 _15859_ ( .A1(_07157_ ), .A2(_07309_ ), .ZN(_07847_ ) );
AOI21_X1 _15860_ ( .A(_06727_ ), .B1(_06661_ ), .B2(_06662_ ), .ZN(_07848_ ) );
OAI21_X1 _15861_ ( .A(_07848_ ), .B1(_06662_ ), .B2(_06661_ ), .ZN(_07849_ ) );
OAI21_X1 _15862_ ( .A(_07153_ ), .B1(_06876_ ), .B2(_02774_ ), .ZN(_07850_ ) );
AOI22_X1 _15863_ ( .A1(_05152_ ), .A2(_07410_ ), .B1(_07505_ ), .B2(_06652_ ), .ZN(_07851_ ) );
AND4_X1 _15864_ ( .A1(_07847_ ), .A2(_07849_ ), .A3(_07850_ ), .A4(_07851_ ), .ZN(_07852_ ) );
NAND3_X1 _15865_ ( .A1(_07845_ ), .A2(_07846_ ), .A3(_07852_ ), .ZN(_07853_ ) );
AOI21_X1 _15866_ ( .A(_07835_ ), .B1(_07853_ ), .B2(_06941_ ), .ZN(_07854_ ) );
OAI21_X1 _15867_ ( .A(_07279_ ), .B1(_05426_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07855_ ) );
OAI21_X1 _15868_ ( .A(_07830_ ), .B1(_07854_ ), .B2(_07855_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
OR3_X1 _15869_ ( .A1(_05453_ ), .A2(_05455_ ), .A3(_06359_ ), .ZN(_07856_ ) );
OR3_X1 _15870_ ( .A1(_07516_ ), .A2(_05371_ ), .A3(_04537_ ), .ZN(_07857_ ) );
OAI21_X1 _15871_ ( .A(_04537_ ), .B1(_07516_ ), .B2(_05371_ ), .ZN(_07858_ ) );
AND3_X1 _15872_ ( .A1(_07857_ ), .A2(_07182_ ), .A3(_07858_ ), .ZN(_07859_ ) );
OAI22_X1 _15873_ ( .A1(_05460_ ), .A2(_07195_ ), .B1(_03119_ ), .B2(_07196_ ), .ZN(_07860_ ) );
OAI21_X1 _15874_ ( .A(_06645_ ), .B1(_07859_ ), .B2(_07860_ ), .ZN(_07861_ ) );
NAND2_X1 _15875_ ( .A1(_07861_ ), .A2(_05605_ ), .ZN(_07862_ ) );
OAI21_X1 _15876_ ( .A(_05101_ ), .B1(_07465_ ), .B2(_07468_ ), .ZN(_07863_ ) );
INV_X1 _15877_ ( .A(_07863_ ), .ZN(_07864_ ) );
OAI21_X1 _15878_ ( .A(_05095_ ), .B1(_07864_ ), .B2(_07471_ ), .ZN(_07865_ ) );
OAI211_X1 _15879_ ( .A(_07863_ ), .B(_05096_ ), .C1(_05100_ ), .C2(_05314_ ), .ZN(_07866_ ) );
NAND3_X1 _15880_ ( .A1(_07865_ ), .A2(_07219_ ), .A3(_07866_ ), .ZN(_07867_ ) );
NAND2_X1 _15881_ ( .A1(_05095_ ), .A2(_07410_ ), .ZN(_07868_ ) );
NAND3_X1 _15882_ ( .A1(_05093_ ), .A2(_03118_ ), .A3(_07505_ ), .ZN(_07869_ ) );
OAI21_X1 _15883_ ( .A(_07153_ ), .B1(_05093_ ), .B2(_03118_ ), .ZN(_07870_ ) );
AND3_X1 _15884_ ( .A1(_07868_ ), .A2(_07869_ ), .A3(_07870_ ), .ZN(_07871_ ) );
AND2_X1 _15885_ ( .A1(_07394_ ), .A2(_06853_ ), .ZN(_07872_ ) );
AOI21_X1 _15886_ ( .A(_07872_ ), .B1(_07127_ ), .B2(_06785_ ), .ZN(_07873_ ) );
OAI211_X1 _15887_ ( .A(_06961_ ), .B(_06786_ ), .C1(_06806_ ), .C2(_06808_ ), .ZN(_07874_ ) );
AOI21_X1 _15888_ ( .A(_07063_ ), .B1(_07873_ ), .B2(_07874_ ), .ZN(_07875_ ) );
AOI21_X1 _15889_ ( .A(_07875_ ), .B1(_07121_ ), .B2(_07872_ ), .ZN(_07876_ ) );
OAI21_X1 _15890_ ( .A(_06902_ ), .B1(_06894_ ), .B2(_06901_ ), .ZN(_07877_ ) );
OAI211_X1 _15891_ ( .A(_07074_ ), .B(_06882_ ), .C1(_03063_ ), .C2(_06799_ ), .ZN(_07878_ ) );
NAND2_X1 _15892_ ( .A1(_07073_ ), .A2(_06844_ ), .ZN(_07879_ ) );
OAI211_X1 _15893_ ( .A(_07878_ ), .B(_06887_ ), .C1(_06882_ ), .C2(_07879_ ), .ZN(_07880_ ) );
OAI21_X1 _15894_ ( .A(_06895_ ), .B1(_06832_ ), .B2(_06817_ ), .ZN(_07881_ ) );
OAI21_X1 _15895_ ( .A(_06882_ ), .B1(_06837_ ), .B2(_06833_ ), .ZN(_07882_ ) );
AND2_X1 _15896_ ( .A1(_07881_ ), .A2(_07882_ ), .ZN(_07883_ ) );
OAI211_X1 _15897_ ( .A(_07880_ ), .B(_07096_ ), .C1(_06872_ ), .C2(_07883_ ), .ZN(_07884_ ) );
NAND3_X1 _15898_ ( .A1(_07877_ ), .A2(_07884_ ), .A3(_06854_ ), .ZN(_07885_ ) );
AND2_X1 _15899_ ( .A1(_07885_ ), .A2(_05332_ ), .ZN(_07886_ ) );
OAI21_X1 _15900_ ( .A(_07886_ ), .B1(_06926_ ), .B2(_07402_ ), .ZN(_07887_ ) );
AND2_X1 _15901_ ( .A1(_07876_ ), .A2(_07887_ ), .ZN(_07888_ ) );
NAND3_X1 _15902_ ( .A1(_07867_ ), .A2(_07871_ ), .A3(_07888_ ), .ZN(_07889_ ) );
AOI21_X1 _15903_ ( .A(_07862_ ), .B1(_07889_ ), .B2(_06941_ ), .ZN(_07890_ ) );
OAI21_X1 _15904_ ( .A(_07279_ ), .B1(_05446_ ), .B2(_06056_ ), .ZN(_07891_ ) );
OAI21_X1 _15905_ ( .A(_07856_ ), .B1(_07890_ ), .B2(_07891_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
OR2_X1 _15906_ ( .A1(_05938_ ), .A2(_06349_ ), .ZN(_07892_ ) );
OAI21_X1 _15907_ ( .A(_07182_ ), .B1(_05067_ ), .B2(_04998_ ), .ZN(_07893_ ) );
OAI22_X1 _15908_ ( .A1(_05354_ ), .A2(_07893_ ), .B1(_02705_ ), .B2(_07196_ ), .ZN(_07894_ ) );
AOI21_X1 _15909_ ( .A(_07894_ ), .B1(_05927_ ), .B2(_06637_ ), .ZN(_07895_ ) );
OAI21_X1 _15910_ ( .A(_05605_ ), .B1(_07895_ ), .B2(_06647_ ), .ZN(_07896_ ) );
NAND3_X1 _15911_ ( .A1(_07209_ ), .A2(_06905_ ), .A3(_07214_ ), .ZN(_07897_ ) );
OAI21_X1 _15912_ ( .A(_06869_ ), .B1(_06910_ ), .B2(_06915_ ), .ZN(_07898_ ) );
OAI211_X1 _15913_ ( .A(_07898_ ), .B(_06914_ ), .C1(_07804_ ), .C2(_06895_ ), .ZN(_07899_ ) );
NAND3_X1 _15914_ ( .A1(_07745_ ), .A2(_07746_ ), .A3(_06805_ ), .ZN(_07900_ ) );
NAND3_X1 _15915_ ( .A1(_07899_ ), .A2(_06874_ ), .A3(_07900_ ), .ZN(_07901_ ) );
OAI211_X1 _15916_ ( .A(_06857_ ), .B(_07901_ ), .C1(_07617_ ), .C2(_07141_ ), .ZN(_07902_ ) );
AOI21_X1 _15917_ ( .A(_07361_ ), .B1(_07897_ ), .B2(_07902_ ), .ZN(_07903_ ) );
NAND4_X1 _15918_ ( .A1(_07567_ ), .A2(_06802_ ), .A3(_06808_ ), .A4(_07291_ ), .ZN(_07904_ ) );
NAND3_X1 _15919_ ( .A1(_07904_ ), .A2(_07902_ ), .A3(_07897_ ), .ZN(_07905_ ) );
AOI221_X4 _15920_ ( .A(_07903_ ), .B1(_07224_ ), .B2(_07309_ ), .C1(_07905_ ), .C2(_06732_ ), .ZN(_07906_ ) );
OAI21_X1 _15921_ ( .A(_07219_ ), .B1(_05157_ ), .B2(_06656_ ), .ZN(_07907_ ) );
OR2_X1 _15922_ ( .A1(_07907_ ), .A2(_06660_ ), .ZN(_07908_ ) );
AOI22_X1 _15923_ ( .A1(_05157_ ), .A2(_07410_ ), .B1(_06659_ ), .B2(_07153_ ), .ZN(_07909_ ) );
NAND2_X1 _15924_ ( .A1(_06657_ ), .A2(_07505_ ), .ZN(_07910_ ) );
AND2_X1 _15925_ ( .A1(_07909_ ), .A2(_07910_ ), .ZN(_07911_ ) );
NAND3_X1 _15926_ ( .A1(_07906_ ), .A2(_07908_ ), .A3(_07911_ ), .ZN(_07912_ ) );
AOI21_X1 _15927_ ( .A(_07896_ ), .B1(_07912_ ), .B2(_06941_ ), .ZN(_07913_ ) );
OAI21_X1 _15928_ ( .A(_07279_ ), .B1(_05535_ ), .B2(\ID_EX_pc [1] ), .ZN(_07914_ ) );
OAI21_X1 _15929_ ( .A(_07892_ ), .B1(_07913_ ), .B2(_07914_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
OR2_X1 _15930_ ( .A1(_06544_ ), .A2(_06349_ ), .ZN(_07915_ ) );
OAI21_X1 _15931_ ( .A(_05327_ ), .B1(_05313_ ), .B2(_05085_ ), .ZN(_07916_ ) );
AOI211_X1 _15932_ ( .A(_05312_ ), .B(_07916_ ), .C1(_05316_ ), .C2(_05090_ ), .ZN(_07917_ ) );
AND2_X1 _15933_ ( .A1(_05310_ ), .A2(_07917_ ), .ZN(_07918_ ) );
NAND4_X1 _15934_ ( .A1(_06789_ ), .A2(_06798_ ), .A3(_05171_ ), .A4(_06746_ ), .ZN(_07919_ ) );
NAND3_X1 _15935_ ( .A1(_07254_ ), .A2(_06905_ ), .A3(_07257_ ), .ZN(_07920_ ) );
NAND3_X1 _15936_ ( .A1(_07649_ ), .A2(_07650_ ), .A3(_06851_ ), .ZN(_07921_ ) );
OAI21_X1 _15937_ ( .A(_06831_ ), .B1(_07033_ ), .B2(_07030_ ), .ZN(_07922_ ) );
AOI21_X1 _15938_ ( .A(_07029_ ), .B1(_05158_ ), .B2(_06799_ ), .ZN(_07923_ ) );
OAI21_X1 _15939_ ( .A(_07922_ ), .B1(_07923_ ), .B2(_06864_ ), .ZN(_07924_ ) );
MUX2_X1 _15940_ ( .A(_07924_ ), .B(_07777_ ), .S(_06811_ ), .Z(_07925_ ) );
OAI211_X1 _15941_ ( .A(_06857_ ), .B(_07921_ ), .C1(_07925_ ), .C2(_06918_ ), .ZN(_07926_ ) );
NAND2_X1 _15942_ ( .A1(_07920_ ), .A2(_07926_ ), .ZN(_07927_ ) );
AOI21_X1 _15943_ ( .A(_07062_ ), .B1(_07919_ ), .B2(_07927_ ), .ZN(_07928_ ) );
AND3_X1 _15944_ ( .A1(_07920_ ), .A2(_07926_ ), .A3(_06927_ ), .ZN(_07929_ ) );
AND3_X1 _15945_ ( .A1(_07270_ ), .A2(_06875_ ), .A3(_07309_ ), .ZN(_07930_ ) );
NOR4_X1 _15946_ ( .A1(_07918_ ), .A2(_07928_ ), .A3(_07929_ ), .A4(_07930_ ), .ZN(_07931_ ) );
OAI21_X1 _15947_ ( .A(_06726_ ), .B1(_05161_ ), .B2(_07026_ ), .ZN(_07932_ ) );
OAI21_X1 _15948_ ( .A(_06922_ ), .B1(_05161_ ), .B2(_07026_ ), .ZN(_07933_ ) );
NAND3_X1 _15949_ ( .A1(_06963_ ), .A2(_05044_ ), .A3(_05073_ ), .ZN(_07934_ ) );
OAI21_X1 _15950_ ( .A(_05323_ ), .B1(_06963_ ), .B2(_05044_ ), .ZN(_07935_ ) );
AND3_X1 _15951_ ( .A1(_07933_ ), .A2(_07934_ ), .A3(_07935_ ), .ZN(_07936_ ) );
AND3_X1 _15952_ ( .A1(_07931_ ), .A2(_07932_ ), .A3(_07936_ ), .ZN(_07937_ ) );
NOR2_X1 _15953_ ( .A1(_07937_ ), .A2(_06939_ ), .ZN(_07938_ ) );
NAND3_X1 _15954_ ( .A1(_05310_ ), .A2(_05317_ ), .A3(_06937_ ), .ZN(_07939_ ) );
AOI21_X1 _15955_ ( .A(_06933_ ), .B1(_05067_ ), .B2(_05068_ ), .ZN(_07940_ ) );
AOI221_X4 _15956_ ( .A(_07940_ ), .B1(\ID_EX_imm [0] ), .B2(_06639_ ), .C1(_05965_ ), .C2(_06636_ ), .ZN(_07941_ ) );
AOI21_X1 _15957_ ( .A(_06647_ ), .B1(_07939_ ), .B2(_07941_ ), .ZN(_07942_ ) );
NOR3_X1 _15958_ ( .A1(_07938_ ), .A2(_05431_ ), .A3(_07942_ ), .ZN(_07943_ ) );
OAI21_X1 _15959_ ( .A(_07279_ ), .B1(_05535_ ), .B2(\ID_EX_pc [0] ), .ZN(_07944_ ) );
OAI21_X1 _15960_ ( .A(_07915_ ), .B1(_07943_ ), .B2(_07944_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
NAND2_X1 _15961_ ( .A1(_05754_ ), .A2(_06401_ ), .ZN(_07945_ ) );
NAND3_X1 _15962_ ( .A1(_07513_ ), .A2(_07515_ ), .A3(_05406_ ), .ZN(_07946_ ) );
NAND3_X1 _15963_ ( .A1(_07517_ ), .A2(_06632_ ), .A3(_07946_ ), .ZN(_07947_ ) );
AOI22_X1 _15964_ ( .A1(_05743_ ), .A2(_06636_ ), .B1(\ID_EX_imm [28] ), .B2(_06950_ ), .ZN(_07948_ ) );
AOI21_X1 _15965_ ( .A(_06646_ ), .B1(_07947_ ), .B2(_07948_ ), .ZN(_07949_ ) );
OR2_X1 _15966_ ( .A1(_07949_ ), .A2(_05430_ ), .ZN(_07950_ ) );
OR3_X1 _15967_ ( .A1(_07465_ ), .A2(_05101_ ), .A3(_07468_ ), .ZN(_07951_ ) );
NAND3_X1 _15968_ ( .A1(_07951_ ), .A2(_07219_ ), .A3(_07863_ ), .ZN(_07952_ ) );
AOI21_X1 _15969_ ( .A(_05333_ ), .B1(_07436_ ), .B2(_06906_ ), .ZN(_07953_ ) );
OR3_X1 _15970_ ( .A1(_06975_ ), .A2(_06979_ ), .A3(_06895_ ), .ZN(_07954_ ) );
OR3_X1 _15971_ ( .A1(_06978_ ), .A2(_06972_ ), .A3(_06882_ ), .ZN(_07955_ ) );
AOI21_X1 _15972_ ( .A(_07551_ ), .B1(_07954_ ), .B2(_07955_ ), .ZN(_07956_ ) );
NOR2_X1 _15973_ ( .A1(_06971_ ), .A2(_06967_ ), .ZN(_07957_ ) );
MUX2_X1 _15974_ ( .A(_07957_ ), .B(_07491_ ), .S(_06895_ ), .Z(_07958_ ) );
AOI211_X1 _15975_ ( .A(_07618_ ), .B(_07956_ ), .C1(_07551_ ), .C2(_07958_ ), .ZN(_07959_ ) );
NOR3_X1 _15976_ ( .A1(_07002_ ), .A2(_07008_ ), .A3(_07401_ ), .ZN(_07960_ ) );
OAI21_X1 _15977_ ( .A(_06926_ ), .B1(_07959_ ), .B2(_07960_ ), .ZN(_07961_ ) );
NAND2_X1 _15978_ ( .A1(_07953_ ), .A2(_07961_ ), .ZN(_07962_ ) );
AND3_X1 _15979_ ( .A1(_06990_ ), .A2(_06744_ ), .A3(_06841_ ), .ZN(_07963_ ) );
AND2_X1 _15980_ ( .A1(_07963_ ), .A2(_06853_ ), .ZN(_07964_ ) );
OR3_X1 _15981_ ( .A1(_07065_ ), .A2(_07478_ ), .A3(_07964_ ), .ZN(_07965_ ) );
AND3_X1 _15982_ ( .A1(_06961_ ), .A2(_06807_ ), .A3(_06964_ ), .ZN(_07966_ ) );
OAI21_X1 _15983_ ( .A(_07966_ ), .B1(_07127_ ), .B2(_06786_ ), .ZN(_07967_ ) );
INV_X1 _15984_ ( .A(_07967_ ), .ZN(_07968_ ) );
OAI21_X1 _15985_ ( .A(_06732_ ), .B1(_07965_ ), .B2(_07968_ ), .ZN(_07969_ ) );
NAND3_X1 _15986_ ( .A1(_07963_ ), .A2(_06926_ ), .A3(_07121_ ), .ZN(_07970_ ) );
OAI21_X1 _15987_ ( .A(_07153_ ), .B1(_05099_ ), .B2(_03095_ ), .ZN(_07971_ ) );
AOI22_X1 _15988_ ( .A1(_05101_ ), .A2(_06922_ ), .B1(_07505_ ), .B2(_07471_ ), .ZN(_07972_ ) );
AND4_X1 _15989_ ( .A1(_07969_ ), .A2(_07970_ ), .A3(_07971_ ), .A4(_07972_ ), .ZN(_07973_ ) );
NAND3_X1 _15990_ ( .A1(_07952_ ), .A2(_07962_ ), .A3(_07973_ ), .ZN(_07974_ ) );
AOI21_X1 _15991_ ( .A(_07950_ ), .B1(_07974_ ), .B2(_06941_ ), .ZN(_07975_ ) );
OAI21_X1 _15992_ ( .A(_06360_ ), .B1(_05742_ ), .B2(_05963_ ), .ZN(_07976_ ) );
OAI21_X1 _15993_ ( .A(_07945_ ), .B1(_07975_ ), .B2(_07976_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _15994_ ( .A1(_05960_ ), .A2(_06401_ ), .ZN(_07977_ ) );
NAND3_X1 _15995_ ( .A1(_07512_ ), .A2(_04653_ ), .A3(_04675_ ), .ZN(_07978_ ) );
NAND2_X1 _15996_ ( .A1(_07978_ ), .A2(_05404_ ), .ZN(_07979_ ) );
AND2_X1 _15997_ ( .A1(_07979_ ), .A2(_04606_ ), .ZN(_07980_ ) );
OR3_X1 _15998_ ( .A1(_07980_ ), .A2(_04629_ ), .A3(_05399_ ), .ZN(_07981_ ) );
OAI21_X1 _15999_ ( .A(_04629_ ), .B1(_07980_ ), .B2(_05399_ ), .ZN(_07982_ ) );
AND3_X1 _16000_ ( .A1(_07981_ ), .A2(_07182_ ), .A3(_07982_ ), .ZN(_07983_ ) );
OAI22_X1 _16001_ ( .A1(_05950_ ), .A2(_07195_ ), .B1(_02349_ ), .B2(_07196_ ), .ZN(_07984_ ) );
OAI21_X1 _16002_ ( .A(_06645_ ), .B1(_07983_ ), .B2(_07984_ ), .ZN(_07985_ ) );
NAND2_X1 _16003_ ( .A1(_07985_ ), .A2(_05605_ ), .ZN(_07986_ ) );
AOI21_X1 _16004_ ( .A(_07451_ ), .B1(_07462_ ), .B2(_07464_ ), .ZN(_07987_ ) );
INV_X1 _16005_ ( .A(_07987_ ), .ZN(_07988_ ) );
INV_X1 _16006_ ( .A(_05283_ ), .ZN(_07989_ ) );
AOI21_X1 _16007_ ( .A(_05278_ ), .B1(_07988_ ), .B2(_07989_ ), .ZN(_07990_ ) );
NOR3_X1 _16008_ ( .A1(_07987_ ), .A2(_05305_ ), .A3(_05283_ ), .ZN(_07991_ ) );
OAI21_X1 _16009_ ( .A(_07219_ ), .B1(_07990_ ), .B2(_07991_ ), .ZN(_07992_ ) );
AND2_X1 _16010_ ( .A1(_05278_ ), .A2(_07410_ ), .ZN(_07993_ ) );
NOR3_X1 _16011_ ( .A1(_05277_ ), .A2(_05307_ ), .A3(_07234_ ), .ZN(_07994_ ) );
AOI21_X1 _16012_ ( .A(_06930_ ), .B1(_05277_ ), .B2(_05307_ ), .ZN(_07995_ ) );
NOR3_X1 _16013_ ( .A1(_07993_ ), .A2(_07994_ ), .A3(_07995_ ), .ZN(_00340_ ) );
OAI21_X1 _16014_ ( .A(_06831_ ), .B1(_06896_ ), .B2(_06838_ ), .ZN(_00341_ ) );
OAI21_X1 _16015_ ( .A(_07032_ ), .B1(_06837_ ), .B2(_06833_ ), .ZN(_00342_ ) );
NAND2_X1 _16016_ ( .A1(_00341_ ), .A2(_00342_ ), .ZN(_00343_ ) );
OAI21_X1 _16017_ ( .A(_06875_ ), .B1(_00343_ ), .B2(_07551_ ), .ZN(_00344_ ) );
OR3_X1 _16018_ ( .A1(_06832_ ), .A2(_06817_ ), .A3(_06895_ ), .ZN(_00345_ ) );
OAI211_X1 _16019_ ( .A(_07074_ ), .B(_06895_ ), .C1(_03063_ ), .C2(_06799_ ), .ZN(_00346_ ) );
AOI21_X1 _16020_ ( .A(_06876_ ), .B1(_00345_ ), .B2(_00346_ ), .ZN(_00347_ ) );
OAI21_X1 _16021_ ( .A(_07309_ ), .B1(_00344_ ), .B2(_00347_ ), .ZN(_00348_ ) );
AOI21_X1 _16022_ ( .A(_00348_ ), .B1(_07618_ ), .B2(_07115_ ), .ZN(_00349_ ) );
INV_X1 _16023_ ( .A(_07065_ ), .ZN(_00350_ ) );
INV_X1 _16024_ ( .A(_07478_ ), .ZN(_00351_ ) );
AND2_X1 _16025_ ( .A1(_07079_ ), .A2(_06874_ ), .ZN(_00352_ ) );
NAND2_X1 _16026_ ( .A1(_00352_ ), .A2(_07038_ ), .ZN(_00353_ ) );
OAI211_X1 _16027_ ( .A(_06782_ ), .B(_07082_ ), .C1(_06783_ ), .C2(_06786_ ), .ZN(_00354_ ) );
NAND4_X1 _16028_ ( .A1(_00350_ ), .A2(_00351_ ), .A3(_00353_ ), .A4(_00354_ ), .ZN(_00355_ ) );
NAND2_X1 _16029_ ( .A1(_00355_ ), .A2(_06732_ ), .ZN(_00356_ ) );
OAI21_X1 _16030_ ( .A(_00356_ ), .B1(_07361_ ), .B2(_00353_ ), .ZN(_00357_ ) );
NOR2_X1 _16031_ ( .A1(_07038_ ), .A2(_05333_ ), .ZN(_00358_ ) );
AOI211_X1 _16032_ ( .A(_00349_ ), .B(_00357_ ), .C1(_07553_ ), .C2(_00358_ ), .ZN(_00359_ ) );
NAND3_X1 _16033_ ( .A1(_07992_ ), .A2(_00340_ ), .A3(_00359_ ), .ZN(_00360_ ) );
AOI21_X1 _16034_ ( .A(_07986_ ), .B1(_00360_ ), .B2(_06941_ ), .ZN(_00361_ ) );
OAI21_X1 _16035_ ( .A(_06360_ ), .B1(_05944_ ), .B2(_05963_ ), .ZN(_00362_ ) );
OAI21_X1 _16036_ ( .A(_07977_ ), .B1(_00361_ ), .B2(_00362_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
OAI21_X1 _16037_ ( .A(_06467_ ), .B1(_06571_ ), .B2(_06574_ ), .ZN(_00363_ ) );
AOI21_X1 _16038_ ( .A(_07051_ ), .B1(_07979_ ), .B2(_04606_ ), .ZN(_00364_ ) );
OAI21_X1 _16039_ ( .A(_00364_ ), .B1(_04606_ ), .B2(_07979_ ), .ZN(_00365_ ) );
NAND3_X1 _16040_ ( .A1(_05995_ ), .A2(_05947_ ), .A3(_06637_ ), .ZN(_00366_ ) );
NAND3_X1 _16041_ ( .A1(_06638_ ), .A2(\ID_EX_imm [26] ), .A3(_06635_ ), .ZN(_00367_ ) );
AND3_X1 _16042_ ( .A1(_00365_ ), .A2(_00366_ ), .A3(_00367_ ), .ZN(_00368_ ) );
OAI21_X1 _16043_ ( .A(_05605_ ), .B1(_00368_ ), .B2(_06647_ ), .ZN(_00369_ ) );
NAND3_X1 _16044_ ( .A1(_07462_ ), .A2(_07451_ ), .A3(_07464_ ), .ZN(_00370_ ) );
NAND3_X1 _16045_ ( .A1(_07988_ ), .A2(_07219_ ), .A3(_00370_ ), .ZN(_00371_ ) );
OAI22_X1 _16046_ ( .A1(_07989_ ), .A2(_07234_ ), .B1(_05284_ ), .B2(_06930_ ), .ZN(_00372_ ) );
AOI21_X1 _16047_ ( .A(_00372_ ), .B1(_05285_ ), .B2(_07410_ ), .ZN(_00373_ ) );
OAI21_X1 _16048_ ( .A(_06875_ ), .B1(_07497_ ), .B2(_07551_ ), .ZN(_00374_ ) );
AND3_X1 _16049_ ( .A1(_07488_ ), .A2(_07489_ ), .A3(_06872_ ), .ZN(_00375_ ) );
OAI21_X1 _16050_ ( .A(_07309_ ), .B1(_00374_ ), .B2(_00375_ ), .ZN(_00376_ ) );
AOI21_X1 _16051_ ( .A(_00376_ ), .B1(_07172_ ), .B2(_07618_ ), .ZN(_00377_ ) );
NOR2_X1 _16052_ ( .A1(_07568_ ), .A2(_07128_ ), .ZN(_00378_ ) );
AND4_X1 _16053_ ( .A1(_06808_ ), .A2(_06789_ ), .A3(_06798_ ), .A4(_06786_ ), .ZN(_00379_ ) );
INV_X1 _16054_ ( .A(_00379_ ), .ZN(_00380_ ) );
NOR2_X1 _16055_ ( .A1(_07147_ ), .A2(_06918_ ), .ZN(_00381_ ) );
NAND2_X1 _16056_ ( .A1(_00381_ ), .A2(_06857_ ), .ZN(_00382_ ) );
INV_X1 _16057_ ( .A(_07127_ ), .ZN(_00383_ ) );
OAI211_X1 _16058_ ( .A(_00380_ ), .B(_00382_ ), .C1(_00383_ ), .C2(_06788_ ), .ZN(_00384_ ) );
OAI21_X1 _16059_ ( .A(_06732_ ), .B1(_00378_ ), .B2(_00384_ ), .ZN(_00385_ ) );
OAI21_X1 _16060_ ( .A(_00385_ ), .B1(_07361_ ), .B2(_00382_ ), .ZN(_00386_ ) );
AOI211_X1 _16061_ ( .A(_00377_ ), .B(_00386_ ), .C1(_07590_ ), .C2(_00358_ ), .ZN(_00387_ ) );
NAND3_X1 _16062_ ( .A1(_00371_ ), .A2(_00373_ ), .A3(_00387_ ), .ZN(_00388_ ) );
AOI21_X1 _16063_ ( .A(_00369_ ), .B1(_00388_ ), .B2(_06941_ ), .ZN(_00389_ ) );
OAI21_X1 _16064_ ( .A(_06360_ ), .B1(_05994_ ), .B2(_05963_ ), .ZN(_00390_ ) );
OAI21_X1 _16065_ ( .A(_00363_ ), .B1(_00389_ ), .B2(_00390_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
NAND2_X1 _16066_ ( .A1(_06019_ ), .A2(_06401_ ), .ZN(_00391_ ) );
INV_X1 _16067_ ( .A(_05403_ ), .ZN(_00392_ ) );
INV_X1 _16068_ ( .A(_04675_ ), .ZN(_00393_ ) );
OAI21_X1 _16069_ ( .A(_00392_ ), .B1(_07511_ ), .B2(_00393_ ), .ZN(_00394_ ) );
AND2_X1 _16070_ ( .A1(_00394_ ), .A2(_04653_ ), .ZN(_00395_ ) );
OAI21_X1 _16071_ ( .A(_06631_ ), .B1(_00394_ ), .B2(_04653_ ), .ZN(_00396_ ) );
OR2_X1 _16072_ ( .A1(_00395_ ), .A2(_00396_ ), .ZN(_00397_ ) );
AOI22_X1 _16073_ ( .A1(_06010_ ), .A2(_06636_ ), .B1(\ID_EX_imm [25] ), .B2(_06950_ ), .ZN(_00398_ ) );
AOI21_X1 _16074_ ( .A(_06646_ ), .B1(_00397_ ), .B2(_00398_ ), .ZN(_00399_ ) );
OR2_X1 _16075_ ( .A1(_00399_ ), .A2(_05430_ ), .ZN(_00400_ ) );
INV_X1 _16076_ ( .A(_05294_ ), .ZN(_00401_ ) );
AOI21_X1 _16077_ ( .A(_00401_ ), .B1(_07453_ ), .B2(_07459_ ), .ZN(_00402_ ) );
OR3_X1 _16078_ ( .A1(_00402_ ), .A2(_05292_ ), .A3(_05300_ ), .ZN(_00403_ ) );
OAI21_X1 _16079_ ( .A(_05300_ ), .B1(_00402_ ), .B2(_05292_ ), .ZN(_00404_ ) );
AND3_X1 _16080_ ( .A1(_00403_ ), .A2(_06726_ ), .A3(_00404_ ), .ZN(_00405_ ) );
AOI22_X1 _16081_ ( .A1(_05300_ ), .A2(_07410_ ), .B1(_07463_ ), .B2(_05323_ ), .ZN(_00406_ ) );
NAND3_X1 _16082_ ( .A1(_06774_ ), .A2(_03039_ ), .A3(_07505_ ), .ZN(_00407_ ) );
NAND2_X1 _16083_ ( .A1(_00406_ ), .A2(_00407_ ), .ZN(_00408_ ) );
NOR2_X1 _16084_ ( .A1(_07208_ ), .A2(_06918_ ), .ZN(_00409_ ) );
AND3_X1 _16085_ ( .A1(_00409_ ), .A2(_07038_ ), .A3(_06927_ ), .ZN(_00410_ ) );
NAND2_X1 _16086_ ( .A1(_00409_ ), .A2(_07038_ ), .ZN(_00411_ ) );
OAI211_X1 _16087_ ( .A(_07479_ ), .B(_00411_ ), .C1(_07609_ ), .C2(_07128_ ), .ZN(_00412_ ) );
AOI21_X1 _16088_ ( .A(_00410_ ), .B1(_00412_ ), .B2(_06732_ ), .ZN(_00413_ ) );
NAND2_X1 _16089_ ( .A1(_07228_ ), .A2(_07401_ ), .ZN(_00414_ ) );
OAI211_X1 _16090_ ( .A(_00414_ ), .B(_00358_ ), .C1(_07401_ ), .C2(_07223_ ), .ZN(_00415_ ) );
AND3_X1 _16091_ ( .A1(_06897_ ), .A2(_06900_ ), .A3(_06805_ ), .ZN(_00416_ ) );
AOI21_X1 _16092_ ( .A(_00416_ ), .B1(_07883_ ), .B2(_07551_ ), .ZN(_00417_ ) );
MUX2_X1 _16093_ ( .A(_00417_ ), .B(_07231_ ), .S(_06919_ ), .Z(_00418_ ) );
OAI211_X1 _16094_ ( .A(_00413_ ), .B(_00415_ ), .C1(_07364_ ), .C2(_00418_ ), .ZN(_00419_ ) );
OR3_X1 _16095_ ( .A1(_00405_ ), .A2(_00408_ ), .A3(_00419_ ), .ZN(_00420_ ) );
AOI21_X1 _16096_ ( .A(_00400_ ), .B1(_00420_ ), .B2(_06941_ ), .ZN(_00421_ ) );
OAI21_X1 _16097_ ( .A(_06360_ ), .B1(_06007_ ), .B2(_05963_ ), .ZN(_00422_ ) );
OAI21_X1 _16098_ ( .A(_00391_ ), .B1(_00421_ ), .B2(_00422_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND3_X1 _16099_ ( .A1(_06027_ ), .A2(_06033_ ), .A3(_06467_ ), .ZN(_00423_ ) );
OAI21_X1 _16100_ ( .A(_07182_ ), .B1(_07511_ ), .B2(_00393_ ), .ZN(_00424_ ) );
AOI21_X1 _16101_ ( .A(_00424_ ), .B1(_00393_ ), .B2(_07511_ ), .ZN(_00425_ ) );
AND2_X1 _16102_ ( .A1(_06023_ ), .A2(_06949_ ), .ZN(_00426_ ) );
AND3_X1 _16103_ ( .A1(_06638_ ), .A2(\ID_EX_imm [24] ), .A3(_06635_ ), .ZN(_00427_ ) );
NOR3_X1 _16104_ ( .A1(_00425_ ), .A2(_00426_ ), .A3(_00427_ ), .ZN(_00428_ ) );
OAI21_X1 _16105_ ( .A(_05605_ ), .B1(_00428_ ), .B2(_06647_ ), .ZN(_00429_ ) );
NOR2_X1 _16106_ ( .A1(_00402_ ), .A2(_06954_ ), .ZN(_00430_ ) );
OAI21_X1 _16107_ ( .A(_00430_ ), .B1(_05294_ ), .B2(_07461_ ), .ZN(_00431_ ) );
AND4_X1 _16108_ ( .A1(_07643_ ), .A2(_06789_ ), .A3(_06798_ ), .A4(_06786_ ), .ZN(_00432_ ) );
AND3_X1 _16109_ ( .A1(_07255_ ), .A2(_07256_ ), .A3(_07096_ ), .ZN(_00433_ ) );
AND2_X1 _16110_ ( .A1(_00433_ ), .A2(_06858_ ), .ZN(_00434_ ) );
OR2_X1 _16111_ ( .A1(_00432_ ), .A2(_00434_ ), .ZN(_00435_ ) );
OAI21_X1 _16112_ ( .A(_06959_ ), .B1(_00435_ ), .B2(_07065_ ), .ZN(_00436_ ) );
NAND3_X1 _16113_ ( .A1(_00433_ ), .A2(_06926_ ), .A3(_06928_ ), .ZN(_00437_ ) );
OR3_X1 _16114_ ( .A1(_07263_ ), .A2(_07264_ ), .A3(_06875_ ), .ZN(_00438_ ) );
AND3_X1 _16115_ ( .A1(_07954_ ), .A2(_07955_ ), .A3(_06872_ ), .ZN(_00439_ ) );
AOI21_X1 _16116_ ( .A(_07551_ ), .B1(_07004_ ), .B2(_07007_ ), .ZN(_00440_ ) );
OAI21_X1 _16117_ ( .A(_07401_ ), .B1(_00439_ ), .B2(_00440_ ), .ZN(_00441_ ) );
NAND3_X1 _16118_ ( .A1(_00438_ ), .A2(_07309_ ), .A3(_00441_ ), .ZN(_00442_ ) );
NAND2_X1 _16119_ ( .A1(_00437_ ), .A2(_00442_ ), .ZN(_00443_ ) );
AND3_X1 _16120_ ( .A1(_07659_ ), .A2(_07660_ ), .A3(_00358_ ), .ZN(_00444_ ) );
NOR3_X1 _16121_ ( .A1(_05290_ ), .A2(_05291_ ), .A3(_07234_ ), .ZN(_00445_ ) );
OAI22_X1 _16122_ ( .A1(_00401_ ), .A2(_05331_ ), .B1(_05293_ ), .B2(_06930_ ), .ZN(_00446_ ) );
NOR4_X1 _16123_ ( .A1(_00443_ ), .A2(_00444_ ), .A3(_00445_ ), .A4(_00446_ ), .ZN(_00447_ ) );
NAND3_X1 _16124_ ( .A1(_00431_ ), .A2(_00436_ ), .A3(_00447_ ), .ZN(_00448_ ) );
AOI21_X1 _16125_ ( .A(_00429_ ), .B1(_00448_ ), .B2(_06941_ ), .ZN(_00449_ ) );
NAND2_X1 _16126_ ( .A1(_06025_ ), .A2(_05648_ ), .ZN(_00450_ ) );
NAND2_X1 _16127_ ( .A1(_00450_ ), .A2(_06522_ ), .ZN(_00451_ ) );
OAI21_X1 _16128_ ( .A(_00423_ ), .B1(_00449_ ), .B2(_00451_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
OR2_X1 _16129_ ( .A1(_06599_ ), .A2(_06349_ ), .ZN(_00452_ ) );
NOR4_X1 _16130_ ( .A1(_06625_ ), .A2(_06626_ ), .A3(_05389_ ), .A4(_05390_ ), .ZN(_00453_ ) );
OAI21_X1 _16131_ ( .A(_04419_ ), .B1(_00453_ ), .B2(_05393_ ), .ZN(_00454_ ) );
NAND2_X1 _16132_ ( .A1(_04418_ ), .A2(_02373_ ), .ZN(_00455_ ) );
AND2_X1 _16133_ ( .A1(_00454_ ), .A2(_00455_ ), .ZN(_00456_ ) );
XNOR2_X1 _16134_ ( .A(_00456_ ), .B(_04442_ ), .ZN(_00457_ ) );
NAND2_X1 _16135_ ( .A1(_00457_ ), .A2(_06632_ ), .ZN(_00458_ ) );
AOI22_X1 _16136_ ( .A1(_06042_ ), .A2(_06637_ ), .B1(\ID_EX_imm [23] ), .B2(_06640_ ), .ZN(_00459_ ) );
AOI21_X1 _16137_ ( .A(_06647_ ), .B1(_00458_ ), .B2(_00459_ ), .ZN(_00460_ ) );
INV_X1 _16138_ ( .A(_05234_ ), .ZN(_00461_ ) );
NAND2_X1 _16139_ ( .A1(_06957_ ), .A2(_07452_ ), .ZN(_00462_ ) );
AOI21_X1 _16140_ ( .A(_06923_ ), .B1(_05243_ ), .B2(_06722_ ), .ZN(_00463_ ) );
AOI21_X1 _16141_ ( .A(_00461_ ), .B1(_00462_ ), .B2(_00463_ ), .ZN(_00464_ ) );
OR3_X1 _16142_ ( .A1(_00464_ ), .A2(_05230_ ), .A3(_07457_ ), .ZN(_00465_ ) );
OAI21_X1 _16143_ ( .A(_05230_ ), .B1(_00464_ ), .B2(_07457_ ), .ZN(_00466_ ) );
NAND3_X1 _16144_ ( .A1(_00465_ ), .A2(_07219_ ), .A3(_00466_ ), .ZN(_00467_ ) );
OAI21_X1 _16145_ ( .A(_07687_ ), .B1(_06874_ ), .B2(_07303_ ), .ZN(_00468_ ) );
NAND2_X1 _16146_ ( .A1(_00468_ ), .A2(_07038_ ), .ZN(_00469_ ) );
AOI21_X1 _16147_ ( .A(_07062_ ), .B1(_07479_ ), .B2(_00469_ ), .ZN(_00470_ ) );
AND3_X1 _16148_ ( .A1(_07313_ ), .A2(_07314_ ), .A3(_06851_ ), .ZN(_00471_ ) );
NAND2_X1 _16149_ ( .A1(_07111_ ), .A2(_06811_ ), .ZN(_00472_ ) );
NAND2_X1 _16150_ ( .A1(_00343_ ), .A2(_06841_ ), .ZN(_00473_ ) );
AND3_X1 _16151_ ( .A1(_00472_ ), .A2(_07140_ ), .A3(_00473_ ), .ZN(_00474_ ) );
OAI21_X1 _16152_ ( .A(_06857_ ), .B1(_00471_ ), .B2(_00474_ ), .ZN(_00475_ ) );
OR3_X1 _16153_ ( .A1(_07311_ ), .A2(_06853_ ), .A3(_06851_ ), .ZN(_00476_ ) );
AOI21_X1 _16154_ ( .A(_05333_ ), .B1(_00475_ ), .B2(_00476_ ), .ZN(_00477_ ) );
AND3_X1 _16155_ ( .A1(_00468_ ), .A2(_06857_ ), .A3(_06927_ ), .ZN(_00478_ ) );
OR3_X1 _16156_ ( .A1(_00470_ ), .A2(_00477_ ), .A3(_00478_ ), .ZN(_00479_ ) );
AND2_X1 _16157_ ( .A1(_05230_ ), .A2(_06922_ ), .ZN(_00480_ ) );
NOR3_X1 _16158_ ( .A1(_05229_ ), .A2(_04420_ ), .A3(_07234_ ), .ZN(_00481_ ) );
AOI21_X1 _16159_ ( .A(_06930_ ), .B1(_05229_ ), .B2(_04420_ ), .ZN(_00482_ ) );
NOR4_X1 _16160_ ( .A1(_00479_ ), .A2(_00480_ ), .A3(_00481_ ), .A4(_00482_ ), .ZN(_00483_ ) );
AOI21_X1 _16161_ ( .A(_06939_ ), .B1(_00467_ ), .B2(_00483_ ), .ZN(_00484_ ) );
NOR3_X1 _16162_ ( .A1(_00460_ ), .A2(_00484_ ), .A3(_05431_ ), .ZN(_00485_ ) );
NAND2_X1 _16163_ ( .A1(_06045_ ), .A2(_05648_ ), .ZN(_00486_ ) );
NAND2_X1 _16164_ ( .A1(_00486_ ), .A2(_06522_ ), .ZN(_00487_ ) );
OAI21_X1 _16165_ ( .A(_00452_ ), .B1(_00485_ ), .B2(_00487_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
OR3_X1 _16166_ ( .A1(_00453_ ), .A2(_04419_ ), .A3(_05393_ ), .ZN(_00488_ ) );
NAND3_X1 _16167_ ( .A1(_00488_ ), .A2(_07182_ ), .A3(_00454_ ), .ZN(_00489_ ) );
AOI22_X1 _16168_ ( .A1(_06068_ ), .A2(_06636_ ), .B1(\ID_EX_imm [22] ), .B2(_06639_ ), .ZN(_00490_ ) );
AOI21_X1 _16169_ ( .A(_06646_ ), .B1(_00489_ ), .B2(_00490_ ), .ZN(_00491_ ) );
AND3_X1 _16170_ ( .A1(_00462_ ), .A2(_00461_ ), .A3(_00463_ ), .ZN(_00492_ ) );
OR3_X1 _16171_ ( .A1(_00492_ ), .A2(_00464_ ), .A3(_06727_ ), .ZN(_00493_ ) );
OR2_X1 _16172_ ( .A1(_07716_ ), .A2(_07717_ ), .ZN(_00494_ ) );
AND2_X1 _16173_ ( .A1(_00494_ ), .A2(_05186_ ), .ZN(_00495_ ) );
AOI22_X1 _16174_ ( .A1(_00495_ ), .A2(_06928_ ), .B1(_07505_ ), .B2(_07457_ ), .ZN(_00496_ ) );
AND4_X1 _16175_ ( .A1(_06808_ ), .A2(_06782_ ), .A3(_06786_ ), .A4(_07346_ ), .ZN(_00497_ ) );
OR3_X1 _16176_ ( .A1(_00497_ ), .A2(_07065_ ), .A3(_00495_ ), .ZN(_00498_ ) );
NAND2_X1 _16177_ ( .A1(_00498_ ), .A2(_06732_ ), .ZN(_00499_ ) );
AOI21_X1 _16178_ ( .A(_05333_ ), .B1(_07730_ ), .B2(_06905_ ), .ZN(_00500_ ) );
NOR3_X1 _16179_ ( .A1(_07368_ ), .A2(_07369_ ), .A3(_06874_ ), .ZN(_00501_ ) );
AOI21_X1 _16180_ ( .A(_06851_ ), .B1(_07498_ ), .B2(_07499_ ), .ZN(_00502_ ) );
OAI21_X1 _16181_ ( .A(_06857_ ), .B1(_00501_ ), .B2(_00502_ ), .ZN(_00503_ ) );
NAND2_X1 _16182_ ( .A1(_00500_ ), .A2(_00503_ ), .ZN(_00504_ ) );
NAND2_X1 _16183_ ( .A1(_05234_ ), .A2(_06922_ ), .ZN(_00505_ ) );
OAI21_X1 _16184_ ( .A(_05323_ ), .B1(_05233_ ), .B2(_02373_ ), .ZN(_00506_ ) );
AND4_X1 _16185_ ( .A1(_00499_ ), .A2(_00504_ ), .A3(_00505_ ), .A4(_00506_ ), .ZN(_00507_ ) );
NAND3_X1 _16186_ ( .A1(_00493_ ), .A2(_00496_ ), .A3(_00507_ ), .ZN(_00508_ ) );
AOI211_X1 _16187_ ( .A(_05430_ ), .B(_00491_ ), .C1(_00508_ ), .C2(_06940_ ), .ZN(_00509_ ) );
AND2_X1 _16188_ ( .A1(_06066_ ), .A2(_05430_ ), .ZN(_00510_ ) );
OR3_X1 _16189_ ( .A1(_00509_ ), .A2(_06353_ ), .A3(_00510_ ), .ZN(_00511_ ) );
NAND2_X1 _16190_ ( .A1(_06065_ ), .A2(_06354_ ), .ZN(_00512_ ) );
NAND2_X1 _16191_ ( .A1(_00511_ ), .A2(_00512_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
NAND2_X1 _16192_ ( .A1(_06104_ ), .A2(_06401_ ), .ZN(_00513_ ) );
AND2_X1 _16193_ ( .A1(_06983_ ), .A2(_05080_ ), .ZN(_00514_ ) );
OR3_X1 _16194_ ( .A1(_07475_ ), .A2(_05089_ ), .A3(_00514_ ), .ZN(_00515_ ) );
OAI21_X1 _16195_ ( .A(_05089_ ), .B1(_07475_ ), .B2(_00514_ ), .ZN(_00516_ ) );
NAND3_X1 _16196_ ( .A1(_00515_ ), .A2(_07219_ ), .A3(_00516_ ), .ZN(_00517_ ) );
NAND2_X1 _16197_ ( .A1(_06746_ ), .A2(_03150_ ), .ZN(_00518_ ) );
AOI21_X1 _16198_ ( .A(_07063_ ), .B1(_06784_ ), .B2(_00518_ ), .ZN(_00519_ ) );
NAND3_X1 _16199_ ( .A1(_00472_ ), .A2(_07618_ ), .A3(_00473_ ), .ZN(_00520_ ) );
NAND3_X1 _16200_ ( .A1(_00345_ ), .A2(_06876_ ), .A3(_00346_ ), .ZN(_00521_ ) );
OAI211_X1 _16201_ ( .A(_06895_ ), .B(_06845_ ), .C1(_06963_ ), .C2(_03150_ ), .ZN(_00522_ ) );
OAI211_X1 _16202_ ( .A(_07551_ ), .B(_00522_ ), .C1(_07879_ ), .C2(_06895_ ), .ZN(_00523_ ) );
NAND3_X1 _16203_ ( .A1(_00521_ ), .A2(_00523_ ), .A3(_07401_ ), .ZN(_00524_ ) );
AOI21_X1 _16204_ ( .A(_07364_ ), .B1(_00520_ ), .B2(_00524_ ), .ZN(_00525_ ) );
AND3_X1 _16205_ ( .A1(_06746_ ), .A2(_03150_ ), .A3(_06927_ ), .ZN(_00526_ ) );
AOI221_X4 _16206_ ( .A(_00526_ ), .B1(_05086_ ), .B2(_05323_ ), .C1(_05089_ ), .C2(_05330_ ), .ZN(_00527_ ) );
OAI21_X1 _16207_ ( .A(_00358_ ), .B1(_07312_ ), .B2(_07315_ ), .ZN(_00528_ ) );
OR2_X1 _16208_ ( .A1(_05087_ ), .A2(_07234_ ), .ZN(_00529_ ) );
NAND3_X1 _16209_ ( .A1(_00527_ ), .A2(_00528_ ), .A3(_00529_ ), .ZN(_00530_ ) );
NOR3_X1 _16210_ ( .A1(_00519_ ), .A2(_00525_ ), .A3(_00530_ ), .ZN(_00531_ ) );
AOI21_X1 _16211_ ( .A(_06939_ ), .B1(_00517_ ), .B2(_00531_ ), .ZN(_00532_ ) );
AOI21_X1 _16212_ ( .A(_05408_ ), .B1(_07518_ ), .B2(_04583_ ), .ZN(_00533_ ) );
XNOR2_X1 _16213_ ( .A(_00533_ ), .B(_04560_ ), .ZN(_00534_ ) );
AOI22_X1 _16214_ ( .A1(_00534_ ), .A2(_06632_ ), .B1(\ID_EX_imm [31] ), .B2(_06640_ ), .ZN(_00535_ ) );
OR2_X1 _16215_ ( .A1(_06097_ ), .A2(_07195_ ), .ZN(_00536_ ) );
AOI21_X1 _16216_ ( .A(_06647_ ), .B1(_00535_ ), .B2(_00536_ ), .ZN(_00537_ ) );
NOR3_X1 _16217_ ( .A1(_00532_ ), .A2(_00537_ ), .A3(_05431_ ), .ZN(_00538_ ) );
OAI21_X1 _16218_ ( .A(_06360_ ), .B1(_06109_ ), .B2(_05963_ ), .ZN(_00539_ ) );
OAI21_X1 _16219_ ( .A(_00513_ ), .B1(_00538_ ), .B2(_00539_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
AND3_X1 _16220_ ( .A1(_04024_ ), .A2(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .A3(_03221_ ), .ZN(\myexu.rst_logic_$_OR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__B_Y ) );
AND3_X1 _16221_ ( .A1(\myexu.state_$_ANDNOT__B_Y ), .A2(_03239_ ), .A3(_04029_ ), .ZN(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ) );
AOI21_X1 _16222_ ( .A(_02222_ ), .B1(_02160_ ), .B2(_02229_ ), .ZN(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16223_ ( .A(IDU_ready_IFU ), .ZN(_00540_ ) );
NAND2_X1 _16224_ ( .A1(_00540_ ), .A2(IDU_valid_EXU ), .ZN(_00541_ ) );
OAI21_X1 _16225_ ( .A(_00541_ ), .B1(_03389_ ), .B2(_03447_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16226_ ( .A1(_03388_ ), .A2(_03447_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16227_ ( .A1(_03388_ ), .A2(_03447_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16228_ ( .A(_03443_ ), .ZN(_00542_ ) );
NOR4_X1 _16229_ ( .A1(_03388_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03223_ ), .A4(_00542_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16230_ ( .A1(_03788_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03223_ ), .A4(_03442_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16231_ ( .A(_03971_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16232_ ( .A(_00541_ ), .B1(_00542_ ), .B2(_00540_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16233_ ( .A1(_03443_ ), .A2(_00540_ ), .B1(_06134_ ), .B2(_04014_ ), .ZN(_00543_ ) );
INV_X1 _16234_ ( .A(loaduse_clear ), .ZN(_00544_ ) );
AOI221_X4 _16235_ ( .A(_00543_ ), .B1(\myidu.state [2] ), .B2(_00544_ ), .C1(_03387_ ), .C2(_03971_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
OR3_X1 _16236_ ( .A1(_03223_ ), .A2(_04014_ ), .A3(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_00545_ ) );
NAND3_X1 _16237_ ( .A1(_03452_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_00546_ ) );
AOI21_X1 _16238_ ( .A(_03498_ ), .B1(_03514_ ), .B2(_03218_ ), .ZN(_00547_ ) );
AND4_X1 _16239_ ( .A1(_03523_ ), .A2(_03473_ ), .A3(_03333_ ), .A4(_03522_ ), .ZN(_00548_ ) );
AOI21_X1 _16240_ ( .A(_03506_ ), .B1(_00548_ ), .B2(_03381_ ), .ZN(_00549_ ) );
OR2_X1 _16241_ ( .A1(_00547_ ), .A2(_00549_ ), .ZN(_00550_ ) );
NAND3_X1 _16242_ ( .A1(_03443_ ), .A2(IDU_ready_IFU ), .A3(_03222_ ), .ZN(_00551_ ) );
OAI211_X1 _16243_ ( .A(_00545_ ), .B(_00546_ ), .C1(_00550_ ), .C2(_00551_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16244_ ( .A(_03452_ ), .B(_04027_ ), .C1(_03443_ ), .C2(_00540_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _16245_ ( .A(_03444_ ), .B(_03452_ ), .C1(_00549_ ), .C2(_00547_ ), .ZN(_00552_ ) );
NAND3_X1 _16246_ ( .A1(_03452_ ), .A2(\myidu.state [2] ), .A3(_00544_ ), .ZN(_00553_ ) );
NAND2_X1 _16247_ ( .A1(_00552_ ), .A2(_00553_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16248_ ( .A1(_03440_ ), .A2(IDU_ready_IFU ), .ZN(_00554_ ) );
OAI21_X1 _16249_ ( .A(_01586_ ), .B1(_03440_ ), .B2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00555_ ) );
INV_X1 _16250_ ( .A(\myifu.state [0] ), .ZN(_00556_ ) );
AOI211_X1 _16251_ ( .A(_00554_ ), .B(_00555_ ), .C1(_00556_ ), .C2(_03440_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
CLKBUF_X2 _16252_ ( .A(_06207_ ), .Z(_00557_ ) );
OR3_X1 _16253_ ( .A1(_02055_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00558_ ) );
OAI21_X1 _16254_ ( .A(_00558_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06208_ ), .ZN(_00559_ ) );
MUX2_X1 _16255_ ( .A(\io_master_rdata [31] ), .B(_00559_ ), .S(_02174_ ), .Z(_00560_ ) );
AND2_X1 _16256_ ( .A1(_00560_ ), .A2(_02176_ ), .ZN(\myifu.data_in [31] ) );
NAND2_X1 _16257_ ( .A1(_02175_ ), .A2(\io_master_rdata [30] ), .ZN(_00561_ ) );
NAND2_X1 _16258_ ( .A1(_06210_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_00562_ ) );
OAI211_X1 _16259_ ( .A(_02174_ ), .B(_00562_ ), .C1(_01760_ ), .C2(_06210_ ), .ZN(_00563_ ) );
AOI21_X1 _16260_ ( .A(_06179_ ), .B1(_00561_ ), .B2(_00563_ ), .ZN(\myifu.data_in [30] ) );
OR3_X1 _16261_ ( .A1(_02055_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06207_ ), .ZN(_00564_ ) );
OAI211_X1 _16262_ ( .A(_02118_ ), .B(_00564_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06208_ ), .ZN(_00565_ ) );
OAI21_X2 _16263_ ( .A(_00565_ ), .B1(\io_master_rdata [21] ), .B2(_02119_ ), .ZN(_00566_ ) );
BUF_X4 _16264_ ( .A(_06192_ ), .Z(_00567_ ) );
NOR2_X1 _16265_ ( .A1(_00566_ ), .A2(_00567_ ), .ZN(\myifu.data_in [21] ) );
OR2_X1 _16266_ ( .A1(_02121_ ), .A2(\io_master_rdata [20] ), .ZN(_00568_ ) );
CLKBUF_X2 _16267_ ( .A(_00557_ ), .Z(_00569_ ) );
OR3_X1 _16268_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00570_ ) );
OAI211_X1 _16269_ ( .A(_02121_ ), .B(_00570_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06210_ ), .ZN(_00571_ ) );
AND3_X1 _16270_ ( .A1(_00568_ ), .A2(_00571_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [20] ) );
OR2_X1 _16271_ ( .A1(_02120_ ), .A2(\io_master_rdata [19] ), .ZN(_00572_ ) );
OR3_X1 _16272_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00573_ ) );
OAI211_X1 _16273_ ( .A(_02121_ ), .B(_00573_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06210_ ), .ZN(_00574_ ) );
AND3_X1 _16274_ ( .A1(_00572_ ), .A2(_00574_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [19] ) );
BUF_X4 _16275_ ( .A(_02119_ ), .Z(_00575_ ) );
OR3_X1 _16276_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00576_ ) );
OAI211_X1 _16277_ ( .A(_00575_ ), .B(_00576_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06209_ ), .ZN(_00577_ ) );
OAI21_X1 _16278_ ( .A(_00577_ ), .B1(\io_master_rdata [18] ), .B2(_00575_ ), .ZN(_00578_ ) );
NOR2_X1 _16279_ ( .A1(_00578_ ), .A2(_00567_ ), .ZN(\myifu.data_in [18] ) );
OR2_X1 _16280_ ( .A1(_02120_ ), .A2(\io_master_rdata [17] ), .ZN(_00579_ ) );
OR3_X1 _16281_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00580_ ) );
OAI211_X1 _16282_ ( .A(_02121_ ), .B(_00580_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06210_ ), .ZN(_00581_ ) );
AND3_X1 _16283_ ( .A1(_00579_ ), .A2(_00581_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [17] ) );
OR3_X1 _16284_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00582_ ) );
OAI211_X1 _16285_ ( .A(_00575_ ), .B(_00582_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06209_ ), .ZN(_00583_ ) );
OAI21_X1 _16286_ ( .A(_00583_ ), .B1(\io_master_rdata [16] ), .B2(_00575_ ), .ZN(_00584_ ) );
NOR2_X1 _16287_ ( .A1(_00584_ ), .A2(_00567_ ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16288_ ( .A1(_02055_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06207_ ), .ZN(_00585_ ) );
OAI211_X1 _16289_ ( .A(_02119_ ), .B(_00585_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06208_ ), .ZN(_00586_ ) );
OAI21_X1 _16290_ ( .A(_00586_ ), .B1(\io_master_rdata [15] ), .B2(_02119_ ), .ZN(_00587_ ) );
NOR2_X1 _16291_ ( .A1(_00587_ ), .A2(_00567_ ), .ZN(\myifu.data_in [15] ) );
OR2_X1 _16292_ ( .A1(_02121_ ), .A2(\io_master_rdata [14] ), .ZN(_00588_ ) );
BUF_X2 _16293_ ( .A(_02120_ ), .Z(_00589_ ) );
CLKBUF_X2 _16294_ ( .A(_00569_ ), .Z(_00590_ ) );
OR3_X1 _16295_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00591_ ) );
OAI211_X1 _16296_ ( .A(_00589_ ), .B(_00591_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00592_ ) );
AND3_X1 _16297_ ( .A1(_00588_ ), .A2(_00592_ ), .A3(_02176_ ), .ZN(\myifu.data_in [14] ) );
OR3_X1 _16298_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00593_ ) );
OAI21_X1 _16299_ ( .A(_00593_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06209_ ), .ZN(_00594_ ) );
MUX2_X1 _16300_ ( .A(\io_master_rdata [13] ), .B(_00594_ ), .S(_02174_ ), .Z(_00595_ ) );
AND2_X1 _16301_ ( .A1(_00595_ ), .A2(_02176_ ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _16302_ ( .A1(_00589_ ), .A2(\io_master_rdata [12] ), .ZN(_00596_ ) );
OR3_X1 _16303_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00597_ ) );
OAI211_X1 _16304_ ( .A(_00589_ ), .B(_00597_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00598_ ) );
AND3_X1 _16305_ ( .A1(_00596_ ), .A2(_00598_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [12] ) );
OR3_X1 _16306_ ( .A1(_02055_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_06207_ ), .ZN(_00599_ ) );
OAI211_X1 _16307_ ( .A(_02118_ ), .B(_00599_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06208_ ), .ZN(_00600_ ) );
OAI21_X2 _16308_ ( .A(_00600_ ), .B1(\io_master_rdata [29] ), .B2(_02119_ ), .ZN(_00601_ ) );
NOR2_X1 _16309_ ( .A1(_00601_ ), .A2(_00567_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16310_ ( .A1(_00589_ ), .A2(\io_master_rdata [11] ), .ZN(_00602_ ) );
OR3_X1 _16311_ ( .A1(_02125_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00603_ ) );
OAI211_X1 _16312_ ( .A(_00589_ ), .B(_00603_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00604_ ) );
AND3_X1 _16313_ ( .A1(_00602_ ), .A2(_00604_ ), .A3(_02176_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16314_ ( .A1(_02120_ ), .A2(\io_master_rdata [10] ), .ZN(_00605_ ) );
OR3_X1 _16315_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00606_ ) );
OAI211_X1 _16316_ ( .A(_02120_ ), .B(_00606_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06210_ ), .ZN(_00607_ ) );
AND3_X1 _16317_ ( .A1(_00605_ ), .A2(_00607_ ), .A3(_02176_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16318_ ( .A1(_02122_ ), .A2(\io_master_rdata [9] ), .ZN(_00608_ ) );
OR3_X1 _16319_ ( .A1(_02125_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00609_ ) );
OAI211_X1 _16320_ ( .A(_02122_ ), .B(_00609_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00610_ ) );
AND3_X1 _16321_ ( .A1(_00608_ ), .A2(_00610_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16322_ ( .A1(_02120_ ), .A2(\io_master_rdata [8] ), .ZN(_00611_ ) );
OR3_X1 _16323_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00612_ ) );
OAI211_X1 _16324_ ( .A(_02120_ ), .B(_00612_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06209_ ), .ZN(_00613_ ) );
AND3_X1 _16325_ ( .A1(_00611_ ), .A2(_00613_ ), .A3(_02176_ ), .ZN(\myifu.data_in [8] ) );
OR3_X1 _16326_ ( .A1(_02055_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00614_ ) );
OAI21_X1 _16327_ ( .A(_00614_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_06208_ ), .ZN(_00615_ ) );
MUX2_X1 _16328_ ( .A(\io_master_rdata [7] ), .B(_00615_ ), .S(_02174_ ), .Z(_00616_ ) );
AND2_X1 _16329_ ( .A1(_00616_ ), .A2(_02176_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16330_ ( .A1(_02125_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00617_ ) );
OAI211_X1 _16331_ ( .A(_02122_ ), .B(_00617_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00618_ ) );
OAI21_X1 _16332_ ( .A(_00618_ ), .B1(\io_master_rdata [6] ), .B2(_02122_ ), .ZN(_00619_ ) );
NOR2_X1 _16333_ ( .A1(_00619_ ), .A2(_06178_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16334_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00620_ ) );
OAI211_X1 _16335_ ( .A(_00575_ ), .B(_00620_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06209_ ), .ZN(_00621_ ) );
OAI21_X1 _16336_ ( .A(_00621_ ), .B1(\io_master_rdata [5] ), .B2(_00575_ ), .ZN(_00622_ ) );
NOR2_X1 _16337_ ( .A1(_00622_ ), .A2(_00567_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16338_ ( .A1(_02125_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00623_ ) );
OAI211_X1 _16339_ ( .A(_00589_ ), .B(_00623_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00624_ ) );
OAI21_X1 _16340_ ( .A(_00624_ ), .B1(\io_master_rdata [4] ), .B2(_02122_ ), .ZN(_00625_ ) );
NOR2_X1 _16341_ ( .A1(_00625_ ), .A2(_00567_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16342_ ( .A1(_02125_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00626_ ) );
OAI211_X1 _16343_ ( .A(_00589_ ), .B(_00626_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00627_ ) );
OAI21_X1 _16344_ ( .A(_00627_ ), .B1(\io_master_rdata [3] ), .B2(_02122_ ), .ZN(_00628_ ) );
NOR2_X1 _16345_ ( .A1(_00628_ ), .A2(_00567_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16346_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00629_ ) );
OAI211_X1 _16347_ ( .A(_02119_ ), .B(_00629_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06209_ ), .ZN(_00630_ ) );
OAI21_X1 _16348_ ( .A(_00630_ ), .B1(\io_master_rdata [2] ), .B2(_00575_ ), .ZN(_00631_ ) );
NOR2_X1 _16349_ ( .A1(_00631_ ), .A2(_00567_ ), .ZN(\myifu.data_in [2] ) );
OR2_X1 _16350_ ( .A1(_02121_ ), .A2(\io_master_rdata [28] ), .ZN(_00632_ ) );
OR3_X1 _16351_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00633_ ) );
OAI211_X1 _16352_ ( .A(_02121_ ), .B(_00633_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06210_ ), .ZN(_00634_ ) );
AND3_X1 _16353_ ( .A1(_00632_ ), .A2(_00634_ ), .A3(_02125_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16354_ ( .A1(_02125_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00635_ ) );
OAI211_X1 _16355_ ( .A(_00589_ ), .B(_00635_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00636_ ) );
OAI21_X1 _16356_ ( .A(_00636_ ), .B1(\io_master_rdata [1] ), .B2(_02122_ ), .ZN(_00637_ ) );
NOR2_X1 _16357_ ( .A1(_00637_ ), .A2(_00567_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16358_ ( .A1(_02123_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00557_ ), .ZN(_00638_ ) );
OAI211_X1 _16359_ ( .A(_02119_ ), .B(_00638_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(_06209_ ), .ZN(_00639_ ) );
OAI21_X1 _16360_ ( .A(_00639_ ), .B1(\io_master_rdata [0] ), .B2(_00575_ ), .ZN(_00640_ ) );
NOR2_X1 _16361_ ( .A1(_00640_ ), .A2(_06179_ ), .ZN(\myifu.data_in [0] ) );
OR2_X1 _16362_ ( .A1(_02121_ ), .A2(\io_master_rdata [27] ), .ZN(_00641_ ) );
OR3_X1 _16363_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00642_ ) );
OAI211_X1 _16364_ ( .A(_00589_ ), .B(_00642_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06210_ ), .ZN(_00643_ ) );
AND3_X1 _16365_ ( .A1(_00641_ ), .A2(_00643_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [27] ) );
OR3_X1 _16366_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00644_ ) );
OAI211_X1 _16367_ ( .A(_00575_ ), .B(_00644_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06209_ ), .ZN(_00645_ ) );
OAI21_X1 _16368_ ( .A(_00645_ ), .B1(\io_master_rdata [26] ), .B2(_02120_ ), .ZN(_00646_ ) );
NOR2_X1 _16369_ ( .A1(_00646_ ), .A2(_06178_ ), .ZN(\myifu.data_in [26] ) );
OR2_X1 _16370_ ( .A1(_02122_ ), .A2(\io_master_rdata [25] ), .ZN(_00647_ ) );
OR3_X1 _16371_ ( .A1(_02125_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00648_ ) );
OAI211_X1 _16372_ ( .A(_02122_ ), .B(_00648_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00649_ ) );
AND3_X1 _16373_ ( .A1(_00647_ ), .A2(_00649_ ), .A3(_02176_ ), .ZN(\myifu.data_in [25] ) );
OR3_X1 _16374_ ( .A1(_02123_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00569_ ), .ZN(_00650_ ) );
OAI211_X1 _16375_ ( .A(_00575_ ), .B(_00650_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06209_ ), .ZN(_00651_ ) );
OAI21_X1 _16376_ ( .A(_00651_ ), .B1(\io_master_rdata [24] ), .B2(_02120_ ), .ZN(_00652_ ) );
NOR2_X1 _16377_ ( .A1(_00652_ ), .A2(_06179_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16378_ ( .A1(_02055_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00557_ ), .ZN(_00653_ ) );
OAI211_X2 _16379_ ( .A(_02119_ ), .B(_00653_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06208_ ), .ZN(_00654_ ) );
OAI21_X2 _16380_ ( .A(_00654_ ), .B1(\io_master_rdata [23] ), .B2(_02119_ ), .ZN(_00655_ ) );
NOR2_X1 _16381_ ( .A1(_00655_ ), .A2(_06179_ ), .ZN(\myifu.data_in [23] ) );
OR2_X1 _16382_ ( .A1(_02121_ ), .A2(\io_master_rdata [22] ), .ZN(_00656_ ) );
OR3_X1 _16383_ ( .A1(_02124_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00590_ ), .ZN(_00657_ ) );
OAI211_X1 _16384_ ( .A(_00589_ ), .B(_00657_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_06210_ ), .ZN(_00658_ ) );
AND3_X1 _16385_ ( .A1(_00656_ ), .A2(_00658_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16386_ ( .A(_00278_ ), .ZN(_00659_ ) );
NAND2_X1 _16387_ ( .A1(_00659_ ), .A2(_02162_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16388_ ( .A1(_06141_ ), .A2(fanout_net_9 ), .ZN(_00660_ ) );
INV_X1 _16389_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00661_ ) );
OAI21_X1 _16390_ ( .A(_02162_ ), .B1(_00660_ ), .B2(_00661_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16391_ ( .A1(_06144_ ), .A2(fanout_net_13 ), .ZN(_00662_ ) );
OAI21_X1 _16392_ ( .A(_02162_ ), .B1(_00662_ ), .B2(_00661_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16393_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .ZN(_00663_ ) );
OAI21_X1 _16394_ ( .A(_02162_ ), .B1(_00663_ ), .B2(_00661_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
AND2_X1 _16395_ ( .A1(_03299_ ), .A2(_03294_ ), .ZN(_00664_ ) );
INV_X1 _16396_ ( .A(_00664_ ), .ZN(_00665_ ) );
OAI21_X1 _16397_ ( .A(\IF_ID_inst [8] ), .B1(_00665_ ), .B2(_03521_ ), .ZN(_00666_ ) );
NOR4_X1 _16398_ ( .A1(_03465_ ), .A2(_03228_ ), .A3(_03469_ ), .A4(_03306_ ), .ZN(_00667_ ) );
AND2_X2 _16399_ ( .A1(_03523_ ), .A2(_03522_ ), .ZN(_00668_ ) );
INV_X1 _16400_ ( .A(_03310_ ), .ZN(_00669_ ) );
AND2_X1 _16401_ ( .A1(_00668_ ), .A2(_00669_ ), .ZN(_00670_ ) );
NAND3_X1 _16402_ ( .A1(_00667_ ), .A2(_00670_ ), .A3(_03542_ ), .ZN(_00671_ ) );
AND2_X1 _16403_ ( .A1(_00671_ ), .A2(_03635_ ), .ZN(_00672_ ) );
OAI221_X1 _16404_ ( .A(_00666_ ), .B1(_03449_ ), .B2(_03219_ ), .C1(_00672_ ), .C2(_03226_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
AND2_X1 _16405_ ( .A1(_03306_ ), .A2(\IF_ID_inst [31] ), .ZN(_00673_ ) );
INV_X1 _16406_ ( .A(_00673_ ), .ZN(_00674_ ) );
OAI221_X1 _16407_ ( .A(_00674_ ), .B1(_03514_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C1(_00670_ ), .C2(_03220_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
NOR2_X1 _16408_ ( .A1(_03514_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00675_ ) );
AOI21_X1 _16409_ ( .A(_03220_ ), .B1(_03523_ ), .B2(_03522_ ), .ZN(_00676_ ) );
NOR2_X1 _16410_ ( .A1(_00675_ ), .A2(_00676_ ), .ZN(_00677_ ) );
BUF_X4 _16411_ ( .A(_00677_ ), .Z(_00678_ ) );
BUF_X4 _16412_ ( .A(_00674_ ), .Z(_00679_ ) );
BUF_X4 _16413_ ( .A(_00669_ ), .Z(_00680_ ) );
OAI211_X1 _16414_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03225_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI211_X1 _16415_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03226_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI211_X1 _16416_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03229_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
OAI21_X1 _16417_ ( .A(\IF_ID_inst [31] ), .B1(_00665_ ), .B2(_03521_ ), .ZN(_00681_ ) );
BUF_X2 _16418_ ( .A(_03514_ ), .Z(_00682_ ) );
OAI221_X1 _16419_ ( .A(_00681_ ), .B1(_03301_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI221_X1 _16420_ ( .A(_00681_ ), .B1(_03318_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI221_X1 _16421_ ( .A(_00681_ ), .B1(_03319_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16422_ ( .A(_00681_ ), .B1(_03449_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _16423_ ( .A(_00681_ ), .B1(_03312_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16424_ ( .A(_00681_ ), .B1(_03323_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16425_ ( .A(_00681_ ), .B1(_03291_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16426_ ( .A(_00681_ ), .B1(_03213_ ), .B2(_03311_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI211_X1 _16427_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03230_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
AOI22_X1 _16428_ ( .A1(_00665_ ), .A2(\IF_ID_inst [31] ), .B1(\IF_ID_inst [7] ), .B2(_03521_ ), .ZN(_00683_ ) );
OAI221_X1 _16429_ ( .A(_00683_ ), .B1(_03229_ ), .B2(_03635_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_03514_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16430_ ( .A(_03687_ ), .ZN(_00684_ ) );
OAI221_X1 _16431_ ( .A(_00684_ ), .B1(_03225_ ), .B2(_00668_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
OAI221_X1 _16432_ ( .A(_03692_ ), .B1(_03230_ ), .B2(_00668_ ), .C1(_00682_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
INV_X1 _16433_ ( .A(_03649_ ), .ZN(_00685_ ) );
OAI221_X1 _16434_ ( .A(_00685_ ), .B1(_03231_ ), .B2(_00668_ ), .C1(_03514_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
INV_X1 _16435_ ( .A(_03602_ ), .ZN(_00686_ ) );
OAI221_X1 _16436_ ( .A(_00686_ ), .B1(_03232_ ), .B2(_00668_ ), .C1(_03514_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16437_ ( .A(_03612_ ), .ZN(_00687_ ) );
OAI221_X1 _16438_ ( .A(_00687_ ), .B1(_03234_ ), .B2(_00668_ ), .C1(_03514_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16439_ ( .A(_03608_ ), .ZN(_00688_ ) );
OAI221_X1 _16440_ ( .A(_00688_ ), .B1(_03235_ ), .B2(_00668_ ), .C1(_03514_ ), .C2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI211_X1 _16441_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03231_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI211_X1 _16442_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03232_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI211_X1 _16443_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03234_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI211_X1 _16444_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03235_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI211_X1 _16445_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03236_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI211_X1 _16446_ ( .A(_00678_ ), .B(_00679_ ), .C1(_03237_ ), .C2(_00680_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI211_X1 _16447_ ( .A(_00677_ ), .B(_00674_ ), .C1(_03238_ ), .C2(_00669_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16448_ ( .A(\IF_ID_inst [11] ), .B1(_00665_ ), .B2(_03521_ ), .ZN(_00689_ ) );
OAI221_X1 _16449_ ( .A(_00689_ ), .B1(_03301_ ), .B2(_03218_ ), .C1(_00672_ ), .C2(_03236_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16450_ ( .A(\IF_ID_inst [10] ), .B1(_00665_ ), .B2(_03521_ ), .ZN(_00690_ ) );
OAI221_X1 _16451_ ( .A(_00690_ ), .B1(_03318_ ), .B2(_03218_ ), .C1(_00672_ ), .C2(_03237_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16452_ ( .A(\IF_ID_inst [9] ), .B1(_00665_ ), .B2(_03521_ ), .ZN(_00691_ ) );
OAI221_X1 _16453_ ( .A(_00691_ ), .B1(_03319_ ), .B2(_03218_ ), .C1(_00672_ ), .C2(_03238_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16454_ ( .A1(_03523_ ), .A2(_03240_ ), .ZN(_00692_ ) );
OAI221_X1 _16455_ ( .A(_00692_ ), .B1(_03312_ ), .B2(_03218_ ), .C1(_00671_ ), .C2(_03229_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
AND3_X1 _16456_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00693_ ) );
CLKBUF_X2 _16457_ ( .A(_03426_ ), .Z(_00694_ ) );
AND3_X1 _16458_ ( .A1(_00694_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00695_ ) );
BUF_X4 _16459_ ( .A(_06137_ ), .Z(_00696_ ) );
AOI211_X1 _16460_ ( .A(_00693_ ), .B(_00695_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_00696_ ), .ZN(_00697_ ) );
NAND2_X2 _16461_ ( .A1(_00661_ ), .A2(\IF_ID_pc [2] ), .ZN(_00698_ ) );
BUF_X4 _16462_ ( .A(_00698_ ), .Z(_00699_ ) );
NAND2_X2 _16463_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00700_ ) );
BUF_X4 _16464_ ( .A(_00700_ ), .Z(_00701_ ) );
BUF_X4 _16465_ ( .A(_06143_ ), .Z(_00702_ ) );
NAND3_X1 _16466_ ( .A1(_00702_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00703_ ) );
NAND4_X1 _16467_ ( .A1(_00697_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00703_ ), .ZN(_00704_ ) );
NOR2_X1 _16468_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00705_ ) );
BUF_X4 _16469_ ( .A(_00705_ ), .Z(_00706_ ) );
BUF_X4 _16470_ ( .A(_06139_ ), .Z(_00707_ ) );
NAND3_X1 _16471_ ( .A1(_00707_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00708_ ) );
NAND3_X1 _16472_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00709_ ) );
AND2_X1 _16473_ ( .A1(_00708_ ), .A2(_00709_ ), .ZN(_00710_ ) );
NAND2_X1 _16474_ ( .A1(_00698_ ), .A2(_00700_ ), .ZN(_00711_ ) );
BUF_X4 _16475_ ( .A(_00711_ ), .Z(_00712_ ) );
BUF_X4 _16476_ ( .A(_06143_ ), .Z(_00713_ ) );
NAND3_X1 _16477_ ( .A1(_00713_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00714_ ) );
BUF_X4 _16478_ ( .A(_06140_ ), .Z(_00715_ ) );
BUF_X4 _16479_ ( .A(_06142_ ), .Z(_00716_ ) );
NAND3_X1 _16480_ ( .A1(_00715_ ), .A2(_00716_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00717_ ) );
NAND4_X1 _16481_ ( .A1(_00710_ ), .A2(_00712_ ), .A3(_00714_ ), .A4(_00717_ ), .ZN(_00718_ ) );
NAND3_X1 _16482_ ( .A1(_00704_ ), .A2(_00706_ ), .A3(_00718_ ), .ZN(_00719_ ) );
AOI21_X1 _16483_ ( .A(\IF_ID_pc [1] ), .B1(_03956_ ), .B2(\IF_ID_pc [2] ), .ZN(_00720_ ) );
INV_X1 _16484_ ( .A(_00720_ ), .ZN(_00721_ ) );
OAI21_X1 _16485_ ( .A(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .B1(_03956_ ), .B2(\IF_ID_pc [2] ), .ZN(_00722_ ) );
NOR2_X1 _16486_ ( .A1(_00721_ ), .A2(_00722_ ), .ZN(_00723_ ) );
AND2_X2 _16487_ ( .A1(_03966_ ), .A2(_00723_ ), .ZN(_00724_ ) );
INV_X1 _16488_ ( .A(_00724_ ), .ZN(_00725_ ) );
BUF_X2 _16489_ ( .A(_00725_ ), .Z(_00726_ ) );
NOR2_X1 _16490_ ( .A1(_00726_ ), .A2(\myifu.data_in [8] ), .ZN(_00727_ ) );
BUF_X4 _16491_ ( .A(_00724_ ), .Z(_00728_ ) );
OAI21_X1 _16492_ ( .A(\myifu.state [2] ), .B1(_00728_ ), .B2(_03621_ ), .ZN(_00729_ ) );
OAI21_X1 _16493_ ( .A(_00719_ ), .B1(_00727_ ), .B2(_00729_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16494_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00730_ ) );
AND3_X1 _16495_ ( .A1(_00694_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00731_ ) );
AOI211_X1 _16496_ ( .A(_00730_ ), .B(_00731_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00696_ ), .ZN(_00732_ ) );
NAND3_X1 _16497_ ( .A1(_00702_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00733_ ) );
NAND4_X1 _16498_ ( .A1(_00732_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00733_ ), .ZN(_00734_ ) );
BUF_X4 _16499_ ( .A(_00705_ ), .Z(_00735_ ) );
NAND3_X1 _16500_ ( .A1(_00707_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00736_ ) );
NAND3_X1 _16501_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00737_ ) );
AND2_X1 _16502_ ( .A1(_00736_ ), .A2(_00737_ ), .ZN(_00738_ ) );
NAND3_X1 _16503_ ( .A1(_00713_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00739_ ) );
NAND3_X1 _16504_ ( .A1(_00715_ ), .A2(_00716_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00740_ ) );
NAND4_X1 _16505_ ( .A1(_00738_ ), .A2(_00712_ ), .A3(_00739_ ), .A4(_00740_ ), .ZN(_00741_ ) );
NAND3_X1 _16506_ ( .A1(_00734_ ), .A2(_00735_ ), .A3(_00741_ ), .ZN(_00742_ ) );
NOR2_X1 _16507_ ( .A1(_00726_ ), .A2(\myifu.data_in [31] ), .ZN(_00743_ ) );
OAI21_X1 _16508_ ( .A(\myifu.state [2] ), .B1(_00728_ ), .B2(_03530_ ), .ZN(_00744_ ) );
OAI21_X1 _16509_ ( .A(_00742_ ), .B1(_00743_ ), .B2(_00744_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
AND2_X1 _16510_ ( .A1(_00561_ ), .A2(_00563_ ), .ZN(_00745_ ) );
OAI211_X1 _16511_ ( .A(_03966_ ), .B(_00723_ ), .C1(_02087_ ), .C2(_00745_ ), .ZN(_00746_ ) );
OAI211_X1 _16512_ ( .A(_00746_ ), .B(\myifu.state [2] ), .C1(_00728_ ), .C2(_03688_ ), .ZN(_00747_ ) );
AND3_X1 _16513_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00748_ ) );
AND3_X1 _16514_ ( .A1(_06140_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00749_ ) );
AOI211_X1 _16515_ ( .A(_00748_ ), .B(_00749_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_06138_ ), .ZN(_00750_ ) );
BUF_X2 _16516_ ( .A(_00698_ ), .Z(_00751_ ) );
BUF_X4 _16517_ ( .A(_00700_ ), .Z(_00752_ ) );
NAND3_X1 _16518_ ( .A1(_06144_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00753_ ) );
NAND4_X1 _16519_ ( .A1(_00750_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00753_ ), .ZN(_00754_ ) );
BUF_X4 _16520_ ( .A(_00705_ ), .Z(_00755_ ) );
BUF_X4 _16521_ ( .A(_06139_ ), .Z(_00756_ ) );
NAND3_X1 _16522_ ( .A1(_00756_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00757_ ) );
NAND3_X1 _16523_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00758_ ) );
AND2_X1 _16524_ ( .A1(_00757_ ), .A2(_00758_ ), .ZN(_00759_ ) );
BUF_X2 _16525_ ( .A(_00711_ ), .Z(_00760_ ) );
BUF_X4 _16526_ ( .A(_06143_ ), .Z(_00761_ ) );
NAND3_X1 _16527_ ( .A1(_00761_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00762_ ) );
BUF_X4 _16528_ ( .A(_06143_ ), .Z(_00763_ ) );
NAND3_X1 _16529_ ( .A1(_06141_ ), .A2(_00763_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00764_ ) );
NAND4_X1 _16530_ ( .A1(_00759_ ), .A2(_00760_ ), .A3(_00762_ ), .A4(_00764_ ), .ZN(_00765_ ) );
NAND3_X1 _16531_ ( .A1(_00754_ ), .A2(_00755_ ), .A3(_00765_ ), .ZN(_00766_ ) );
NAND2_X1 _16532_ ( .A1(_00747_ ), .A2(_00766_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
INV_X1 _16533_ ( .A(\myifu.state [2] ), .ZN(_00767_ ) );
BUF_X4 _16534_ ( .A(_00767_ ), .Z(_00768_ ) );
BUF_X4 _16535_ ( .A(_00725_ ), .Z(_00769_ ) );
AOI21_X1 _16536_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00770_ ) );
BUF_X4 _16537_ ( .A(_00724_ ), .Z(_00771_ ) );
OAI21_X1 _16538_ ( .A(_00771_ ), .B1(_00566_ ), .B2(_06192_ ), .ZN(_00772_ ) );
NAND2_X1 _16539_ ( .A1(_00770_ ), .A2(_00772_ ), .ZN(_00773_ ) );
AND3_X1 _16540_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00774_ ) );
AND3_X1 _16541_ ( .A1(_06140_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00775_ ) );
AOI211_X1 _16542_ ( .A(_00774_ ), .B(_00775_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_06138_ ), .ZN(_00776_ ) );
NAND3_X1 _16543_ ( .A1(_06144_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00777_ ) );
NAND4_X1 _16544_ ( .A1(_00776_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00777_ ), .ZN(_00778_ ) );
NAND3_X1 _16545_ ( .A1(_00756_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00779_ ) );
NAND3_X1 _16546_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00780_ ) );
AND2_X1 _16547_ ( .A1(_00779_ ), .A2(_00780_ ), .ZN(_00781_ ) );
NAND3_X1 _16548_ ( .A1(_00761_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00782_ ) );
NAND3_X1 _16549_ ( .A1(_06141_ ), .A2(_00763_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00783_ ) );
NAND4_X1 _16550_ ( .A1(_00781_ ), .A2(_00760_ ), .A3(_00782_ ), .A4(_00783_ ), .ZN(_00784_ ) );
NAND3_X1 _16551_ ( .A1(_00778_ ), .A2(_00755_ ), .A3(_00784_ ), .ZN(_00785_ ) );
NAND2_X1 _16552_ ( .A1(_00773_ ), .A2(_00785_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
AOI21_X1 _16553_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00786_ ) );
NAND2_X1 _16554_ ( .A1(_00568_ ), .A2(_00571_ ), .ZN(_00787_ ) );
OAI21_X1 _16555_ ( .A(_00771_ ), .B1(_00787_ ), .B2(_06192_ ), .ZN(_00788_ ) );
NAND2_X1 _16556_ ( .A1(_00786_ ), .A2(_00788_ ), .ZN(_00789_ ) );
AND3_X1 _16557_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00790_ ) );
AND3_X1 _16558_ ( .A1(_06140_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00791_ ) );
AOI211_X1 _16559_ ( .A(_00790_ ), .B(_00791_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_06138_ ), .ZN(_00792_ ) );
NAND3_X1 _16560_ ( .A1(_06144_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00793_ ) );
NAND4_X1 _16561_ ( .A1(_00792_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00793_ ), .ZN(_00794_ ) );
NAND3_X1 _16562_ ( .A1(_00756_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00795_ ) );
NAND3_X1 _16563_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00796_ ) );
AND2_X1 _16564_ ( .A1(_00795_ ), .A2(_00796_ ), .ZN(_00797_ ) );
NAND3_X1 _16565_ ( .A1(_00761_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00798_ ) );
NAND3_X1 _16566_ ( .A1(_06141_ ), .A2(_00763_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00799_ ) );
NAND4_X1 _16567_ ( .A1(_00797_ ), .A2(_00760_ ), .A3(_00798_ ), .A4(_00799_ ), .ZN(_00800_ ) );
NAND3_X1 _16568_ ( .A1(_00794_ ), .A2(_00755_ ), .A3(_00800_ ), .ZN(_00801_ ) );
NAND2_X1 _16569_ ( .A1(_00789_ ), .A2(_00801_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
AOI21_X1 _16570_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00802_ ) );
NAND2_X1 _16571_ ( .A1(_00572_ ), .A2(_00574_ ), .ZN(_00803_ ) );
BUF_X4 _16572_ ( .A(_02087_ ), .Z(_00804_ ) );
OAI21_X1 _16573_ ( .A(_00771_ ), .B1(_00803_ ), .B2(_00804_ ), .ZN(_00805_ ) );
NAND2_X1 _16574_ ( .A1(_00802_ ), .A2(_00805_ ), .ZN(_00806_ ) );
AND3_X1 _16575_ ( .A1(fanout_net_13 ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00807_ ) );
AND3_X1 _16576_ ( .A1(_06140_ ), .A2(fanout_net_9 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00808_ ) );
AOI211_X1 _16577_ ( .A(_00807_ ), .B(_00808_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_06138_ ), .ZN(_00809_ ) );
NAND3_X1 _16578_ ( .A1(_06144_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00810_ ) );
NAND4_X1 _16579_ ( .A1(_00809_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00810_ ), .ZN(_00811_ ) );
BUF_X4 _16580_ ( .A(_06139_ ), .Z(_00812_ ) );
NAND3_X1 _16581_ ( .A1(_00812_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00813_ ) );
NAND3_X1 _16582_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00814_ ) );
AND2_X1 _16583_ ( .A1(_00813_ ), .A2(_00814_ ), .ZN(_00815_ ) );
BUF_X4 _16584_ ( .A(_00711_ ), .Z(_00816_ ) );
BUF_X4 _16585_ ( .A(_00816_ ), .Z(_00817_ ) );
NAND3_X1 _16586_ ( .A1(_00761_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00818_ ) );
NAND3_X1 _16587_ ( .A1(_06141_ ), .A2(_00763_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00819_ ) );
NAND4_X1 _16588_ ( .A1(_00815_ ), .A2(_00817_ ), .A3(_00818_ ), .A4(_00819_ ), .ZN(_00820_ ) );
NAND3_X1 _16589_ ( .A1(_00811_ ), .A2(_00755_ ), .A3(_00820_ ), .ZN(_00821_ ) );
NAND2_X1 _16590_ ( .A1(_00806_ ), .A2(_00821_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
AND3_X1 _16591_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00822_ ) );
AND3_X1 _16592_ ( .A1(_00694_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00823_ ) );
AOI211_X1 _16593_ ( .A(_00822_ ), .B(_00823_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_00696_ ), .ZN(_00824_ ) );
NAND3_X1 _16594_ ( .A1(_00702_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00825_ ) );
NAND4_X1 _16595_ ( .A1(_00824_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00825_ ), .ZN(_00826_ ) );
NAND3_X1 _16596_ ( .A1(_00707_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00827_ ) );
NAND3_X1 _16597_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00828_ ) );
AND2_X1 _16598_ ( .A1(_00827_ ), .A2(_00828_ ), .ZN(_00829_ ) );
NAND3_X1 _16599_ ( .A1(_00713_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00830_ ) );
BUF_X4 _16600_ ( .A(_06143_ ), .Z(_00831_ ) );
NAND3_X1 _16601_ ( .A1(_00715_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00832_ ) );
NAND4_X1 _16602_ ( .A1(_00829_ ), .A2(_00712_ ), .A3(_00830_ ), .A4(_00832_ ), .ZN(_00833_ ) );
NAND3_X1 _16603_ ( .A1(_00826_ ), .A2(_00735_ ), .A3(_00833_ ), .ZN(_00834_ ) );
BUF_X4 _16604_ ( .A(_00724_ ), .Z(_00835_ ) );
OAI21_X1 _16605_ ( .A(_00835_ ), .B1(_00578_ ), .B2(_06178_ ), .ZN(_00836_ ) );
NAND2_X1 _16606_ ( .A1(_00836_ ), .A2(\myifu.state [2] ), .ZN(_00837_ ) );
CLKBUF_X2 _16607_ ( .A(_00725_ ), .Z(_00838_ ) );
AND2_X1 _16608_ ( .A1(_00838_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00839_ ) );
OAI21_X1 _16609_ ( .A(_00834_ ), .B1(_00837_ ), .B2(_00839_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
AOI21_X1 _16610_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00840_ ) );
NAND2_X1 _16611_ ( .A1(_00579_ ), .A2(_00581_ ), .ZN(_00841_ ) );
OAI21_X1 _16612_ ( .A(_00771_ ), .B1(_00841_ ), .B2(_00804_ ), .ZN(_00842_ ) );
NAND2_X1 _16613_ ( .A1(_00840_ ), .A2(_00842_ ), .ZN(_00843_ ) );
AND3_X1 _16614_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00844_ ) );
AND3_X1 _16615_ ( .A1(_06140_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00845_ ) );
AOI211_X1 _16616_ ( .A(_00844_ ), .B(_00845_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_06138_ ), .ZN(_00846_ ) );
NAND3_X1 _16617_ ( .A1(_06144_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00847_ ) );
NAND4_X1 _16618_ ( .A1(_00846_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00847_ ), .ZN(_00848_ ) );
NAND3_X1 _16619_ ( .A1(_00812_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00849_ ) );
NAND3_X1 _16620_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00850_ ) );
AND2_X1 _16621_ ( .A1(_00849_ ), .A2(_00850_ ), .ZN(_00851_ ) );
NAND3_X1 _16622_ ( .A1(_00761_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00852_ ) );
BUF_X4 _16623_ ( .A(_06143_ ), .Z(_00853_ ) );
NAND3_X1 _16624_ ( .A1(_06141_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00854_ ) );
NAND4_X1 _16625_ ( .A1(_00851_ ), .A2(_00817_ ), .A3(_00852_ ), .A4(_00854_ ), .ZN(_00855_ ) );
NAND3_X1 _16626_ ( .A1(_00848_ ), .A2(_00755_ ), .A3(_00855_ ), .ZN(_00856_ ) );
NAND2_X1 _16627_ ( .A1(_00843_ ), .A2(_00856_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
AND3_X1 _16628_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00857_ ) );
AND3_X1 _16629_ ( .A1(_00694_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00858_ ) );
AOI211_X1 _16630_ ( .A(_00857_ ), .B(_00858_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_00696_ ), .ZN(_00859_ ) );
NAND3_X1 _16631_ ( .A1(_00702_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00860_ ) );
NAND4_X1 _16632_ ( .A1(_00859_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00860_ ), .ZN(_00861_ ) );
NAND3_X1 _16633_ ( .A1(_00707_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00862_ ) );
NAND3_X1 _16634_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00863_ ) );
AND2_X1 _16635_ ( .A1(_00862_ ), .A2(_00863_ ), .ZN(_00864_ ) );
NAND3_X1 _16636_ ( .A1(_00713_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00865_ ) );
NAND3_X1 _16637_ ( .A1(_00715_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00866_ ) );
NAND4_X1 _16638_ ( .A1(_00864_ ), .A2(_00712_ ), .A3(_00865_ ), .A4(_00866_ ), .ZN(_00867_ ) );
NAND3_X1 _16639_ ( .A1(_00861_ ), .A2(_00735_ ), .A3(_00867_ ), .ZN(_00868_ ) );
OAI21_X1 _16640_ ( .A(_00835_ ), .B1(_00584_ ), .B2(_06178_ ), .ZN(_00869_ ) );
NAND2_X1 _16641_ ( .A1(_00869_ ), .A2(\myifu.state [2] ), .ZN(_00870_ ) );
AND2_X1 _16642_ ( .A1(_00838_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00871_ ) );
OAI21_X1 _16643_ ( .A(_00868_ ), .B1(_00870_ ), .B2(_00871_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
AOI21_X1 _16644_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00872_ ) );
OAI21_X1 _16645_ ( .A(_00771_ ), .B1(_00587_ ), .B2(_00804_ ), .ZN(_00873_ ) );
NAND2_X1 _16646_ ( .A1(_00872_ ), .A2(_00873_ ), .ZN(_00874_ ) );
AND3_X1 _16647_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00875_ ) );
AND3_X1 _16648_ ( .A1(_06140_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00876_ ) );
AOI211_X1 _16649_ ( .A(_00875_ ), .B(_00876_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_06138_ ), .ZN(_00877_ ) );
BUF_X4 _16650_ ( .A(_06143_ ), .Z(_00878_ ) );
NAND3_X1 _16651_ ( .A1(_00878_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00879_ ) );
NAND4_X1 _16652_ ( .A1(_00877_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00879_ ), .ZN(_00880_ ) );
NAND3_X1 _16653_ ( .A1(_00812_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00881_ ) );
NAND3_X1 _16654_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00882_ ) );
AND2_X1 _16655_ ( .A1(_00881_ ), .A2(_00882_ ), .ZN(_00883_ ) );
NAND3_X1 _16656_ ( .A1(_00761_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00884_ ) );
BUF_X4 _16657_ ( .A(_06139_ ), .Z(_00885_ ) );
BUF_X4 _16658_ ( .A(_00885_ ), .Z(_00886_ ) );
NAND3_X1 _16659_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00887_ ) );
NAND4_X1 _16660_ ( .A1(_00883_ ), .A2(_00817_ ), .A3(_00884_ ), .A4(_00887_ ), .ZN(_00888_ ) );
NAND3_X1 _16661_ ( .A1(_00880_ ), .A2(_00755_ ), .A3(_00888_ ), .ZN(_00889_ ) );
NAND2_X1 _16662_ ( .A1(_00874_ ), .A2(_00889_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
AND3_X1 _16663_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00890_ ) );
AND3_X1 _16664_ ( .A1(_00694_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00891_ ) );
AOI211_X1 _16665_ ( .A(_00890_ ), .B(_00891_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_00696_ ), .ZN(_00892_ ) );
NAND3_X1 _16666_ ( .A1(_00702_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00893_ ) );
NAND4_X1 _16667_ ( .A1(_00892_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00893_ ), .ZN(_00894_ ) );
NAND3_X1 _16668_ ( .A1(_00885_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00895_ ) );
NAND3_X1 _16669_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00896_ ) );
AND2_X1 _16670_ ( .A1(_00895_ ), .A2(_00896_ ), .ZN(_00897_ ) );
NAND3_X1 _16671_ ( .A1(_00713_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00898_ ) );
NAND3_X1 _16672_ ( .A1(_00715_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00899_ ) );
NAND4_X1 _16673_ ( .A1(_00897_ ), .A2(_00816_ ), .A3(_00898_ ), .A4(_00899_ ), .ZN(_00900_ ) );
NAND3_X1 _16674_ ( .A1(_00894_ ), .A2(_00735_ ), .A3(_00900_ ), .ZN(_00901_ ) );
AND2_X1 _16675_ ( .A1(_00726_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00902_ ) );
OAI21_X1 _16676_ ( .A(\myifu.state [2] ), .B1(_00726_ ), .B2(\myifu.data_in [14] ), .ZN(_00903_ ) );
OAI21_X1 _16677_ ( .A(_00901_ ), .B1(_00902_ ), .B2(_00903_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
AND3_X1 _16678_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00904_ ) );
AND3_X1 _16679_ ( .A1(_00694_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00905_ ) );
AOI211_X1 _16680_ ( .A(_00904_ ), .B(_00905_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_00696_ ), .ZN(_00906_ ) );
NAND3_X1 _16681_ ( .A1(_00702_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00907_ ) );
NAND4_X1 _16682_ ( .A1(_00906_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00907_ ), .ZN(_00908_ ) );
NAND3_X1 _16683_ ( .A1(_00885_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00909_ ) );
NAND3_X1 _16684_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00910_ ) );
AND2_X1 _16685_ ( .A1(_00909_ ), .A2(_00910_ ), .ZN(_00911_ ) );
NAND3_X1 _16686_ ( .A1(_00716_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_00912_ ) );
NAND3_X1 _16687_ ( .A1(_00715_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_00913_ ) );
NAND4_X1 _16688_ ( .A1(_00911_ ), .A2(_00816_ ), .A3(_00912_ ), .A4(_00913_ ), .ZN(_00914_ ) );
NAND3_X1 _16689_ ( .A1(_00908_ ), .A2(_00735_ ), .A3(_00914_ ), .ZN(_00915_ ) );
AND2_X1 _16690_ ( .A1(_00726_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00916_ ) );
OAI21_X1 _16691_ ( .A(\myifu.state [2] ), .B1(_00726_ ), .B2(\myifu.data_in [13] ), .ZN(_00917_ ) );
OAI21_X1 _16692_ ( .A(_00915_ ), .B1(_00916_ ), .B2(_00917_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
AOI21_X1 _16693_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00918_ ) );
NAND2_X1 _16694_ ( .A1(_00596_ ), .A2(_00598_ ), .ZN(_00919_ ) );
OAI21_X1 _16695_ ( .A(_00771_ ), .B1(_00919_ ), .B2(_00804_ ), .ZN(_00920_ ) );
NAND2_X1 _16696_ ( .A1(_00918_ ), .A2(_00920_ ), .ZN(_00921_ ) );
AND3_X1 _16697_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_00922_ ) );
AND3_X1 _16698_ ( .A1(_06140_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_00923_ ) );
BUF_X4 _16699_ ( .A(_06137_ ), .Z(_00924_ ) );
AOI211_X1 _16700_ ( .A(_00922_ ), .B(_00923_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_00924_ ), .ZN(_00925_ ) );
NAND3_X1 _16701_ ( .A1(_00878_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_00926_ ) );
NAND4_X1 _16702_ ( .A1(_00925_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00926_ ), .ZN(_00927_ ) );
NAND3_X1 _16703_ ( .A1(_00812_ ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_00928_ ) );
NAND3_X1 _16704_ ( .A1(fanout_net_14 ), .A2(fanout_net_10 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_00929_ ) );
AND2_X1 _16705_ ( .A1(_00928_ ), .A2(_00929_ ), .ZN(_00930_ ) );
BUF_X4 _16706_ ( .A(_06143_ ), .Z(_00931_ ) );
NAND3_X1 _16707_ ( .A1(_00931_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_00932_ ) );
NAND3_X1 _16708_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_00933_ ) );
NAND4_X1 _16709_ ( .A1(_00930_ ), .A2(_00817_ ), .A3(_00932_ ), .A4(_00933_ ), .ZN(_00934_ ) );
NAND3_X1 _16710_ ( .A1(_00927_ ), .A2(_00755_ ), .A3(_00934_ ), .ZN(_00935_ ) );
NAND2_X1 _16711_ ( .A1(_00921_ ), .A2(_00935_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
OAI21_X1 _16712_ ( .A(_00835_ ), .B1(_00601_ ), .B2(_06178_ ), .ZN(_00936_ ) );
OAI211_X1 _16713_ ( .A(_00936_ ), .B(\myifu.state [2] ), .C1(_00728_ ), .C2(_03694_ ), .ZN(_00937_ ) );
AND3_X1 _16714_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_00938_ ) );
AND3_X1 _16715_ ( .A1(_06140_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_00939_ ) );
AOI211_X1 _16716_ ( .A(_00938_ ), .B(_00939_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_00924_ ), .ZN(_00940_ ) );
NAND3_X1 _16717_ ( .A1(_00878_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_00941_ ) );
NAND4_X1 _16718_ ( .A1(_00940_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00941_ ), .ZN(_00942_ ) );
NAND3_X1 _16719_ ( .A1(_00812_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_00943_ ) );
NAND3_X1 _16720_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_00944_ ) );
AND2_X1 _16721_ ( .A1(_00943_ ), .A2(_00944_ ), .ZN(_00945_ ) );
NAND3_X1 _16722_ ( .A1(_00931_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_00946_ ) );
NAND3_X1 _16723_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_00947_ ) );
NAND4_X1 _16724_ ( .A1(_00945_ ), .A2(_00817_ ), .A3(_00946_ ), .A4(_00947_ ), .ZN(_00948_ ) );
NAND3_X1 _16725_ ( .A1(_00942_ ), .A2(_00755_ ), .A3(_00948_ ), .ZN(_00949_ ) );
NAND2_X1 _16726_ ( .A1(_00937_ ), .A2(_00949_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16727_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_00950_ ) );
AND3_X1 _16728_ ( .A1(_00694_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_00951_ ) );
AOI211_X1 _16729_ ( .A(_00950_ ), .B(_00951_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_00696_ ), .ZN(_00952_ ) );
NAND3_X1 _16730_ ( .A1(_00702_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_00953_ ) );
NAND4_X1 _16731_ ( .A1(_00952_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00953_ ), .ZN(_00954_ ) );
NAND3_X1 _16732_ ( .A1(_00885_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_00955_ ) );
NAND3_X1 _16733_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_00956_ ) );
AND2_X1 _16734_ ( .A1(_00955_ ), .A2(_00956_ ), .ZN(_00957_ ) );
NAND3_X1 _16735_ ( .A1(_00716_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_00958_ ) );
NAND3_X1 _16736_ ( .A1(_00756_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_00959_ ) );
NAND4_X1 _16737_ ( .A1(_00957_ ), .A2(_00816_ ), .A3(_00958_ ), .A4(_00959_ ), .ZN(_00960_ ) );
NAND3_X1 _16738_ ( .A1(_00954_ ), .A2(_00735_ ), .A3(_00960_ ), .ZN(_00961_ ) );
NOR2_X1 _16739_ ( .A1(_00726_ ), .A2(\myifu.data_in [11] ), .ZN(_00962_ ) );
OAI21_X1 _16740_ ( .A(\myifu.state [2] ), .B1(_00728_ ), .B2(_03633_ ), .ZN(_00963_ ) );
OAI21_X1 _16741_ ( .A(_00961_ ), .B1(_00962_ ), .B2(_00963_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
AND3_X1 _16742_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_00964_ ) );
AND3_X1 _16743_ ( .A1(_00694_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_00965_ ) );
AOI211_X1 _16744_ ( .A(_00964_ ), .B(_00965_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_06137_ ), .ZN(_00966_ ) );
NAND3_X1 _16745_ ( .A1(_00763_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_00967_ ) );
NAND4_X1 _16746_ ( .A1(_00966_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00967_ ), .ZN(_00968_ ) );
NAND3_X1 _16747_ ( .A1(_00885_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_00969_ ) );
NAND3_X1 _16748_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_00970_ ) );
AND2_X1 _16749_ ( .A1(_00969_ ), .A2(_00970_ ), .ZN(_00971_ ) );
NAND3_X1 _16750_ ( .A1(_00716_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_00972_ ) );
NAND3_X1 _16751_ ( .A1(_00756_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_00973_ ) );
NAND4_X1 _16752_ ( .A1(_00971_ ), .A2(_00816_ ), .A3(_00972_ ), .A4(_00973_ ), .ZN(_00974_ ) );
NAND3_X1 _16753_ ( .A1(_00968_ ), .A2(_00735_ ), .A3(_00974_ ), .ZN(_00975_ ) );
NOR2_X1 _16754_ ( .A1(_00726_ ), .A2(\myifu.data_in [10] ), .ZN(_00976_ ) );
OAI21_X1 _16755_ ( .A(\myifu.state [2] ), .B1(_00728_ ), .B2(_03629_ ), .ZN(_00977_ ) );
OAI21_X1 _16756_ ( .A(_00975_ ), .B1(_00976_ ), .B2(_00977_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
NAND2_X1 _16757_ ( .A1(_00608_ ), .A2(_00610_ ), .ZN(_00978_ ) );
OAI21_X1 _16758_ ( .A(_00724_ ), .B1(_00978_ ), .B2(_06178_ ), .ZN(_00979_ ) );
OAI211_X1 _16759_ ( .A(_00979_ ), .B(\myifu.state [2] ), .C1(_00728_ ), .C2(_03617_ ), .ZN(_00980_ ) );
AND3_X1 _16760_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_00981_ ) );
CLKBUF_X2 _16761_ ( .A(_06139_ ), .Z(_00982_ ) );
AND3_X1 _16762_ ( .A1(_00982_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_00983_ ) );
AOI211_X1 _16763_ ( .A(_00981_ ), .B(_00983_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_00924_ ), .ZN(_00984_ ) );
NAND3_X1 _16764_ ( .A1(_00878_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_00985_ ) );
NAND4_X1 _16765_ ( .A1(_00984_ ), .A2(_00751_ ), .A3(_00752_ ), .A4(_00985_ ), .ZN(_00986_ ) );
NAND3_X1 _16766_ ( .A1(_00812_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_00987_ ) );
NAND3_X1 _16767_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_00988_ ) );
AND2_X1 _16768_ ( .A1(_00987_ ), .A2(_00988_ ), .ZN(_00989_ ) );
NAND3_X1 _16769_ ( .A1(_00931_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_00990_ ) );
NAND3_X1 _16770_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_00991_ ) );
NAND4_X1 _16771_ ( .A1(_00989_ ), .A2(_00817_ ), .A3(_00990_ ), .A4(_00991_ ), .ZN(_00992_ ) );
NAND3_X1 _16772_ ( .A1(_00986_ ), .A2(_00755_ ), .A3(_00992_ ), .ZN(_00993_ ) );
NAND2_X1 _16773_ ( .A1(_00980_ ), .A2(_00993_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
AND3_X1 _16774_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_00994_ ) );
AND3_X1 _16775_ ( .A1(_00694_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_00995_ ) );
AOI211_X1 _16776_ ( .A(_00994_ ), .B(_00995_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_06137_ ), .ZN(_00996_ ) );
NAND3_X1 _16777_ ( .A1(_00763_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_00997_ ) );
NAND4_X1 _16778_ ( .A1(_00996_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_00997_ ), .ZN(_00998_ ) );
NAND3_X1 _16779_ ( .A1(_00885_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_00999_ ) );
NAND3_X1 _16780_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_01000_ ) );
AND2_X1 _16781_ ( .A1(_00999_ ), .A2(_01000_ ), .ZN(_01001_ ) );
NAND3_X1 _16782_ ( .A1(_00716_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_01002_ ) );
NAND3_X1 _16783_ ( .A1(_00756_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_01003_ ) );
NAND4_X1 _16784_ ( .A1(_01001_ ), .A2(_00816_ ), .A3(_01002_ ), .A4(_01003_ ), .ZN(_01004_ ) );
NAND3_X1 _16785_ ( .A1(_00998_ ), .A2(_00735_ ), .A3(_01004_ ), .ZN(_01005_ ) );
NOR4_X1 _16786_ ( .A1(\myifu.data_in [7] ), .A2(_03967_ ), .A3(_00722_ ), .A4(_00721_ ), .ZN(_01006_ ) );
OAI21_X1 _16787_ ( .A(\myifu.state [2] ), .B1(_00728_ ), .B2(_03678_ ), .ZN(_01007_ ) );
OAI21_X1 _16788_ ( .A(_01005_ ), .B1(_01006_ ), .B2(_01007_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AND3_X1 _16789_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_01008_ ) );
AND3_X1 _16790_ ( .A1(_06139_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_01009_ ) );
AOI211_X1 _16791_ ( .A(_01008_ ), .B(_01009_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_06137_ ), .ZN(_01010_ ) );
NAND3_X1 _16792_ ( .A1(_00763_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_01011_ ) );
NAND4_X1 _16793_ ( .A1(_01010_ ), .A2(_00699_ ), .A3(_00701_ ), .A4(_01011_ ), .ZN(_01012_ ) );
NAND3_X1 _16794_ ( .A1(_00885_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_01013_ ) );
NAND3_X1 _16795_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_01014_ ) );
AND2_X1 _16796_ ( .A1(_01013_ ), .A2(_01014_ ), .ZN(_01015_ ) );
NAND3_X1 _16797_ ( .A1(_00716_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_01016_ ) );
NAND3_X1 _16798_ ( .A1(_00756_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_01017_ ) );
NAND4_X1 _16799_ ( .A1(_01015_ ), .A2(_00816_ ), .A3(_01016_ ), .A4(_01017_ ), .ZN(_01018_ ) );
NAND3_X1 _16800_ ( .A1(_01012_ ), .A2(_00735_ ), .A3(_01018_ ), .ZN(_01019_ ) );
NOR2_X1 _16801_ ( .A1(\myifu.data_in [6] ), .A2(_00726_ ), .ZN(_01020_ ) );
OAI21_X1 _16802_ ( .A(\myifu.state [2] ), .B1(_00771_ ), .B2(_03302_ ), .ZN(_01021_ ) );
OAI21_X1 _16803_ ( .A(_01019_ ), .B1(_01020_ ), .B2(_01021_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
AOI21_X1 _16804_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01022_ ) );
OAI21_X1 _16805_ ( .A(_00771_ ), .B1(_00622_ ), .B2(_00804_ ), .ZN(_01023_ ) );
NAND2_X1 _16806_ ( .A1(_01022_ ), .A2(_01023_ ), .ZN(_01024_ ) );
AND3_X1 _16807_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_01025_ ) );
AND3_X1 _16808_ ( .A1(_00982_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_01026_ ) );
AOI211_X1 _16809_ ( .A(_01025_ ), .B(_01026_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00924_ ), .ZN(_01027_ ) );
BUF_X4 _16810_ ( .A(_00698_ ), .Z(_01028_ ) );
BUF_X4 _16811_ ( .A(_00700_ ), .Z(_01029_ ) );
NAND3_X1 _16812_ ( .A1(_00878_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_01030_ ) );
NAND4_X1 _16813_ ( .A1(_01027_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01030_ ), .ZN(_01031_ ) );
NAND3_X1 _16814_ ( .A1(_00812_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_01032_ ) );
NAND3_X1 _16815_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_01033_ ) );
AND2_X1 _16816_ ( .A1(_01032_ ), .A2(_01033_ ), .ZN(_01034_ ) );
NAND3_X1 _16817_ ( .A1(_00931_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_01035_ ) );
NAND3_X1 _16818_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_01036_ ) );
NAND4_X1 _16819_ ( .A1(_01034_ ), .A2(_00817_ ), .A3(_01035_ ), .A4(_01036_ ), .ZN(_01037_ ) );
NAND3_X1 _16820_ ( .A1(_01031_ ), .A2(_00755_ ), .A3(_01037_ ), .ZN(_01038_ ) );
NAND2_X1 _16821_ ( .A1(_01024_ ), .A2(_01038_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
AOI21_X1 _16822_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01039_ ) );
OAI21_X1 _16823_ ( .A(_00771_ ), .B1(_00625_ ), .B2(_00804_ ), .ZN(_01040_ ) );
NAND2_X1 _16824_ ( .A1(_01039_ ), .A2(_01040_ ), .ZN(_01041_ ) );
AND3_X1 _16825_ ( .A1(fanout_net_15 ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_01042_ ) );
AND3_X1 _16826_ ( .A1(_00982_ ), .A2(fanout_net_11 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_01043_ ) );
AOI211_X1 _16827_ ( .A(_01042_ ), .B(_01043_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00924_ ), .ZN(_01044_ ) );
NAND3_X1 _16828_ ( .A1(_00878_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_01045_ ) );
NAND4_X1 _16829_ ( .A1(_01044_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01045_ ), .ZN(_01046_ ) );
NAND3_X1 _16830_ ( .A1(_00812_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_01047_ ) );
NAND3_X1 _16831_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_01048_ ) );
AND2_X1 _16832_ ( .A1(_01047_ ), .A2(_01048_ ), .ZN(_01049_ ) );
NAND3_X1 _16833_ ( .A1(_00931_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_01050_ ) );
NAND3_X1 _16834_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_01051_ ) );
NAND4_X1 _16835_ ( .A1(_01049_ ), .A2(_00817_ ), .A3(_01050_ ), .A4(_01051_ ), .ZN(_01052_ ) );
NAND3_X1 _16836_ ( .A1(_01046_ ), .A2(_00706_ ), .A3(_01052_ ), .ZN(_01053_ ) );
NAND2_X1 _16837_ ( .A1(_01041_ ), .A2(_01053_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _16838_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01054_ ) );
OAI21_X1 _16839_ ( .A(_00835_ ), .B1(_00628_ ), .B2(_00804_ ), .ZN(_01055_ ) );
NAND2_X1 _16840_ ( .A1(_01054_ ), .A2(_01055_ ), .ZN(_01056_ ) );
AND3_X1 _16841_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_01057_ ) );
AND3_X1 _16842_ ( .A1(_00982_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_01058_ ) );
AOI211_X1 _16843_ ( .A(_01057_ ), .B(_01058_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00924_ ), .ZN(_01059_ ) );
NAND3_X1 _16844_ ( .A1(_00878_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_01060_ ) );
NAND4_X1 _16845_ ( .A1(_01059_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01060_ ), .ZN(_01061_ ) );
NAND3_X1 _16846_ ( .A1(_00812_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_01062_ ) );
NAND3_X1 _16847_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_01063_ ) );
AND2_X1 _16848_ ( .A1(_01062_ ), .A2(_01063_ ), .ZN(_01064_ ) );
NAND3_X1 _16849_ ( .A1(_00931_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_01065_ ) );
NAND3_X1 _16850_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_01066_ ) );
NAND4_X1 _16851_ ( .A1(_01064_ ), .A2(_00817_ ), .A3(_01065_ ), .A4(_01066_ ), .ZN(_01067_ ) );
NAND3_X1 _16852_ ( .A1(_01061_ ), .A2(_00706_ ), .A3(_01067_ ), .ZN(_01068_ ) );
NAND2_X1 _16853_ ( .A1(_01056_ ), .A2(_01068_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
AOI21_X1 _16854_ ( .A(_00768_ ), .B1(_00769_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01069_ ) );
OAI21_X1 _16855_ ( .A(_00835_ ), .B1(_00631_ ), .B2(_00804_ ), .ZN(_01070_ ) );
NAND2_X1 _16856_ ( .A1(_01069_ ), .A2(_01070_ ), .ZN(_01071_ ) );
AND3_X1 _16857_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_01072_ ) );
AND3_X1 _16858_ ( .A1(_00982_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_01073_ ) );
AOI211_X1 _16859_ ( .A(_01072_ ), .B(_01073_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_00924_ ), .ZN(_01074_ ) );
NAND3_X1 _16860_ ( .A1(_00878_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_01075_ ) );
NAND4_X1 _16861_ ( .A1(_01074_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01075_ ), .ZN(_01076_ ) );
NAND3_X1 _16862_ ( .A1(_00812_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_01077_ ) );
NAND3_X1 _16863_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_01078_ ) );
AND2_X1 _16864_ ( .A1(_01077_ ), .A2(_01078_ ), .ZN(_01079_ ) );
NAND3_X1 _16865_ ( .A1(_00931_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_01080_ ) );
NAND3_X1 _16866_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_01081_ ) );
NAND4_X1 _16867_ ( .A1(_01079_ ), .A2(_00817_ ), .A3(_01080_ ), .A4(_01081_ ), .ZN(_01082_ ) );
NAND3_X1 _16868_ ( .A1(_01076_ ), .A2(_00706_ ), .A3(_01082_ ), .ZN(_01083_ ) );
NAND2_X1 _16869_ ( .A1(_01071_ ), .A2(_01083_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
AOI21_X1 _16870_ ( .A(_00767_ ), .B1(_00838_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01084_ ) );
OAI21_X1 _16871_ ( .A(_00835_ ), .B1(_00637_ ), .B2(_00804_ ), .ZN(_01085_ ) );
NAND2_X1 _16872_ ( .A1(_01084_ ), .A2(_01085_ ), .ZN(_01086_ ) );
AND3_X1 _16873_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_01087_ ) );
AND3_X1 _16874_ ( .A1(_00982_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_01088_ ) );
AOI211_X1 _16875_ ( .A(_01087_ ), .B(_01088_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_00924_ ), .ZN(_01089_ ) );
NAND3_X1 _16876_ ( .A1(_00878_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_01090_ ) );
NAND4_X1 _16877_ ( .A1(_01089_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01090_ ), .ZN(_01091_ ) );
NAND3_X1 _16878_ ( .A1(_00707_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_01092_ ) );
NAND3_X1 _16879_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_01093_ ) );
AND2_X1 _16880_ ( .A1(_01092_ ), .A2(_01093_ ), .ZN(_01094_ ) );
NAND3_X1 _16881_ ( .A1(_00931_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_01095_ ) );
NAND3_X1 _16882_ ( .A1(_00886_ ), .A2(_00853_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_01096_ ) );
NAND4_X1 _16883_ ( .A1(_01094_ ), .A2(_00712_ ), .A3(_01095_ ), .A4(_01096_ ), .ZN(_01097_ ) );
NAND3_X1 _16884_ ( .A1(_01091_ ), .A2(_00706_ ), .A3(_01097_ ), .ZN(_01098_ ) );
NAND2_X1 _16885_ ( .A1(_01086_ ), .A2(_01098_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
OR2_X1 _16886_ ( .A1(_00838_ ), .A2(\myifu.data_in [28] ), .ZN(_01099_ ) );
OAI211_X1 _16887_ ( .A(_01099_ ), .B(\myifu.state [2] ), .C1(_00728_ ), .C2(_03650_ ), .ZN(_01100_ ) );
AND3_X1 _16888_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_01101_ ) );
AND3_X1 _16889_ ( .A1(_00982_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01102_ ) );
AOI211_X1 _16890_ ( .A(_01101_ ), .B(_01102_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00924_ ), .ZN(_01103_ ) );
NAND3_X1 _16891_ ( .A1(_00878_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01104_ ) );
NAND4_X1 _16892_ ( .A1(_01103_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01104_ ), .ZN(_01105_ ) );
NAND3_X1 _16893_ ( .A1(_00707_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01106_ ) );
NAND3_X1 _16894_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01107_ ) );
AND2_X1 _16895_ ( .A1(_01106_ ), .A2(_01107_ ), .ZN(_01108_ ) );
NAND3_X1 _16896_ ( .A1(_00931_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01109_ ) );
NAND3_X1 _16897_ ( .A1(_00886_ ), .A2(_00713_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01110_ ) );
NAND4_X1 _16898_ ( .A1(_01108_ ), .A2(_00712_ ), .A3(_01109_ ), .A4(_01110_ ), .ZN(_01111_ ) );
NAND3_X1 _16899_ ( .A1(_01105_ ), .A2(_00706_ ), .A3(_01111_ ), .ZN(_01112_ ) );
NAND2_X1 _16900_ ( .A1(_01100_ ), .A2(_01112_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
AND3_X1 _16901_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01113_ ) );
AND3_X1 _16902_ ( .A1(_06139_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01114_ ) );
AOI211_X1 _16903_ ( .A(_01113_ ), .B(_01114_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_06137_ ), .ZN(_01115_ ) );
NAND3_X1 _16904_ ( .A1(_00763_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01116_ ) );
NAND4_X1 _16905_ ( .A1(_01115_ ), .A2(_00698_ ), .A3(_00700_ ), .A4(_01116_ ), .ZN(_01117_ ) );
NAND3_X1 _16906_ ( .A1(_00885_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01118_ ) );
NAND3_X1 _16907_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01119_ ) );
AND2_X1 _16908_ ( .A1(_01118_ ), .A2(_01119_ ), .ZN(_01120_ ) );
NAND3_X1 _16909_ ( .A1(_00716_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01121_ ) );
NAND3_X1 _16910_ ( .A1(_00756_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01122_ ) );
NAND4_X1 _16911_ ( .A1(_01120_ ), .A2(_00816_ ), .A3(_01121_ ), .A4(_01122_ ), .ZN(_01123_ ) );
NAND3_X1 _16912_ ( .A1(_01117_ ), .A2(_00735_ ), .A3(_01123_ ), .ZN(_01124_ ) );
OAI21_X1 _16913_ ( .A(_00835_ ), .B1(_00640_ ), .B2(_06178_ ), .ZN(_01125_ ) );
NAND2_X1 _16914_ ( .A1(_01125_ ), .A2(\myifu.state [2] ), .ZN(_01126_ ) );
AND2_X1 _16915_ ( .A1(_00838_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01127_ ) );
OAI21_X1 _16916_ ( .A(_01124_ ), .B1(_01126_ ), .B2(_01127_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
NAND2_X1 _16917_ ( .A1(_00641_ ), .A2(_00643_ ), .ZN(_01128_ ) );
OAI21_X1 _16918_ ( .A(_00724_ ), .B1(_01128_ ), .B2(_02087_ ), .ZN(_01129_ ) );
OAI211_X1 _16919_ ( .A(_01129_ ), .B(\myifu.state [2] ), .C1(_00728_ ), .C2(_03603_ ), .ZN(_01130_ ) );
AND3_X1 _16920_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01131_ ) );
AND3_X1 _16921_ ( .A1(_00982_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01132_ ) );
AOI211_X1 _16922_ ( .A(_01131_ ), .B(_01132_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00924_ ), .ZN(_01133_ ) );
NAND3_X1 _16923_ ( .A1(_00761_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01134_ ) );
NAND4_X1 _16924_ ( .A1(_01133_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01134_ ), .ZN(_01135_ ) );
NAND3_X1 _16925_ ( .A1(_00707_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01136_ ) );
NAND3_X1 _16926_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01137_ ) );
AND2_X1 _16927_ ( .A1(_01136_ ), .A2(_01137_ ), .ZN(_01138_ ) );
NAND3_X1 _16928_ ( .A1(_00931_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01139_ ) );
NAND3_X1 _16929_ ( .A1(_00715_ ), .A2(_00713_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01140_ ) );
NAND4_X1 _16930_ ( .A1(_01138_ ), .A2(_00712_ ), .A3(_01139_ ), .A4(_01140_ ), .ZN(_01141_ ) );
NAND3_X1 _16931_ ( .A1(_01135_ ), .A2(_00706_ ), .A3(_01141_ ), .ZN(_01142_ ) );
NAND2_X1 _16932_ ( .A1(_01130_ ), .A2(_01142_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
AND3_X1 _16933_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01143_ ) );
AND3_X1 _16934_ ( .A1(_06139_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01144_ ) );
AOI211_X1 _16935_ ( .A(_01143_ ), .B(_01144_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_06137_ ), .ZN(_01145_ ) );
NAND3_X1 _16936_ ( .A1(_00763_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01146_ ) );
NAND4_X1 _16937_ ( .A1(_01145_ ), .A2(_00698_ ), .A3(_00700_ ), .A4(_01146_ ), .ZN(_01147_ ) );
NAND3_X1 _16938_ ( .A1(_00885_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01148_ ) );
NAND3_X1 _16939_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01149_ ) );
AND2_X1 _16940_ ( .A1(_01148_ ), .A2(_01149_ ), .ZN(_01150_ ) );
NAND3_X1 _16941_ ( .A1(_00716_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01151_ ) );
NAND3_X1 _16942_ ( .A1(_00756_ ), .A2(_00831_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01152_ ) );
NAND4_X1 _16943_ ( .A1(_01150_ ), .A2(_00816_ ), .A3(_01151_ ), .A4(_01152_ ), .ZN(_01153_ ) );
NAND3_X1 _16944_ ( .A1(_01147_ ), .A2(_00705_ ), .A3(_01153_ ), .ZN(_01154_ ) );
NOR2_X1 _16945_ ( .A1(\myifu.data_in [26] ), .A2(_00726_ ), .ZN(_01155_ ) );
OAI21_X1 _16946_ ( .A(\myifu.state [2] ), .B1(_00771_ ), .B2(_03613_ ), .ZN(_01156_ ) );
OAI21_X1 _16947_ ( .A(_01154_ ), .B1(_01155_ ), .B2(_01156_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
OR2_X1 _16948_ ( .A1(_00838_ ), .A2(\myifu.data_in [25] ), .ZN(_01157_ ) );
AOI21_X1 _16949_ ( .A(_00767_ ), .B1(_00838_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_01158_ ) );
NAND2_X1 _16950_ ( .A1(_01157_ ), .A2(_01158_ ), .ZN(_01159_ ) );
AND3_X1 _16951_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01160_ ) );
AND3_X1 _16952_ ( .A1(_00982_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01161_ ) );
AOI211_X1 _16953_ ( .A(_01160_ ), .B(_01161_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_00696_ ), .ZN(_01162_ ) );
NAND3_X1 _16954_ ( .A1(_00761_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01163_ ) );
NAND4_X1 _16955_ ( .A1(_01162_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01163_ ), .ZN(_01164_ ) );
NAND3_X1 _16956_ ( .A1(_00707_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01165_ ) );
NAND3_X1 _16957_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01166_ ) );
AND2_X1 _16958_ ( .A1(_01165_ ), .A2(_01166_ ), .ZN(_01167_ ) );
NAND3_X1 _16959_ ( .A1(_00702_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01168_ ) );
NAND3_X1 _16960_ ( .A1(_00715_ ), .A2(_00713_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01169_ ) );
NAND4_X1 _16961_ ( .A1(_01167_ ), .A2(_00712_ ), .A3(_01168_ ), .A4(_01169_ ), .ZN(_01170_ ) );
NAND3_X1 _16962_ ( .A1(_01164_ ), .A2(_00706_ ), .A3(_01170_ ), .ZN(_01171_ ) );
NAND2_X1 _16963_ ( .A1(_01159_ ), .A2(_01171_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
AND3_X1 _16964_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01172_ ) );
AND3_X1 _16965_ ( .A1(_06139_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01173_ ) );
AOI211_X1 _16966_ ( .A(_01172_ ), .B(_01173_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_06137_ ), .ZN(_01174_ ) );
NAND3_X1 _16967_ ( .A1(_00763_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01175_ ) );
NAND4_X1 _16968_ ( .A1(_01174_ ), .A2(_00698_ ), .A3(_00700_ ), .A4(_01175_ ), .ZN(_01176_ ) );
NAND3_X1 _16969_ ( .A1(_00885_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01177_ ) );
NAND3_X1 _16970_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01178_ ) );
AND2_X1 _16971_ ( .A1(_01177_ ), .A2(_01178_ ), .ZN(_01179_ ) );
NAND3_X1 _16972_ ( .A1(_00716_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01180_ ) );
NAND3_X1 _16973_ ( .A1(_00756_ ), .A2(_06143_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01181_ ) );
NAND4_X1 _16974_ ( .A1(_01179_ ), .A2(_00816_ ), .A3(_01180_ ), .A4(_01181_ ), .ZN(_01182_ ) );
NAND3_X1 _16975_ ( .A1(_01176_ ), .A2(_00705_ ), .A3(_01182_ ), .ZN(_01183_ ) );
OAI21_X1 _16976_ ( .A(_00835_ ), .B1(_00652_ ), .B2(_06178_ ), .ZN(_01184_ ) );
NAND2_X1 _16977_ ( .A1(_01184_ ), .A2(\myifu.state [2] ), .ZN(_01185_ ) );
AND2_X1 _16978_ ( .A1(_00838_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01186_ ) );
OAI21_X1 _16979_ ( .A(_01183_ ), .B1(_01185_ ), .B2(_01186_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
AOI21_X1 _16980_ ( .A(_00767_ ), .B1(_00838_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01187_ ) );
OAI21_X1 _16981_ ( .A(_00835_ ), .B1(_00655_ ), .B2(_00804_ ), .ZN(_01188_ ) );
NAND2_X1 _16982_ ( .A1(_01187_ ), .A2(_01188_ ), .ZN(_01189_ ) );
AND3_X1 _16983_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01190_ ) );
AND3_X1 _16984_ ( .A1(_00982_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01191_ ) );
AOI211_X1 _16985_ ( .A(_01190_ ), .B(_01191_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_00696_ ), .ZN(_01192_ ) );
NAND3_X1 _16986_ ( .A1(_00761_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01193_ ) );
NAND4_X1 _16987_ ( .A1(_01192_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01193_ ), .ZN(_01194_ ) );
NAND3_X1 _16988_ ( .A1(_00707_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01195_ ) );
NAND3_X1 _16989_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01196_ ) );
AND2_X1 _16990_ ( .A1(_01195_ ), .A2(_01196_ ), .ZN(_01197_ ) );
NAND3_X1 _16991_ ( .A1(_00702_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01198_ ) );
NAND3_X1 _16992_ ( .A1(_00715_ ), .A2(_00713_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01199_ ) );
NAND4_X1 _16993_ ( .A1(_01197_ ), .A2(_00712_ ), .A3(_01198_ ), .A4(_01199_ ), .ZN(_01200_ ) );
NAND3_X1 _16994_ ( .A1(_01194_ ), .A2(_00706_ ), .A3(_01200_ ), .ZN(_01201_ ) );
NAND2_X1 _16995_ ( .A1(_01189_ ), .A2(_01201_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
AOI21_X1 _16996_ ( .A(_00767_ ), .B1(_00838_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_01202_ ) );
NAND2_X1 _16997_ ( .A1(_00656_ ), .A2(_00658_ ), .ZN(_01203_ ) );
OAI21_X1 _16998_ ( .A(_00835_ ), .B1(_01203_ ), .B2(_06178_ ), .ZN(_01204_ ) );
NAND2_X1 _16999_ ( .A1(_01202_ ), .A2(_01204_ ), .ZN(_01205_ ) );
AND3_X1 _17000_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01206_ ) );
AND3_X1 _17001_ ( .A1(_00694_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01207_ ) );
AOI211_X1 _17002_ ( .A(_01206_ ), .B(_01207_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_00696_ ), .ZN(_01208_ ) );
NAND3_X1 _17003_ ( .A1(_00761_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01209_ ) );
NAND4_X1 _17004_ ( .A1(_01208_ ), .A2(_01028_ ), .A3(_01029_ ), .A4(_01209_ ), .ZN(_01210_ ) );
NAND3_X1 _17005_ ( .A1(_00707_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01211_ ) );
NAND3_X1 _17006_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01212_ ) );
AND2_X1 _17007_ ( .A1(_01211_ ), .A2(_01212_ ), .ZN(_01213_ ) );
NAND3_X1 _17008_ ( .A1(_00702_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01214_ ) );
NAND3_X1 _17009_ ( .A1(_00715_ ), .A2(_00713_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01215_ ) );
NAND4_X1 _17010_ ( .A1(_01213_ ), .A2(_00712_ ), .A3(_01214_ ), .A4(_01215_ ), .ZN(_01216_ ) );
NAND3_X1 _17011_ ( .A1(_01210_ ), .A2(_00706_ ), .A3(_01216_ ), .ZN(_01217_ ) );
NAND2_X1 _17012_ ( .A1(_01205_ ), .A2(_01217_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI211_X1 _17013_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_03440_ ), .C1(_03780_ ), .C2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17014_ ( .A(_03968_ ), .ZN(_01218_ ) );
NAND4_X1 _17015_ ( .A1(_03965_ ), .A2(_03960_ ), .A3(\myifu.state [2] ), .A4(_01218_ ), .ZN(_01219_ ) );
NOR2_X1 _17016_ ( .A1(_02050_ ), .A2(_00556_ ), .ZN(_01220_ ) );
INV_X1 _17017_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01221_ ) );
AOI21_X1 _17018_ ( .A(_00554_ ), .B1(_01220_ ), .B2(_01221_ ), .ZN(_01222_ ) );
AOI21_X1 _17019_ ( .A(reset ), .B1(_01219_ ), .B2(_01222_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _17020_ ( .A1(_06127_ ), .A2(_02087_ ), .ZN(_01223_ ) );
AND3_X1 _17021_ ( .A1(_01964_ ), .A2(_02012_ ), .A3(_02049_ ), .ZN(_01224_ ) );
NOR4_X1 _17022_ ( .A1(_01223_ ), .A2(\myidu.stall_quest_fencei ), .A3(_00556_ ), .A4(_01224_ ), .ZN(_01225_ ) );
AND2_X1 _17023_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01226_ ) );
OR4_X1 _17024_ ( .A1(reset ), .A2(_01225_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A4(_01226_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _17025_ ( .A(_01587_ ), .B(\myifu.state [2] ), .C1(_03967_ ), .C2(_03968_ ), .ZN(_01227_ ) );
NAND2_X1 _17026_ ( .A1(_01223_ ), .A2(_02163_ ), .ZN(_01228_ ) );
NAND2_X1 _17027_ ( .A1(_01227_ ), .A2(_01228_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _17028_ ( .A1(_03965_ ), .A2(_03960_ ), .A3(\myifu.state [2] ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17029_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01229_ ) );
NOR3_X1 _17030_ ( .A1(_01229_ ), .A2(_00662_ ), .A3(_00760_ ), .ZN(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ) );
NOR3_X1 _17031_ ( .A1(_01229_ ), .A2(_00663_ ), .A3(_00760_ ), .ZN(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ) );
AND4_X1 _17032_ ( .A1(\IF_ID_pc [4] ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00760_ ), .ZN(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ) );
AND4_X1 _17033_ ( .A1(\IF_ID_pc [4] ), .A2(_06136_ ), .A3(_06144_ ), .A4(_00760_ ), .ZN(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ) );
NOR3_X1 _17034_ ( .A1(_01229_ ), .A2(_00660_ ), .A3(_00760_ ), .ZN(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ) );
AND4_X1 _17035_ ( .A1(_06141_ ), .A2(_06136_ ), .A3(\IF_ID_pc [3] ), .A4(_00760_ ), .ZN(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _17036_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06138_ ), .A3(_00760_ ), .ZN(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ) );
AND4_X1 _17037_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06138_ ), .A3(_00751_ ), .A4(_00752_ ), .ZN(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ) );
AND3_X1 _17038_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_06141_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ) );
AND3_X1 _17039_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_06144_ ), .ZN(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ) );
AND3_X1 _17040_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ) );
AND3_X1 _17041_ ( .A1(_02162_ ), .A2(_06138_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ) );
OR2_X1 _17042_ ( .A1(_01223_ ), .A2(_00556_ ), .ZN(_01230_ ) );
AND2_X1 _17043_ ( .A1(_02012_ ), .A2(_02049_ ), .ZN(_01231_ ) );
NAND3_X1 _17044_ ( .A1(_01231_ ), .A2(_01964_ ), .A3(\myifu.state [0] ), .ZN(_01232_ ) );
NOR3_X1 _17045_ ( .A1(_03441_ ), .A2(_00554_ ), .A3(_01226_ ), .ZN(_01233_ ) );
NAND3_X1 _17046_ ( .A1(_00556_ ), .A2(_03440_ ), .A3(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01234_ ) );
NAND4_X1 _17047_ ( .A1(_01230_ ), .A2(_01232_ ), .A3(_01233_ ), .A4(_01234_ ), .ZN(_01235_ ) );
AND2_X1 _17048_ ( .A1(_03966_ ), .A2(_01218_ ), .ZN(_01236_ ) );
INV_X1 _17049_ ( .A(_01236_ ), .ZN(_01237_ ) );
AOI21_X1 _17050_ ( .A(_01235_ ), .B1(_02052_ ), .B2(_01237_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
NOR3_X1 _17051_ ( .A1(_03788_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03442_ ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
INV_X1 _17052_ ( .A(_03272_ ), .ZN(_01238_ ) );
AOI211_X1 _17053_ ( .A(_00540_ ), .B(_00542_ ), .C1(_03219_ ), .C2(_01238_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
NAND3_X1 _17054_ ( .A1(_01233_ ), .A2(_01587_ ), .A3(_01234_ ), .ZN(_01239_ ) );
AOI21_X1 _17055_ ( .A(_01239_ ), .B1(_02050_ ), .B2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND3_X1 _17056_ ( .A1(_03960_ ), .A2(fanout_net_45 ), .A3(_06232_ ), .ZN(_01240_ ) );
INV_X1 _17057_ ( .A(fanout_net_45 ), .ZN(_01241_ ) );
BUF_X4 _17058_ ( .A(_01241_ ), .Z(_01242_ ) );
AOI21_X1 _17059_ ( .A(_01240_ ), .B1(_01242_ ), .B2(\mylsu.state [0] ), .ZN(_01243_ ) );
AOI21_X1 _17060_ ( .A(_01243_ ), .B1(\mylsu.state [0] ), .B2(_06134_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ) );
AOI211_X1 _17061_ ( .A(_04031_ ), .B(_01243_ ), .C1(\mylsu.state [0] ), .C2(_06134_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
AND2_X1 _17062_ ( .A1(\myexu.rst_logic_$_OR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__B_Y ), .A2(_02134_ ), .ZN(_01244_ ) );
AND2_X1 _17063_ ( .A1(_02147_ ), .A2(_01244_ ), .ZN(_01245_ ) );
INV_X1 _17064_ ( .A(_01245_ ), .ZN(_01246_ ) );
OAI22_X1 _17065_ ( .A1(_06132_ ), .A2(_01246_ ), .B1(_06233_ ), .B2(_06163_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _17066_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01247_ ) );
OR4_X1 _17067_ ( .A1(_06134_ ), .A2(_02151_ ), .A3(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ), .A4(_01247_ ), .ZN(_01248_ ) );
NOR4_X1 _17068_ ( .A1(_02152_ ), .A2(_02158_ ), .A3(_04031_ ), .A4(_01248_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
INV_X1 _17069_ ( .A(_02158_ ), .ZN(_01249_ ) );
AND2_X1 _17070_ ( .A1(io_master_wready ), .A2(io_master_awready ), .ZN(_01250_ ) );
NOR2_X1 _17071_ ( .A1(_03982_ ), .A2(_01250_ ), .ZN(_01251_ ) );
AND4_X1 _17072_ ( .A1(io_master_awready ), .A2(_06214_ ), .A3(_04026_ ), .A4(_01251_ ), .ZN(_01252_ ) );
OAI211_X1 _17073_ ( .A(_01249_ ), .B(_01252_ ), .C1(_02129_ ), .C2(_02151_ ), .ZN(_01253_ ) );
NAND3_X1 _17074_ ( .A1(_04029_ ), .A2(\mylsu.state [2] ), .A3(_06121_ ), .ZN(_01254_ ) );
OAI21_X1 _17075_ ( .A(_01253_ ), .B1(io_master_wready ), .B2(_01254_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
AND3_X1 _17076_ ( .A1(_02149_ ), .A2(\mylsu.state [0] ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_01255_ ) );
AND2_X1 _17077_ ( .A1(_06145_ ), .A2(_01255_ ), .ZN(_01256_ ) );
INV_X1 _17078_ ( .A(_02152_ ), .ZN(_01257_ ) );
NAND4_X1 _17079_ ( .A1(_01256_ ), .A2(_01257_ ), .A3(_01249_ ), .A4(_01250_ ), .ZN(_01258_ ) );
NAND3_X1 _17080_ ( .A1(_04026_ ), .A2(\mylsu.state [2] ), .A3(io_master_wready ), .ZN(_01259_ ) );
NAND3_X1 _17081_ ( .A1(_04026_ ), .A2(\mylsu.state [4] ), .A3(io_master_awready ), .ZN(_01260_ ) );
NAND3_X1 _17082_ ( .A1(_06228_ ), .A2(\mylsu.state [1] ), .A3(_04026_ ), .ZN(_01261_ ) );
NAND4_X1 _17083_ ( .A1(_01258_ ), .A2(_01259_ ), .A3(_01260_ ), .A4(_01261_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
OAI21_X1 _17084_ ( .A(_01245_ ), .B1(_06127_ ), .B2(_06169_ ), .ZN(_01262_ ) );
NAND3_X1 _17085_ ( .A1(_03960_ ), .A2(_00319_ ), .A3(_06232_ ), .ZN(_01263_ ) );
NAND4_X1 _17086_ ( .A1(_01255_ ), .A2(EXU_valid_LSU ), .A3(_04026_ ), .A4(_01247_ ), .ZN(_01264_ ) );
OAI21_X1 _17087_ ( .A(_01264_ ), .B1(_02129_ ), .B2(_02151_ ), .ZN(_01265_ ) );
OR4_X1 _17088_ ( .A1(\EX_LS_dest_csreg_mem [28] ), .A2(_02128_ ), .A3(_01256_ ), .A4(_02151_ ), .ZN(_01266_ ) );
NAND3_X1 _17089_ ( .A1(_01265_ ), .A2(_01266_ ), .A3(_01249_ ), .ZN(_01267_ ) );
AND3_X1 _17090_ ( .A1(_02158_ ), .A2(_06145_ ), .A3(_01255_ ), .ZN(_01268_ ) );
AOI21_X1 _17091_ ( .A(_04031_ ), .B1(\mylsu.state [0] ), .B2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_01269_ ) );
NAND3_X1 _17092_ ( .A1(_02151_ ), .A2(_02132_ ), .A3(\myexu.rst_logic_$_OR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__B_Y ), .ZN(_01270_ ) );
OAI211_X1 _17093_ ( .A(_01269_ ), .B(_01270_ ), .C1(_06228_ ), .C2(_06221_ ), .ZN(_01271_ ) );
AOI211_X1 _17094_ ( .A(_01268_ ), .B(_01271_ ), .C1(_02218_ ), .C2(_01244_ ), .ZN(_01272_ ) );
NAND4_X1 _17095_ ( .A1(_01262_ ), .A2(_01263_ ), .A3(_01267_ ), .A4(_01272_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND3_X1 _17096_ ( .A1(_04026_ ), .A2(\mylsu.state [4] ), .A3(_06122_ ), .ZN(_01273_ ) );
AND4_X1 _17097_ ( .A1(\mylsu.state [0] ), .A2(_02149_ ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .A4(_06122_ ), .ZN(_01274_ ) );
NAND3_X1 _17098_ ( .A1(_01274_ ), .A2(io_master_wready ), .A3(_04026_ ), .ZN(_01275_ ) );
OR3_X1 _17099_ ( .A1(_01275_ ), .A2(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A3(_03982_ ), .ZN(_01276_ ) );
OAI21_X1 _17100_ ( .A(_01273_ ), .B1(_02220_ ), .B2(_01276_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
AOI21_X1 _17101_ ( .A(\EX_LS_pc [21] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01277_ ) );
NAND3_X1 _17102_ ( .A1(_03988_ ), .A2(\EX_LS_flag [2] ), .A3(\EX_LS_result_csreg_mem [21] ), .ZN(_01278_ ) );
OAI211_X1 _17103_ ( .A(_03984_ ), .B(_01278_ ), .C1(_02183_ ), .C2(_03976_ ), .ZN(_01279_ ) );
AOI21_X1 _17104_ ( .A(_01279_ ), .B1(_02220_ ), .B2(_06148_ ), .ZN(_01280_ ) );
NOR2_X1 _17105_ ( .A1(_01277_ ), .A2(_01280_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _17106_ ( .A(\LS_WB_wdata_csreg [20] ), .B(\EX_LS_result_csreg_mem [20] ), .S(_03976_ ), .Z(_01281_ ) );
INV_X1 _17107_ ( .A(_03983_ ), .ZN(_01282_ ) );
OR2_X1 _17108_ ( .A1(_03973_ ), .A2(_01282_ ), .ZN(_01283_ ) );
BUF_X4 _17109_ ( .A(_01283_ ), .Z(_01284_ ) );
BUF_X4 _17110_ ( .A(_01284_ ), .Z(_01285_ ) );
MUX2_X1 _17111_ ( .A(_01281_ ), .B(\EX_LS_pc [20] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
OAI22_X1 _17112_ ( .A1(_06165_ ), .A2(_02185_ ), .B1(_04010_ ), .B2(_06254_ ), .ZN(_01286_ ) );
MUX2_X1 _17113_ ( .A(_01286_ ), .B(\EX_LS_pc [19] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
AOI21_X1 _17114_ ( .A(\EX_LS_pc [18] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01287_ ) );
MUX2_X1 _17115_ ( .A(\LS_WB_wdata_csreg [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_02233_ ), .Z(_01288_ ) );
NOR3_X1 _17116_ ( .A1(_03973_ ), .A2(_01282_ ), .A3(_01288_ ), .ZN(_01289_ ) );
NOR2_X1 _17117_ ( .A1(_01287_ ), .A2(_01289_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
OAI22_X1 _17118_ ( .A1(_06165_ ), .A2(_02187_ ), .B1(_04010_ ), .B2(_05592_ ), .ZN(_01290_ ) );
MUX2_X1 _17119_ ( .A(_01290_ ), .B(\EX_LS_pc [17] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
OAI22_X1 _17120_ ( .A1(_06165_ ), .A2(_02188_ ), .B1(_04010_ ), .B2(_05613_ ), .ZN(_01291_ ) );
MUX2_X1 _17121_ ( .A(_01291_ ), .B(\EX_LS_pc [16] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
AOI21_X1 _17122_ ( .A(\EX_LS_pc [15] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01292_ ) );
BUF_X4 _17123_ ( .A(_02234_ ), .Z(_01293_ ) );
OAI21_X1 _17124_ ( .A(_03984_ ), .B1(_01293_ ), .B2(_06268_ ), .ZN(_01294_ ) );
BUF_X4 _17125_ ( .A(_02234_ ), .Z(_01295_ ) );
AOI221_X4 _17126_ ( .A(_01294_ ), .B1(\LS_WB_wdata_csreg [15] ), .B2(_01295_ ), .C1(_02220_ ), .C2(_06148_ ), .ZN(_01296_ ) );
NOR2_X1 _17127_ ( .A1(_01292_ ), .A2(_01296_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _17128_ ( .A(\EX_LS_pc [14] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01297_ ) );
OAI21_X1 _17129_ ( .A(_03983_ ), .B1(_01293_ ), .B2(_05659_ ), .ZN(_01298_ ) );
AOI221_X4 _17130_ ( .A(_01298_ ), .B1(\LS_WB_wdata_csreg [14] ), .B2(_01295_ ), .C1(_02220_ ), .C2(_06148_ ), .ZN(_01299_ ) );
NOR2_X1 _17131_ ( .A1(_01297_ ), .A2(_01299_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
OAI22_X1 _17132_ ( .A1(_06165_ ), .A2(_02191_ ), .B1(_04010_ ), .B2(_05678_ ), .ZN(_01300_ ) );
MUX2_X1 _17133_ ( .A(_01300_ ), .B(\EX_LS_pc [13] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
OAI22_X1 _17134_ ( .A1(_06165_ ), .A2(_02192_ ), .B1(_04010_ ), .B2(_05705_ ), .ZN(_01301_ ) );
MUX2_X1 _17135_ ( .A(_01301_ ), .B(\EX_LS_pc [12] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _17136_ ( .A(\EX_LS_pc [30] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01302_ ) );
MUX2_X1 _17137_ ( .A(\LS_WB_wdata_csreg [30] ), .B(\EX_LS_result_csreg_mem [30] ), .S(_02233_ ), .Z(_01303_ ) );
NOR3_X1 _17138_ ( .A1(_03973_ ), .A2(_01282_ ), .A3(_01303_ ), .ZN(_01304_ ) );
NOR2_X1 _17139_ ( .A1(_01302_ ), .A2(_01304_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
OAI22_X1 _17140_ ( .A1(_06165_ ), .A2(_02194_ ), .B1(_04010_ ), .B2(_05729_ ), .ZN(_01305_ ) );
MUX2_X1 _17141_ ( .A(_01305_ ), .B(\EX_LS_pc [11] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
AOI221_X4 _17142_ ( .A(_01284_ ), .B1(\LS_WB_wdata_csreg [10] ), .B2(_01295_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [10] ), .ZN(_01306_ ) );
AOI21_X1 _17143_ ( .A(\EX_LS_pc [10] ), .B1(_03974_ ), .B2(_03984_ ), .ZN(_01307_ ) );
NOR2_X1 _17144_ ( .A1(_01306_ ), .A2(_01307_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
AOI221_X4 _17145_ ( .A(_01284_ ), .B1(\LS_WB_wdata_csreg [9] ), .B2(_01295_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [9] ), .ZN(_01308_ ) );
AOI21_X1 _17146_ ( .A(\EX_LS_pc [9] ), .B1(_03974_ ), .B2(_03984_ ), .ZN(_01309_ ) );
NOR2_X1 _17147_ ( .A1(_01308_ ), .A2(_01309_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
OAI22_X1 _17148_ ( .A1(_06165_ ), .A2(_02197_ ), .B1(_04010_ ), .B2(_05804_ ), .ZN(_01310_ ) );
MUX2_X1 _17149_ ( .A(_01310_ ), .B(\EX_LS_pc [8] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
AOI21_X1 _17150_ ( .A(\EX_LS_pc [7] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01311_ ) );
OAI21_X1 _17151_ ( .A(_03983_ ), .B1(_01293_ ), .B2(_06247_ ), .ZN(_01312_ ) );
AOI221_X4 _17152_ ( .A(_01312_ ), .B1(\LS_WB_wdata_csreg [7] ), .B2(_01295_ ), .C1(_02220_ ), .C2(_06148_ ), .ZN(_01313_ ) );
NOR2_X1 _17153_ ( .A1(_01311_ ), .A2(_01313_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _17154_ ( .A1(_06165_ ), .A2(_02199_ ), .B1(_04010_ ), .B2(_05840_ ), .ZN(_01314_ ) );
MUX2_X1 _17155_ ( .A(_01314_ ), .B(\EX_LS_pc [6] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
OAI22_X1 _17156_ ( .A1(_06165_ ), .A2(_02200_ ), .B1(_04010_ ), .B2(_05858_ ), .ZN(_01315_ ) );
MUX2_X1 _17157_ ( .A(_01315_ ), .B(\EX_LS_pc [5] ), .S(_01285_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
AOI21_X1 _17158_ ( .A(\EX_LS_pc [4] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01316_ ) );
OAI21_X1 _17159_ ( .A(_03983_ ), .B1(_01293_ ), .B2(_05885_ ), .ZN(_01317_ ) );
AOI221_X4 _17160_ ( .A(_01317_ ), .B1(\LS_WB_wdata_csreg [4] ), .B2(_01295_ ), .C1(_02220_ ), .C2(_06148_ ), .ZN(_01318_ ) );
NOR2_X1 _17161_ ( .A1(_01316_ ), .A2(_01318_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
OAI22_X1 _17162_ ( .A1(_03976_ ), .A2(_02202_ ), .B1(_03978_ ), .B2(_05898_ ), .ZN(_01319_ ) );
MUX2_X1 _17163_ ( .A(_01319_ ), .B(\EX_LS_pc [3] ), .S(_01284_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
OAI22_X1 _17164_ ( .A1(_03976_ ), .A2(_02203_ ), .B1(_03978_ ), .B2(_06238_ ), .ZN(_01320_ ) );
MUX2_X1 _17165_ ( .A(_01320_ ), .B(\EX_LS_pc [2] ), .S(_01284_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
OAI22_X1 _17166_ ( .A1(_03976_ ), .A2(_02193_ ), .B1(_03978_ ), .B2(_05454_ ), .ZN(_01321_ ) );
MUX2_X1 _17167_ ( .A(_01321_ ), .B(\EX_LS_pc [29] ), .S(_01284_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
AOI21_X1 _17168_ ( .A(\EX_LS_pc [1] ), .B1(_03975_ ), .B2(_03985_ ), .ZN(_01322_ ) );
OAI21_X1 _17169_ ( .A(_03983_ ), .B1(_01293_ ), .B2(_06239_ ), .ZN(_01323_ ) );
AOI221_X4 _17170_ ( .A(_01323_ ), .B1(\LS_WB_wdata_csreg [1] ), .B2(_01293_ ), .C1(_02220_ ), .C2(_06148_ ), .ZN(_01324_ ) );
NOR2_X1 _17171_ ( .A1(_01322_ ), .A2(_01324_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
OAI22_X1 _17172_ ( .A1(_03976_ ), .A2(_02206_ ), .B1(_03978_ ), .B2(_06240_ ), .ZN(_01325_ ) );
MUX2_X1 _17173_ ( .A(_01325_ ), .B(\EX_LS_pc [0] ), .S(_01284_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
OAI22_X1 _17174_ ( .A1(_03976_ ), .A2(_02204_ ), .B1(_03978_ ), .B2(_05746_ ), .ZN(_01326_ ) );
MUX2_X1 _17175_ ( .A(_01326_ ), .B(\EX_LS_pc [28] ), .S(_01284_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _17176_ ( .A(\EX_LS_pc [27] ), .B1(_03974_ ), .B2(_03985_ ), .ZN(_01327_ ) );
OAI21_X1 _17177_ ( .A(_03983_ ), .B1(_01293_ ), .B2(_05952_ ), .ZN(_01328_ ) );
AOI221_X4 _17178_ ( .A(_01328_ ), .B1(\LS_WB_wdata_csreg [27] ), .B2(_01293_ ), .C1(_02220_ ), .C2(_06148_ ), .ZN(_01329_ ) );
NOR2_X1 _17179_ ( .A1(_01327_ ), .A2(_01329_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
AOI221_X4 _17180_ ( .A(_01284_ ), .B1(\LS_WB_wdata_csreg [26] ), .B2(_01295_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [26] ), .ZN(_01330_ ) );
AOI21_X1 _17181_ ( .A(\EX_LS_pc [26] ), .B1(_03974_ ), .B2(_03984_ ), .ZN(_01331_ ) );
NOR2_X1 _17182_ ( .A1(_01330_ ), .A2(_01331_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI221_X4 _17183_ ( .A(_01283_ ), .B1(\LS_WB_wdata_csreg [25] ), .B2(_01295_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [25] ), .ZN(_01332_ ) );
AOI21_X1 _17184_ ( .A(\EX_LS_pc [25] ), .B1(_03974_ ), .B2(_03984_ ), .ZN(_01333_ ) );
NOR2_X1 _17185_ ( .A1(_01332_ ), .A2(_01333_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
AOI221_X4 _17186_ ( .A(_01283_ ), .B1(\LS_WB_wdata_csreg [24] ), .B2(_01295_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [24] ), .ZN(_01334_ ) );
AOI21_X1 _17187_ ( .A(\EX_LS_pc [24] ), .B1(_03974_ ), .B2(_03984_ ), .ZN(_01335_ ) );
NOR2_X1 _17188_ ( .A1(_01334_ ), .A2(_01335_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _17189_ ( .A(\EX_LS_pc [23] ), .B1(_03974_ ), .B2(_03984_ ), .ZN(_01336_ ) );
OAI21_X1 _17190_ ( .A(_03983_ ), .B1(_01293_ ), .B2(_06267_ ), .ZN(_01337_ ) );
AOI221_X4 _17191_ ( .A(_01337_ ), .B1(\LS_WB_wdata_csreg [23] ), .B2(_01293_ ), .C1(_02219_ ), .C2(_06148_ ), .ZN(_01338_ ) );
NOR2_X1 _17192_ ( .A1(_01336_ ), .A2(_01338_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
OAI22_X1 _17193_ ( .A1(_03976_ ), .A2(_02212_ ), .B1(_03978_ ), .B2(_06057_ ), .ZN(_01339_ ) );
MUX2_X1 _17194_ ( .A(_01339_ ), .B(\EX_LS_pc [22] ), .S(_01284_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
AOI221_X4 _17195_ ( .A(_01283_ ), .B1(\LS_WB_wdata_csreg [31] ), .B2(_01295_ ), .C1(\EX_LS_flag [2] ), .C2(\EX_LS_result_csreg_mem [31] ), .ZN(_01340_ ) );
AOI21_X1 _17196_ ( .A(\EX_LS_pc [31] ), .B1(_03974_ ), .B2(_03984_ ), .ZN(_01341_ ) );
NOR2_X1 _17197_ ( .A1(_01340_ ), .A2(_01341_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
INV_X1 _17198_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01342_ ) );
AND2_X1 _17199_ ( .A1(_01342_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01343_ ) );
INV_X1 _17200_ ( .A(\mylsu.typ_tmp [1] ), .ZN(_01344_ ) );
AND2_X1 _17201_ ( .A1(_01343_ ), .A2(_01344_ ), .ZN(_01345_ ) );
BUF_X2 _17202_ ( .A(_01345_ ), .Z(_01346_ ) );
NAND2_X1 _17203_ ( .A1(_01344_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01347_ ) );
NOR2_X1 _17204_ ( .A1(_01347_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01348_ ) );
OR2_X1 _17205_ ( .A1(_01346_ ), .A2(_01348_ ), .ZN(_01349_ ) );
NOR2_X2 _17206_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01350_ ) );
INV_X1 _17207_ ( .A(_01350_ ), .ZN(_01351_ ) );
OR3_X1 _17208_ ( .A1(_00587_ ), .A2(_06128_ ), .A3(_01351_ ), .ZN(_01352_ ) );
NAND3_X1 _17209_ ( .A1(_00560_ ), .A2(_02076_ ), .A3(_01351_ ), .ZN(_01353_ ) );
NAND2_X1 _17210_ ( .A1(_01352_ ), .A2(_01353_ ), .ZN(_01354_ ) );
AND2_X1 _17211_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01355_ ) );
AND2_X1 _17212_ ( .A1(_01355_ ), .A2(_01342_ ), .ZN(_01356_ ) );
BUF_X4 _17213_ ( .A(_01356_ ), .Z(_01357_ ) );
INV_X1 _17214_ ( .A(_01357_ ), .ZN(_01358_ ) );
NOR2_X2 _17215_ ( .A1(_01354_ ), .A2(_01358_ ), .ZN(_01359_ ) );
BUF_X4 _17216_ ( .A(_01355_ ), .Z(_01360_ ) );
INV_X1 _17217_ ( .A(_01360_ ), .ZN(_01361_ ) );
OR2_X2 _17218_ ( .A1(_00566_ ), .A2(_06128_ ), .ZN(_01362_ ) );
AOI211_X1 _17219_ ( .A(_01349_ ), .B(_01359_ ), .C1(_01361_ ), .C2(_01362_ ), .ZN(_01363_ ) );
OAI21_X1 _17220_ ( .A(_01363_ ), .B1(_01342_ ), .B2(_01361_ ), .ZN(_01364_ ) );
INV_X1 _17221_ ( .A(_01346_ ), .ZN(_01365_ ) );
BUF_X4 _17222_ ( .A(_01365_ ), .Z(_01366_ ) );
NOR2_X2 _17223_ ( .A1(_00587_ ), .A2(_06129_ ), .ZN(_01367_ ) );
NOR2_X1 _17224_ ( .A1(_06174_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01368_ ) );
NOR2_X1 _17225_ ( .A1(_00655_ ), .A2(_06128_ ), .ZN(_01369_ ) );
NOR2_X1 _17226_ ( .A1(_06170_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01370_ ) );
AOI22_X1 _17227_ ( .A1(_01367_ ), .A2(_01368_ ), .B1(_01369_ ), .B2(_01370_ ), .ZN(_01371_ ) );
NAND3_X1 _17228_ ( .A1(_00616_ ), .A2(_06211_ ), .A3(_01350_ ), .ZN(_01372_ ) );
NAND4_X1 _17229_ ( .A1(_00560_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_02076_ ), .ZN(_01373_ ) );
AND3_X4 _17230_ ( .A1(_01371_ ), .A2(_01372_ ), .A3(_01373_ ), .ZN(_01374_ ) );
BUF_X4 _17231_ ( .A(_01374_ ), .Z(_01375_ ) );
OAI21_X1 _17232_ ( .A(_01364_ ), .B1(_01366_ ), .B2(_01375_ ), .ZN(_01376_ ) );
MUX2_X1 _17233_ ( .A(\EX_LS_result_reg [21] ), .B(_01376_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
NOR2_X2 _17234_ ( .A1(_01359_ ), .A2(_01349_ ), .ZN(_01377_ ) );
BUF_X4 _17235_ ( .A(_01377_ ), .Z(_01378_ ) );
BUF_X4 _17236_ ( .A(_01357_ ), .Z(_01379_ ) );
NAND3_X1 _17237_ ( .A1(_00568_ ), .A2(_00571_ ), .A3(\io_master_arid [1] ), .ZN(_01380_ ) );
AND2_X1 _17238_ ( .A1(_01360_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01381_ ) );
BUF_X4 _17239_ ( .A(_01381_ ), .Z(_01382_ ) );
NOR2_X1 _17240_ ( .A1(_01380_ ), .A2(_01382_ ), .ZN(_01383_ ) );
OAI21_X1 _17241_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01383_ ), .ZN(_01384_ ) );
OAI21_X1 _17242_ ( .A(_01384_ ), .B1(_01366_ ), .B2(_01375_ ), .ZN(_01385_ ) );
MUX2_X1 _17243_ ( .A(\EX_LS_result_reg [20] ), .B(_01385_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _17244_ ( .A1(_00572_ ), .A2(_00574_ ), .A3(_06211_ ), .ZN(_01386_ ) );
NOR2_X1 _17245_ ( .A1(_01386_ ), .A2(_01382_ ), .ZN(_01387_ ) );
OAI21_X1 _17246_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01387_ ), .ZN(_01388_ ) );
BUF_X4 _17247_ ( .A(_01374_ ), .Z(_01389_ ) );
OAI21_X1 _17248_ ( .A(_01388_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01390_ ) );
MUX2_X1 _17249_ ( .A(\EX_LS_result_reg [19] ), .B(_01390_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
NOR3_X1 _17250_ ( .A1(_00578_ ), .A2(_06131_ ), .A3(_01360_ ), .ZN(_01391_ ) );
OAI21_X1 _17251_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01391_ ), .ZN(_01392_ ) );
OAI21_X1 _17252_ ( .A(_01392_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01393_ ) );
MUX2_X1 _17253_ ( .A(\EX_LS_result_reg [18] ), .B(_01393_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
NAND3_X1 _17254_ ( .A1(_00579_ ), .A2(_00581_ ), .A3(_06211_ ), .ZN(_01394_ ) );
NOR2_X1 _17255_ ( .A1(_01394_ ), .A2(_01382_ ), .ZN(_01395_ ) );
OAI21_X1 _17256_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01395_ ), .ZN(_01396_ ) );
OAI21_X1 _17257_ ( .A(_01396_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01397_ ) );
MUX2_X1 _17258_ ( .A(\EX_LS_result_reg [17] ), .B(_01397_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
NOR3_X1 _17259_ ( .A1(_00584_ ), .A2(_06131_ ), .A3(_01360_ ), .ZN(_01398_ ) );
OAI21_X1 _17260_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01398_ ), .ZN(_01399_ ) );
OAI21_X1 _17261_ ( .A(_01399_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01400_ ) );
MUX2_X1 _17262_ ( .A(\EX_LS_result_reg [16] ), .B(_01400_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
NOR3_X1 _17263_ ( .A1(_01346_ ), .A2(_01360_ ), .A3(_01348_ ), .ZN(_01401_ ) );
NAND2_X1 _17264_ ( .A1(_01367_ ), .A2(_01401_ ), .ZN(_01402_ ) );
NAND2_X1 _17265_ ( .A1(_01354_ ), .A2(_01360_ ), .ZN(_01403_ ) );
BUF_X4 _17266_ ( .A(_01365_ ), .Z(_01404_ ) );
OAI211_X1 _17267_ ( .A(_01402_ ), .B(_01403_ ), .C1(_01375_ ), .C2(_01404_ ), .ZN(_01405_ ) );
MUX2_X1 _17268_ ( .A(\EX_LS_result_reg [15] ), .B(_01405_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
NOR2_X1 _17269_ ( .A1(_01361_ ), .A2(_01350_ ), .ZN(_01406_ ) );
NOR2_X1 _17270_ ( .A1(_06130_ ), .A2(_01406_ ), .ZN(_01407_ ) );
INV_X1 _17271_ ( .A(_01349_ ), .ZN(_01408_ ) );
AND2_X1 _17272_ ( .A1(_01407_ ), .A2(_01408_ ), .ZN(_01409_ ) );
AND3_X1 _17273_ ( .A1(_00588_ ), .A2(_00592_ ), .A3(_01409_ ), .ZN(_01410_ ) );
NOR2_X1 _17274_ ( .A1(_00745_ ), .A2(_06131_ ), .ZN(_01411_ ) );
AOI21_X1 _17275_ ( .A(_01410_ ), .B1(_01411_ ), .B2(_01406_ ), .ZN(_01412_ ) );
OAI21_X1 _17276_ ( .A(_01412_ ), .B1(_01375_ ), .B2(_01404_ ), .ZN(_01413_ ) );
MUX2_X1 _17277_ ( .A(\EX_LS_result_reg [14] ), .B(_01413_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
NAND2_X1 _17278_ ( .A1(_00595_ ), .A2(_06211_ ), .ZN(_01414_ ) );
NOR2_X1 _17279_ ( .A1(_00601_ ), .A2(_06128_ ), .ZN(_01415_ ) );
INV_X1 _17280_ ( .A(_01415_ ), .ZN(_01416_ ) );
MUX2_X1 _17281_ ( .A(_01414_ ), .B(_01416_ ), .S(_01406_ ), .Z(_01417_ ) );
OAI22_X1 _17282_ ( .A1(_01375_ ), .A2(_01404_ ), .B1(_01349_ ), .B2(_01417_ ), .ZN(_01418_ ) );
MUX2_X1 _17283_ ( .A(\EX_LS_result_reg [13] ), .B(_01418_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
AND4_X1 _17284_ ( .A1(\io_master_arid [1] ), .A2(_00632_ ), .A3(_00634_ ), .A4(_01406_ ), .ZN(_01419_ ) );
AND3_X1 _17285_ ( .A1(_00596_ ), .A2(_00598_ ), .A3(_01407_ ), .ZN(_01420_ ) );
OAI21_X1 _17286_ ( .A(_01408_ ), .B1(_01419_ ), .B2(_01420_ ), .ZN(_01421_ ) );
OAI21_X1 _17287_ ( .A(_01421_ ), .B1(_01375_ ), .B2(_01404_ ), .ZN(_01422_ ) );
MUX2_X1 _17288_ ( .A(\EX_LS_result_reg [12] ), .B(_01422_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
AOI211_X1 _17289_ ( .A(_06130_ ), .B(_01382_ ), .C1(_00561_ ), .C2(_00563_ ), .ZN(_01423_ ) );
OAI21_X1 _17290_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01423_ ), .ZN(_01424_ ) );
OAI21_X1 _17291_ ( .A(_01424_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01425_ ) );
MUX2_X1 _17292_ ( .A(\EX_LS_result_reg [30] ), .B(_01425_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
AND4_X1 _17293_ ( .A1(\io_master_arid [1] ), .A2(_00641_ ), .A3(_00643_ ), .A4(_01406_ ), .ZN(_01426_ ) );
AND3_X1 _17294_ ( .A1(_00602_ ), .A2(_00604_ ), .A3(_01407_ ), .ZN(_01427_ ) );
OAI21_X1 _17295_ ( .A(_01408_ ), .B1(_01426_ ), .B2(_01427_ ), .ZN(_01428_ ) );
OAI21_X1 _17296_ ( .A(_01428_ ), .B1(_01375_ ), .B2(_01404_ ), .ZN(_01429_ ) );
MUX2_X1 _17297_ ( .A(\EX_LS_result_reg [11] ), .B(_01429_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
NAND3_X1 _17298_ ( .A1(_00605_ ), .A2(_00607_ ), .A3(_01409_ ), .ZN(_01430_ ) );
NOR2_X1 _17299_ ( .A1(_00646_ ), .A2(_06169_ ), .ZN(_01431_ ) );
NAND2_X1 _17300_ ( .A1(_01431_ ), .A2(_01406_ ), .ZN(_01432_ ) );
OAI211_X1 _17301_ ( .A(_01430_ ), .B(_01432_ ), .C1(_01375_ ), .C2(_01404_ ), .ZN(_01433_ ) );
MUX2_X1 _17302_ ( .A(\EX_LS_result_reg [10] ), .B(_01433_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
NAND3_X1 _17303_ ( .A1(_00608_ ), .A2(_00610_ ), .A3(_01409_ ), .ZN(_01434_ ) );
NAND4_X1 _17304_ ( .A1(_00647_ ), .A2(_00649_ ), .A3(\io_master_arid [1] ), .A4(_01406_ ), .ZN(_01435_ ) );
OAI211_X1 _17305_ ( .A(_01434_ ), .B(_01435_ ), .C1(_01375_ ), .C2(_01365_ ), .ZN(_01436_ ) );
MUX2_X1 _17306_ ( .A(\EX_LS_result_reg [9] ), .B(_01436_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NAND3_X1 _17307_ ( .A1(_00611_ ), .A2(_00613_ ), .A3(_01409_ ), .ZN(_01437_ ) );
NOR2_X1 _17308_ ( .A1(_00652_ ), .A2(_06131_ ), .ZN(_01438_ ) );
NAND2_X1 _17309_ ( .A1(_01438_ ), .A2(_01406_ ), .ZN(_01439_ ) );
OAI211_X1 _17310_ ( .A(_01437_ ), .B(_01439_ ), .C1(_01375_ ), .C2(_01365_ ), .ZN(_01440_ ) );
MUX2_X1 _17311_ ( .A(\EX_LS_result_reg [8] ), .B(_01440_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
OR3_X4 _17312_ ( .A1(_01374_ ), .A2(\mylsu.typ_tmp [2] ), .A3(_01347_ ), .ZN(_01441_ ) );
AND2_X1 _17313_ ( .A1(_00616_ ), .A2(_06211_ ), .ZN(_01442_ ) );
MUX2_X1 _17314_ ( .A(_01442_ ), .B(_01369_ ), .S(_01406_ ), .Z(_01443_ ) );
OAI21_X1 _17315_ ( .A(_01443_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01347_ ), .ZN(_01444_ ) );
AOI21_X1 _17316_ ( .A(_01346_ ), .B1(_01441_ ), .B2(_01444_ ), .ZN(_01445_ ) );
NOR2_X1 _17317_ ( .A1(_01374_ ), .A2(_01365_ ), .ZN(_01446_ ) );
OR2_X2 _17318_ ( .A1(_01445_ ), .A2(_01446_ ), .ZN(_01447_ ) );
MUX2_X2 _17319_ ( .A(\EX_LS_result_reg [7] ), .B(_01447_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _17320_ ( .A1(_01242_ ), .A2(\EX_LS_result_reg [6] ), .ZN(_01448_ ) );
NOR2_X1 _17321_ ( .A1(_01401_ ), .A2(_01350_ ), .ZN(_01449_ ) );
INV_X1 _17322_ ( .A(_01449_ ), .ZN(_01450_ ) );
AND2_X1 _17323_ ( .A1(_01349_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01451_ ) );
NOR2_X1 _17324_ ( .A1(_01450_ ), .A2(_01451_ ), .ZN(_01452_ ) );
AOI211_X1 _17325_ ( .A(_01242_ ), .B(_06169_ ), .C1(_01203_ ), .C2(_01452_ ), .ZN(_01453_ ) );
NAND2_X1 _17326_ ( .A1(_00619_ ), .A2(_01450_ ), .ZN(_01454_ ) );
NAND2_X1 _17327_ ( .A1(_01453_ ), .A2(_01454_ ), .ZN(_01455_ ) );
NAND3_X1 _17328_ ( .A1(_00588_ ), .A2(_00592_ ), .A3(_06170_ ), .ZN(_01456_ ) );
OR2_X1 _17329_ ( .A1(_00745_ ), .A2(_06170_ ), .ZN(_01457_ ) );
AND3_X1 _17330_ ( .A1(_01456_ ), .A2(_01451_ ), .A3(_01457_ ), .ZN(_01458_ ) );
OAI21_X1 _17331_ ( .A(_01448_ ), .B1(_01455_ ), .B2(_01458_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _17332_ ( .A(_01416_ ), .B(_01362_ ), .S(_01370_ ), .Z(_01459_ ) );
MUX2_X1 _17333_ ( .A(_01459_ ), .B(_01414_ ), .S(_01368_ ), .Z(_01460_ ) );
NOR2_X2 _17334_ ( .A1(_01460_ ), .A2(_01350_ ), .ZN(_01461_ ) );
NOR3_X2 _17335_ ( .A1(_00622_ ), .A2(_06129_ ), .A3(_01351_ ), .ZN(_01462_ ) );
OAI21_X1 _17336_ ( .A(_01346_ ), .B1(_01461_ ), .B2(_01462_ ), .ZN(_01463_ ) );
OAI21_X1 _17337_ ( .A(_01348_ ), .B1(_01461_ ), .B2(_01462_ ), .ZN(_01464_ ) );
NOR3_X1 _17338_ ( .A1(_00566_ ), .A2(_06130_ ), .A3(_01350_ ), .ZN(_01465_ ) );
OAI21_X1 _17339_ ( .A(_01382_ ), .B1(_01465_ ), .B2(_01462_ ), .ZN(_01466_ ) );
OR3_X1 _17340_ ( .A1(_00622_ ), .A2(_06130_ ), .A3(_01382_ ), .ZN(_01467_ ) );
AOI21_X1 _17341_ ( .A(_01357_ ), .B1(_01466_ ), .B2(_01467_ ), .ZN(_01468_ ) );
INV_X1 _17342_ ( .A(_01465_ ), .ZN(_01469_ ) );
INV_X1 _17343_ ( .A(_01462_ ), .ZN(_01470_ ) );
AOI21_X1 _17344_ ( .A(_01358_ ), .B1(_01469_ ), .B2(_01470_ ), .ZN(_01471_ ) );
OAI22_X1 _17345_ ( .A1(_01468_ ), .A2(_01471_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01347_ ), .ZN(_01472_ ) );
AND2_X2 _17346_ ( .A1(_01464_ ), .A2(_01472_ ), .ZN(_01473_ ) );
OAI21_X1 _17347_ ( .A(_01463_ ), .B1(_01473_ ), .B2(_01346_ ), .ZN(_01474_ ) );
MUX2_X1 _17348_ ( .A(\EX_LS_result_reg [5] ), .B(_01474_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
AOI221_X4 _17349_ ( .A(_01242_ ), .B1(_00787_ ), .B2(_01452_ ), .C1(_00625_ ), .C2(_01450_ ), .ZN(_01475_ ) );
AND3_X1 _17350_ ( .A1(_00632_ ), .A2(_00634_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01476_ ) );
OAI21_X1 _17351_ ( .A(_01451_ ), .B1(_00919_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01477_ ) );
OAI211_X1 _17352_ ( .A(_01475_ ), .B(\io_master_arid [1] ), .C1(_01476_ ), .C2(_01477_ ), .ZN(_01478_ ) );
NAND2_X1 _17353_ ( .A1(_01242_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_01479_ ) );
NAND2_X1 _17354_ ( .A1(_01478_ ), .A2(_01479_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
AOI221_X4 _17355_ ( .A(_01241_ ), .B1(_00803_ ), .B2(_01452_ ), .C1(_00628_ ), .C2(_01450_ ), .ZN(_01480_ ) );
AND3_X1 _17356_ ( .A1(_00641_ ), .A2(_00643_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01481_ ) );
NAND3_X1 _17357_ ( .A1(_00602_ ), .A2(_00604_ ), .A3(_06170_ ), .ZN(_01482_ ) );
NAND2_X1 _17358_ ( .A1(_01482_ ), .A2(_01451_ ), .ZN(_01483_ ) );
OAI211_X1 _17359_ ( .A(_01480_ ), .B(\io_master_arid [1] ), .C1(_01481_ ), .C2(_01483_ ), .ZN(_01484_ ) );
NAND2_X1 _17360_ ( .A1(_01242_ ), .A2(\EX_LS_result_reg [3] ), .ZN(_01485_ ) );
NAND2_X1 _17361_ ( .A1(_01484_ ), .A2(_01485_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
NOR4_X1 _17362_ ( .A1(_00578_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(_06170_ ), .A4(_06129_ ), .ZN(_01486_ ) );
NOR3_X1 _17363_ ( .A1(_00646_ ), .A2(_06129_ ), .A3(_01370_ ), .ZN(_01487_ ) );
OAI22_X1 _17364_ ( .A1(_01486_ ), .A2(_01487_ ), .B1(_06174_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01488_ ) );
NAND4_X1 _17365_ ( .A1(_00605_ ), .A2(_00607_ ), .A3(_06211_ ), .A4(_01368_ ), .ZN(_01489_ ) );
AOI21_X1 _17366_ ( .A(_01350_ ), .B1(_01488_ ), .B2(_01489_ ), .ZN(_01490_ ) );
NOR3_X1 _17367_ ( .A1(_00631_ ), .A2(_06129_ ), .A3(_01351_ ), .ZN(_01491_ ) );
OAI21_X1 _17368_ ( .A(_01346_ ), .B1(_01490_ ), .B2(_01491_ ), .ZN(_01492_ ) );
OAI21_X1 _17369_ ( .A(_01348_ ), .B1(_01490_ ), .B2(_01491_ ), .ZN(_01493_ ) );
NOR3_X1 _17370_ ( .A1(_00578_ ), .A2(_06130_ ), .A3(_01350_ ), .ZN(_01494_ ) );
OAI21_X1 _17371_ ( .A(_01382_ ), .B1(_01494_ ), .B2(_01491_ ), .ZN(_01495_ ) );
OR3_X1 _17372_ ( .A1(_00631_ ), .A2(_06130_ ), .A3(_01381_ ), .ZN(_01496_ ) );
AOI21_X1 _17373_ ( .A(_01357_ ), .B1(_01495_ ), .B2(_01496_ ), .ZN(_01497_ ) );
INV_X1 _17374_ ( .A(_01494_ ), .ZN(_01498_ ) );
INV_X1 _17375_ ( .A(_01491_ ), .ZN(_01499_ ) );
AOI21_X1 _17376_ ( .A(_01358_ ), .B1(_01498_ ), .B2(_01499_ ), .ZN(_01500_ ) );
OAI22_X1 _17377_ ( .A1(_01497_ ), .A2(_01500_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01347_ ), .ZN(_01501_ ) );
AND2_X1 _17378_ ( .A1(_01493_ ), .A2(_01501_ ), .ZN(_01502_ ) );
OAI21_X1 _17379_ ( .A(_01492_ ), .B1(_01502_ ), .B2(_01346_ ), .ZN(_01503_ ) );
MUX2_X1 _17380_ ( .A(\EX_LS_result_reg [2] ), .B(_01503_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
NOR3_X1 _17381_ ( .A1(_00601_ ), .A2(_06131_ ), .A3(_01360_ ), .ZN(_01504_ ) );
OAI21_X1 _17382_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01504_ ), .ZN(_01505_ ) );
OAI21_X1 _17383_ ( .A(_01505_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01506_ ) );
MUX2_X1 _17384_ ( .A(\EX_LS_result_reg [29] ), .B(_01506_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
AOI221_X4 _17385_ ( .A(_01241_ ), .B1(_00841_ ), .B2(_01452_ ), .C1(_00637_ ), .C2(_01450_ ), .ZN(_01507_ ) );
AND3_X1 _17386_ ( .A1(_00647_ ), .A2(_00649_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01508_ ) );
OAI21_X1 _17387_ ( .A(_01451_ ), .B1(_00978_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01509_ ) );
OAI211_X1 _17388_ ( .A(_01507_ ), .B(\io_master_arid [1] ), .C1(_01508_ ), .C2(_01509_ ), .ZN(_01510_ ) );
NAND2_X1 _17389_ ( .A1(_01242_ ), .A2(\EX_LS_result_reg [1] ), .ZN(_01511_ ) );
NAND2_X1 _17390_ ( .A1(_01510_ ), .A2(_01511_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
NOR4_X1 _17391_ ( .A1(_00584_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(_06170_ ), .A4(_06129_ ), .ZN(_01512_ ) );
NOR3_X1 _17392_ ( .A1(_00652_ ), .A2(_06129_ ), .A3(_01370_ ), .ZN(_01513_ ) );
OAI22_X1 _17393_ ( .A1(_01512_ ), .A2(_01513_ ), .B1(_06174_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01514_ ) );
NAND4_X1 _17394_ ( .A1(_00611_ ), .A2(_00613_ ), .A3(_06211_ ), .A4(_01368_ ), .ZN(_01515_ ) );
AOI21_X1 _17395_ ( .A(_01350_ ), .B1(_01514_ ), .B2(_01515_ ), .ZN(_01516_ ) );
NOR3_X1 _17396_ ( .A1(_00640_ ), .A2(_06129_ ), .A3(_01351_ ), .ZN(_01517_ ) );
OAI21_X1 _17397_ ( .A(_01346_ ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01518_ ) );
OAI21_X1 _17398_ ( .A(_01348_ ), .B1(_01516_ ), .B2(_01517_ ), .ZN(_01519_ ) );
NOR3_X1 _17399_ ( .A1(_00584_ ), .A2(_06129_ ), .A3(_01350_ ), .ZN(_01520_ ) );
OAI21_X1 _17400_ ( .A(_01382_ ), .B1(_01520_ ), .B2(_01517_ ), .ZN(_01521_ ) );
OR3_X1 _17401_ ( .A1(_00640_ ), .A2(_06130_ ), .A3(_01381_ ), .ZN(_01522_ ) );
AOI21_X1 _17402_ ( .A(_01357_ ), .B1(_01521_ ), .B2(_01522_ ), .ZN(_01523_ ) );
INV_X1 _17403_ ( .A(_01520_ ), .ZN(_01524_ ) );
INV_X1 _17404_ ( .A(_01517_ ), .ZN(_01525_ ) );
AOI21_X1 _17405_ ( .A(_01358_ ), .B1(_01524_ ), .B2(_01525_ ), .ZN(_01526_ ) );
OAI22_X1 _17406_ ( .A1(_01523_ ), .A2(_01526_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01347_ ), .ZN(_01527_ ) );
AND2_X1 _17407_ ( .A1(_01519_ ), .A2(_01527_ ), .ZN(_01528_ ) );
OAI21_X1 _17408_ ( .A(_01518_ ), .B1(_01528_ ), .B2(_01346_ ), .ZN(_01529_ ) );
MUX2_X1 _17409_ ( .A(\EX_LS_result_reg [0] ), .B(_01529_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
AND4_X1 _17410_ ( .A1(_06211_ ), .A2(_00632_ ), .A3(_00634_ ), .A4(_01361_ ), .ZN(_01530_ ) );
OAI21_X1 _17411_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01530_ ), .ZN(_01531_ ) );
OAI21_X1 _17412_ ( .A(_01531_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01532_ ) );
MUX2_X1 _17413_ ( .A(\EX_LS_result_reg [28] ), .B(_01532_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
NOR2_X1 _17414_ ( .A1(_01446_ ), .A2(_01242_ ), .ZN(_01533_ ) );
NOR3_X1 _17415_ ( .A1(_01128_ ), .A2(_06169_ ), .A3(_01382_ ), .ZN(_01534_ ) );
OAI21_X1 _17416_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01534_ ), .ZN(_01535_ ) );
AOI22_X1 _17417_ ( .A1(_01533_ ), .A2(_01535_ ), .B1(_01242_ ), .B2(_04607_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
NOR3_X1 _17418_ ( .A1(_00646_ ), .A2(_06131_ ), .A3(_01360_ ), .ZN(_01536_ ) );
OAI21_X1 _17419_ ( .A(_01377_ ), .B1(_01357_ ), .B2(_01536_ ), .ZN(_01537_ ) );
OAI21_X1 _17420_ ( .A(_01537_ ), .B1(_01366_ ), .B2(_01389_ ), .ZN(_01538_ ) );
MUX2_X1 _17421_ ( .A(\EX_LS_result_reg [26] ), .B(_01538_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
AND4_X1 _17422_ ( .A1(\io_master_arid [1] ), .A2(_00647_ ), .A3(_00649_ ), .A4(_01361_ ), .ZN(_01539_ ) );
OAI21_X1 _17423_ ( .A(_01378_ ), .B1(_01379_ ), .B2(_01539_ ), .ZN(_01540_ ) );
AOI22_X1 _17424_ ( .A1(_01533_ ), .A2(_01540_ ), .B1(_01242_ ), .B2(_04631_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
NOR3_X1 _17425_ ( .A1(_00652_ ), .A2(_06131_ ), .A3(_01360_ ), .ZN(_01541_ ) );
OAI21_X1 _17426_ ( .A(_01377_ ), .B1(_01357_ ), .B2(_01541_ ), .ZN(_01542_ ) );
OAI21_X1 _17427_ ( .A(_01542_ ), .B1(_01404_ ), .B2(_01389_ ), .ZN(_01543_ ) );
MUX2_X1 _17428_ ( .A(\EX_LS_result_reg [24] ), .B(_01543_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _17429_ ( .A1(_00655_ ), .A2(_06131_ ), .A3(_01360_ ), .ZN(_01544_ ) );
OAI21_X1 _17430_ ( .A(_01377_ ), .B1(_01357_ ), .B2(_01544_ ), .ZN(_01545_ ) );
OAI21_X1 _17431_ ( .A(_01545_ ), .B1(_01404_ ), .B2(_01389_ ), .ZN(_01546_ ) );
MUX2_X1 _17432_ ( .A(\EX_LS_result_reg [23] ), .B(_01546_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _17433_ ( .A1(_01203_ ), .A2(_06131_ ), .A3(_01382_ ), .ZN(_01547_ ) );
OAI21_X1 _17434_ ( .A(_01377_ ), .B1(_01357_ ), .B2(_01547_ ), .ZN(_01548_ ) );
OAI21_X1 _17435_ ( .A(_01548_ ), .B1(_01404_ ), .B2(_01374_ ), .ZN(_01549_ ) );
MUX2_X1 _17436_ ( .A(\EX_LS_result_reg [22] ), .B(_01549_ ), .S(fanout_net_45 ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17437_ ( .A1(_00560_ ), .A2(\io_master_arid [1] ), .A3(_01361_ ), .ZN(_01550_ ) );
OAI21_X1 _17438_ ( .A(_01377_ ), .B1(_01357_ ), .B2(_01550_ ), .ZN(_01551_ ) );
OAI21_X1 _17439_ ( .A(_01551_ ), .B1(_01404_ ), .B2(_01374_ ), .ZN(_01552_ ) );
MUX2_X1 _17440_ ( .A(\EX_LS_result_reg [31] ), .B(_01552_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17441_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(\LS_WB_waddr_reg [2] ), .ZN(_01553_ ) );
INV_X1 _17442_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01554_ ) );
INV_X1 _17443_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01555_ ) );
NAND3_X1 _17444_ ( .A1(_01553_ ), .A2(_01554_ ), .A3(_01555_ ), .ZN(_01556_ ) );
AND2_X1 _17445_ ( .A1(_01585_ ), .A2(LS_WB_wen_reg ), .ZN(_01557_ ) );
NAND2_X1 _17446_ ( .A1(_01556_ ), .A2(_01557_ ), .ZN(_01558_ ) );
BUF_X4 _17447_ ( .A(_01558_ ), .Z(_01559_ ) );
INV_X1 _17448_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01560_ ) );
INV_X1 _17449_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01561_ ) );
AOI21_X1 _17450_ ( .A(_01559_ ), .B1(_01560_ ), .B2(_01561_ ), .ZN(_01562_ ) );
NOR4_X1 _17451_ ( .A1(_01562_ ), .A2(_01554_ ), .A3(_01555_ ), .A4(_01559_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
AOI21_X1 _17452_ ( .A(_01559_ ), .B1(_01554_ ), .B2(_01555_ ), .ZN(_01563_ ) );
NOR2_X1 _17453_ ( .A1(_01558_ ), .A2(_01560_ ), .ZN(_01564_ ) );
NOR4_X1 _17454_ ( .A1(_01563_ ), .A2(_01564_ ), .A3(_01561_ ), .A4(_01559_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
NOR2_X1 _17455_ ( .A1(_01558_ ), .A2(_01554_ ), .ZN(_01565_ ) );
AND4_X1 _17456_ ( .A1(_01561_ ), .A2(_01565_ ), .A3(_01564_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
NOR2_X1 _17457_ ( .A1(_01559_ ), .A2(_01561_ ), .ZN(_01566_ ) );
NOR4_X1 _17458_ ( .A1(_01563_ ), .A2(_01566_ ), .A3(_01560_ ), .A4(_01559_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
NOR2_X1 _17459_ ( .A1(_01559_ ), .A2(_01555_ ), .ZN(_01567_ ) );
AND4_X1 _17460_ ( .A1(_01561_ ), .A2(_01567_ ), .A3(_01564_ ), .A4(_01554_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
CLKBUF_X1 _17461_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
NOR4_X1 _17462_ ( .A1(_01562_ ), .A2(_01565_ ), .A3(_01555_ ), .A4(_01559_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
AND4_X1 _17463_ ( .A1(_01560_ ), .A2(_01567_ ), .A3(_01566_ ), .A4(_01554_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17464_ ( .A1(_01560_ ), .A2(_01565_ ), .A3(_01566_ ), .A4(_01555_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
AND4_X1 _17465_ ( .A1(_01560_ ), .A2(_01565_ ), .A3(_01566_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
NOR4_X1 _17466_ ( .A1(_01563_ ), .A2(_01560_ ), .A3(_01561_ ), .A4(_01559_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17467_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01567_ ), .A3(_01564_ ), .A4(_01554_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17468_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01565_ ), .A3(_01564_ ), .A4(_01555_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17469_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01567_ ), .A3(_01564_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
AND4_X1 _17470_ ( .A1(_01561_ ), .A2(_01565_ ), .A3(_01564_ ), .A4(_01555_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
NOR4_X1 _17471_ ( .A1(_01562_ ), .A2(_01567_ ), .A3(_01554_ ), .A4(_01559_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17472_ ( .A1(_02053_ ), .A2(_01748_ ), .A3(_02060_ ), .ZN(_01568_ ) );
NAND2_X1 _17473_ ( .A1(_01568_ ), .A2(_01748_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17474_ ( .A(reset ), .B(_02053_ ), .C1(_02054_ ), .C2(_06205_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17475_ ( .A(_01556_ ), .Z(_01569_ ) );
CLKBUF_X2 _17476_ ( .A(_01557_ ), .Z(_01570_ ) );
AND3_X1 _17477_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17478_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17479_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17480_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17481_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17482_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17483_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17484_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17485_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17486_ ( .A1(_01569_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01570_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17487_ ( .A(_01556_ ), .Z(_01571_ ) );
CLKBUF_X2 _17488_ ( .A(_01557_ ), .Z(_01572_ ) );
AND3_X1 _17489_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17490_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17491_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17492_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17493_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17494_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17495_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17496_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17497_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17498_ ( .A1(_01571_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01572_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17499_ ( .A(_01556_ ), .Z(_01573_ ) );
CLKBUF_X2 _17500_ ( .A(_01557_ ), .Z(_01574_ ) );
AND3_X1 _17501_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17502_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17503_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17504_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17505_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17506_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17507_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17508_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17509_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17510_ ( .A1(_01573_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01574_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17511_ ( .A1(_01556_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01557_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17512_ ( .A1(_01556_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01557_ ), .ZN(\myreg.Reg[1]_$_DFFE_PP__Q_D ) );
AND3_X1 _17513_ ( .A1(_01748_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17514_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01575_ ) );
AND2_X1 _17515_ ( .A1(_01575_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01576_ ) );
INV_X1 _17516_ ( .A(_01576_ ), .ZN(_01577_ ) );
NOR2_X1 _17517_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01578_ ) );
OAI211_X1 _17518_ ( .A(_01586_ ), .B(\mysc.state [0] ), .C1(_01577_ ), .C2(_01578_ ), .ZN(_01579_ ) );
INV_X1 _17519_ ( .A(_01579_ ), .ZN(_01580_ ) );
OR3_X1 _17520_ ( .A1(_01580_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17521_ ( .A1(_01577_ ), .A2(reset ), .A3(_01578_ ), .ZN(_01581_ ) );
NAND2_X1 _17522_ ( .A1(_01581_ ), .A2(\mysc.state [0] ), .ZN(_01582_ ) );
OR3_X1 _17523_ ( .A1(_04013_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01583_ ) );
NAND2_X1 _17524_ ( .A1(_01582_ ), .A2(_01583_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17525_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07996_ ) );
CLKGATE_X1 _17526_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_07997_ ) );
CLKGATE_X1 _17527_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07998_ ) );
CLKGATE_X1 _17528_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07999_ ) );
CLKGATE_X1 _17529_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_08000_ ) );
CLKGATE_X1 _17530_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_08001_ ) );
CLKGATE_X1 _17531_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_08002_ ) );
CLKGATE_X1 _17532_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_08003_ ) );
CLKGATE_X1 _17533_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_08004_ ) );
CLKGATE_X1 _17534_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_08005_ ) );
CLKGATE_X1 _17535_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_08006_ ) );
CLKGATE_X1 _17536_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_08007_ ) );
CLKGATE_X1 _17537_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_08008_ ) );
CLKGATE_X1 _17538_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_08009_ ) );
CLKGATE_X1 _17539_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_08010_ ) );
CLKGATE_X1 _17540_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_08011_ ) );
CLKGATE_X1 _17541_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_08012_ ) );
CLKGATE_X1 _17542_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08013_ ) );
CLKGATE_X1 _17543_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_08014_ ) );
CLKGATE_X1 _17544_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PN0P__Q_E ), .GCK(_08015_ ) );
CLKGATE_X1 _17545_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PN0P__Q_E ), .GCK(_08016_ ) );
CLKGATE_X1 _17546_ ( .CK(clock ), .E(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_08017_ ) );
CLKGATE_X1 _17547_ ( .CK(clock ), .E(\myexu.rst_logic_$_OR__B_A_$_ANDNOT__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__A_B_$_ANDNOT__B_Y ), .GCK(_08018_ ) );
CLKGATE_X1 _17548_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_08019_ ) );
CLKGATE_X1 _17549_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_08020_ ) );
CLKGATE_X1 _17550_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_08021_ ) );
CLKGATE_X1 _17551_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_08022_ ) );
CLKGATE_X1 _17552_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_08023_ ) );
CLKGATE_X1 _17553_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_08024_ ) );
CLKGATE_X1 _17554_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_08025_ ) );
CLKGATE_X1 _17555_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_08026_ ) );
CLKGATE_X1 _17556_ ( .CK(clock ), .E(\myifu.myicache.tag[3]_$_DFFE_PP__Q_E ), .GCK(_08027_ ) );
CLKGATE_X1 _17557_ ( .CK(clock ), .E(\myifu.myicache.tag[2]_$_DFFE_PP__Q_E ), .GCK(_08028_ ) );
CLKGATE_X1 _17558_ ( .CK(clock ), .E(\myifu.myicache.tag[1]_$_DFFE_PP__Q_E ), .GCK(_08029_ ) );
CLKGATE_X1 _17559_ ( .CK(clock ), .E(\myifu.myicache.tag[0]_$_DFFE_PP__Q_E ), .GCK(_08030_ ) );
CLKGATE_X1 _17560_ ( .CK(clock ), .E(\myifu.myicache.data[7]_$_DFFE_PP__Q_E ), .GCK(_08031_ ) );
CLKGATE_X1 _17561_ ( .CK(clock ), .E(\myifu.myicache.data[6]_$_DFFE_PP__Q_E ), .GCK(_08032_ ) );
CLKGATE_X1 _17562_ ( .CK(clock ), .E(\myifu.myicache.data[5]_$_DFFE_PP__Q_E ), .GCK(_08033_ ) );
CLKGATE_X1 _17563_ ( .CK(clock ), .E(\myifu.myicache.data[4]_$_DFFE_PP__Q_E ), .GCK(_08034_ ) );
CLKGATE_X1 _17564_ ( .CK(clock ), .E(\myifu.myicache.data[3]_$_DFFE_PP__Q_E ), .GCK(_08035_ ) );
CLKGATE_X1 _17565_ ( .CK(clock ), .E(\myifu.myicache.data[2]_$_DFFE_PP__Q_E ), .GCK(_08036_ ) );
CLKGATE_X1 _17566_ ( .CK(clock ), .E(\myifu.myicache.data[1]_$_DFFE_PP__Q_E ), .GCK(_08037_ ) );
CLKGATE_X1 _17567_ ( .CK(clock ), .E(\myifu.myicache.data[0]_$_DFFE_PP__Q_E ), .GCK(_08038_ ) );
CLKGATE_X1 _17568_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_08039_ ) );
CLKGATE_X1 _17569_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_08040_ ) );
CLKGATE_X1 _17570_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_08041_ ) );
CLKGATE_X1 _17571_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_08042_ ) );
CLKGATE_X1 _17572_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_08043_ ) );
CLKGATE_X1 _17573_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08044_ ) );
CLKGATE_X1 _17574_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08045_ ) );
CLKGATE_X1 _17575_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08046_ ) );
CLKGATE_X1 _17576_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_08047_ ) );
CLKGATE_X1 _17577_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08048_ ) );
CLKGATE_X1 _17578_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_08049_ ) );
CLKGATE_X1 _17579_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_08050_ ) );
CLKGATE_X1 _17580_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_08051_ ) );
CLKGATE_X1 _17581_ ( .CK(clock ), .E(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_S_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08052_ ) );
CLKGATE_X1 _17582_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y ), .GCK(_08053_ ) );
CLKGATE_X1 _17583_ ( .CK(clock ), .E(\myexu.state_$_ANDNOT__B_Y_$_AND__A_Y ), .GCK(_08054_ ) );
CLKGATE_X1 _17584_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_08055_ ) );
CLKGATE_X1 _17585_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_08056_ ) );
CLKGATE_X1 _17586_ ( .CK(clock ), .E(\mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_E ), .GCK(_08057_ ) );
CLKGATE_X1 _17587_ ( .CK(clock ), .E(\mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_E ), .GCK(_08058_ ) );
CLKGATE_X1 _17588_ ( .CK(clock ), .E(\mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_E ), .GCK(_08059_ ) );
CLKGATE_X1 _17589_ ( .CK(clock ), .E(\mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_E ), .GCK(_08060_ ) );
LOGIC1_X1 _17590_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17591_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00064_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00065_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08389_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08388_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08387_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08386_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08385_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08384_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08383_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08382_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08381_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08380_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08379_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08378_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08377_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08376_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08375_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08374_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08373_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08372_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08371_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08370_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08369_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08368_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08367_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08366_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08365_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08364_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08363_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08362_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08361_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08360_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08359_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08060_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08358_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08059_ ), .Q(\mtvec [31] ), .QN(_08357_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08059_ ), .Q(\mtvec [30] ), .QN(_08356_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08059_ ), .Q(\mtvec [21] ), .QN(_08355_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08059_ ), .Q(\mtvec [20] ), .QN(_08354_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08059_ ), .Q(\mtvec [19] ), .QN(_08353_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08059_ ), .Q(\mtvec [18] ), .QN(_08352_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08059_ ), .Q(\mtvec [17] ), .QN(_08351_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08059_ ), .Q(\mtvec [16] ), .QN(_08350_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08059_ ), .Q(\mtvec [15] ), .QN(_08349_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08059_ ), .Q(\mtvec [14] ), .QN(_08348_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08059_ ), .Q(\mtvec [13] ), .QN(_08347_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08059_ ), .Q(\mtvec [12] ), .QN(_08346_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08059_ ), .Q(\mtvec [29] ), .QN(_08345_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08059_ ), .Q(\mtvec [11] ), .QN(_08344_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08059_ ), .Q(\mtvec [10] ), .QN(_08343_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08059_ ), .Q(\mtvec [9] ), .QN(_08342_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08059_ ), .Q(\mtvec [8] ), .QN(_08341_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08059_ ), .Q(\mtvec [7] ), .QN(_08340_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08059_ ), .Q(\mtvec [6] ), .QN(_08339_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08059_ ), .Q(\mtvec [5] ), .QN(_08338_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08059_ ), .Q(\mtvec [4] ), .QN(_08337_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08059_ ), .Q(\mtvec [3] ), .QN(_08336_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08059_ ), .Q(\mtvec [2] ), .QN(_08335_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08059_ ), .Q(\mtvec [28] ), .QN(_08334_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08059_ ), .Q(\mtvec [1] ), .QN(_08333_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08059_ ), .Q(\mtvec [0] ), .QN(_08332_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08059_ ), .Q(\mtvec [27] ), .QN(_08331_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08059_ ), .Q(\mtvec [26] ), .QN(_08330_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08059_ ), .Q(\mtvec [25] ), .QN(_08329_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08059_ ), .Q(\mtvec [24] ), .QN(_08328_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08059_ ), .Q(\mtvec [23] ), .QN(_08327_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08059_ ), .Q(\mtvec [22] ), .QN(_08326_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q ( .D(_00000_ ), .CK(_08058_ ), .Q(\mepc [31] ), .QN(_08325_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_1 ( .D(_00066_ ), .CK(_08058_ ), .Q(\mepc [30] ), .QN(_08324_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_10 ( .D(_00067_ ), .CK(_08058_ ), .Q(\mepc [21] ), .QN(_08323_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_11 ( .D(_00068_ ), .CK(_08058_ ), .Q(\mepc [20] ), .QN(_08322_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_12 ( .D(_00069_ ), .CK(_08058_ ), .Q(\mepc [19] ), .QN(_08321_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_13 ( .D(_00070_ ), .CK(_08058_ ), .Q(\mepc [18] ), .QN(_08320_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_14 ( .D(_00071_ ), .CK(_08058_ ), .Q(\mepc [17] ), .QN(_08319_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_15 ( .D(_00072_ ), .CK(_08058_ ), .Q(\mepc [16] ), .QN(_08318_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_16 ( .D(_00073_ ), .CK(_08058_ ), .Q(\mepc [15] ), .QN(_08317_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_17 ( .D(_00074_ ), .CK(_08058_ ), .Q(\mepc [14] ), .QN(_08316_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_18 ( .D(_00075_ ), .CK(_08058_ ), .Q(\mepc [13] ), .QN(_08315_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_19 ( .D(_00076_ ), .CK(_08058_ ), .Q(\mepc [12] ), .QN(_08314_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_2 ( .D(_00077_ ), .CK(_08058_ ), .Q(\mepc [29] ), .QN(_08313_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_20 ( .D(_00078_ ), .CK(_08058_ ), .Q(\mepc [11] ), .QN(_08312_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_21 ( .D(_00079_ ), .CK(_08058_ ), .Q(\mepc [10] ), .QN(_08311_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_22 ( .D(_00080_ ), .CK(_08058_ ), .Q(\mepc [9] ), .QN(_08310_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_23 ( .D(_00081_ ), .CK(_08058_ ), .Q(\mepc [8] ), .QN(_08309_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_24 ( .D(_00082_ ), .CK(_08058_ ), .Q(\mepc [7] ), .QN(_08308_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_25 ( .D(_00083_ ), .CK(_08058_ ), .Q(\mepc [6] ), .QN(_08307_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_26 ( .D(_00084_ ), .CK(_08058_ ), .Q(\mepc [5] ), .QN(_08306_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_27 ( .D(_00085_ ), .CK(_08058_ ), .Q(\mepc [4] ), .QN(_08305_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_28 ( .D(_00086_ ), .CK(_08058_ ), .Q(\mepc [3] ), .QN(_08304_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_29 ( .D(_00087_ ), .CK(_08058_ ), .Q(\mepc [2] ), .QN(_08303_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_3 ( .D(_00088_ ), .CK(_08058_ ), .Q(\mepc [28] ), .QN(_08302_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_30 ( .D(_00089_ ), .CK(_08058_ ), .Q(\mepc [1] ), .QN(_08301_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_31 ( .D(_00090_ ), .CK(_08058_ ), .Q(\mepc [0] ), .QN(_08300_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_4 ( .D(_00091_ ), .CK(_08058_ ), .Q(\mepc [27] ), .QN(_08299_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_5 ( .D(_00092_ ), .CK(_08058_ ), .Q(\mepc [26] ), .QN(_08298_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_6 ( .D(_00093_ ), .CK(_08058_ ), .Q(\mepc [25] ), .QN(_08297_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_7 ( .D(_00094_ ), .CK(_08058_ ), .Q(\mepc [24] ), .QN(_08296_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_8 ( .D(_00095_ ), .CK(_08058_ ), .Q(\mepc [23] ), .QN(_08295_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_SDFFE_PP0P__Q_9 ( .D(_00096_ ), .CK(_08058_ ), .Q(\mepc [22] ), .QN(_08294_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q ( .D(_00097_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08293_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_1 ( .D(_00098_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08292_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_10 ( .D(_00099_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08291_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_11 ( .D(_00100_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08290_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_12 ( .D(_00101_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08289_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_13 ( .D(_00102_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08288_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_14 ( .D(_00103_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08287_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_15 ( .D(_00104_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08286_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_16 ( .D(_00105_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08285_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_17 ( .D(_00106_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08284_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_18 ( .D(_00107_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08283_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_19 ( .D(_00108_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08282_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_2 ( .D(_00109_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08281_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_20 ( .D(_00110_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08280_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_21 ( .D(_00111_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08279_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_22 ( .D(_00112_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08278_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_23 ( .D(_00113_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08277_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_24 ( .D(_00114_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08276_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_25 ( .D(_00115_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08275_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_26 ( .D(_00116_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08274_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_27 ( .D(_00117_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08273_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_28 ( .D(_00118_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08272_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_29 ( .D(_00119_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08271_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_3 ( .D(_00120_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08270_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_30 ( .D(_00121_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08269_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_31 ( .D(_00122_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08268_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_4 ( .D(_00123_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08267_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_5 ( .D(_00124_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08266_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_6 ( .D(_00125_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08265_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_7 ( .D(_00126_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08264_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_8 ( .D(_00127_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08263_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFE_PP0P__Q_9 ( .D(_00128_ ), .CK(_08057_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08390_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PP0__Q ( .D(_00129_ ), .CK(clock ), .Q(excp_written ), .QN(_08391_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08262_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08392_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08393_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08394_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08395_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08396_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08397_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08398_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08399_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08400_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08401_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08402_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08403_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08404_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08405_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08406_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08407_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08408_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08409_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08410_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08411_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08412_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08413_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08414_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08415_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08416_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08417_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08418_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08419_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08420_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08421_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_08056_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08261_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00130_ ), .CK(_08055_ ), .Q(\myec.state [1] ), .QN(_08260_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00131_ ), .CK(_08055_ ), .Q(\myec.state [0] ), .QN(_08422_ ) );
DFF_X1 \myexu.check_quest_$_SDFF_PN0__Q ( .D(_00132_ ), .CK(clock ), .Q(check_quest ), .QN(_08423_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08259_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08424_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08425_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08426_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08427_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08428_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08429_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08430_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08431_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08432_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08433_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08258_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00133_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08257_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00134_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08256_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00135_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08255_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00136_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08254_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00137_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08253_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00138_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08252_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00139_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08251_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00140_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08250_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00141_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08249_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00142_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08248_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00143_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08247_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00144_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08246_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00145_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08245_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00146_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08244_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00147_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08243_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00148_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08242_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00149_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08241_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00150_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08240_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00151_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08239_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00152_ ), .CK(_08054_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08238_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q ( .D(_00153_ ), .CK(_08053_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08237_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_1 ( .D(_00154_ ), .CK(_08053_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08236_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_2 ( .D(_00155_ ), .CK(_08053_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08235_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_3 ( .D(_00156_ ), .CK(_08053_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08234_ ) );
DFF_X1 \myexu.dest_reg_$_SDFFE_PN0P__Q_4 ( .D(_00157_ ), .CK(_08053_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08233_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q ( .D(_00158_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [30] ), .QN(_08232_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_1 ( .D(_00159_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [29] ), .QN(_08231_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_10 ( .D(_00160_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [20] ), .QN(_08230_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_11 ( .D(_00161_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [19] ), .QN(_08229_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_12 ( .D(_00162_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [18] ), .QN(_08228_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_13 ( .D(_00163_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [17] ), .QN(_08227_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_14 ( .D(_00164_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [16] ), .QN(_08226_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_15 ( .D(_00165_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [15] ), .QN(_08225_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_16 ( .D(_00166_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [14] ), .QN(_08224_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_17 ( .D(_00167_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [13] ), .QN(_08223_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_18 ( .D(_00168_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [12] ), .QN(_08222_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_19 ( .D(_00169_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [11] ), .QN(_08221_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_2 ( .D(_00170_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [28] ), .QN(_08220_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_20 ( .D(_00171_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [10] ), .QN(_08219_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_21 ( .D(_00172_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [9] ), .QN(_08218_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_22 ( .D(_00173_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [8] ), .QN(_08217_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_23 ( .D(_00174_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [7] ), .QN(_08216_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_24 ( .D(_00175_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [6] ), .QN(_08215_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_25 ( .D(_00176_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [5] ), .QN(_08214_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_26 ( .D(_00177_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [4] ), .QN(_08213_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_27 ( .D(_00178_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [3] ), .QN(_08212_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_28 ( .D(_00179_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [2] ), .QN(_08211_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_29 ( .D(_00180_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [1] ), .QN(_08210_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_3 ( .D(_00181_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [27] ), .QN(_08209_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_30 ( .D(_00182_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [0] ), .QN(_08208_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_4 ( .D(_00183_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [26] ), .QN(_08207_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_5 ( .D(_00184_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [25] ), .QN(_08206_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_6 ( .D(_00185_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [24] ), .QN(_08205_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_7 ( .D(_00186_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [23] ), .QN(_08204_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_8 ( .D(_00187_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [22] ), .QN(_08203_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN0P__Q_9 ( .D(_00188_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [21] ), .QN(_08202_ ) );
DFF_X1 \myexu.pc_jump_$_SDFFE_PN1P__Q ( .D(_00189_ ), .CK(_08052_ ), .Q(\myexu.pc_jump [31] ), .QN(_08201_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q ( .D(_00190_ ), .CK(_08053_ ), .Q(\EX_LS_pc [31] ), .QN(_08200_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_1 ( .D(_00191_ ), .CK(_08053_ ), .Q(\EX_LS_pc [30] ), .QN(_08199_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_10 ( .D(_00192_ ), .CK(_08053_ ), .Q(\EX_LS_pc [21] ), .QN(_08198_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_11 ( .D(_00193_ ), .CK(_08053_ ), .Q(\EX_LS_pc [20] ), .QN(_08197_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_12 ( .D(_00194_ ), .CK(_08053_ ), .Q(\EX_LS_pc [19] ), .QN(_08196_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_13 ( .D(_00195_ ), .CK(_08053_ ), .Q(\EX_LS_pc [18] ), .QN(_08195_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_14 ( .D(_00196_ ), .CK(_08053_ ), .Q(\EX_LS_pc [17] ), .QN(_08194_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_15 ( .D(_00197_ ), .CK(_08053_ ), .Q(\EX_LS_pc [16] ), .QN(_08193_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_16 ( .D(_00198_ ), .CK(_08053_ ), .Q(\EX_LS_pc [15] ), .QN(_08192_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_17 ( .D(_00199_ ), .CK(_08053_ ), .Q(\EX_LS_pc [14] ), .QN(_08191_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_18 ( .D(_00200_ ), .CK(_08053_ ), .Q(\EX_LS_pc [13] ), .QN(_08190_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_19 ( .D(_00201_ ), .CK(_08053_ ), .Q(\EX_LS_pc [12] ), .QN(_08189_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_2 ( .D(_00202_ ), .CK(_08053_ ), .Q(\EX_LS_pc [29] ), .QN(_08188_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_20 ( .D(_00203_ ), .CK(_08053_ ), .Q(\EX_LS_pc [11] ), .QN(_08187_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_21 ( .D(_00204_ ), .CK(_08053_ ), .Q(\EX_LS_pc [10] ), .QN(_08186_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_22 ( .D(_00205_ ), .CK(_08053_ ), .Q(\EX_LS_pc [9] ), .QN(_08185_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_23 ( .D(_00206_ ), .CK(_08053_ ), .Q(\EX_LS_pc [8] ), .QN(_08184_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_24 ( .D(_00207_ ), .CK(_08053_ ), .Q(\EX_LS_pc [7] ), .QN(_08183_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_25 ( .D(_00208_ ), .CK(_08053_ ), .Q(\EX_LS_pc [6] ), .QN(_08182_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_26 ( .D(_00209_ ), .CK(_08053_ ), .Q(\EX_LS_pc [5] ), .QN(_08181_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_27 ( .D(_00210_ ), .CK(_08053_ ), .Q(\EX_LS_pc [4] ), .QN(_08180_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_28 ( .D(_00211_ ), .CK(_08053_ ), .Q(\EX_LS_pc [3] ), .QN(_08179_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_29 ( .D(_00212_ ), .CK(_08053_ ), .Q(\EX_LS_pc [2] ), .QN(_08178_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_3 ( .D(_00213_ ), .CK(_08053_ ), .Q(\EX_LS_pc [28] ), .QN(_08177_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_30 ( .D(_00214_ ), .CK(_08053_ ), .Q(\EX_LS_pc [1] ), .QN(_08176_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_31 ( .D(_00215_ ), .CK(_08053_ ), .Q(\EX_LS_pc [0] ), .QN(_08175_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_4 ( .D(_00216_ ), .CK(_08053_ ), .Q(\EX_LS_pc [27] ), .QN(_08174_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_5 ( .D(_00217_ ), .CK(_08053_ ), .Q(\EX_LS_pc [26] ), .QN(_08173_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_6 ( .D(_00218_ ), .CK(_08053_ ), .Q(\EX_LS_pc [25] ), .QN(_08172_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_7 ( .D(_00219_ ), .CK(_08053_ ), .Q(\EX_LS_pc [24] ), .QN(_08171_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_8 ( .D(_00220_ ), .CK(_08053_ ), .Q(\EX_LS_pc [23] ), .QN(_08170_ ) );
DFF_X1 \myexu.pc_out_$_SDFFE_PN0P__Q_9 ( .D(_00221_ ), .CK(_08053_ ), .Q(\EX_LS_pc [22] ), .QN(_08434_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08435_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08436_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08437_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08438_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08439_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08440_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08441_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08442_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08443_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08444_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08445_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08446_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08447_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08448_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08449_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08450_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08451_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08452_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08453_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08454_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08455_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08456_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08457_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08458_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08459_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08460_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08461_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08462_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08463_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08464_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08465_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_08054_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08466_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_08054_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.state_$_SDFF_PN0__Q ( .D(_00223_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PN0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q ( .D(_00222_ ), .CK(_08053_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_1 ( .D(_00224_ ), .CK(_08053_ ), .Q(\EX_LS_flag [1] ), .QN(_08169_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_2 ( .D(_00225_ ), .CK(_08053_ ), .Q(\EX_LS_flag [0] ), .QN(_08168_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_3 ( .D(_00226_ ), .CK(_08053_ ), .Q(\EX_LS_typ [4] ), .QN(_08167_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_4 ( .D(_00227_ ), .CK(_08053_ ), .Q(\EX_LS_typ [3] ), .QN(_08166_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_5 ( .D(_00228_ ), .CK(_08053_ ), .Q(\EX_LS_typ [2] ), .QN(_08165_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_6 ( .D(_00229_ ), .CK(_08053_ ), .Q(\EX_LS_typ [1] ), .QN(_08164_ ) );
DFF_X1 \myexu.typ_out_$_SDFFE_PN0P__Q_7 ( .D(_00230_ ), .CK(_08053_ ), .Q(\EX_LS_typ [0] ), .QN(_08163_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00231_ ), .CK(_08051_ ), .Q(\ID_EX_csr [11] ), .QN(_08162_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00232_ ), .CK(_08051_ ), .Q(\ID_EX_csr [10] ), .QN(_08161_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00233_ ), .CK(_08051_ ), .Q(\ID_EX_csr [1] ), .QN(_08160_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00234_ ), .CK(_08051_ ), .Q(\ID_EX_csr [0] ), .QN(_08159_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00235_ ), .CK(_08051_ ), .Q(\ID_EX_csr [9] ), .QN(_08158_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00236_ ), .CK(_08051_ ), .Q(\ID_EX_csr [8] ), .QN(_08157_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00237_ ), .CK(_08051_ ), .Q(\ID_EX_csr [7] ), .QN(_08156_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00238_ ), .CK(_08051_ ), .Q(\ID_EX_csr [6] ), .QN(_08155_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00239_ ), .CK(_08051_ ), .Q(\ID_EX_csr [5] ), .QN(_08154_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00240_ ), .CK(_08051_ ), .Q(\ID_EX_csr [4] ), .QN(_08153_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00241_ ), .CK(_08051_ ), .Q(\ID_EX_csr [3] ), .QN(_08152_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00242_ ), .CK(_08051_ ), .Q(\ID_EX_csr [2] ), .QN(_08151_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00243_ ), .CK(_08050_ ), .Q(exception_quest_IDU ), .QN(_08150_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00244_ ), .CK(_08049_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_08048_ ), .Q(\ID_EX_imm [31] ), .QN(_08467_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_08048_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_08048_ ), .Q(\ID_EX_imm [21] ), .QN(_08468_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_08048_ ), .Q(\ID_EX_imm [20] ), .QN(_08469_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_08048_ ), .Q(\ID_EX_imm [19] ), .QN(_08470_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_08048_ ), .Q(\ID_EX_imm [18] ), .QN(_08471_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_08048_ ), .Q(\ID_EX_imm [17] ), .QN(_08472_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_08048_ ), .Q(\ID_EX_imm [16] ), .QN(_08473_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_08048_ ), .Q(\ID_EX_imm [15] ), .QN(_08474_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_08048_ ), .Q(\ID_EX_imm [14] ), .QN(_08475_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_08048_ ), .Q(\ID_EX_imm [13] ), .QN(_08476_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_08048_ ), .Q(\ID_EX_imm [12] ), .QN(_08477_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_08048_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_1_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_08048_ ), .Q(\ID_EX_imm [11] ), .QN(_08478_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_08048_ ), .Q(\ID_EX_imm [10] ), .QN(_08479_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_08048_ ), .Q(\ID_EX_imm [9] ), .QN(_08480_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_08048_ ), .Q(\ID_EX_imm [8] ), .QN(_08481_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_08048_ ), .Q(\ID_EX_imm [7] ), .QN(_08482_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_08048_ ), .Q(\ID_EX_imm [6] ), .QN(_08483_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_08048_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_08048_ ), .Q(\ID_EX_imm [4] ), .QN(_08484_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_08048_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_08048_ ), .Q(\ID_EX_imm [2] ), .QN(_08485_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_08048_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_08048_ ), .Q(\ID_EX_imm [1] ), .QN(_08486_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_08048_ ), .Q(\ID_EX_imm [0] ), .QN(_08487_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_08048_ ), .Q(\ID_EX_imm [27] ), .QN(_08488_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_08048_ ), .Q(\ID_EX_imm [26] ), .QN(_08489_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_08048_ ), .Q(\ID_EX_imm [25] ), .QN(_08490_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_08048_ ), .Q(\ID_EX_imm [24] ), .QN(_08491_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_08048_ ), .Q(\ID_EX_imm [23] ), .QN(_08492_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__B_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_08048_ ), .Q(\ID_EX_imm [22] ), .QN(_08493_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08047_ ), .Q(\ID_EX_pc [31] ), .QN(_08494_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08047_ ), .Q(\ID_EX_pc [30] ), .QN(_08495_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08047_ ), .Q(\ID_EX_pc [21] ), .QN(_08496_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08047_ ), .Q(\ID_EX_pc [20] ), .QN(_08497_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08047_ ), .Q(\ID_EX_pc [19] ), .QN(_08498_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08047_ ), .Q(\ID_EX_pc [18] ), .QN(_08499_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08047_ ), .Q(\ID_EX_pc [17] ), .QN(_08500_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08047_ ), .Q(\ID_EX_pc [16] ), .QN(_08501_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08047_ ), .Q(\ID_EX_pc [15] ), .QN(_08502_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08047_ ), .Q(\ID_EX_pc [14] ), .QN(_08503_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08047_ ), .Q(\ID_EX_pc [13] ), .QN(_08504_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08047_ ), .Q(\ID_EX_pc [12] ), .QN(_08505_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08047_ ), .Q(\ID_EX_pc [29] ), .QN(_08506_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08047_ ), .Q(\ID_EX_pc [11] ), .QN(_08507_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08047_ ), .Q(\ID_EX_pc [10] ), .QN(_08508_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08047_ ), .Q(\ID_EX_pc [9] ), .QN(_08509_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08047_ ), .Q(\ID_EX_pc [8] ), .QN(_08510_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08047_ ), .Q(\ID_EX_pc [7] ), .QN(_08511_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08047_ ), .Q(\ID_EX_pc [6] ), .QN(_08512_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08047_ ), .Q(\ID_EX_pc [5] ), .QN(_08513_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_08047_ ), .Q(\ID_EX_pc [4] ), .QN(_08514_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_08047_ ), .Q(\ID_EX_pc [3] ), .QN(_08515_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_08047_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08047_ ), .Q(\ID_EX_pc [28] ), .QN(_08516_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_08047_ ), .Q(\ID_EX_pc [1] ), .QN(_08517_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_08047_ ), .Q(\ID_EX_pc [0] ), .QN(_08518_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08047_ ), .Q(\ID_EX_pc [27] ), .QN(_08519_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08047_ ), .Q(\ID_EX_pc [26] ), .QN(_08520_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08047_ ), .Q(\ID_EX_pc [25] ), .QN(_08521_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08047_ ), .Q(\ID_EX_pc [24] ), .QN(_08522_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08047_ ), .Q(\ID_EX_pc [23] ), .QN(_08523_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08047_ ), .Q(\ID_EX_pc [22] ), .QN(_08149_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00245_ ), .CK(_08046_ ), .Q(\ID_EX_rd [4] ), .QN(_08148_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00246_ ), .CK(_08046_ ), .Q(\ID_EX_rd [3] ), .QN(_08147_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00247_ ), .CK(_08046_ ), .Q(\ID_EX_rd [2] ), .QN(_08146_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00248_ ), .CK(_08046_ ), .Q(\ID_EX_rd [1] ), .QN(_08145_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00249_ ), .CK(_08046_ ), .Q(\ID_EX_rd [0] ), .QN(_08144_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00250_ ), .CK(_08045_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08143_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00251_ ), .CK(_08045_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08142_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00253_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08140_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00252_ ), .CK(_08045_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08141_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00255_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08138_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00254_ ), .CK(_08045_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08139_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00257_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08136_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00256_ ), .CK(_08045_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08137_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00259_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08134_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00258_ ), .CK(_08044_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08135_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00260_ ), .CK(_08044_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08133_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00262_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08131_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00261_ ), .CK(_08044_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08132_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00264_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08129_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00263_ ), .CK(_08044_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08130_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00266_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08127_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00265_ ), .CK(_08044_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08128_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00268_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08125_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00267_ ), .CK(_08043_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08126_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00269_ ), .CK(_08042_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08124_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08525_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00270_ ), .CK(_08041_ ), .Q(\ID_EX_typ [7] ), .QN(_08524_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00271_ ), .CK(_08041_ ), .Q(\ID_EX_typ [6] ), .QN(_08123_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00272_ ), .CK(_08041_ ), .Q(\ID_EX_typ [5] ), .QN(_08122_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00273_ ), .CK(_08041_ ), .Q(\ID_EX_typ [4] ), .QN(\myexu.check_quest_$_SDFF_PN0__Q_D_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00274_ ), .CK(_08041_ ), .Q(\ID_EX_typ [3] ), .QN(_08121_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00275_ ), .CK(_08041_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00276_ ), .CK(_08041_ ), .Q(\ID_EX_typ [1] ), .QN(_08120_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00277_ ), .CK(_08041_ ), .Q(\ID_EX_typ [0] ), .QN(_08526_ ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_08040_ ), .Q(check_assert ), .QN(_08527_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_08039_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_08039_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_08039_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_08039_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_08039_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_08039_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_08039_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_08039_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_08039_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_08039_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_08039_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_08039_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_08039_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_08039_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_08039_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_08039_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_08039_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_08039_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_08039_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_08039_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_08039_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_08039_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_08039_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_08039_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_08039_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_08039_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_08039_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_08039_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_08039_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_08039_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_08039_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_08039_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08528_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08529_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08530_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08531_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08532_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08533_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08534_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08535_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08536_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08537_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08538_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08539_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08540_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08541_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08542_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08543_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08544_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08545_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08546_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08547_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08548_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08549_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08550_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08551_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08552_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08553_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08554_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08555_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08556_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08557_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08558_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08038_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08559_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08560_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08561_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08562_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08563_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08564_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08565_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08566_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08567_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08037_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08036_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08035_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08034_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08033_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08032_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_08031_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08800_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08801_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08802_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08803_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08804_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08805_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08806_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08807_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08808_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08809_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08030_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08810_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08811_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08812_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08813_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08814_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08815_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08816_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08817_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08818_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08819_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08820_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08821_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08822_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08823_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08824_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08825_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08826_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08827_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08828_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08829_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08830_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08831_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08832_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08833_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08834_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08835_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08836_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08029_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08837_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08838_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08839_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08840_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08841_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08842_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08843_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08844_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08845_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08846_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08847_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08848_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08849_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08850_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08851_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08852_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08853_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08854_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08855_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08856_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08857_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08858_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08859_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08860_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08861_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08862_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08863_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08028_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08864_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08865_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08866_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08867_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08868_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08869_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08870_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08871_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08872_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08873_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08874_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08875_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08876_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08877_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08878_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08879_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08880_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08881_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08882_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08883_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08884_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08885_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08886_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08887_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08888_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08889_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08890_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_08027_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08119_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00278_ ), .CK(_08026_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08118_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00279_ ), .CK(_08025_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08117_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00280_ ), .CK(_08024_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08891_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_08023_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08116_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00281_ ), .CK(_08022_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00282_ ), .CK(_08021_ ), .Q(\IF_ID_pc [30] ), .QN(_08115_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00283_ ), .CK(_08021_ ), .Q(\IF_ID_pc [21] ), .QN(_08114_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00284_ ), .CK(_08021_ ), .Q(\IF_ID_pc [20] ), .QN(_08113_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00285_ ), .CK(_08021_ ), .Q(\IF_ID_pc [19] ), .QN(_08112_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00286_ ), .CK(_08021_ ), .Q(\IF_ID_pc [18] ), .QN(_08111_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00287_ ), .CK(_08021_ ), .Q(\IF_ID_pc [17] ), .QN(_08110_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00288_ ), .CK(_08021_ ), .Q(\IF_ID_pc [16] ), .QN(_08109_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00289_ ), .CK(_08021_ ), .Q(\IF_ID_pc [15] ), .QN(_08108_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00290_ ), .CK(_08021_ ), .Q(\IF_ID_pc [14] ), .QN(_08107_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00291_ ), .CK(_08021_ ), .Q(\IF_ID_pc [13] ), .QN(_08106_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00292_ ), .CK(_08021_ ), .Q(\IF_ID_pc [12] ), .QN(_08105_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00293_ ), .CK(_08021_ ), .Q(\IF_ID_pc [29] ), .QN(_08104_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00294_ ), .CK(_08021_ ), .Q(\IF_ID_pc [11] ), .QN(_08103_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00295_ ), .CK(_08021_ ), .Q(\IF_ID_pc [10] ), .QN(_08102_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00296_ ), .CK(_08021_ ), .Q(\IF_ID_pc [9] ), .QN(_08101_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00297_ ), .CK(_08021_ ), .Q(\IF_ID_pc [8] ), .QN(_08100_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00298_ ), .CK(_08021_ ), .Q(\IF_ID_pc [7] ), .QN(_08099_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00299_ ), .CK(_08021_ ), .Q(\IF_ID_pc [6] ), .QN(_08098_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00300_ ), .CK(_08021_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00301_ ), .CK(_08021_ ), .Q(\IF_ID_pc [4] ), .QN(_08097_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00303_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08096_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00302_ ), .CK(_08021_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00305_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08094_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00304_ ), .CK(_08021_ ), .Q(\IF_ID_pc [2] ), .QN(_08095_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00306_ ), .CK(_08021_ ), .Q(\IF_ID_pc [28] ), .QN(_08093_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00307_ ), .CK(_08021_ ), .Q(\IF_ID_pc [1] ), .QN(_08092_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00308_ ), .CK(_08021_ ), .Q(\IF_ID_pc [27] ), .QN(_08091_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00309_ ), .CK(_08021_ ), .Q(\IF_ID_pc [26] ), .QN(_08090_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00310_ ), .CK(_08021_ ), .Q(\IF_ID_pc [25] ), .QN(_08089_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00311_ ), .CK(_08021_ ), .Q(\IF_ID_pc [24] ), .QN(_08088_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00312_ ), .CK(_08021_ ), .Q(\IF_ID_pc [23] ), .QN(_08087_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00313_ ), .CK(_08021_ ), .Q(\IF_ID_pc [22] ), .QN(_08086_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00314_ ), .CK(_08021_ ), .Q(\IF_ID_pc [31] ), .QN(_08085_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08893_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08084_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00315_ ), .CK(_08020_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08892_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00317_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00316_ ), .CK(_08019_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08083_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08894_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08895_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08896_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08897_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08898_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08899_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08900_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08901_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08902_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08903_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08904_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08905_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08906_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08907_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08908_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08909_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08910_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08911_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08912_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08913_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08914_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08915_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08916_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08917_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08918_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08919_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08920_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08921_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08922_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08923_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08924_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08018_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08925_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08926_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08927_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08928_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08929_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08930_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08931_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08932_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08933_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08934_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08935_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08936_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08937_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08938_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08939_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08940_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08941_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08942_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08943_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08944_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08945_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08946_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08947_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08948_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08949_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08950_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08951_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08952_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08953_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08954_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08955_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08956_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_08017_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08082_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PN0P__Q ( .D(_00318_ ), .CK(_08016_ ), .Q(LS_WB_pc ), .QN(_08081_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PN0P__Q ( .D(_00319_ ), .CK(_08015_ ), .Q(\mylsu.previous_load_done ), .QN(_08957_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08958_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08959_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08960_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(\mylsu.state_$_DFF_P__Q_1_D_$_OR__Y_A_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__Y_B_$_OR__Y_B_$_NAND__A_Y_$_NOR__A_Y_$_ANDNOT__A_B_$_OR__Y_B ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_08018_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_08018_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08961_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_08018_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08080_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00320_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08079_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00321_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08078_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00322_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08077_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00323_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08076_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00324_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08075_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00325_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_08074_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00326_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_08073_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00327_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_08072_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00328_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_08071_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00329_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_08070_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00330_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_08069_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00331_ ), .CK(_08018_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08962_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_08018_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08963_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_08018_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08964_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_08018_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08965_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_08018_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08966_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08967_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08968_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08969_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08970_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08971_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08972_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08973_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08974_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08975_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08976_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08977_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08978_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08979_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08980_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08981_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08982_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08983_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08984_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08985_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08986_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08987_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08988_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08989_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08990_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08991_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08992_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08993_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08994_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08995_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08996_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08997_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_08018_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08998_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08999_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_09000_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_09001_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_09002_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_09003_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_09004_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_09005_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_09006_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_09007_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_09008_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_09009_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_09010_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_09011_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_09012_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_09013_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_09014_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_09015_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_09016_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_09017_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_09018_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_09019_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_09020_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_09021_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_09022_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_09023_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_09024_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_09025_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_09026_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_09027_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_09028_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_09029_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_08014_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_08068_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q ( .D(_00332_ ), .CK(_08013_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_08067_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_1 ( .D(_00333_ ), .CK(_08013_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_08066_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_2 ( .D(_00334_ ), .CK(_08013_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_08065_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_3 ( .D(_00335_ ), .CK(_08013_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_08064_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_4 ( .D(_00336_ ), .CK(_08013_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_08063_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PN0P__Q_5 ( .D(_00337_ ), .CK(_08013_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_08062_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PN0P__Q ( .D(_00338_ ), .CK(_08013_ ), .Q(LS_WB_wen_reg ), .QN(_09030_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_09031_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_09032_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08012_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08011_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08010_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08009_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08008_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08007_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08006_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08005_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08004_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08003_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08002_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08001_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_08000_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07999_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07998_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_1_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_10_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_10_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_11_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_11_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_12_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_12_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_13_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_13_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_14_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_14_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_15_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_16_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_15_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_17_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_16_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_18_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_17_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_19_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_2_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_20_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_18_A_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_21_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_22_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_23_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_22_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_24_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_25_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.pc_jump_$_SDFFE_PN0P__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_26_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_27_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_28_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_29_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_3_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_2_A_$_ANDNOT__Y_A_$_OR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_30_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_31_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_4_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_5_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_6_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_7_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_8_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_8_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[1]_$_DFFE_PP__Q_9_D ), .CK(_07997_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_XOR__Y_9_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00339_ ), .CK(_07996_ ), .Q(loaduse_clear ), .QN(_09033_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_09034_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_09035_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_08061_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\EX_LS_dest_csreg_mem [1] ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(fanout_net_39 ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(fanout_net_39 ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(fanout_net_39 ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(fanout_net_39 ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(fanout_net_39 ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(fanout_net_39 ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_44 ) );
BUF_X8 fanout_buf_45 ( .A(\mylsu.state [3] ), .Z(fanout_net_45 ) );

endmodule
