
module ysyx_23060229_multiplier(

);


endmodule
