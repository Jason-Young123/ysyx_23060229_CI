//Generate the verilog at 2025-09-29T17:35:26 by iSTA.
module ysyx_23060229 (
clock,
reset,
io_interrupt,
io_master_awready,
io_master_awvalid,
io_master_wready,
io_master_wvalid,
io_master_wlast,
io_master_bready,
io_master_bvalid,
io_master_arready,
io_master_arvalid,
io_master_rready,
io_master_rvalid,
io_master_rlast,
io_slave_awready,
io_slave_awvalid,
io_slave_wready,
io_slave_wvalid,
io_slave_wlast,
io_slave_bready,
io_slave_bvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_rready,
io_slave_rvalid,
io_slave_rlast,
io_master_awaddr,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_awburst,
io_master_wdata,
io_master_wstrb,
io_master_bresp,
io_master_bid,
io_master_araddr,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_arburst,
io_master_rresp,
io_master_rdata,
io_master_rid,
io_slave_awaddr,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_awburst,
io_slave_wdata,
io_slave_wstrb,
io_slave_bresp,
io_slave_bid,
io_slave_araddr,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_arburst,
io_slave_rresp,
io_slave_rdata,
io_slave_rid
);

input clock ;
input reset ;
input io_interrupt ;
input io_master_awready ;
output io_master_awvalid ;
input io_master_wready ;
output io_master_wvalid ;
output io_master_wlast ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_arready ;
output io_master_arvalid ;
output io_master_rready ;
input io_master_rvalid ;
input io_master_rlast ;
output io_slave_awready ;
input io_slave_awvalid ;
output io_slave_wready ;
input io_slave_wvalid ;
input io_slave_wlast ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
input io_slave_rready ;
output io_slave_rvalid ;
output io_slave_rlast ;
output [31:0] io_master_awaddr ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
output [1:0] io_master_awburst ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [1:0] io_master_bresp ;
input [3:0] io_master_bid ;
output [31:0] io_master_araddr ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [1:0] io_master_arburst ;
input [1:0] io_master_rresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [31:0] io_slave_awaddr ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
input [1:0] io_slave_awburst ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;
output [1:0] io_slave_bresp ;
output [3:0] io_slave_bid ;
input [31:0] io_slave_araddr ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [1:0] io_slave_arburst ;
output [1:0] io_slave_rresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;

wire clock ;
wire reset ;
wire io_interrupt ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_master_wlast ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_rlast ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire io_slave_wlast ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_rlast ;
wire _00000_ ;
wire _00001_ ;
wire _00002_ ;
wire _00003_ ;
wire _00004_ ;
wire _00005_ ;
wire _00006_ ;
wire _00007_ ;
wire _00008_ ;
wire _00009_ ;
wire _00010_ ;
wire _00011_ ;
wire _00012_ ;
wire _00013_ ;
wire _00014_ ;
wire _00015_ ;
wire _00016_ ;
wire _00017_ ;
wire _00018_ ;
wire _00019_ ;
wire _00020_ ;
wire _00021_ ;
wire _00022_ ;
wire _00023_ ;
wire _00024_ ;
wire _00025_ ;
wire _00026_ ;
wire _00027_ ;
wire _00028_ ;
wire _00029_ ;
wire _00030_ ;
wire _00031_ ;
wire _00032_ ;
wire _00033_ ;
wire _00034_ ;
wire _00035_ ;
wire _00036_ ;
wire _00037_ ;
wire _00038_ ;
wire _00039_ ;
wire _00040_ ;
wire _00041_ ;
wire _00042_ ;
wire _00043_ ;
wire _00044_ ;
wire _00045_ ;
wire _00046_ ;
wire _00047_ ;
wire _00048_ ;
wire _00049_ ;
wire _00050_ ;
wire _00051_ ;
wire _00052_ ;
wire _00053_ ;
wire _00054_ ;
wire _00055_ ;
wire _00056_ ;
wire _00057_ ;
wire _00058_ ;
wire _00059_ ;
wire _00060_ ;
wire _00061_ ;
wire _00062_ ;
wire _00063_ ;
wire _00064_ ;
wire _00065_ ;
wire _00066_ ;
wire _00067_ ;
wire _00068_ ;
wire _00069_ ;
wire _00070_ ;
wire _00071_ ;
wire _00072_ ;
wire _00073_ ;
wire _00074_ ;
wire _00075_ ;
wire _00076_ ;
wire _00077_ ;
wire _00078_ ;
wire _00079_ ;
wire _00080_ ;
wire _00081_ ;
wire _00082_ ;
wire _00083_ ;
wire _00084_ ;
wire _00085_ ;
wire _00086_ ;
wire _00087_ ;
wire _00088_ ;
wire _00089_ ;
wire _00090_ ;
wire _00091_ ;
wire _00092_ ;
wire _00093_ ;
wire _00094_ ;
wire _00095_ ;
wire _00096_ ;
wire _00097_ ;
wire _00098_ ;
wire _00099_ ;
wire _00100_ ;
wire _00101_ ;
wire _00102_ ;
wire _00103_ ;
wire _00104_ ;
wire _00105_ ;
wire _00106_ ;
wire _00107_ ;
wire _00108_ ;
wire _00109_ ;
wire _00110_ ;
wire _00111_ ;
wire _00112_ ;
wire _00113_ ;
wire _00114_ ;
wire _00115_ ;
wire _00116_ ;
wire _00117_ ;
wire _00118_ ;
wire _00119_ ;
wire _00120_ ;
wire _00121_ ;
wire _00122_ ;
wire _00123_ ;
wire _00124_ ;
wire _00125_ ;
wire _00126_ ;
wire _00127_ ;
wire _00128_ ;
wire _00129_ ;
wire _00130_ ;
wire _00131_ ;
wire _00132_ ;
wire _00133_ ;
wire _00134_ ;
wire _00135_ ;
wire _00136_ ;
wire _00137_ ;
wire _00138_ ;
wire _00139_ ;
wire _00140_ ;
wire _00141_ ;
wire _00142_ ;
wire _00143_ ;
wire _00144_ ;
wire _00145_ ;
wire _00146_ ;
wire _00147_ ;
wire _00148_ ;
wire _00149_ ;
wire _00150_ ;
wire _00151_ ;
wire _00152_ ;
wire _00153_ ;
wire _00154_ ;
wire _00155_ ;
wire _00156_ ;
wire _00157_ ;
wire _00158_ ;
wire _00159_ ;
wire _00160_ ;
wire _00161_ ;
wire _00162_ ;
wire _00163_ ;
wire _00164_ ;
wire _00165_ ;
wire _00166_ ;
wire _00167_ ;
wire _00168_ ;
wire _00169_ ;
wire _00170_ ;
wire _00171_ ;
wire _00172_ ;
wire _00173_ ;
wire _00174_ ;
wire _00175_ ;
wire _00176_ ;
wire _00177_ ;
wire _00178_ ;
wire _00179_ ;
wire _00180_ ;
wire _00181_ ;
wire _00182_ ;
wire _00183_ ;
wire _00184_ ;
wire _00185_ ;
wire _00186_ ;
wire _00187_ ;
wire _00188_ ;
wire _00189_ ;
wire _00190_ ;
wire _00191_ ;
wire _00192_ ;
wire _00193_ ;
wire _00194_ ;
wire _00195_ ;
wire _00196_ ;
wire _00197_ ;
wire _00198_ ;
wire _00199_ ;
wire _00200_ ;
wire _00201_ ;
wire _00202_ ;
wire _00203_ ;
wire _00204_ ;
wire _00205_ ;
wire _00206_ ;
wire _00207_ ;
wire _00208_ ;
wire _00209_ ;
wire _00210_ ;
wire _00211_ ;
wire _00212_ ;
wire _00213_ ;
wire _00214_ ;
wire _00215_ ;
wire _00216_ ;
wire _00217_ ;
wire _00218_ ;
wire _00219_ ;
wire _00220_ ;
wire _00221_ ;
wire _00222_ ;
wire _00223_ ;
wire _00224_ ;
wire _00225_ ;
wire _00226_ ;
wire _00227_ ;
wire _00228_ ;
wire _00229_ ;
wire _00230_ ;
wire _00231_ ;
wire _00232_ ;
wire _00233_ ;
wire _00234_ ;
wire _00235_ ;
wire _00236_ ;
wire _00237_ ;
wire _00238_ ;
wire _00239_ ;
wire _00240_ ;
wire _00241_ ;
wire _00242_ ;
wire _00243_ ;
wire _00244_ ;
wire _00245_ ;
wire _00246_ ;
wire _00247_ ;
wire _00248_ ;
wire _00249_ ;
wire _00250_ ;
wire _00251_ ;
wire _00252_ ;
wire _00253_ ;
wire _00254_ ;
wire _00255_ ;
wire _00256_ ;
wire _00257_ ;
wire _00258_ ;
wire _00259_ ;
wire _00260_ ;
wire _00261_ ;
wire _00262_ ;
wire _00263_ ;
wire _00264_ ;
wire _00265_ ;
wire _00266_ ;
wire _00267_ ;
wire _00268_ ;
wire _00269_ ;
wire _00270_ ;
wire _00271_ ;
wire _00272_ ;
wire _00273_ ;
wire _00274_ ;
wire _00275_ ;
wire _00276_ ;
wire _00277_ ;
wire _00278_ ;
wire _00279_ ;
wire _00280_ ;
wire _00281_ ;
wire _00282_ ;
wire _00283_ ;
wire _00284_ ;
wire _00285_ ;
wire _00286_ ;
wire _00287_ ;
wire _00288_ ;
wire _00289_ ;
wire _00290_ ;
wire _00291_ ;
wire _00292_ ;
wire _00293_ ;
wire _00294_ ;
wire _00295_ ;
wire _00296_ ;
wire _00297_ ;
wire _00298_ ;
wire _00299_ ;
wire _00300_ ;
wire _00301_ ;
wire _00302_ ;
wire _00303_ ;
wire _00304_ ;
wire _00305_ ;
wire _00306_ ;
wire _00307_ ;
wire _00308_ ;
wire _00309_ ;
wire _00310_ ;
wire _00311_ ;
wire _00312_ ;
wire _00313_ ;
wire _00314_ ;
wire _00315_ ;
wire _00316_ ;
wire _00317_ ;
wire _00318_ ;
wire _00319_ ;
wire _00320_ ;
wire _00321_ ;
wire _00322_ ;
wire _00323_ ;
wire _00324_ ;
wire _00325_ ;
wire _00326_ ;
wire _00327_ ;
wire _00328_ ;
wire _00329_ ;
wire _00330_ ;
wire _00331_ ;
wire _00332_ ;
wire _00333_ ;
wire _00334_ ;
wire _00335_ ;
wire _00336_ ;
wire _00337_ ;
wire _00338_ ;
wire _00339_ ;
wire _00340_ ;
wire _00341_ ;
wire _00342_ ;
wire _00343_ ;
wire _00344_ ;
wire _00345_ ;
wire _00346_ ;
wire _00347_ ;
wire _00348_ ;
wire _00349_ ;
wire _00350_ ;
wire _00351_ ;
wire _00352_ ;
wire _00353_ ;
wire _00354_ ;
wire _00355_ ;
wire _00356_ ;
wire _00357_ ;
wire _00358_ ;
wire _00359_ ;
wire _00360_ ;
wire _00361_ ;
wire _00362_ ;
wire _00363_ ;
wire _00364_ ;
wire _00365_ ;
wire _00366_ ;
wire _00367_ ;
wire _00368_ ;
wire _00369_ ;
wire _00370_ ;
wire _00371_ ;
wire _00372_ ;
wire _00373_ ;
wire _00374_ ;
wire _00375_ ;
wire _00376_ ;
wire _00377_ ;
wire _00378_ ;
wire _00379_ ;
wire _00380_ ;
wire _00381_ ;
wire _00382_ ;
wire _00383_ ;
wire _00384_ ;
wire _00385_ ;
wire _00386_ ;
wire _00387_ ;
wire _00388_ ;
wire _00389_ ;
wire _00390_ ;
wire _00391_ ;
wire _00392_ ;
wire _00393_ ;
wire _00394_ ;
wire _00395_ ;
wire _00396_ ;
wire _00397_ ;
wire _00398_ ;
wire _00399_ ;
wire _00400_ ;
wire _00401_ ;
wire _00402_ ;
wire _00403_ ;
wire _00404_ ;
wire _00405_ ;
wire _00406_ ;
wire _00407_ ;
wire _00408_ ;
wire _00409_ ;
wire _00410_ ;
wire _00411_ ;
wire _00412_ ;
wire _00413_ ;
wire _00414_ ;
wire _00415_ ;
wire _00416_ ;
wire _00417_ ;
wire _00418_ ;
wire _00419_ ;
wire _00420_ ;
wire _00421_ ;
wire _00422_ ;
wire _00423_ ;
wire _00424_ ;
wire _00425_ ;
wire _00426_ ;
wire _00427_ ;
wire _00428_ ;
wire _00429_ ;
wire _00430_ ;
wire _00431_ ;
wire _00432_ ;
wire _00433_ ;
wire _00434_ ;
wire _00435_ ;
wire _00436_ ;
wire _00437_ ;
wire _00438_ ;
wire _00439_ ;
wire _00440_ ;
wire _00441_ ;
wire _00442_ ;
wire _00443_ ;
wire _00444_ ;
wire _00445_ ;
wire _00446_ ;
wire _00447_ ;
wire _00448_ ;
wire _00449_ ;
wire _00450_ ;
wire _00451_ ;
wire _00452_ ;
wire _00453_ ;
wire _00454_ ;
wire _00455_ ;
wire _00456_ ;
wire _00457_ ;
wire _00458_ ;
wire _00459_ ;
wire _00460_ ;
wire _00461_ ;
wire _00462_ ;
wire _00463_ ;
wire _00464_ ;
wire _00465_ ;
wire _00466_ ;
wire _00467_ ;
wire _00468_ ;
wire _00469_ ;
wire _00470_ ;
wire _00471_ ;
wire _00472_ ;
wire _00473_ ;
wire _00474_ ;
wire _00475_ ;
wire _00476_ ;
wire _00477_ ;
wire _00478_ ;
wire _00479_ ;
wire _00480_ ;
wire _00481_ ;
wire _00482_ ;
wire _00483_ ;
wire _00484_ ;
wire _00485_ ;
wire _00486_ ;
wire _00487_ ;
wire _00488_ ;
wire _00489_ ;
wire _00490_ ;
wire _00491_ ;
wire _00492_ ;
wire _00493_ ;
wire _00494_ ;
wire _00495_ ;
wire _00496_ ;
wire _00497_ ;
wire _00498_ ;
wire _00499_ ;
wire _00500_ ;
wire _00501_ ;
wire _00502_ ;
wire _00503_ ;
wire _00504_ ;
wire _00505_ ;
wire _00506_ ;
wire _00507_ ;
wire _00508_ ;
wire _00509_ ;
wire _00510_ ;
wire _00511_ ;
wire _00512_ ;
wire _00513_ ;
wire _00514_ ;
wire _00515_ ;
wire _00516_ ;
wire _00517_ ;
wire _00518_ ;
wire _00519_ ;
wire _00520_ ;
wire _00521_ ;
wire _00522_ ;
wire _00523_ ;
wire _00524_ ;
wire _00525_ ;
wire _00526_ ;
wire _00527_ ;
wire _00528_ ;
wire _00529_ ;
wire _00530_ ;
wire _00531_ ;
wire _00532_ ;
wire _00533_ ;
wire _00534_ ;
wire _00535_ ;
wire _00536_ ;
wire _00537_ ;
wire _00538_ ;
wire _00539_ ;
wire _00540_ ;
wire _00541_ ;
wire _00542_ ;
wire _00543_ ;
wire _00544_ ;
wire _00545_ ;
wire _00546_ ;
wire _00547_ ;
wire _00548_ ;
wire _00549_ ;
wire _00550_ ;
wire _00551_ ;
wire _00552_ ;
wire _00553_ ;
wire _00554_ ;
wire _00555_ ;
wire _00556_ ;
wire _00557_ ;
wire _00558_ ;
wire _00559_ ;
wire _00560_ ;
wire _00561_ ;
wire _00562_ ;
wire _00563_ ;
wire _00564_ ;
wire _00565_ ;
wire _00566_ ;
wire _00567_ ;
wire _00568_ ;
wire _00569_ ;
wire _00570_ ;
wire _00571_ ;
wire _00572_ ;
wire _00573_ ;
wire _00574_ ;
wire _00575_ ;
wire _00576_ ;
wire _00577_ ;
wire _00578_ ;
wire _00579_ ;
wire _00580_ ;
wire _00581_ ;
wire _00582_ ;
wire _00583_ ;
wire _00584_ ;
wire _00585_ ;
wire _00586_ ;
wire _00587_ ;
wire _00588_ ;
wire _00589_ ;
wire _00590_ ;
wire _00591_ ;
wire _00592_ ;
wire _00593_ ;
wire _00594_ ;
wire _00595_ ;
wire _00596_ ;
wire _00597_ ;
wire _00598_ ;
wire _00599_ ;
wire _00600_ ;
wire _00601_ ;
wire _00602_ ;
wire _00603_ ;
wire _00604_ ;
wire _00605_ ;
wire _00606_ ;
wire _00607_ ;
wire _00608_ ;
wire _00609_ ;
wire _00610_ ;
wire _00611_ ;
wire _00612_ ;
wire _00613_ ;
wire _00614_ ;
wire _00615_ ;
wire _00616_ ;
wire _00617_ ;
wire _00618_ ;
wire _00619_ ;
wire _00620_ ;
wire _00621_ ;
wire _00622_ ;
wire _00623_ ;
wire _00624_ ;
wire _00625_ ;
wire _00626_ ;
wire _00627_ ;
wire _00628_ ;
wire _00629_ ;
wire _00630_ ;
wire _00631_ ;
wire _00632_ ;
wire _00633_ ;
wire _00634_ ;
wire _00635_ ;
wire _00636_ ;
wire _00637_ ;
wire _00638_ ;
wire _00639_ ;
wire _00640_ ;
wire _00641_ ;
wire _00642_ ;
wire _00643_ ;
wire _00644_ ;
wire _00645_ ;
wire _00646_ ;
wire _00647_ ;
wire _00648_ ;
wire _00649_ ;
wire _00650_ ;
wire _00651_ ;
wire _00652_ ;
wire _00653_ ;
wire _00654_ ;
wire _00655_ ;
wire _00656_ ;
wire _00657_ ;
wire _00658_ ;
wire _00659_ ;
wire _00660_ ;
wire _00661_ ;
wire _00662_ ;
wire _00663_ ;
wire _00664_ ;
wire _00665_ ;
wire _00666_ ;
wire _00667_ ;
wire _00668_ ;
wire _00669_ ;
wire _00670_ ;
wire _00671_ ;
wire _00672_ ;
wire _00673_ ;
wire _00674_ ;
wire _00675_ ;
wire _00676_ ;
wire _00677_ ;
wire _00678_ ;
wire _00679_ ;
wire _00680_ ;
wire _00681_ ;
wire _00682_ ;
wire _00683_ ;
wire _00684_ ;
wire _00685_ ;
wire _00686_ ;
wire _00687_ ;
wire _00688_ ;
wire _00689_ ;
wire _00690_ ;
wire _00691_ ;
wire _00692_ ;
wire _00693_ ;
wire _00694_ ;
wire _00695_ ;
wire _00696_ ;
wire _00697_ ;
wire _00698_ ;
wire _00699_ ;
wire _00700_ ;
wire _00701_ ;
wire _00702_ ;
wire _00703_ ;
wire _00704_ ;
wire _00705_ ;
wire _00706_ ;
wire _00707_ ;
wire _00708_ ;
wire _00709_ ;
wire _00710_ ;
wire _00711_ ;
wire _00712_ ;
wire _00713_ ;
wire _00714_ ;
wire _00715_ ;
wire _00716_ ;
wire _00717_ ;
wire _00718_ ;
wire _00719_ ;
wire _00720_ ;
wire _00721_ ;
wire _00722_ ;
wire _00723_ ;
wire _00724_ ;
wire _00725_ ;
wire _00726_ ;
wire _00727_ ;
wire _00728_ ;
wire _00729_ ;
wire _00730_ ;
wire _00731_ ;
wire _00732_ ;
wire _00733_ ;
wire _00734_ ;
wire _00735_ ;
wire _00736_ ;
wire _00737_ ;
wire _00738_ ;
wire _00739_ ;
wire _00740_ ;
wire _00741_ ;
wire _00742_ ;
wire _00743_ ;
wire _00744_ ;
wire _00745_ ;
wire _00746_ ;
wire _00747_ ;
wire _00748_ ;
wire _00749_ ;
wire _00750_ ;
wire _00751_ ;
wire _00752_ ;
wire _00753_ ;
wire _00754_ ;
wire _00755_ ;
wire _00756_ ;
wire _00757_ ;
wire _00758_ ;
wire _00759_ ;
wire _00760_ ;
wire _00761_ ;
wire _00762_ ;
wire _00763_ ;
wire _00764_ ;
wire _00765_ ;
wire _00766_ ;
wire _00767_ ;
wire _00768_ ;
wire _00769_ ;
wire _00770_ ;
wire _00771_ ;
wire _00772_ ;
wire _00773_ ;
wire _00774_ ;
wire _00775_ ;
wire _00776_ ;
wire _00777_ ;
wire _00778_ ;
wire _00779_ ;
wire _00780_ ;
wire _00781_ ;
wire _00782_ ;
wire _00783_ ;
wire _00784_ ;
wire _00785_ ;
wire _00786_ ;
wire _00787_ ;
wire _00788_ ;
wire _00789_ ;
wire _00790_ ;
wire _00791_ ;
wire _00792_ ;
wire _00793_ ;
wire _00794_ ;
wire _00795_ ;
wire _00796_ ;
wire _00797_ ;
wire _00798_ ;
wire _00799_ ;
wire _00800_ ;
wire _00801_ ;
wire _00802_ ;
wire _00803_ ;
wire _00804_ ;
wire _00805_ ;
wire _00806_ ;
wire _00807_ ;
wire _00808_ ;
wire _00809_ ;
wire _00810_ ;
wire _00811_ ;
wire _00812_ ;
wire _00813_ ;
wire _00814_ ;
wire _00815_ ;
wire _00816_ ;
wire _00817_ ;
wire _00818_ ;
wire _00819_ ;
wire _00820_ ;
wire _00821_ ;
wire _00822_ ;
wire _00823_ ;
wire _00824_ ;
wire _00825_ ;
wire _00826_ ;
wire _00827_ ;
wire _00828_ ;
wire _00829_ ;
wire _00830_ ;
wire _00831_ ;
wire _00832_ ;
wire _00833_ ;
wire _00834_ ;
wire _00835_ ;
wire _00836_ ;
wire _00837_ ;
wire _00838_ ;
wire _00839_ ;
wire _00840_ ;
wire _00841_ ;
wire _00842_ ;
wire _00843_ ;
wire _00844_ ;
wire _00845_ ;
wire _00846_ ;
wire _00847_ ;
wire _00848_ ;
wire _00849_ ;
wire _00850_ ;
wire _00851_ ;
wire _00852_ ;
wire _00853_ ;
wire _00854_ ;
wire _00855_ ;
wire _00856_ ;
wire _00857_ ;
wire _00858_ ;
wire _00859_ ;
wire _00860_ ;
wire _00861_ ;
wire _00862_ ;
wire _00863_ ;
wire _00864_ ;
wire _00865_ ;
wire _00866_ ;
wire _00867_ ;
wire _00868_ ;
wire _00869_ ;
wire _00870_ ;
wire _00871_ ;
wire _00872_ ;
wire _00873_ ;
wire _00874_ ;
wire _00875_ ;
wire _00876_ ;
wire _00877_ ;
wire _00878_ ;
wire _00879_ ;
wire _00880_ ;
wire _00881_ ;
wire _00882_ ;
wire _00883_ ;
wire _00884_ ;
wire _00885_ ;
wire _00886_ ;
wire _00887_ ;
wire _00888_ ;
wire _00889_ ;
wire _00890_ ;
wire _00891_ ;
wire _00892_ ;
wire _00893_ ;
wire _00894_ ;
wire _00895_ ;
wire _00896_ ;
wire _00897_ ;
wire _00898_ ;
wire _00899_ ;
wire _00900_ ;
wire _00901_ ;
wire _00902_ ;
wire _00903_ ;
wire _00904_ ;
wire _00905_ ;
wire _00906_ ;
wire _00907_ ;
wire _00908_ ;
wire _00909_ ;
wire _00910_ ;
wire _00911_ ;
wire _00912_ ;
wire _00913_ ;
wire _00914_ ;
wire _00915_ ;
wire _00916_ ;
wire _00917_ ;
wire _00918_ ;
wire _00919_ ;
wire _00920_ ;
wire _00921_ ;
wire _00922_ ;
wire _00923_ ;
wire _00924_ ;
wire _00925_ ;
wire _00926_ ;
wire _00927_ ;
wire _00928_ ;
wire _00929_ ;
wire _00930_ ;
wire _00931_ ;
wire _00932_ ;
wire _00933_ ;
wire _00934_ ;
wire _00935_ ;
wire _00936_ ;
wire _00937_ ;
wire _00938_ ;
wire _00939_ ;
wire _00940_ ;
wire _00941_ ;
wire _00942_ ;
wire _00943_ ;
wire _00944_ ;
wire _00945_ ;
wire _00946_ ;
wire _00947_ ;
wire _00948_ ;
wire _00949_ ;
wire _00950_ ;
wire _00951_ ;
wire _00952_ ;
wire _00953_ ;
wire _00954_ ;
wire _00955_ ;
wire _00956_ ;
wire _00957_ ;
wire _00958_ ;
wire _00959_ ;
wire _00960_ ;
wire _00961_ ;
wire _00962_ ;
wire _00963_ ;
wire _00964_ ;
wire _00965_ ;
wire _00966_ ;
wire _00967_ ;
wire _00968_ ;
wire _00969_ ;
wire _00970_ ;
wire _00971_ ;
wire _00972_ ;
wire _00973_ ;
wire _00974_ ;
wire _00975_ ;
wire _00976_ ;
wire _00977_ ;
wire _00978_ ;
wire _00979_ ;
wire _00980_ ;
wire _00981_ ;
wire _00982_ ;
wire _00983_ ;
wire _00984_ ;
wire _00985_ ;
wire _00986_ ;
wire _00987_ ;
wire _00988_ ;
wire _00989_ ;
wire _00990_ ;
wire _00991_ ;
wire _00992_ ;
wire _00993_ ;
wire _00994_ ;
wire _00995_ ;
wire _00996_ ;
wire _00997_ ;
wire _00998_ ;
wire _00999_ ;
wire _01000_ ;
wire _01001_ ;
wire _01002_ ;
wire _01003_ ;
wire _01004_ ;
wire _01005_ ;
wire _01006_ ;
wire _01007_ ;
wire _01008_ ;
wire _01009_ ;
wire _01010_ ;
wire _01011_ ;
wire _01012_ ;
wire _01013_ ;
wire _01014_ ;
wire _01015_ ;
wire _01016_ ;
wire _01017_ ;
wire _01018_ ;
wire _01019_ ;
wire _01020_ ;
wire _01021_ ;
wire _01022_ ;
wire _01023_ ;
wire _01024_ ;
wire _01025_ ;
wire _01026_ ;
wire _01027_ ;
wire _01028_ ;
wire _01029_ ;
wire _01030_ ;
wire _01031_ ;
wire _01032_ ;
wire _01033_ ;
wire _01034_ ;
wire _01035_ ;
wire _01036_ ;
wire _01037_ ;
wire _01038_ ;
wire _01039_ ;
wire _01040_ ;
wire _01041_ ;
wire _01042_ ;
wire _01043_ ;
wire _01044_ ;
wire _01045_ ;
wire _01046_ ;
wire _01047_ ;
wire _01048_ ;
wire _01049_ ;
wire _01050_ ;
wire _01051_ ;
wire _01052_ ;
wire _01053_ ;
wire _01054_ ;
wire _01055_ ;
wire _01056_ ;
wire _01057_ ;
wire _01058_ ;
wire _01059_ ;
wire _01060_ ;
wire _01061_ ;
wire _01062_ ;
wire _01063_ ;
wire _01064_ ;
wire _01065_ ;
wire _01066_ ;
wire _01067_ ;
wire _01068_ ;
wire _01069_ ;
wire _01070_ ;
wire _01071_ ;
wire _01072_ ;
wire _01073_ ;
wire _01074_ ;
wire _01075_ ;
wire _01076_ ;
wire _01077_ ;
wire _01078_ ;
wire _01079_ ;
wire _01080_ ;
wire _01081_ ;
wire _01082_ ;
wire _01083_ ;
wire _01084_ ;
wire _01085_ ;
wire _01086_ ;
wire _01087_ ;
wire _01088_ ;
wire _01089_ ;
wire _01090_ ;
wire _01091_ ;
wire _01092_ ;
wire _01093_ ;
wire _01094_ ;
wire _01095_ ;
wire _01096_ ;
wire _01097_ ;
wire _01098_ ;
wire _01099_ ;
wire _01100_ ;
wire _01101_ ;
wire _01102_ ;
wire _01103_ ;
wire _01104_ ;
wire _01105_ ;
wire _01106_ ;
wire _01107_ ;
wire _01108_ ;
wire _01109_ ;
wire _01110_ ;
wire _01111_ ;
wire _01112_ ;
wire _01113_ ;
wire _01114_ ;
wire _01115_ ;
wire _01116_ ;
wire _01117_ ;
wire _01118_ ;
wire _01119_ ;
wire _01120_ ;
wire _01121_ ;
wire _01122_ ;
wire _01123_ ;
wire _01124_ ;
wire _01125_ ;
wire _01126_ ;
wire _01127_ ;
wire _01128_ ;
wire _01129_ ;
wire _01130_ ;
wire _01131_ ;
wire _01132_ ;
wire _01133_ ;
wire _01134_ ;
wire _01135_ ;
wire _01136_ ;
wire _01137_ ;
wire _01138_ ;
wire _01139_ ;
wire _01140_ ;
wire _01141_ ;
wire _01142_ ;
wire _01143_ ;
wire _01144_ ;
wire _01145_ ;
wire _01146_ ;
wire _01147_ ;
wire _01148_ ;
wire _01149_ ;
wire _01150_ ;
wire _01151_ ;
wire _01152_ ;
wire _01153_ ;
wire _01154_ ;
wire _01155_ ;
wire _01156_ ;
wire _01157_ ;
wire _01158_ ;
wire _01159_ ;
wire _01160_ ;
wire _01161_ ;
wire _01162_ ;
wire _01163_ ;
wire _01164_ ;
wire _01165_ ;
wire _01166_ ;
wire _01167_ ;
wire _01168_ ;
wire _01169_ ;
wire _01170_ ;
wire _01171_ ;
wire _01172_ ;
wire _01173_ ;
wire _01174_ ;
wire _01175_ ;
wire _01176_ ;
wire _01177_ ;
wire _01178_ ;
wire _01179_ ;
wire _01180_ ;
wire _01181_ ;
wire _01182_ ;
wire _01183_ ;
wire _01184_ ;
wire _01185_ ;
wire _01186_ ;
wire _01187_ ;
wire _01188_ ;
wire _01189_ ;
wire _01190_ ;
wire _01191_ ;
wire _01192_ ;
wire _01193_ ;
wire _01194_ ;
wire _01195_ ;
wire _01196_ ;
wire _01197_ ;
wire _01198_ ;
wire _01199_ ;
wire _01200_ ;
wire _01201_ ;
wire _01202_ ;
wire _01203_ ;
wire _01204_ ;
wire _01205_ ;
wire _01206_ ;
wire _01207_ ;
wire _01208_ ;
wire _01209_ ;
wire _01210_ ;
wire _01211_ ;
wire _01212_ ;
wire _01213_ ;
wire _01214_ ;
wire _01215_ ;
wire _01216_ ;
wire _01217_ ;
wire _01218_ ;
wire _01219_ ;
wire _01220_ ;
wire _01221_ ;
wire _01222_ ;
wire _01223_ ;
wire _01224_ ;
wire _01225_ ;
wire _01226_ ;
wire _01227_ ;
wire _01228_ ;
wire _01229_ ;
wire _01230_ ;
wire _01231_ ;
wire _01232_ ;
wire _01233_ ;
wire _01234_ ;
wire _01235_ ;
wire _01236_ ;
wire _01237_ ;
wire _01238_ ;
wire _01239_ ;
wire _01240_ ;
wire _01241_ ;
wire _01242_ ;
wire _01243_ ;
wire _01244_ ;
wire _01245_ ;
wire _01246_ ;
wire _01247_ ;
wire _01248_ ;
wire _01249_ ;
wire _01250_ ;
wire _01251_ ;
wire _01252_ ;
wire _01253_ ;
wire _01254_ ;
wire _01255_ ;
wire _01256_ ;
wire _01257_ ;
wire _01258_ ;
wire _01259_ ;
wire _01260_ ;
wire _01261_ ;
wire _01262_ ;
wire _01263_ ;
wire _01264_ ;
wire _01265_ ;
wire _01266_ ;
wire _01267_ ;
wire _01268_ ;
wire _01269_ ;
wire _01270_ ;
wire _01271_ ;
wire _01272_ ;
wire _01273_ ;
wire _01274_ ;
wire _01275_ ;
wire _01276_ ;
wire _01277_ ;
wire _01278_ ;
wire _01279_ ;
wire _01280_ ;
wire _01281_ ;
wire _01282_ ;
wire _01283_ ;
wire _01284_ ;
wire _01285_ ;
wire _01286_ ;
wire _01287_ ;
wire _01288_ ;
wire _01289_ ;
wire _01290_ ;
wire _01291_ ;
wire _01292_ ;
wire _01293_ ;
wire _01294_ ;
wire _01295_ ;
wire _01296_ ;
wire _01297_ ;
wire _01298_ ;
wire _01299_ ;
wire _01300_ ;
wire _01301_ ;
wire _01302_ ;
wire _01303_ ;
wire _01304_ ;
wire _01305_ ;
wire _01306_ ;
wire _01307_ ;
wire _01308_ ;
wire _01309_ ;
wire _01310_ ;
wire _01311_ ;
wire _01312_ ;
wire _01313_ ;
wire _01314_ ;
wire _01315_ ;
wire _01316_ ;
wire _01317_ ;
wire _01318_ ;
wire _01319_ ;
wire _01320_ ;
wire _01321_ ;
wire _01322_ ;
wire _01323_ ;
wire _01324_ ;
wire _01325_ ;
wire _01326_ ;
wire _01327_ ;
wire _01328_ ;
wire _01329_ ;
wire _01330_ ;
wire _01331_ ;
wire _01332_ ;
wire _01333_ ;
wire _01334_ ;
wire _01335_ ;
wire _01336_ ;
wire _01337_ ;
wire _01338_ ;
wire _01339_ ;
wire _01340_ ;
wire _01341_ ;
wire _01342_ ;
wire _01343_ ;
wire _01344_ ;
wire _01345_ ;
wire _01346_ ;
wire _01347_ ;
wire _01348_ ;
wire _01349_ ;
wire _01350_ ;
wire _01351_ ;
wire _01352_ ;
wire _01353_ ;
wire _01354_ ;
wire _01355_ ;
wire _01356_ ;
wire _01357_ ;
wire _01358_ ;
wire _01359_ ;
wire _01360_ ;
wire _01361_ ;
wire _01362_ ;
wire _01363_ ;
wire _01364_ ;
wire _01365_ ;
wire _01366_ ;
wire _01367_ ;
wire _01368_ ;
wire _01369_ ;
wire _01370_ ;
wire _01371_ ;
wire _01372_ ;
wire _01373_ ;
wire _01374_ ;
wire _01375_ ;
wire _01376_ ;
wire _01377_ ;
wire _01378_ ;
wire _01379_ ;
wire _01380_ ;
wire _01381_ ;
wire _01382_ ;
wire _01383_ ;
wire _01384_ ;
wire _01385_ ;
wire _01386_ ;
wire _01387_ ;
wire _01388_ ;
wire _01389_ ;
wire _01390_ ;
wire _01391_ ;
wire _01392_ ;
wire _01393_ ;
wire _01394_ ;
wire _01395_ ;
wire _01396_ ;
wire _01397_ ;
wire _01398_ ;
wire _01399_ ;
wire _01400_ ;
wire _01401_ ;
wire _01402_ ;
wire _01403_ ;
wire _01404_ ;
wire _01405_ ;
wire _01406_ ;
wire _01407_ ;
wire _01408_ ;
wire _01409_ ;
wire _01410_ ;
wire _01411_ ;
wire _01412_ ;
wire _01413_ ;
wire _01414_ ;
wire _01415_ ;
wire _01416_ ;
wire _01417_ ;
wire _01418_ ;
wire _01419_ ;
wire _01420_ ;
wire _01421_ ;
wire _01422_ ;
wire _01423_ ;
wire _01424_ ;
wire _01425_ ;
wire _01426_ ;
wire _01427_ ;
wire _01428_ ;
wire _01429_ ;
wire _01430_ ;
wire _01431_ ;
wire _01432_ ;
wire _01433_ ;
wire _01434_ ;
wire _01435_ ;
wire _01436_ ;
wire _01437_ ;
wire _01438_ ;
wire _01439_ ;
wire _01440_ ;
wire _01441_ ;
wire _01442_ ;
wire _01443_ ;
wire _01444_ ;
wire _01445_ ;
wire _01446_ ;
wire _01447_ ;
wire _01448_ ;
wire _01449_ ;
wire _01450_ ;
wire _01451_ ;
wire _01452_ ;
wire _01453_ ;
wire _01454_ ;
wire _01455_ ;
wire _01456_ ;
wire _01457_ ;
wire _01458_ ;
wire _01459_ ;
wire _01460_ ;
wire _01461_ ;
wire _01462_ ;
wire _01463_ ;
wire _01464_ ;
wire _01465_ ;
wire _01466_ ;
wire _01467_ ;
wire _01468_ ;
wire _01469_ ;
wire _01470_ ;
wire _01471_ ;
wire _01472_ ;
wire _01473_ ;
wire _01474_ ;
wire _01475_ ;
wire _01476_ ;
wire _01477_ ;
wire _01478_ ;
wire _01479_ ;
wire _01480_ ;
wire _01481_ ;
wire _01482_ ;
wire _01483_ ;
wire _01484_ ;
wire _01485_ ;
wire _01486_ ;
wire _01487_ ;
wire _01488_ ;
wire _01489_ ;
wire _01490_ ;
wire _01491_ ;
wire _01492_ ;
wire _01493_ ;
wire _01494_ ;
wire _01495_ ;
wire _01496_ ;
wire _01497_ ;
wire _01498_ ;
wire _01499_ ;
wire _01500_ ;
wire _01501_ ;
wire _01502_ ;
wire _01503_ ;
wire _01504_ ;
wire _01505_ ;
wire _01506_ ;
wire _01507_ ;
wire _01508_ ;
wire _01509_ ;
wire _01510_ ;
wire _01511_ ;
wire _01512_ ;
wire _01513_ ;
wire _01514_ ;
wire _01515_ ;
wire _01516_ ;
wire _01517_ ;
wire _01518_ ;
wire _01519_ ;
wire _01520_ ;
wire _01521_ ;
wire _01522_ ;
wire _01523_ ;
wire _01524_ ;
wire _01525_ ;
wire _01526_ ;
wire _01527_ ;
wire _01528_ ;
wire _01529_ ;
wire _01530_ ;
wire _01531_ ;
wire _01532_ ;
wire _01533_ ;
wire _01534_ ;
wire _01535_ ;
wire _01536_ ;
wire _01537_ ;
wire _01538_ ;
wire _01539_ ;
wire _01540_ ;
wire _01541_ ;
wire _01542_ ;
wire _01543_ ;
wire _01544_ ;
wire _01545_ ;
wire _01546_ ;
wire _01547_ ;
wire _01548_ ;
wire _01549_ ;
wire _01550_ ;
wire _01551_ ;
wire _01552_ ;
wire _01553_ ;
wire _01554_ ;
wire _01555_ ;
wire _01556_ ;
wire _01557_ ;
wire _01558_ ;
wire _01559_ ;
wire _01560_ ;
wire _01561_ ;
wire _01562_ ;
wire _01563_ ;
wire _01564_ ;
wire _01565_ ;
wire _01566_ ;
wire _01567_ ;
wire _01568_ ;
wire _01569_ ;
wire _01570_ ;
wire _01571_ ;
wire _01572_ ;
wire _01573_ ;
wire _01574_ ;
wire _01575_ ;
wire _01576_ ;
wire _01577_ ;
wire _01578_ ;
wire _01579_ ;
wire _01580_ ;
wire _01581_ ;
wire _01582_ ;
wire _01583_ ;
wire _01584_ ;
wire _01585_ ;
wire _01586_ ;
wire _01587_ ;
wire _01588_ ;
wire _01589_ ;
wire _01590_ ;
wire _01591_ ;
wire _01592_ ;
wire _01593_ ;
wire _01594_ ;
wire _01595_ ;
wire _01596_ ;
wire _01597_ ;
wire _01598_ ;
wire _01599_ ;
wire _01600_ ;
wire _01601_ ;
wire _01602_ ;
wire _01603_ ;
wire _01604_ ;
wire _01605_ ;
wire _01606_ ;
wire _01607_ ;
wire _01608_ ;
wire _01609_ ;
wire _01610_ ;
wire _01611_ ;
wire _01612_ ;
wire _01613_ ;
wire _01614_ ;
wire _01615_ ;
wire _01616_ ;
wire _01617_ ;
wire _01618_ ;
wire _01619_ ;
wire _01620_ ;
wire _01621_ ;
wire _01622_ ;
wire _01623_ ;
wire _01624_ ;
wire _01625_ ;
wire _01626_ ;
wire _01627_ ;
wire _01628_ ;
wire _01629_ ;
wire _01630_ ;
wire _01631_ ;
wire _01632_ ;
wire _01633_ ;
wire _01634_ ;
wire _01635_ ;
wire _01636_ ;
wire _01637_ ;
wire _01638_ ;
wire _01639_ ;
wire _01640_ ;
wire _01641_ ;
wire _01642_ ;
wire _01643_ ;
wire _01644_ ;
wire _01645_ ;
wire _01646_ ;
wire _01647_ ;
wire _01648_ ;
wire _01649_ ;
wire _01650_ ;
wire _01651_ ;
wire _01652_ ;
wire _01653_ ;
wire _01654_ ;
wire _01655_ ;
wire _01656_ ;
wire _01657_ ;
wire _01658_ ;
wire _01659_ ;
wire _01660_ ;
wire _01661_ ;
wire _01662_ ;
wire _01663_ ;
wire _01664_ ;
wire _01665_ ;
wire _01666_ ;
wire _01667_ ;
wire _01668_ ;
wire _01669_ ;
wire _01670_ ;
wire _01671_ ;
wire _01672_ ;
wire _01673_ ;
wire _01674_ ;
wire _01675_ ;
wire _01676_ ;
wire _01677_ ;
wire _01678_ ;
wire _01679_ ;
wire _01680_ ;
wire _01681_ ;
wire _01682_ ;
wire _01683_ ;
wire _01684_ ;
wire _01685_ ;
wire _01686_ ;
wire _01687_ ;
wire _01688_ ;
wire _01689_ ;
wire _01690_ ;
wire _01691_ ;
wire _01692_ ;
wire _01693_ ;
wire _01694_ ;
wire _01695_ ;
wire _01696_ ;
wire _01697_ ;
wire _01698_ ;
wire _01699_ ;
wire _01700_ ;
wire _01701_ ;
wire _01702_ ;
wire _01703_ ;
wire _01704_ ;
wire _01705_ ;
wire _01706_ ;
wire _01707_ ;
wire _01708_ ;
wire _01709_ ;
wire _01710_ ;
wire _01711_ ;
wire _01712_ ;
wire _01713_ ;
wire _01714_ ;
wire _01715_ ;
wire _01716_ ;
wire _01717_ ;
wire _01718_ ;
wire _01719_ ;
wire _01720_ ;
wire _01721_ ;
wire _01722_ ;
wire _01723_ ;
wire _01724_ ;
wire _01725_ ;
wire _01726_ ;
wire _01727_ ;
wire _01728_ ;
wire _01729_ ;
wire _01730_ ;
wire _01731_ ;
wire _01732_ ;
wire _01733_ ;
wire _01734_ ;
wire _01735_ ;
wire _01736_ ;
wire _01737_ ;
wire _01738_ ;
wire _01739_ ;
wire _01740_ ;
wire _01741_ ;
wire _01742_ ;
wire _01743_ ;
wire _01744_ ;
wire _01745_ ;
wire _01746_ ;
wire _01747_ ;
wire _01748_ ;
wire _01749_ ;
wire _01750_ ;
wire _01751_ ;
wire _01752_ ;
wire _01753_ ;
wire _01754_ ;
wire _01755_ ;
wire _01756_ ;
wire _01757_ ;
wire _01758_ ;
wire _01759_ ;
wire _01760_ ;
wire _01761_ ;
wire _01762_ ;
wire _01763_ ;
wire _01764_ ;
wire _01765_ ;
wire _01766_ ;
wire _01767_ ;
wire _01768_ ;
wire _01769_ ;
wire _01770_ ;
wire _01771_ ;
wire _01772_ ;
wire _01773_ ;
wire _01774_ ;
wire _01775_ ;
wire _01776_ ;
wire _01777_ ;
wire _01778_ ;
wire _01779_ ;
wire _01780_ ;
wire _01781_ ;
wire _01782_ ;
wire _01783_ ;
wire _01784_ ;
wire _01785_ ;
wire _01786_ ;
wire _01787_ ;
wire _01788_ ;
wire _01789_ ;
wire _01790_ ;
wire _01791_ ;
wire _01792_ ;
wire _01793_ ;
wire _01794_ ;
wire _01795_ ;
wire _01796_ ;
wire _01797_ ;
wire _01798_ ;
wire _01799_ ;
wire _01800_ ;
wire _01801_ ;
wire _01802_ ;
wire _01803_ ;
wire _01804_ ;
wire _01805_ ;
wire _01806_ ;
wire _01807_ ;
wire _01808_ ;
wire _01809_ ;
wire _01810_ ;
wire _01811_ ;
wire _01812_ ;
wire _01813_ ;
wire _01814_ ;
wire _01815_ ;
wire _01816_ ;
wire _01817_ ;
wire _01818_ ;
wire _01819_ ;
wire _01820_ ;
wire _01821_ ;
wire _01822_ ;
wire _01823_ ;
wire _01824_ ;
wire _01825_ ;
wire _01826_ ;
wire _01827_ ;
wire _01828_ ;
wire _01829_ ;
wire _01830_ ;
wire _01831_ ;
wire _01832_ ;
wire _01833_ ;
wire _01834_ ;
wire _01835_ ;
wire _01836_ ;
wire _01837_ ;
wire _01838_ ;
wire _01839_ ;
wire _01840_ ;
wire _01841_ ;
wire _01842_ ;
wire _01843_ ;
wire _01844_ ;
wire _01845_ ;
wire _01846_ ;
wire _01847_ ;
wire _01848_ ;
wire _01849_ ;
wire _01850_ ;
wire _01851_ ;
wire _01852_ ;
wire _01853_ ;
wire _01854_ ;
wire _01855_ ;
wire _01856_ ;
wire _01857_ ;
wire _01858_ ;
wire _01859_ ;
wire _01860_ ;
wire _01861_ ;
wire _01862_ ;
wire _01863_ ;
wire _01864_ ;
wire _01865_ ;
wire _01866_ ;
wire _01867_ ;
wire _01868_ ;
wire _01869_ ;
wire _01870_ ;
wire _01871_ ;
wire _01872_ ;
wire _01873_ ;
wire _01874_ ;
wire _01875_ ;
wire _01876_ ;
wire _01877_ ;
wire _01878_ ;
wire _01879_ ;
wire _01880_ ;
wire _01881_ ;
wire _01882_ ;
wire _01883_ ;
wire _01884_ ;
wire _01885_ ;
wire _01886_ ;
wire _01887_ ;
wire _01888_ ;
wire _01889_ ;
wire _01890_ ;
wire _01891_ ;
wire _01892_ ;
wire _01893_ ;
wire _01894_ ;
wire _01895_ ;
wire _01896_ ;
wire _01897_ ;
wire _01898_ ;
wire _01899_ ;
wire _01900_ ;
wire _01901_ ;
wire _01902_ ;
wire _01903_ ;
wire _01904_ ;
wire _01905_ ;
wire _01906_ ;
wire _01907_ ;
wire _01908_ ;
wire _01909_ ;
wire _01910_ ;
wire _01911_ ;
wire _01912_ ;
wire _01913_ ;
wire _01914_ ;
wire _01915_ ;
wire _01916_ ;
wire _01917_ ;
wire _01918_ ;
wire _01919_ ;
wire _01920_ ;
wire _01921_ ;
wire _01922_ ;
wire _01923_ ;
wire _01924_ ;
wire _01925_ ;
wire _01926_ ;
wire _01927_ ;
wire _01928_ ;
wire _01929_ ;
wire _01930_ ;
wire _01931_ ;
wire _01932_ ;
wire _01933_ ;
wire _01934_ ;
wire _01935_ ;
wire _01936_ ;
wire _01937_ ;
wire _01938_ ;
wire _01939_ ;
wire _01940_ ;
wire _01941_ ;
wire _01942_ ;
wire _01943_ ;
wire _01944_ ;
wire _01945_ ;
wire _01946_ ;
wire _01947_ ;
wire _01948_ ;
wire _01949_ ;
wire _01950_ ;
wire _01951_ ;
wire _01952_ ;
wire _01953_ ;
wire _01954_ ;
wire _01955_ ;
wire _01956_ ;
wire _01957_ ;
wire _01958_ ;
wire _01959_ ;
wire _01960_ ;
wire _01961_ ;
wire _01962_ ;
wire _01963_ ;
wire _01964_ ;
wire _01965_ ;
wire _01966_ ;
wire _01967_ ;
wire _01968_ ;
wire _01969_ ;
wire _01970_ ;
wire _01971_ ;
wire _01972_ ;
wire _01973_ ;
wire _01974_ ;
wire _01975_ ;
wire _01976_ ;
wire _01977_ ;
wire _01978_ ;
wire _01979_ ;
wire _01980_ ;
wire _01981_ ;
wire _01982_ ;
wire _01983_ ;
wire _01984_ ;
wire _01985_ ;
wire _01986_ ;
wire _01987_ ;
wire _01988_ ;
wire _01989_ ;
wire _01990_ ;
wire _01991_ ;
wire _01992_ ;
wire _01993_ ;
wire _01994_ ;
wire _01995_ ;
wire _01996_ ;
wire _01997_ ;
wire _01998_ ;
wire _01999_ ;
wire _02000_ ;
wire _02001_ ;
wire _02002_ ;
wire _02003_ ;
wire _02004_ ;
wire _02005_ ;
wire _02006_ ;
wire _02007_ ;
wire _02008_ ;
wire _02009_ ;
wire _02010_ ;
wire _02011_ ;
wire _02012_ ;
wire _02013_ ;
wire _02014_ ;
wire _02015_ ;
wire _02016_ ;
wire _02017_ ;
wire _02018_ ;
wire _02019_ ;
wire _02020_ ;
wire _02021_ ;
wire _02022_ ;
wire _02023_ ;
wire _02024_ ;
wire _02025_ ;
wire _02026_ ;
wire _02027_ ;
wire _02028_ ;
wire _02029_ ;
wire _02030_ ;
wire _02031_ ;
wire _02032_ ;
wire _02033_ ;
wire _02034_ ;
wire _02035_ ;
wire _02036_ ;
wire _02037_ ;
wire _02038_ ;
wire _02039_ ;
wire _02040_ ;
wire _02041_ ;
wire _02042_ ;
wire _02043_ ;
wire _02044_ ;
wire _02045_ ;
wire _02046_ ;
wire _02047_ ;
wire _02048_ ;
wire _02049_ ;
wire _02050_ ;
wire _02051_ ;
wire _02052_ ;
wire _02053_ ;
wire _02054_ ;
wire _02055_ ;
wire _02056_ ;
wire _02057_ ;
wire _02058_ ;
wire _02059_ ;
wire _02060_ ;
wire _02061_ ;
wire _02062_ ;
wire _02063_ ;
wire _02064_ ;
wire _02065_ ;
wire _02066_ ;
wire _02067_ ;
wire _02068_ ;
wire _02069_ ;
wire _02070_ ;
wire _02071_ ;
wire _02072_ ;
wire _02073_ ;
wire _02074_ ;
wire _02075_ ;
wire _02076_ ;
wire _02077_ ;
wire _02078_ ;
wire _02079_ ;
wire _02080_ ;
wire _02081_ ;
wire _02082_ ;
wire _02083_ ;
wire _02084_ ;
wire _02085_ ;
wire _02086_ ;
wire _02087_ ;
wire _02088_ ;
wire _02089_ ;
wire _02090_ ;
wire _02091_ ;
wire _02092_ ;
wire _02093_ ;
wire _02094_ ;
wire _02095_ ;
wire _02096_ ;
wire _02097_ ;
wire _02098_ ;
wire _02099_ ;
wire _02100_ ;
wire _02101_ ;
wire _02102_ ;
wire _02103_ ;
wire _02104_ ;
wire _02105_ ;
wire _02106_ ;
wire _02107_ ;
wire _02108_ ;
wire _02109_ ;
wire _02110_ ;
wire _02111_ ;
wire _02112_ ;
wire _02113_ ;
wire _02114_ ;
wire _02115_ ;
wire _02116_ ;
wire _02117_ ;
wire _02118_ ;
wire _02119_ ;
wire _02120_ ;
wire _02121_ ;
wire _02122_ ;
wire _02123_ ;
wire _02124_ ;
wire _02125_ ;
wire _02126_ ;
wire _02127_ ;
wire _02128_ ;
wire _02129_ ;
wire _02130_ ;
wire _02131_ ;
wire _02132_ ;
wire _02133_ ;
wire _02134_ ;
wire _02135_ ;
wire _02136_ ;
wire _02137_ ;
wire _02138_ ;
wire _02139_ ;
wire _02140_ ;
wire _02141_ ;
wire _02142_ ;
wire _02143_ ;
wire _02144_ ;
wire _02145_ ;
wire _02146_ ;
wire _02147_ ;
wire _02148_ ;
wire _02149_ ;
wire _02150_ ;
wire _02151_ ;
wire _02152_ ;
wire _02153_ ;
wire _02154_ ;
wire _02155_ ;
wire _02156_ ;
wire _02157_ ;
wire _02158_ ;
wire _02159_ ;
wire _02160_ ;
wire _02161_ ;
wire _02162_ ;
wire _02163_ ;
wire _02164_ ;
wire _02165_ ;
wire _02166_ ;
wire _02167_ ;
wire _02168_ ;
wire _02169_ ;
wire _02170_ ;
wire _02171_ ;
wire _02172_ ;
wire _02173_ ;
wire _02174_ ;
wire _02175_ ;
wire _02176_ ;
wire _02177_ ;
wire _02178_ ;
wire _02179_ ;
wire _02180_ ;
wire _02181_ ;
wire _02182_ ;
wire _02183_ ;
wire _02184_ ;
wire _02185_ ;
wire _02186_ ;
wire _02187_ ;
wire _02188_ ;
wire _02189_ ;
wire _02190_ ;
wire _02191_ ;
wire _02192_ ;
wire _02193_ ;
wire _02194_ ;
wire _02195_ ;
wire _02196_ ;
wire _02197_ ;
wire _02198_ ;
wire _02199_ ;
wire _02200_ ;
wire _02201_ ;
wire _02202_ ;
wire _02203_ ;
wire _02204_ ;
wire _02205_ ;
wire _02206_ ;
wire _02207_ ;
wire _02208_ ;
wire _02209_ ;
wire _02210_ ;
wire _02211_ ;
wire _02212_ ;
wire _02213_ ;
wire _02214_ ;
wire _02215_ ;
wire _02216_ ;
wire _02217_ ;
wire _02218_ ;
wire _02219_ ;
wire _02220_ ;
wire _02221_ ;
wire _02222_ ;
wire _02223_ ;
wire _02224_ ;
wire _02225_ ;
wire _02226_ ;
wire _02227_ ;
wire _02228_ ;
wire _02229_ ;
wire _02230_ ;
wire _02231_ ;
wire _02232_ ;
wire _02233_ ;
wire _02234_ ;
wire _02235_ ;
wire _02236_ ;
wire _02237_ ;
wire _02238_ ;
wire _02239_ ;
wire _02240_ ;
wire _02241_ ;
wire _02242_ ;
wire _02243_ ;
wire _02244_ ;
wire _02245_ ;
wire _02246_ ;
wire _02247_ ;
wire _02248_ ;
wire _02249_ ;
wire _02250_ ;
wire _02251_ ;
wire _02252_ ;
wire _02253_ ;
wire _02254_ ;
wire _02255_ ;
wire _02256_ ;
wire _02257_ ;
wire _02258_ ;
wire _02259_ ;
wire _02260_ ;
wire _02261_ ;
wire _02262_ ;
wire _02263_ ;
wire _02264_ ;
wire _02265_ ;
wire _02266_ ;
wire _02267_ ;
wire _02268_ ;
wire _02269_ ;
wire _02270_ ;
wire _02271_ ;
wire _02272_ ;
wire _02273_ ;
wire _02274_ ;
wire _02275_ ;
wire _02276_ ;
wire _02277_ ;
wire _02278_ ;
wire _02279_ ;
wire _02280_ ;
wire _02281_ ;
wire _02282_ ;
wire _02283_ ;
wire _02284_ ;
wire _02285_ ;
wire _02286_ ;
wire _02287_ ;
wire _02288_ ;
wire _02289_ ;
wire _02290_ ;
wire _02291_ ;
wire _02292_ ;
wire _02293_ ;
wire _02294_ ;
wire _02295_ ;
wire _02296_ ;
wire _02297_ ;
wire _02298_ ;
wire _02299_ ;
wire _02300_ ;
wire _02301_ ;
wire _02302_ ;
wire _02303_ ;
wire _02304_ ;
wire _02305_ ;
wire _02306_ ;
wire _02307_ ;
wire _02308_ ;
wire _02309_ ;
wire _02310_ ;
wire _02311_ ;
wire _02312_ ;
wire _02313_ ;
wire _02314_ ;
wire _02315_ ;
wire _02316_ ;
wire _02317_ ;
wire _02318_ ;
wire _02319_ ;
wire _02320_ ;
wire _02321_ ;
wire _02322_ ;
wire _02323_ ;
wire _02324_ ;
wire _02325_ ;
wire _02326_ ;
wire _02327_ ;
wire _02328_ ;
wire _02329_ ;
wire _02330_ ;
wire _02331_ ;
wire _02332_ ;
wire _02333_ ;
wire _02334_ ;
wire _02335_ ;
wire _02336_ ;
wire _02337_ ;
wire _02338_ ;
wire _02339_ ;
wire _02340_ ;
wire _02341_ ;
wire _02342_ ;
wire _02343_ ;
wire _02344_ ;
wire _02345_ ;
wire _02346_ ;
wire _02347_ ;
wire _02348_ ;
wire _02349_ ;
wire _02350_ ;
wire _02351_ ;
wire _02352_ ;
wire _02353_ ;
wire _02354_ ;
wire _02355_ ;
wire _02356_ ;
wire _02357_ ;
wire _02358_ ;
wire _02359_ ;
wire _02360_ ;
wire _02361_ ;
wire _02362_ ;
wire _02363_ ;
wire _02364_ ;
wire _02365_ ;
wire _02366_ ;
wire _02367_ ;
wire _02368_ ;
wire _02369_ ;
wire _02370_ ;
wire _02371_ ;
wire _02372_ ;
wire _02373_ ;
wire _02374_ ;
wire _02375_ ;
wire _02376_ ;
wire _02377_ ;
wire _02378_ ;
wire _02379_ ;
wire _02380_ ;
wire _02381_ ;
wire _02382_ ;
wire _02383_ ;
wire _02384_ ;
wire _02385_ ;
wire _02386_ ;
wire _02387_ ;
wire _02388_ ;
wire _02389_ ;
wire _02390_ ;
wire _02391_ ;
wire _02392_ ;
wire _02393_ ;
wire _02394_ ;
wire _02395_ ;
wire _02396_ ;
wire _02397_ ;
wire _02398_ ;
wire _02399_ ;
wire _02400_ ;
wire _02401_ ;
wire _02402_ ;
wire _02403_ ;
wire _02404_ ;
wire _02405_ ;
wire _02406_ ;
wire _02407_ ;
wire _02408_ ;
wire _02409_ ;
wire _02410_ ;
wire _02411_ ;
wire _02412_ ;
wire _02413_ ;
wire _02414_ ;
wire _02415_ ;
wire _02416_ ;
wire _02417_ ;
wire _02418_ ;
wire _02419_ ;
wire _02420_ ;
wire _02421_ ;
wire _02422_ ;
wire _02423_ ;
wire _02424_ ;
wire _02425_ ;
wire _02426_ ;
wire _02427_ ;
wire _02428_ ;
wire _02429_ ;
wire _02430_ ;
wire _02431_ ;
wire _02432_ ;
wire _02433_ ;
wire _02434_ ;
wire _02435_ ;
wire _02436_ ;
wire _02437_ ;
wire _02438_ ;
wire _02439_ ;
wire _02440_ ;
wire _02441_ ;
wire _02442_ ;
wire _02443_ ;
wire _02444_ ;
wire _02445_ ;
wire _02446_ ;
wire _02447_ ;
wire _02448_ ;
wire _02449_ ;
wire _02450_ ;
wire _02451_ ;
wire _02452_ ;
wire _02453_ ;
wire _02454_ ;
wire _02455_ ;
wire _02456_ ;
wire _02457_ ;
wire _02458_ ;
wire _02459_ ;
wire _02460_ ;
wire _02461_ ;
wire _02462_ ;
wire _02463_ ;
wire _02464_ ;
wire _02465_ ;
wire _02466_ ;
wire _02467_ ;
wire _02468_ ;
wire _02469_ ;
wire _02470_ ;
wire _02471_ ;
wire _02472_ ;
wire _02473_ ;
wire _02474_ ;
wire _02475_ ;
wire _02476_ ;
wire _02477_ ;
wire _02478_ ;
wire _02479_ ;
wire _02480_ ;
wire _02481_ ;
wire _02482_ ;
wire _02483_ ;
wire _02484_ ;
wire _02485_ ;
wire _02486_ ;
wire _02487_ ;
wire _02488_ ;
wire _02489_ ;
wire _02490_ ;
wire _02491_ ;
wire _02492_ ;
wire _02493_ ;
wire _02494_ ;
wire _02495_ ;
wire _02496_ ;
wire _02497_ ;
wire _02498_ ;
wire _02499_ ;
wire _02500_ ;
wire _02501_ ;
wire _02502_ ;
wire _02503_ ;
wire _02504_ ;
wire _02505_ ;
wire _02506_ ;
wire _02507_ ;
wire _02508_ ;
wire _02509_ ;
wire _02510_ ;
wire _02511_ ;
wire _02512_ ;
wire _02513_ ;
wire _02514_ ;
wire _02515_ ;
wire _02516_ ;
wire _02517_ ;
wire _02518_ ;
wire _02519_ ;
wire _02520_ ;
wire _02521_ ;
wire _02522_ ;
wire _02523_ ;
wire _02524_ ;
wire _02525_ ;
wire _02526_ ;
wire _02527_ ;
wire _02528_ ;
wire _02529_ ;
wire _02530_ ;
wire _02531_ ;
wire _02532_ ;
wire _02533_ ;
wire _02534_ ;
wire _02535_ ;
wire _02536_ ;
wire _02537_ ;
wire _02538_ ;
wire _02539_ ;
wire _02540_ ;
wire _02541_ ;
wire _02542_ ;
wire _02543_ ;
wire _02544_ ;
wire _02545_ ;
wire _02546_ ;
wire _02547_ ;
wire _02548_ ;
wire _02549_ ;
wire _02550_ ;
wire _02551_ ;
wire _02552_ ;
wire _02553_ ;
wire _02554_ ;
wire _02555_ ;
wire _02556_ ;
wire _02557_ ;
wire _02558_ ;
wire _02559_ ;
wire _02560_ ;
wire _02561_ ;
wire _02562_ ;
wire _02563_ ;
wire _02564_ ;
wire _02565_ ;
wire _02566_ ;
wire _02567_ ;
wire _02568_ ;
wire _02569_ ;
wire _02570_ ;
wire _02571_ ;
wire _02572_ ;
wire _02573_ ;
wire _02574_ ;
wire _02575_ ;
wire _02576_ ;
wire _02577_ ;
wire _02578_ ;
wire _02579_ ;
wire _02580_ ;
wire _02581_ ;
wire _02582_ ;
wire _02583_ ;
wire _02584_ ;
wire _02585_ ;
wire _02586_ ;
wire _02587_ ;
wire _02588_ ;
wire _02589_ ;
wire _02590_ ;
wire _02591_ ;
wire _02592_ ;
wire _02593_ ;
wire _02594_ ;
wire _02595_ ;
wire _02596_ ;
wire _02597_ ;
wire _02598_ ;
wire _02599_ ;
wire _02600_ ;
wire _02601_ ;
wire _02602_ ;
wire _02603_ ;
wire _02604_ ;
wire _02605_ ;
wire _02606_ ;
wire _02607_ ;
wire _02608_ ;
wire _02609_ ;
wire _02610_ ;
wire _02611_ ;
wire _02612_ ;
wire _02613_ ;
wire _02614_ ;
wire _02615_ ;
wire _02616_ ;
wire _02617_ ;
wire _02618_ ;
wire _02619_ ;
wire _02620_ ;
wire _02621_ ;
wire _02622_ ;
wire _02623_ ;
wire _02624_ ;
wire _02625_ ;
wire _02626_ ;
wire _02627_ ;
wire _02628_ ;
wire _02629_ ;
wire _02630_ ;
wire _02631_ ;
wire _02632_ ;
wire _02633_ ;
wire _02634_ ;
wire _02635_ ;
wire _02636_ ;
wire _02637_ ;
wire _02638_ ;
wire _02639_ ;
wire _02640_ ;
wire _02641_ ;
wire _02642_ ;
wire _02643_ ;
wire _02644_ ;
wire _02645_ ;
wire _02646_ ;
wire _02647_ ;
wire _02648_ ;
wire _02649_ ;
wire _02650_ ;
wire _02651_ ;
wire _02652_ ;
wire _02653_ ;
wire _02654_ ;
wire _02655_ ;
wire _02656_ ;
wire _02657_ ;
wire _02658_ ;
wire _02659_ ;
wire _02660_ ;
wire _02661_ ;
wire _02662_ ;
wire _02663_ ;
wire _02664_ ;
wire _02665_ ;
wire _02666_ ;
wire _02667_ ;
wire _02668_ ;
wire _02669_ ;
wire _02670_ ;
wire _02671_ ;
wire _02672_ ;
wire _02673_ ;
wire _02674_ ;
wire _02675_ ;
wire _02676_ ;
wire _02677_ ;
wire _02678_ ;
wire _02679_ ;
wire _02680_ ;
wire _02681_ ;
wire _02682_ ;
wire _02683_ ;
wire _02684_ ;
wire _02685_ ;
wire _02686_ ;
wire _02687_ ;
wire _02688_ ;
wire _02689_ ;
wire _02690_ ;
wire _02691_ ;
wire _02692_ ;
wire _02693_ ;
wire _02694_ ;
wire _02695_ ;
wire _02696_ ;
wire _02697_ ;
wire _02698_ ;
wire _02699_ ;
wire _02700_ ;
wire _02701_ ;
wire _02702_ ;
wire _02703_ ;
wire _02704_ ;
wire _02705_ ;
wire _02706_ ;
wire _02707_ ;
wire _02708_ ;
wire _02709_ ;
wire _02710_ ;
wire _02711_ ;
wire _02712_ ;
wire _02713_ ;
wire _02714_ ;
wire _02715_ ;
wire _02716_ ;
wire _02717_ ;
wire _02718_ ;
wire _02719_ ;
wire _02720_ ;
wire _02721_ ;
wire _02722_ ;
wire _02723_ ;
wire _02724_ ;
wire _02725_ ;
wire _02726_ ;
wire _02727_ ;
wire _02728_ ;
wire _02729_ ;
wire _02730_ ;
wire _02731_ ;
wire _02732_ ;
wire _02733_ ;
wire _02734_ ;
wire _02735_ ;
wire _02736_ ;
wire _02737_ ;
wire _02738_ ;
wire _02739_ ;
wire _02740_ ;
wire _02741_ ;
wire _02742_ ;
wire _02743_ ;
wire _02744_ ;
wire _02745_ ;
wire _02746_ ;
wire _02747_ ;
wire _02748_ ;
wire _02749_ ;
wire _02750_ ;
wire _02751_ ;
wire _02752_ ;
wire _02753_ ;
wire _02754_ ;
wire _02755_ ;
wire _02756_ ;
wire _02757_ ;
wire _02758_ ;
wire _02759_ ;
wire _02760_ ;
wire _02761_ ;
wire _02762_ ;
wire _02763_ ;
wire _02764_ ;
wire _02765_ ;
wire _02766_ ;
wire _02767_ ;
wire _02768_ ;
wire _02769_ ;
wire _02770_ ;
wire _02771_ ;
wire _02772_ ;
wire _02773_ ;
wire _02774_ ;
wire _02775_ ;
wire _02776_ ;
wire _02777_ ;
wire _02778_ ;
wire _02779_ ;
wire _02780_ ;
wire _02781_ ;
wire _02782_ ;
wire _02783_ ;
wire _02784_ ;
wire _02785_ ;
wire _02786_ ;
wire _02787_ ;
wire _02788_ ;
wire _02789_ ;
wire _02790_ ;
wire _02791_ ;
wire _02792_ ;
wire _02793_ ;
wire _02794_ ;
wire _02795_ ;
wire _02796_ ;
wire _02797_ ;
wire _02798_ ;
wire _02799_ ;
wire _02800_ ;
wire _02801_ ;
wire _02802_ ;
wire _02803_ ;
wire _02804_ ;
wire _02805_ ;
wire _02806_ ;
wire _02807_ ;
wire _02808_ ;
wire _02809_ ;
wire _02810_ ;
wire _02811_ ;
wire _02812_ ;
wire _02813_ ;
wire _02814_ ;
wire _02815_ ;
wire _02816_ ;
wire _02817_ ;
wire _02818_ ;
wire _02819_ ;
wire _02820_ ;
wire _02821_ ;
wire _02822_ ;
wire _02823_ ;
wire _02824_ ;
wire _02825_ ;
wire _02826_ ;
wire _02827_ ;
wire _02828_ ;
wire _02829_ ;
wire _02830_ ;
wire _02831_ ;
wire _02832_ ;
wire _02833_ ;
wire _02834_ ;
wire _02835_ ;
wire _02836_ ;
wire _02837_ ;
wire _02838_ ;
wire _02839_ ;
wire _02840_ ;
wire _02841_ ;
wire _02842_ ;
wire _02843_ ;
wire _02844_ ;
wire _02845_ ;
wire _02846_ ;
wire _02847_ ;
wire _02848_ ;
wire _02849_ ;
wire _02850_ ;
wire _02851_ ;
wire _02852_ ;
wire _02853_ ;
wire _02854_ ;
wire _02855_ ;
wire _02856_ ;
wire _02857_ ;
wire _02858_ ;
wire _02859_ ;
wire _02860_ ;
wire _02861_ ;
wire _02862_ ;
wire _02863_ ;
wire _02864_ ;
wire _02865_ ;
wire _02866_ ;
wire _02867_ ;
wire _02868_ ;
wire _02869_ ;
wire _02870_ ;
wire _02871_ ;
wire _02872_ ;
wire _02873_ ;
wire _02874_ ;
wire _02875_ ;
wire _02876_ ;
wire _02877_ ;
wire _02878_ ;
wire _02879_ ;
wire _02880_ ;
wire _02881_ ;
wire _02882_ ;
wire _02883_ ;
wire _02884_ ;
wire _02885_ ;
wire _02886_ ;
wire _02887_ ;
wire _02888_ ;
wire _02889_ ;
wire _02890_ ;
wire _02891_ ;
wire _02892_ ;
wire _02893_ ;
wire _02894_ ;
wire _02895_ ;
wire _02896_ ;
wire _02897_ ;
wire _02898_ ;
wire _02899_ ;
wire _02900_ ;
wire _02901_ ;
wire _02902_ ;
wire _02903_ ;
wire _02904_ ;
wire _02905_ ;
wire _02906_ ;
wire _02907_ ;
wire _02908_ ;
wire _02909_ ;
wire _02910_ ;
wire _02911_ ;
wire _02912_ ;
wire _02913_ ;
wire _02914_ ;
wire _02915_ ;
wire _02916_ ;
wire _02917_ ;
wire _02918_ ;
wire _02919_ ;
wire _02920_ ;
wire _02921_ ;
wire _02922_ ;
wire _02923_ ;
wire _02924_ ;
wire _02925_ ;
wire _02926_ ;
wire _02927_ ;
wire _02928_ ;
wire _02929_ ;
wire _02930_ ;
wire _02931_ ;
wire _02932_ ;
wire _02933_ ;
wire _02934_ ;
wire _02935_ ;
wire _02936_ ;
wire _02937_ ;
wire _02938_ ;
wire _02939_ ;
wire _02940_ ;
wire _02941_ ;
wire _02942_ ;
wire _02943_ ;
wire _02944_ ;
wire _02945_ ;
wire _02946_ ;
wire _02947_ ;
wire _02948_ ;
wire _02949_ ;
wire _02950_ ;
wire _02951_ ;
wire _02952_ ;
wire _02953_ ;
wire _02954_ ;
wire _02955_ ;
wire _02956_ ;
wire _02957_ ;
wire _02958_ ;
wire _02959_ ;
wire _02960_ ;
wire _02961_ ;
wire _02962_ ;
wire _02963_ ;
wire _02964_ ;
wire _02965_ ;
wire _02966_ ;
wire _02967_ ;
wire _02968_ ;
wire _02969_ ;
wire _02970_ ;
wire _02971_ ;
wire _02972_ ;
wire _02973_ ;
wire _02974_ ;
wire _02975_ ;
wire _02976_ ;
wire _02977_ ;
wire _02978_ ;
wire _02979_ ;
wire _02980_ ;
wire _02981_ ;
wire _02982_ ;
wire _02983_ ;
wire _02984_ ;
wire _02985_ ;
wire _02986_ ;
wire _02987_ ;
wire _02988_ ;
wire _02989_ ;
wire _02990_ ;
wire _02991_ ;
wire _02992_ ;
wire _02993_ ;
wire _02994_ ;
wire _02995_ ;
wire _02996_ ;
wire _02997_ ;
wire _02998_ ;
wire _02999_ ;
wire _03000_ ;
wire _03001_ ;
wire _03002_ ;
wire _03003_ ;
wire _03004_ ;
wire _03005_ ;
wire _03006_ ;
wire _03007_ ;
wire _03008_ ;
wire _03009_ ;
wire _03010_ ;
wire _03011_ ;
wire _03012_ ;
wire _03013_ ;
wire _03014_ ;
wire _03015_ ;
wire _03016_ ;
wire _03017_ ;
wire _03018_ ;
wire _03019_ ;
wire _03020_ ;
wire _03021_ ;
wire _03022_ ;
wire _03023_ ;
wire _03024_ ;
wire _03025_ ;
wire _03026_ ;
wire _03027_ ;
wire _03028_ ;
wire _03029_ ;
wire _03030_ ;
wire _03031_ ;
wire _03032_ ;
wire _03033_ ;
wire _03034_ ;
wire _03035_ ;
wire _03036_ ;
wire _03037_ ;
wire _03038_ ;
wire _03039_ ;
wire _03040_ ;
wire _03041_ ;
wire _03042_ ;
wire _03043_ ;
wire _03044_ ;
wire _03045_ ;
wire _03046_ ;
wire _03047_ ;
wire _03048_ ;
wire _03049_ ;
wire _03050_ ;
wire _03051_ ;
wire _03052_ ;
wire _03053_ ;
wire _03054_ ;
wire _03055_ ;
wire _03056_ ;
wire _03057_ ;
wire _03058_ ;
wire _03059_ ;
wire _03060_ ;
wire _03061_ ;
wire _03062_ ;
wire _03063_ ;
wire _03064_ ;
wire _03065_ ;
wire _03066_ ;
wire _03067_ ;
wire _03068_ ;
wire _03069_ ;
wire _03070_ ;
wire _03071_ ;
wire _03072_ ;
wire _03073_ ;
wire _03074_ ;
wire _03075_ ;
wire _03076_ ;
wire _03077_ ;
wire _03078_ ;
wire _03079_ ;
wire _03080_ ;
wire _03081_ ;
wire _03082_ ;
wire _03083_ ;
wire _03084_ ;
wire _03085_ ;
wire _03086_ ;
wire _03087_ ;
wire _03088_ ;
wire _03089_ ;
wire _03090_ ;
wire _03091_ ;
wire _03092_ ;
wire _03093_ ;
wire _03094_ ;
wire _03095_ ;
wire _03096_ ;
wire _03097_ ;
wire _03098_ ;
wire _03099_ ;
wire _03100_ ;
wire _03101_ ;
wire _03102_ ;
wire _03103_ ;
wire _03104_ ;
wire _03105_ ;
wire _03106_ ;
wire _03107_ ;
wire _03108_ ;
wire _03109_ ;
wire _03110_ ;
wire _03111_ ;
wire _03112_ ;
wire _03113_ ;
wire _03114_ ;
wire _03115_ ;
wire _03116_ ;
wire _03117_ ;
wire _03118_ ;
wire _03119_ ;
wire _03120_ ;
wire _03121_ ;
wire _03122_ ;
wire _03123_ ;
wire _03124_ ;
wire _03125_ ;
wire _03126_ ;
wire _03127_ ;
wire _03128_ ;
wire _03129_ ;
wire _03130_ ;
wire _03131_ ;
wire _03132_ ;
wire _03133_ ;
wire _03134_ ;
wire _03135_ ;
wire _03136_ ;
wire _03137_ ;
wire _03138_ ;
wire _03139_ ;
wire _03140_ ;
wire _03141_ ;
wire _03142_ ;
wire _03143_ ;
wire _03144_ ;
wire _03145_ ;
wire _03146_ ;
wire _03147_ ;
wire _03148_ ;
wire _03149_ ;
wire _03150_ ;
wire _03151_ ;
wire _03152_ ;
wire _03153_ ;
wire _03154_ ;
wire _03155_ ;
wire _03156_ ;
wire _03157_ ;
wire _03158_ ;
wire _03159_ ;
wire _03160_ ;
wire _03161_ ;
wire _03162_ ;
wire _03163_ ;
wire _03164_ ;
wire _03165_ ;
wire _03166_ ;
wire _03167_ ;
wire _03168_ ;
wire _03169_ ;
wire _03170_ ;
wire _03171_ ;
wire _03172_ ;
wire _03173_ ;
wire _03174_ ;
wire _03175_ ;
wire _03176_ ;
wire _03177_ ;
wire _03178_ ;
wire _03179_ ;
wire _03180_ ;
wire _03181_ ;
wire _03182_ ;
wire _03183_ ;
wire _03184_ ;
wire _03185_ ;
wire _03186_ ;
wire _03187_ ;
wire _03188_ ;
wire _03189_ ;
wire _03190_ ;
wire _03191_ ;
wire _03192_ ;
wire _03193_ ;
wire _03194_ ;
wire _03195_ ;
wire _03196_ ;
wire _03197_ ;
wire _03198_ ;
wire _03199_ ;
wire _03200_ ;
wire _03201_ ;
wire _03202_ ;
wire _03203_ ;
wire _03204_ ;
wire _03205_ ;
wire _03206_ ;
wire _03207_ ;
wire _03208_ ;
wire _03209_ ;
wire _03210_ ;
wire _03211_ ;
wire _03212_ ;
wire _03213_ ;
wire _03214_ ;
wire _03215_ ;
wire _03216_ ;
wire _03217_ ;
wire _03218_ ;
wire _03219_ ;
wire _03220_ ;
wire _03221_ ;
wire _03222_ ;
wire _03223_ ;
wire _03224_ ;
wire _03225_ ;
wire _03226_ ;
wire _03227_ ;
wire _03228_ ;
wire _03229_ ;
wire _03230_ ;
wire _03231_ ;
wire _03232_ ;
wire _03233_ ;
wire _03234_ ;
wire _03235_ ;
wire _03236_ ;
wire _03237_ ;
wire _03238_ ;
wire _03239_ ;
wire _03240_ ;
wire _03241_ ;
wire _03242_ ;
wire _03243_ ;
wire _03244_ ;
wire _03245_ ;
wire _03246_ ;
wire _03247_ ;
wire _03248_ ;
wire _03249_ ;
wire _03250_ ;
wire _03251_ ;
wire _03252_ ;
wire _03253_ ;
wire _03254_ ;
wire _03255_ ;
wire _03256_ ;
wire _03257_ ;
wire _03258_ ;
wire _03259_ ;
wire _03260_ ;
wire _03261_ ;
wire _03262_ ;
wire _03263_ ;
wire _03264_ ;
wire _03265_ ;
wire _03266_ ;
wire _03267_ ;
wire _03268_ ;
wire _03269_ ;
wire _03270_ ;
wire _03271_ ;
wire _03272_ ;
wire _03273_ ;
wire _03274_ ;
wire _03275_ ;
wire _03276_ ;
wire _03277_ ;
wire _03278_ ;
wire _03279_ ;
wire _03280_ ;
wire _03281_ ;
wire _03282_ ;
wire _03283_ ;
wire _03284_ ;
wire _03285_ ;
wire _03286_ ;
wire _03287_ ;
wire _03288_ ;
wire _03289_ ;
wire _03290_ ;
wire _03291_ ;
wire _03292_ ;
wire _03293_ ;
wire _03294_ ;
wire _03295_ ;
wire _03296_ ;
wire _03297_ ;
wire _03298_ ;
wire _03299_ ;
wire _03300_ ;
wire _03301_ ;
wire _03302_ ;
wire _03303_ ;
wire _03304_ ;
wire _03305_ ;
wire _03306_ ;
wire _03307_ ;
wire _03308_ ;
wire _03309_ ;
wire _03310_ ;
wire _03311_ ;
wire _03312_ ;
wire _03313_ ;
wire _03314_ ;
wire _03315_ ;
wire _03316_ ;
wire _03317_ ;
wire _03318_ ;
wire _03319_ ;
wire _03320_ ;
wire _03321_ ;
wire _03322_ ;
wire _03323_ ;
wire _03324_ ;
wire _03325_ ;
wire _03326_ ;
wire _03327_ ;
wire _03328_ ;
wire _03329_ ;
wire _03330_ ;
wire _03331_ ;
wire _03332_ ;
wire _03333_ ;
wire _03334_ ;
wire _03335_ ;
wire _03336_ ;
wire _03337_ ;
wire _03338_ ;
wire _03339_ ;
wire _03340_ ;
wire _03341_ ;
wire _03342_ ;
wire _03343_ ;
wire _03344_ ;
wire _03345_ ;
wire _03346_ ;
wire _03347_ ;
wire _03348_ ;
wire _03349_ ;
wire _03350_ ;
wire _03351_ ;
wire _03352_ ;
wire _03353_ ;
wire _03354_ ;
wire _03355_ ;
wire _03356_ ;
wire _03357_ ;
wire _03358_ ;
wire _03359_ ;
wire _03360_ ;
wire _03361_ ;
wire _03362_ ;
wire _03363_ ;
wire _03364_ ;
wire _03365_ ;
wire _03366_ ;
wire _03367_ ;
wire _03368_ ;
wire _03369_ ;
wire _03370_ ;
wire _03371_ ;
wire _03372_ ;
wire _03373_ ;
wire _03374_ ;
wire _03375_ ;
wire _03376_ ;
wire _03377_ ;
wire _03378_ ;
wire _03379_ ;
wire _03380_ ;
wire _03381_ ;
wire _03382_ ;
wire _03383_ ;
wire _03384_ ;
wire _03385_ ;
wire _03386_ ;
wire _03387_ ;
wire _03388_ ;
wire _03389_ ;
wire _03390_ ;
wire _03391_ ;
wire _03392_ ;
wire _03393_ ;
wire _03394_ ;
wire _03395_ ;
wire _03396_ ;
wire _03397_ ;
wire _03398_ ;
wire _03399_ ;
wire _03400_ ;
wire _03401_ ;
wire _03402_ ;
wire _03403_ ;
wire _03404_ ;
wire _03405_ ;
wire _03406_ ;
wire _03407_ ;
wire _03408_ ;
wire _03409_ ;
wire _03410_ ;
wire _03411_ ;
wire _03412_ ;
wire _03413_ ;
wire _03414_ ;
wire _03415_ ;
wire _03416_ ;
wire _03417_ ;
wire _03418_ ;
wire _03419_ ;
wire _03420_ ;
wire _03421_ ;
wire _03422_ ;
wire _03423_ ;
wire _03424_ ;
wire _03425_ ;
wire _03426_ ;
wire _03427_ ;
wire _03428_ ;
wire _03429_ ;
wire _03430_ ;
wire _03431_ ;
wire _03432_ ;
wire _03433_ ;
wire _03434_ ;
wire _03435_ ;
wire _03436_ ;
wire _03437_ ;
wire _03438_ ;
wire _03439_ ;
wire _03440_ ;
wire _03441_ ;
wire _03442_ ;
wire _03443_ ;
wire _03444_ ;
wire _03445_ ;
wire _03446_ ;
wire _03447_ ;
wire _03448_ ;
wire _03449_ ;
wire _03450_ ;
wire _03451_ ;
wire _03452_ ;
wire _03453_ ;
wire _03454_ ;
wire _03455_ ;
wire _03456_ ;
wire _03457_ ;
wire _03458_ ;
wire _03459_ ;
wire _03460_ ;
wire _03461_ ;
wire _03462_ ;
wire _03463_ ;
wire _03464_ ;
wire _03465_ ;
wire _03466_ ;
wire _03467_ ;
wire _03468_ ;
wire _03469_ ;
wire _03470_ ;
wire _03471_ ;
wire _03472_ ;
wire _03473_ ;
wire _03474_ ;
wire _03475_ ;
wire _03476_ ;
wire _03477_ ;
wire _03478_ ;
wire _03479_ ;
wire _03480_ ;
wire _03481_ ;
wire _03482_ ;
wire _03483_ ;
wire _03484_ ;
wire _03485_ ;
wire _03486_ ;
wire _03487_ ;
wire _03488_ ;
wire _03489_ ;
wire _03490_ ;
wire _03491_ ;
wire _03492_ ;
wire _03493_ ;
wire _03494_ ;
wire _03495_ ;
wire _03496_ ;
wire _03497_ ;
wire _03498_ ;
wire _03499_ ;
wire _03500_ ;
wire _03501_ ;
wire _03502_ ;
wire _03503_ ;
wire _03504_ ;
wire _03505_ ;
wire _03506_ ;
wire _03507_ ;
wire _03508_ ;
wire _03509_ ;
wire _03510_ ;
wire _03511_ ;
wire _03512_ ;
wire _03513_ ;
wire _03514_ ;
wire _03515_ ;
wire _03516_ ;
wire _03517_ ;
wire _03518_ ;
wire _03519_ ;
wire _03520_ ;
wire _03521_ ;
wire _03522_ ;
wire _03523_ ;
wire _03524_ ;
wire _03525_ ;
wire _03526_ ;
wire _03527_ ;
wire _03528_ ;
wire _03529_ ;
wire _03530_ ;
wire _03531_ ;
wire _03532_ ;
wire _03533_ ;
wire _03534_ ;
wire _03535_ ;
wire _03536_ ;
wire _03537_ ;
wire _03538_ ;
wire _03539_ ;
wire _03540_ ;
wire _03541_ ;
wire _03542_ ;
wire _03543_ ;
wire _03544_ ;
wire _03545_ ;
wire _03546_ ;
wire _03547_ ;
wire _03548_ ;
wire _03549_ ;
wire _03550_ ;
wire _03551_ ;
wire _03552_ ;
wire _03553_ ;
wire _03554_ ;
wire _03555_ ;
wire _03556_ ;
wire _03557_ ;
wire _03558_ ;
wire _03559_ ;
wire _03560_ ;
wire _03561_ ;
wire _03562_ ;
wire _03563_ ;
wire _03564_ ;
wire _03565_ ;
wire _03566_ ;
wire _03567_ ;
wire _03568_ ;
wire _03569_ ;
wire _03570_ ;
wire _03571_ ;
wire _03572_ ;
wire _03573_ ;
wire _03574_ ;
wire _03575_ ;
wire _03576_ ;
wire _03577_ ;
wire _03578_ ;
wire _03579_ ;
wire _03580_ ;
wire _03581_ ;
wire _03582_ ;
wire _03583_ ;
wire _03584_ ;
wire _03585_ ;
wire _03586_ ;
wire _03587_ ;
wire _03588_ ;
wire _03589_ ;
wire _03590_ ;
wire _03591_ ;
wire _03592_ ;
wire _03593_ ;
wire _03594_ ;
wire _03595_ ;
wire _03596_ ;
wire _03597_ ;
wire _03598_ ;
wire _03599_ ;
wire _03600_ ;
wire _03601_ ;
wire _03602_ ;
wire _03603_ ;
wire _03604_ ;
wire _03605_ ;
wire _03606_ ;
wire _03607_ ;
wire _03608_ ;
wire _03609_ ;
wire _03610_ ;
wire _03611_ ;
wire _03612_ ;
wire _03613_ ;
wire _03614_ ;
wire _03615_ ;
wire _03616_ ;
wire _03617_ ;
wire _03618_ ;
wire _03619_ ;
wire _03620_ ;
wire _03621_ ;
wire _03622_ ;
wire _03623_ ;
wire _03624_ ;
wire _03625_ ;
wire _03626_ ;
wire _03627_ ;
wire _03628_ ;
wire _03629_ ;
wire _03630_ ;
wire _03631_ ;
wire _03632_ ;
wire _03633_ ;
wire _03634_ ;
wire _03635_ ;
wire _03636_ ;
wire _03637_ ;
wire _03638_ ;
wire _03639_ ;
wire _03640_ ;
wire _03641_ ;
wire _03642_ ;
wire _03643_ ;
wire _03644_ ;
wire _03645_ ;
wire _03646_ ;
wire _03647_ ;
wire _03648_ ;
wire _03649_ ;
wire _03650_ ;
wire _03651_ ;
wire _03652_ ;
wire _03653_ ;
wire _03654_ ;
wire _03655_ ;
wire _03656_ ;
wire _03657_ ;
wire _03658_ ;
wire _03659_ ;
wire _03660_ ;
wire _03661_ ;
wire _03662_ ;
wire _03663_ ;
wire _03664_ ;
wire _03665_ ;
wire _03666_ ;
wire _03667_ ;
wire _03668_ ;
wire _03669_ ;
wire _03670_ ;
wire _03671_ ;
wire _03672_ ;
wire _03673_ ;
wire _03674_ ;
wire _03675_ ;
wire _03676_ ;
wire _03677_ ;
wire _03678_ ;
wire _03679_ ;
wire _03680_ ;
wire _03681_ ;
wire _03682_ ;
wire _03683_ ;
wire _03684_ ;
wire _03685_ ;
wire _03686_ ;
wire _03687_ ;
wire _03688_ ;
wire _03689_ ;
wire _03690_ ;
wire _03691_ ;
wire _03692_ ;
wire _03693_ ;
wire _03694_ ;
wire _03695_ ;
wire _03696_ ;
wire _03697_ ;
wire _03698_ ;
wire _03699_ ;
wire _03700_ ;
wire _03701_ ;
wire _03702_ ;
wire _03703_ ;
wire _03704_ ;
wire _03705_ ;
wire _03706_ ;
wire _03707_ ;
wire _03708_ ;
wire _03709_ ;
wire _03710_ ;
wire _03711_ ;
wire _03712_ ;
wire _03713_ ;
wire _03714_ ;
wire _03715_ ;
wire _03716_ ;
wire _03717_ ;
wire _03718_ ;
wire _03719_ ;
wire _03720_ ;
wire _03721_ ;
wire _03722_ ;
wire _03723_ ;
wire _03724_ ;
wire _03725_ ;
wire _03726_ ;
wire _03727_ ;
wire _03728_ ;
wire _03729_ ;
wire _03730_ ;
wire _03731_ ;
wire _03732_ ;
wire _03733_ ;
wire _03734_ ;
wire _03735_ ;
wire _03736_ ;
wire _03737_ ;
wire _03738_ ;
wire _03739_ ;
wire _03740_ ;
wire _03741_ ;
wire _03742_ ;
wire _03743_ ;
wire _03744_ ;
wire _03745_ ;
wire _03746_ ;
wire _03747_ ;
wire _03748_ ;
wire _03749_ ;
wire _03750_ ;
wire _03751_ ;
wire _03752_ ;
wire _03753_ ;
wire _03754_ ;
wire _03755_ ;
wire _03756_ ;
wire _03757_ ;
wire _03758_ ;
wire _03759_ ;
wire _03760_ ;
wire _03761_ ;
wire _03762_ ;
wire _03763_ ;
wire _03764_ ;
wire _03765_ ;
wire _03766_ ;
wire _03767_ ;
wire _03768_ ;
wire _03769_ ;
wire _03770_ ;
wire _03771_ ;
wire _03772_ ;
wire _03773_ ;
wire _03774_ ;
wire _03775_ ;
wire _03776_ ;
wire _03777_ ;
wire _03778_ ;
wire _03779_ ;
wire _03780_ ;
wire _03781_ ;
wire _03782_ ;
wire _03783_ ;
wire _03784_ ;
wire _03785_ ;
wire _03786_ ;
wire _03787_ ;
wire _03788_ ;
wire _03789_ ;
wire _03790_ ;
wire _03791_ ;
wire _03792_ ;
wire _03793_ ;
wire _03794_ ;
wire _03795_ ;
wire _03796_ ;
wire _03797_ ;
wire _03798_ ;
wire _03799_ ;
wire _03800_ ;
wire _03801_ ;
wire _03802_ ;
wire _03803_ ;
wire _03804_ ;
wire _03805_ ;
wire _03806_ ;
wire _03807_ ;
wire _03808_ ;
wire _03809_ ;
wire _03810_ ;
wire _03811_ ;
wire _03812_ ;
wire _03813_ ;
wire _03814_ ;
wire _03815_ ;
wire _03816_ ;
wire _03817_ ;
wire _03818_ ;
wire _03819_ ;
wire _03820_ ;
wire _03821_ ;
wire _03822_ ;
wire _03823_ ;
wire _03824_ ;
wire _03825_ ;
wire _03826_ ;
wire _03827_ ;
wire _03828_ ;
wire _03829_ ;
wire _03830_ ;
wire _03831_ ;
wire _03832_ ;
wire _03833_ ;
wire _03834_ ;
wire _03835_ ;
wire _03836_ ;
wire _03837_ ;
wire _03838_ ;
wire _03839_ ;
wire _03840_ ;
wire _03841_ ;
wire _03842_ ;
wire _03843_ ;
wire _03844_ ;
wire _03845_ ;
wire _03846_ ;
wire _03847_ ;
wire _03848_ ;
wire _03849_ ;
wire _03850_ ;
wire _03851_ ;
wire _03852_ ;
wire _03853_ ;
wire _03854_ ;
wire _03855_ ;
wire _03856_ ;
wire _03857_ ;
wire _03858_ ;
wire _03859_ ;
wire _03860_ ;
wire _03861_ ;
wire _03862_ ;
wire _03863_ ;
wire _03864_ ;
wire _03865_ ;
wire _03866_ ;
wire _03867_ ;
wire _03868_ ;
wire _03869_ ;
wire _03870_ ;
wire _03871_ ;
wire _03872_ ;
wire _03873_ ;
wire _03874_ ;
wire _03875_ ;
wire _03876_ ;
wire _03877_ ;
wire _03878_ ;
wire _03879_ ;
wire _03880_ ;
wire _03881_ ;
wire _03882_ ;
wire _03883_ ;
wire _03884_ ;
wire _03885_ ;
wire _03886_ ;
wire _03887_ ;
wire _03888_ ;
wire _03889_ ;
wire _03890_ ;
wire _03891_ ;
wire _03892_ ;
wire _03893_ ;
wire _03894_ ;
wire _03895_ ;
wire _03896_ ;
wire _03897_ ;
wire _03898_ ;
wire _03899_ ;
wire _03900_ ;
wire _03901_ ;
wire _03902_ ;
wire _03903_ ;
wire _03904_ ;
wire _03905_ ;
wire _03906_ ;
wire _03907_ ;
wire _03908_ ;
wire _03909_ ;
wire _03910_ ;
wire _03911_ ;
wire _03912_ ;
wire _03913_ ;
wire _03914_ ;
wire _03915_ ;
wire _03916_ ;
wire _03917_ ;
wire _03918_ ;
wire _03919_ ;
wire _03920_ ;
wire _03921_ ;
wire _03922_ ;
wire _03923_ ;
wire _03924_ ;
wire _03925_ ;
wire _03926_ ;
wire _03927_ ;
wire _03928_ ;
wire _03929_ ;
wire _03930_ ;
wire _03931_ ;
wire _03932_ ;
wire _03933_ ;
wire _03934_ ;
wire _03935_ ;
wire _03936_ ;
wire _03937_ ;
wire _03938_ ;
wire _03939_ ;
wire _03940_ ;
wire _03941_ ;
wire _03942_ ;
wire _03943_ ;
wire _03944_ ;
wire _03945_ ;
wire _03946_ ;
wire _03947_ ;
wire _03948_ ;
wire _03949_ ;
wire _03950_ ;
wire _03951_ ;
wire _03952_ ;
wire _03953_ ;
wire _03954_ ;
wire _03955_ ;
wire _03956_ ;
wire _03957_ ;
wire _03958_ ;
wire _03959_ ;
wire _03960_ ;
wire _03961_ ;
wire _03962_ ;
wire _03963_ ;
wire _03964_ ;
wire _03965_ ;
wire _03966_ ;
wire _03967_ ;
wire _03968_ ;
wire _03969_ ;
wire _03970_ ;
wire _03971_ ;
wire _03972_ ;
wire _03973_ ;
wire _03974_ ;
wire _03975_ ;
wire _03976_ ;
wire _03977_ ;
wire _03978_ ;
wire _03979_ ;
wire _03980_ ;
wire _03981_ ;
wire _03982_ ;
wire _03983_ ;
wire _03984_ ;
wire _03985_ ;
wire _03986_ ;
wire _03987_ ;
wire _03988_ ;
wire _03989_ ;
wire _03990_ ;
wire _03991_ ;
wire _03992_ ;
wire _03993_ ;
wire _03994_ ;
wire _03995_ ;
wire _03996_ ;
wire _03997_ ;
wire _03998_ ;
wire _03999_ ;
wire _04000_ ;
wire _04001_ ;
wire _04002_ ;
wire _04003_ ;
wire _04004_ ;
wire _04005_ ;
wire _04006_ ;
wire _04007_ ;
wire _04008_ ;
wire _04009_ ;
wire _04010_ ;
wire _04011_ ;
wire _04012_ ;
wire _04013_ ;
wire _04014_ ;
wire _04015_ ;
wire _04016_ ;
wire _04017_ ;
wire _04018_ ;
wire _04019_ ;
wire _04020_ ;
wire _04021_ ;
wire _04022_ ;
wire _04023_ ;
wire _04024_ ;
wire _04025_ ;
wire _04026_ ;
wire _04027_ ;
wire _04028_ ;
wire _04029_ ;
wire _04030_ ;
wire _04031_ ;
wire _04032_ ;
wire _04033_ ;
wire _04034_ ;
wire _04035_ ;
wire _04036_ ;
wire _04037_ ;
wire _04038_ ;
wire _04039_ ;
wire _04040_ ;
wire _04041_ ;
wire _04042_ ;
wire _04043_ ;
wire _04044_ ;
wire _04045_ ;
wire _04046_ ;
wire _04047_ ;
wire _04048_ ;
wire _04049_ ;
wire _04050_ ;
wire _04051_ ;
wire _04052_ ;
wire _04053_ ;
wire _04054_ ;
wire _04055_ ;
wire _04056_ ;
wire _04057_ ;
wire _04058_ ;
wire _04059_ ;
wire _04060_ ;
wire _04061_ ;
wire _04062_ ;
wire _04063_ ;
wire _04064_ ;
wire _04065_ ;
wire _04066_ ;
wire _04067_ ;
wire _04068_ ;
wire _04069_ ;
wire _04070_ ;
wire _04071_ ;
wire _04072_ ;
wire _04073_ ;
wire _04074_ ;
wire _04075_ ;
wire _04076_ ;
wire _04077_ ;
wire _04078_ ;
wire _04079_ ;
wire _04080_ ;
wire _04081_ ;
wire _04082_ ;
wire _04083_ ;
wire _04084_ ;
wire _04085_ ;
wire _04086_ ;
wire _04087_ ;
wire _04088_ ;
wire _04089_ ;
wire _04090_ ;
wire _04091_ ;
wire _04092_ ;
wire _04093_ ;
wire _04094_ ;
wire _04095_ ;
wire _04096_ ;
wire _04097_ ;
wire _04098_ ;
wire _04099_ ;
wire _04100_ ;
wire _04101_ ;
wire _04102_ ;
wire _04103_ ;
wire _04104_ ;
wire _04105_ ;
wire _04106_ ;
wire _04107_ ;
wire _04108_ ;
wire _04109_ ;
wire _04110_ ;
wire _04111_ ;
wire _04112_ ;
wire _04113_ ;
wire _04114_ ;
wire _04115_ ;
wire _04116_ ;
wire _04117_ ;
wire _04118_ ;
wire _04119_ ;
wire _04120_ ;
wire _04121_ ;
wire _04122_ ;
wire _04123_ ;
wire _04124_ ;
wire _04125_ ;
wire _04126_ ;
wire _04127_ ;
wire _04128_ ;
wire _04129_ ;
wire _04130_ ;
wire _04131_ ;
wire _04132_ ;
wire _04133_ ;
wire _04134_ ;
wire _04135_ ;
wire _04136_ ;
wire _04137_ ;
wire _04138_ ;
wire _04139_ ;
wire _04140_ ;
wire _04141_ ;
wire _04142_ ;
wire _04143_ ;
wire _04144_ ;
wire _04145_ ;
wire _04146_ ;
wire _04147_ ;
wire _04148_ ;
wire _04149_ ;
wire _04150_ ;
wire _04151_ ;
wire _04152_ ;
wire _04153_ ;
wire _04154_ ;
wire _04155_ ;
wire _04156_ ;
wire _04157_ ;
wire _04158_ ;
wire _04159_ ;
wire _04160_ ;
wire _04161_ ;
wire _04162_ ;
wire _04163_ ;
wire _04164_ ;
wire _04165_ ;
wire _04166_ ;
wire _04167_ ;
wire _04168_ ;
wire _04169_ ;
wire _04170_ ;
wire _04171_ ;
wire _04172_ ;
wire _04173_ ;
wire _04174_ ;
wire _04175_ ;
wire _04176_ ;
wire _04177_ ;
wire _04178_ ;
wire _04179_ ;
wire _04180_ ;
wire _04181_ ;
wire _04182_ ;
wire _04183_ ;
wire _04184_ ;
wire _04185_ ;
wire _04186_ ;
wire _04187_ ;
wire _04188_ ;
wire _04189_ ;
wire _04190_ ;
wire _04191_ ;
wire _04192_ ;
wire _04193_ ;
wire _04194_ ;
wire _04195_ ;
wire _04196_ ;
wire _04197_ ;
wire _04198_ ;
wire _04199_ ;
wire _04200_ ;
wire _04201_ ;
wire _04202_ ;
wire _04203_ ;
wire _04204_ ;
wire _04205_ ;
wire _04206_ ;
wire _04207_ ;
wire _04208_ ;
wire _04209_ ;
wire _04210_ ;
wire _04211_ ;
wire _04212_ ;
wire _04213_ ;
wire _04214_ ;
wire _04215_ ;
wire _04216_ ;
wire _04217_ ;
wire _04218_ ;
wire _04219_ ;
wire _04220_ ;
wire _04221_ ;
wire _04222_ ;
wire _04223_ ;
wire _04224_ ;
wire _04225_ ;
wire _04226_ ;
wire _04227_ ;
wire _04228_ ;
wire _04229_ ;
wire _04230_ ;
wire _04231_ ;
wire _04232_ ;
wire _04233_ ;
wire _04234_ ;
wire _04235_ ;
wire _04236_ ;
wire _04237_ ;
wire _04238_ ;
wire _04239_ ;
wire _04240_ ;
wire _04241_ ;
wire _04242_ ;
wire _04243_ ;
wire _04244_ ;
wire _04245_ ;
wire _04246_ ;
wire _04247_ ;
wire _04248_ ;
wire _04249_ ;
wire _04250_ ;
wire _04251_ ;
wire _04252_ ;
wire _04253_ ;
wire _04254_ ;
wire _04255_ ;
wire _04256_ ;
wire _04257_ ;
wire _04258_ ;
wire _04259_ ;
wire _04260_ ;
wire _04261_ ;
wire _04262_ ;
wire _04263_ ;
wire _04264_ ;
wire _04265_ ;
wire _04266_ ;
wire _04267_ ;
wire _04268_ ;
wire _04269_ ;
wire _04270_ ;
wire _04271_ ;
wire _04272_ ;
wire _04273_ ;
wire _04274_ ;
wire _04275_ ;
wire _04276_ ;
wire _04277_ ;
wire _04278_ ;
wire _04279_ ;
wire _04280_ ;
wire _04281_ ;
wire _04282_ ;
wire _04283_ ;
wire _04284_ ;
wire _04285_ ;
wire _04286_ ;
wire _04287_ ;
wire _04288_ ;
wire _04289_ ;
wire _04290_ ;
wire _04291_ ;
wire _04292_ ;
wire _04293_ ;
wire _04294_ ;
wire _04295_ ;
wire _04296_ ;
wire _04297_ ;
wire _04298_ ;
wire _04299_ ;
wire _04300_ ;
wire _04301_ ;
wire _04302_ ;
wire _04303_ ;
wire _04304_ ;
wire _04305_ ;
wire _04306_ ;
wire _04307_ ;
wire _04308_ ;
wire _04309_ ;
wire _04310_ ;
wire _04311_ ;
wire _04312_ ;
wire _04313_ ;
wire _04314_ ;
wire _04315_ ;
wire _04316_ ;
wire _04317_ ;
wire _04318_ ;
wire _04319_ ;
wire _04320_ ;
wire _04321_ ;
wire _04322_ ;
wire _04323_ ;
wire _04324_ ;
wire _04325_ ;
wire _04326_ ;
wire _04327_ ;
wire _04328_ ;
wire _04329_ ;
wire _04330_ ;
wire _04331_ ;
wire _04332_ ;
wire _04333_ ;
wire _04334_ ;
wire _04335_ ;
wire _04336_ ;
wire _04337_ ;
wire _04338_ ;
wire _04339_ ;
wire _04340_ ;
wire _04341_ ;
wire _04342_ ;
wire _04343_ ;
wire _04344_ ;
wire _04345_ ;
wire _04346_ ;
wire _04347_ ;
wire _04348_ ;
wire _04349_ ;
wire _04350_ ;
wire _04351_ ;
wire _04352_ ;
wire _04353_ ;
wire _04354_ ;
wire _04355_ ;
wire _04356_ ;
wire _04357_ ;
wire _04358_ ;
wire _04359_ ;
wire _04360_ ;
wire _04361_ ;
wire _04362_ ;
wire _04363_ ;
wire _04364_ ;
wire _04365_ ;
wire _04366_ ;
wire _04367_ ;
wire _04368_ ;
wire _04369_ ;
wire _04370_ ;
wire _04371_ ;
wire _04372_ ;
wire _04373_ ;
wire _04374_ ;
wire _04375_ ;
wire _04376_ ;
wire _04377_ ;
wire _04378_ ;
wire _04379_ ;
wire _04380_ ;
wire _04381_ ;
wire _04382_ ;
wire _04383_ ;
wire _04384_ ;
wire _04385_ ;
wire _04386_ ;
wire _04387_ ;
wire _04388_ ;
wire _04389_ ;
wire _04390_ ;
wire _04391_ ;
wire _04392_ ;
wire _04393_ ;
wire _04394_ ;
wire _04395_ ;
wire _04396_ ;
wire _04397_ ;
wire _04398_ ;
wire _04399_ ;
wire _04400_ ;
wire _04401_ ;
wire _04402_ ;
wire _04403_ ;
wire _04404_ ;
wire _04405_ ;
wire _04406_ ;
wire _04407_ ;
wire _04408_ ;
wire _04409_ ;
wire _04410_ ;
wire _04411_ ;
wire _04412_ ;
wire _04413_ ;
wire _04414_ ;
wire _04415_ ;
wire _04416_ ;
wire _04417_ ;
wire _04418_ ;
wire _04419_ ;
wire _04420_ ;
wire _04421_ ;
wire _04422_ ;
wire _04423_ ;
wire _04424_ ;
wire _04425_ ;
wire _04426_ ;
wire _04427_ ;
wire _04428_ ;
wire _04429_ ;
wire _04430_ ;
wire _04431_ ;
wire _04432_ ;
wire _04433_ ;
wire _04434_ ;
wire _04435_ ;
wire _04436_ ;
wire _04437_ ;
wire _04438_ ;
wire _04439_ ;
wire _04440_ ;
wire _04441_ ;
wire _04442_ ;
wire _04443_ ;
wire _04444_ ;
wire _04445_ ;
wire _04446_ ;
wire _04447_ ;
wire _04448_ ;
wire _04449_ ;
wire _04450_ ;
wire _04451_ ;
wire _04452_ ;
wire _04453_ ;
wire _04454_ ;
wire _04455_ ;
wire _04456_ ;
wire _04457_ ;
wire _04458_ ;
wire _04459_ ;
wire _04460_ ;
wire _04461_ ;
wire _04462_ ;
wire _04463_ ;
wire _04464_ ;
wire _04465_ ;
wire _04466_ ;
wire _04467_ ;
wire _04468_ ;
wire _04469_ ;
wire _04470_ ;
wire _04471_ ;
wire _04472_ ;
wire _04473_ ;
wire _04474_ ;
wire _04475_ ;
wire _04476_ ;
wire _04477_ ;
wire _04478_ ;
wire _04479_ ;
wire _04480_ ;
wire _04481_ ;
wire _04482_ ;
wire _04483_ ;
wire _04484_ ;
wire _04485_ ;
wire _04486_ ;
wire _04487_ ;
wire _04488_ ;
wire _04489_ ;
wire _04490_ ;
wire _04491_ ;
wire _04492_ ;
wire _04493_ ;
wire _04494_ ;
wire _04495_ ;
wire _04496_ ;
wire _04497_ ;
wire _04498_ ;
wire _04499_ ;
wire _04500_ ;
wire _04501_ ;
wire _04502_ ;
wire _04503_ ;
wire _04504_ ;
wire _04505_ ;
wire _04506_ ;
wire _04507_ ;
wire _04508_ ;
wire _04509_ ;
wire _04510_ ;
wire _04511_ ;
wire _04512_ ;
wire _04513_ ;
wire _04514_ ;
wire _04515_ ;
wire _04516_ ;
wire _04517_ ;
wire _04518_ ;
wire _04519_ ;
wire _04520_ ;
wire _04521_ ;
wire _04522_ ;
wire _04523_ ;
wire _04524_ ;
wire _04525_ ;
wire _04526_ ;
wire _04527_ ;
wire _04528_ ;
wire _04529_ ;
wire _04530_ ;
wire _04531_ ;
wire _04532_ ;
wire _04533_ ;
wire _04534_ ;
wire _04535_ ;
wire _04536_ ;
wire _04537_ ;
wire _04538_ ;
wire _04539_ ;
wire _04540_ ;
wire _04541_ ;
wire _04542_ ;
wire _04543_ ;
wire _04544_ ;
wire _04545_ ;
wire _04546_ ;
wire _04547_ ;
wire _04548_ ;
wire _04549_ ;
wire _04550_ ;
wire _04551_ ;
wire _04552_ ;
wire _04553_ ;
wire _04554_ ;
wire _04555_ ;
wire _04556_ ;
wire _04557_ ;
wire _04558_ ;
wire _04559_ ;
wire _04560_ ;
wire _04561_ ;
wire _04562_ ;
wire _04563_ ;
wire _04564_ ;
wire _04565_ ;
wire _04566_ ;
wire _04567_ ;
wire _04568_ ;
wire _04569_ ;
wire _04570_ ;
wire _04571_ ;
wire _04572_ ;
wire _04573_ ;
wire _04574_ ;
wire _04575_ ;
wire _04576_ ;
wire _04577_ ;
wire _04578_ ;
wire _04579_ ;
wire _04580_ ;
wire _04581_ ;
wire _04582_ ;
wire _04583_ ;
wire _04584_ ;
wire _04585_ ;
wire _04586_ ;
wire _04587_ ;
wire _04588_ ;
wire _04589_ ;
wire _04590_ ;
wire _04591_ ;
wire _04592_ ;
wire _04593_ ;
wire _04594_ ;
wire _04595_ ;
wire _04596_ ;
wire _04597_ ;
wire _04598_ ;
wire _04599_ ;
wire _04600_ ;
wire _04601_ ;
wire _04602_ ;
wire _04603_ ;
wire _04604_ ;
wire _04605_ ;
wire _04606_ ;
wire _04607_ ;
wire _04608_ ;
wire _04609_ ;
wire _04610_ ;
wire _04611_ ;
wire _04612_ ;
wire _04613_ ;
wire _04614_ ;
wire _04615_ ;
wire _04616_ ;
wire _04617_ ;
wire _04618_ ;
wire _04619_ ;
wire _04620_ ;
wire _04621_ ;
wire _04622_ ;
wire _04623_ ;
wire _04624_ ;
wire _04625_ ;
wire _04626_ ;
wire _04627_ ;
wire _04628_ ;
wire _04629_ ;
wire _04630_ ;
wire _04631_ ;
wire _04632_ ;
wire _04633_ ;
wire _04634_ ;
wire _04635_ ;
wire _04636_ ;
wire _04637_ ;
wire _04638_ ;
wire _04639_ ;
wire _04640_ ;
wire _04641_ ;
wire _04642_ ;
wire _04643_ ;
wire _04644_ ;
wire _04645_ ;
wire _04646_ ;
wire _04647_ ;
wire _04648_ ;
wire _04649_ ;
wire _04650_ ;
wire _04651_ ;
wire _04652_ ;
wire _04653_ ;
wire _04654_ ;
wire _04655_ ;
wire _04656_ ;
wire _04657_ ;
wire _04658_ ;
wire _04659_ ;
wire _04660_ ;
wire _04661_ ;
wire _04662_ ;
wire _04663_ ;
wire _04664_ ;
wire _04665_ ;
wire _04666_ ;
wire _04667_ ;
wire _04668_ ;
wire _04669_ ;
wire _04670_ ;
wire _04671_ ;
wire _04672_ ;
wire _04673_ ;
wire _04674_ ;
wire _04675_ ;
wire _04676_ ;
wire _04677_ ;
wire _04678_ ;
wire _04679_ ;
wire _04680_ ;
wire _04681_ ;
wire _04682_ ;
wire _04683_ ;
wire _04684_ ;
wire _04685_ ;
wire _04686_ ;
wire _04687_ ;
wire _04688_ ;
wire _04689_ ;
wire _04690_ ;
wire _04691_ ;
wire _04692_ ;
wire _04693_ ;
wire _04694_ ;
wire _04695_ ;
wire _04696_ ;
wire _04697_ ;
wire _04698_ ;
wire _04699_ ;
wire _04700_ ;
wire _04701_ ;
wire _04702_ ;
wire _04703_ ;
wire _04704_ ;
wire _04705_ ;
wire _04706_ ;
wire _04707_ ;
wire _04708_ ;
wire _04709_ ;
wire _04710_ ;
wire _04711_ ;
wire _04712_ ;
wire _04713_ ;
wire _04714_ ;
wire _04715_ ;
wire _04716_ ;
wire _04717_ ;
wire _04718_ ;
wire _04719_ ;
wire _04720_ ;
wire _04721_ ;
wire _04722_ ;
wire _04723_ ;
wire _04724_ ;
wire _04725_ ;
wire _04726_ ;
wire _04727_ ;
wire _04728_ ;
wire _04729_ ;
wire _04730_ ;
wire _04731_ ;
wire _04732_ ;
wire _04733_ ;
wire _04734_ ;
wire _04735_ ;
wire _04736_ ;
wire _04737_ ;
wire _04738_ ;
wire _04739_ ;
wire _04740_ ;
wire _04741_ ;
wire _04742_ ;
wire _04743_ ;
wire _04744_ ;
wire _04745_ ;
wire _04746_ ;
wire _04747_ ;
wire _04748_ ;
wire _04749_ ;
wire _04750_ ;
wire _04751_ ;
wire _04752_ ;
wire _04753_ ;
wire _04754_ ;
wire _04755_ ;
wire _04756_ ;
wire _04757_ ;
wire _04758_ ;
wire _04759_ ;
wire _04760_ ;
wire _04761_ ;
wire _04762_ ;
wire _04763_ ;
wire _04764_ ;
wire _04765_ ;
wire _04766_ ;
wire _04767_ ;
wire _04768_ ;
wire _04769_ ;
wire _04770_ ;
wire _04771_ ;
wire _04772_ ;
wire _04773_ ;
wire _04774_ ;
wire _04775_ ;
wire _04776_ ;
wire _04777_ ;
wire _04778_ ;
wire _04779_ ;
wire _04780_ ;
wire _04781_ ;
wire _04782_ ;
wire _04783_ ;
wire _04784_ ;
wire _04785_ ;
wire _04786_ ;
wire _04787_ ;
wire _04788_ ;
wire _04789_ ;
wire _04790_ ;
wire _04791_ ;
wire _04792_ ;
wire _04793_ ;
wire _04794_ ;
wire _04795_ ;
wire _04796_ ;
wire _04797_ ;
wire _04798_ ;
wire _04799_ ;
wire _04800_ ;
wire _04801_ ;
wire _04802_ ;
wire _04803_ ;
wire _04804_ ;
wire _04805_ ;
wire _04806_ ;
wire _04807_ ;
wire _04808_ ;
wire _04809_ ;
wire _04810_ ;
wire _04811_ ;
wire _04812_ ;
wire _04813_ ;
wire _04814_ ;
wire _04815_ ;
wire _04816_ ;
wire _04817_ ;
wire _04818_ ;
wire _04819_ ;
wire _04820_ ;
wire _04821_ ;
wire _04822_ ;
wire _04823_ ;
wire _04824_ ;
wire _04825_ ;
wire _04826_ ;
wire _04827_ ;
wire _04828_ ;
wire _04829_ ;
wire _04830_ ;
wire _04831_ ;
wire _04832_ ;
wire _04833_ ;
wire _04834_ ;
wire _04835_ ;
wire _04836_ ;
wire _04837_ ;
wire _04838_ ;
wire _04839_ ;
wire _04840_ ;
wire _04841_ ;
wire _04842_ ;
wire _04843_ ;
wire _04844_ ;
wire _04845_ ;
wire _04846_ ;
wire _04847_ ;
wire _04848_ ;
wire _04849_ ;
wire _04850_ ;
wire _04851_ ;
wire _04852_ ;
wire _04853_ ;
wire _04854_ ;
wire _04855_ ;
wire _04856_ ;
wire _04857_ ;
wire _04858_ ;
wire _04859_ ;
wire _04860_ ;
wire _04861_ ;
wire _04862_ ;
wire _04863_ ;
wire _04864_ ;
wire _04865_ ;
wire _04866_ ;
wire _04867_ ;
wire _04868_ ;
wire _04869_ ;
wire _04870_ ;
wire _04871_ ;
wire _04872_ ;
wire _04873_ ;
wire _04874_ ;
wire _04875_ ;
wire _04876_ ;
wire _04877_ ;
wire _04878_ ;
wire _04879_ ;
wire _04880_ ;
wire _04881_ ;
wire _04882_ ;
wire _04883_ ;
wire _04884_ ;
wire _04885_ ;
wire _04886_ ;
wire _04887_ ;
wire _04888_ ;
wire _04889_ ;
wire _04890_ ;
wire _04891_ ;
wire _04892_ ;
wire _04893_ ;
wire _04894_ ;
wire _04895_ ;
wire _04896_ ;
wire _04897_ ;
wire _04898_ ;
wire _04899_ ;
wire _04900_ ;
wire _04901_ ;
wire _04902_ ;
wire _04903_ ;
wire _04904_ ;
wire _04905_ ;
wire _04906_ ;
wire _04907_ ;
wire _04908_ ;
wire _04909_ ;
wire _04910_ ;
wire _04911_ ;
wire _04912_ ;
wire _04913_ ;
wire _04914_ ;
wire _04915_ ;
wire _04916_ ;
wire _04917_ ;
wire _04918_ ;
wire _04919_ ;
wire _04920_ ;
wire _04921_ ;
wire _04922_ ;
wire _04923_ ;
wire _04924_ ;
wire _04925_ ;
wire _04926_ ;
wire _04927_ ;
wire _04928_ ;
wire _04929_ ;
wire _04930_ ;
wire _04931_ ;
wire _04932_ ;
wire _04933_ ;
wire _04934_ ;
wire _04935_ ;
wire _04936_ ;
wire _04937_ ;
wire _04938_ ;
wire _04939_ ;
wire _04940_ ;
wire _04941_ ;
wire _04942_ ;
wire _04943_ ;
wire _04944_ ;
wire _04945_ ;
wire _04946_ ;
wire _04947_ ;
wire _04948_ ;
wire _04949_ ;
wire _04950_ ;
wire _04951_ ;
wire _04952_ ;
wire _04953_ ;
wire _04954_ ;
wire _04955_ ;
wire _04956_ ;
wire _04957_ ;
wire _04958_ ;
wire _04959_ ;
wire _04960_ ;
wire _04961_ ;
wire _04962_ ;
wire _04963_ ;
wire _04964_ ;
wire _04965_ ;
wire _04966_ ;
wire _04967_ ;
wire _04968_ ;
wire _04969_ ;
wire _04970_ ;
wire _04971_ ;
wire _04972_ ;
wire _04973_ ;
wire _04974_ ;
wire _04975_ ;
wire _04976_ ;
wire _04977_ ;
wire _04978_ ;
wire _04979_ ;
wire _04980_ ;
wire _04981_ ;
wire _04982_ ;
wire _04983_ ;
wire _04984_ ;
wire _04985_ ;
wire _04986_ ;
wire _04987_ ;
wire _04988_ ;
wire _04989_ ;
wire _04990_ ;
wire _04991_ ;
wire _04992_ ;
wire _04993_ ;
wire _04994_ ;
wire _04995_ ;
wire _04996_ ;
wire _04997_ ;
wire _04998_ ;
wire _04999_ ;
wire _05000_ ;
wire _05001_ ;
wire _05002_ ;
wire _05003_ ;
wire _05004_ ;
wire _05005_ ;
wire _05006_ ;
wire _05007_ ;
wire _05008_ ;
wire _05009_ ;
wire _05010_ ;
wire _05011_ ;
wire _05012_ ;
wire _05013_ ;
wire _05014_ ;
wire _05015_ ;
wire _05016_ ;
wire _05017_ ;
wire _05018_ ;
wire _05019_ ;
wire _05020_ ;
wire _05021_ ;
wire _05022_ ;
wire _05023_ ;
wire _05024_ ;
wire _05025_ ;
wire _05026_ ;
wire _05027_ ;
wire _05028_ ;
wire _05029_ ;
wire _05030_ ;
wire _05031_ ;
wire _05032_ ;
wire _05033_ ;
wire _05034_ ;
wire _05035_ ;
wire _05036_ ;
wire _05037_ ;
wire _05038_ ;
wire _05039_ ;
wire _05040_ ;
wire _05041_ ;
wire _05042_ ;
wire _05043_ ;
wire _05044_ ;
wire _05045_ ;
wire _05046_ ;
wire _05047_ ;
wire _05048_ ;
wire _05049_ ;
wire _05050_ ;
wire _05051_ ;
wire _05052_ ;
wire _05053_ ;
wire _05054_ ;
wire _05055_ ;
wire _05056_ ;
wire _05057_ ;
wire _05058_ ;
wire _05059_ ;
wire _05060_ ;
wire _05061_ ;
wire _05062_ ;
wire _05063_ ;
wire _05064_ ;
wire _05065_ ;
wire _05066_ ;
wire _05067_ ;
wire _05068_ ;
wire _05069_ ;
wire _05070_ ;
wire _05071_ ;
wire _05072_ ;
wire _05073_ ;
wire _05074_ ;
wire _05075_ ;
wire _05076_ ;
wire _05077_ ;
wire _05078_ ;
wire _05079_ ;
wire _05080_ ;
wire _05081_ ;
wire _05082_ ;
wire _05083_ ;
wire _05084_ ;
wire _05085_ ;
wire _05086_ ;
wire _05087_ ;
wire _05088_ ;
wire _05089_ ;
wire _05090_ ;
wire _05091_ ;
wire _05092_ ;
wire _05093_ ;
wire _05094_ ;
wire _05095_ ;
wire _05096_ ;
wire _05097_ ;
wire _05098_ ;
wire _05099_ ;
wire _05100_ ;
wire _05101_ ;
wire _05102_ ;
wire _05103_ ;
wire _05104_ ;
wire _05105_ ;
wire _05106_ ;
wire _05107_ ;
wire _05108_ ;
wire _05109_ ;
wire _05110_ ;
wire _05111_ ;
wire _05112_ ;
wire _05113_ ;
wire _05114_ ;
wire _05115_ ;
wire _05116_ ;
wire _05117_ ;
wire _05118_ ;
wire _05119_ ;
wire _05120_ ;
wire _05121_ ;
wire _05122_ ;
wire _05123_ ;
wire _05124_ ;
wire _05125_ ;
wire _05126_ ;
wire _05127_ ;
wire _05128_ ;
wire _05129_ ;
wire _05130_ ;
wire _05131_ ;
wire _05132_ ;
wire _05133_ ;
wire _05134_ ;
wire _05135_ ;
wire _05136_ ;
wire _05137_ ;
wire _05138_ ;
wire _05139_ ;
wire _05140_ ;
wire _05141_ ;
wire _05142_ ;
wire _05143_ ;
wire _05144_ ;
wire _05145_ ;
wire _05146_ ;
wire _05147_ ;
wire _05148_ ;
wire _05149_ ;
wire _05150_ ;
wire _05151_ ;
wire _05152_ ;
wire _05153_ ;
wire _05154_ ;
wire _05155_ ;
wire _05156_ ;
wire _05157_ ;
wire _05158_ ;
wire _05159_ ;
wire _05160_ ;
wire _05161_ ;
wire _05162_ ;
wire _05163_ ;
wire _05164_ ;
wire _05165_ ;
wire _05166_ ;
wire _05167_ ;
wire _05168_ ;
wire _05169_ ;
wire _05170_ ;
wire _05171_ ;
wire _05172_ ;
wire _05173_ ;
wire _05174_ ;
wire _05175_ ;
wire _05176_ ;
wire _05177_ ;
wire _05178_ ;
wire _05179_ ;
wire _05180_ ;
wire _05181_ ;
wire _05182_ ;
wire _05183_ ;
wire _05184_ ;
wire _05185_ ;
wire _05186_ ;
wire _05187_ ;
wire _05188_ ;
wire _05189_ ;
wire _05190_ ;
wire _05191_ ;
wire _05192_ ;
wire _05193_ ;
wire _05194_ ;
wire _05195_ ;
wire _05196_ ;
wire _05197_ ;
wire _05198_ ;
wire _05199_ ;
wire _05200_ ;
wire _05201_ ;
wire _05202_ ;
wire _05203_ ;
wire _05204_ ;
wire _05205_ ;
wire _05206_ ;
wire _05207_ ;
wire _05208_ ;
wire _05209_ ;
wire _05210_ ;
wire _05211_ ;
wire _05212_ ;
wire _05213_ ;
wire _05214_ ;
wire _05215_ ;
wire _05216_ ;
wire _05217_ ;
wire _05218_ ;
wire _05219_ ;
wire _05220_ ;
wire _05221_ ;
wire _05222_ ;
wire _05223_ ;
wire _05224_ ;
wire _05225_ ;
wire _05226_ ;
wire _05227_ ;
wire _05228_ ;
wire _05229_ ;
wire _05230_ ;
wire _05231_ ;
wire _05232_ ;
wire _05233_ ;
wire _05234_ ;
wire _05235_ ;
wire _05236_ ;
wire _05237_ ;
wire _05238_ ;
wire _05239_ ;
wire _05240_ ;
wire _05241_ ;
wire _05242_ ;
wire _05243_ ;
wire _05244_ ;
wire _05245_ ;
wire _05246_ ;
wire _05247_ ;
wire _05248_ ;
wire _05249_ ;
wire _05250_ ;
wire _05251_ ;
wire _05252_ ;
wire _05253_ ;
wire _05254_ ;
wire _05255_ ;
wire _05256_ ;
wire _05257_ ;
wire _05258_ ;
wire _05259_ ;
wire _05260_ ;
wire _05261_ ;
wire _05262_ ;
wire _05263_ ;
wire _05264_ ;
wire _05265_ ;
wire _05266_ ;
wire _05267_ ;
wire _05268_ ;
wire _05269_ ;
wire _05270_ ;
wire _05271_ ;
wire _05272_ ;
wire _05273_ ;
wire _05274_ ;
wire _05275_ ;
wire _05276_ ;
wire _05277_ ;
wire _05278_ ;
wire _05279_ ;
wire _05280_ ;
wire _05281_ ;
wire _05282_ ;
wire _05283_ ;
wire _05284_ ;
wire _05285_ ;
wire _05286_ ;
wire _05287_ ;
wire _05288_ ;
wire _05289_ ;
wire _05290_ ;
wire _05291_ ;
wire _05292_ ;
wire _05293_ ;
wire _05294_ ;
wire _05295_ ;
wire _05296_ ;
wire _05297_ ;
wire _05298_ ;
wire _05299_ ;
wire _05300_ ;
wire _05301_ ;
wire _05302_ ;
wire _05303_ ;
wire _05304_ ;
wire _05305_ ;
wire _05306_ ;
wire _05307_ ;
wire _05308_ ;
wire _05309_ ;
wire _05310_ ;
wire _05311_ ;
wire _05312_ ;
wire _05313_ ;
wire _05314_ ;
wire _05315_ ;
wire _05316_ ;
wire _05317_ ;
wire _05318_ ;
wire _05319_ ;
wire _05320_ ;
wire _05321_ ;
wire _05322_ ;
wire _05323_ ;
wire _05324_ ;
wire _05325_ ;
wire _05326_ ;
wire _05327_ ;
wire _05328_ ;
wire _05329_ ;
wire _05330_ ;
wire _05331_ ;
wire _05332_ ;
wire _05333_ ;
wire _05334_ ;
wire _05335_ ;
wire _05336_ ;
wire _05337_ ;
wire _05338_ ;
wire _05339_ ;
wire _05340_ ;
wire _05341_ ;
wire _05342_ ;
wire _05343_ ;
wire _05344_ ;
wire _05345_ ;
wire _05346_ ;
wire _05347_ ;
wire _05348_ ;
wire _05349_ ;
wire _05350_ ;
wire _05351_ ;
wire _05352_ ;
wire _05353_ ;
wire _05354_ ;
wire _05355_ ;
wire _05356_ ;
wire _05357_ ;
wire _05358_ ;
wire _05359_ ;
wire _05360_ ;
wire _05361_ ;
wire _05362_ ;
wire _05363_ ;
wire _05364_ ;
wire _05365_ ;
wire _05366_ ;
wire _05367_ ;
wire _05368_ ;
wire _05369_ ;
wire _05370_ ;
wire _05371_ ;
wire _05372_ ;
wire _05373_ ;
wire _05374_ ;
wire _05375_ ;
wire _05376_ ;
wire _05377_ ;
wire _05378_ ;
wire _05379_ ;
wire _05380_ ;
wire _05381_ ;
wire _05382_ ;
wire _05383_ ;
wire _05384_ ;
wire _05385_ ;
wire _05386_ ;
wire _05387_ ;
wire _05388_ ;
wire _05389_ ;
wire _05390_ ;
wire _05391_ ;
wire _05392_ ;
wire _05393_ ;
wire _05394_ ;
wire _05395_ ;
wire _05396_ ;
wire _05397_ ;
wire _05398_ ;
wire _05399_ ;
wire _05400_ ;
wire _05401_ ;
wire _05402_ ;
wire _05403_ ;
wire _05404_ ;
wire _05405_ ;
wire _05406_ ;
wire _05407_ ;
wire _05408_ ;
wire _05409_ ;
wire _05410_ ;
wire _05411_ ;
wire _05412_ ;
wire _05413_ ;
wire _05414_ ;
wire _05415_ ;
wire _05416_ ;
wire _05417_ ;
wire _05418_ ;
wire _05419_ ;
wire _05420_ ;
wire _05421_ ;
wire _05422_ ;
wire _05423_ ;
wire _05424_ ;
wire _05425_ ;
wire _05426_ ;
wire _05427_ ;
wire _05428_ ;
wire _05429_ ;
wire _05430_ ;
wire _05431_ ;
wire _05432_ ;
wire _05433_ ;
wire _05434_ ;
wire _05435_ ;
wire _05436_ ;
wire _05437_ ;
wire _05438_ ;
wire _05439_ ;
wire _05440_ ;
wire _05441_ ;
wire _05442_ ;
wire _05443_ ;
wire _05444_ ;
wire _05445_ ;
wire _05446_ ;
wire _05447_ ;
wire _05448_ ;
wire _05449_ ;
wire _05450_ ;
wire _05451_ ;
wire _05452_ ;
wire _05453_ ;
wire _05454_ ;
wire _05455_ ;
wire _05456_ ;
wire _05457_ ;
wire _05458_ ;
wire _05459_ ;
wire _05460_ ;
wire _05461_ ;
wire _05462_ ;
wire _05463_ ;
wire _05464_ ;
wire _05465_ ;
wire _05466_ ;
wire _05467_ ;
wire _05468_ ;
wire _05469_ ;
wire _05470_ ;
wire _05471_ ;
wire _05472_ ;
wire _05473_ ;
wire _05474_ ;
wire _05475_ ;
wire _05476_ ;
wire _05477_ ;
wire _05478_ ;
wire _05479_ ;
wire _05480_ ;
wire _05481_ ;
wire _05482_ ;
wire _05483_ ;
wire _05484_ ;
wire _05485_ ;
wire _05486_ ;
wire _05487_ ;
wire _05488_ ;
wire _05489_ ;
wire _05490_ ;
wire _05491_ ;
wire _05492_ ;
wire _05493_ ;
wire _05494_ ;
wire _05495_ ;
wire _05496_ ;
wire _05497_ ;
wire _05498_ ;
wire _05499_ ;
wire _05500_ ;
wire _05501_ ;
wire _05502_ ;
wire _05503_ ;
wire _05504_ ;
wire _05505_ ;
wire _05506_ ;
wire _05507_ ;
wire _05508_ ;
wire _05509_ ;
wire _05510_ ;
wire _05511_ ;
wire _05512_ ;
wire _05513_ ;
wire _05514_ ;
wire _05515_ ;
wire _05516_ ;
wire _05517_ ;
wire _05518_ ;
wire _05519_ ;
wire _05520_ ;
wire _05521_ ;
wire _05522_ ;
wire _05523_ ;
wire _05524_ ;
wire _05525_ ;
wire _05526_ ;
wire _05527_ ;
wire _05528_ ;
wire _05529_ ;
wire _05530_ ;
wire _05531_ ;
wire _05532_ ;
wire _05533_ ;
wire _05534_ ;
wire _05535_ ;
wire _05536_ ;
wire _05537_ ;
wire _05538_ ;
wire _05539_ ;
wire _05540_ ;
wire _05541_ ;
wire _05542_ ;
wire _05543_ ;
wire _05544_ ;
wire _05545_ ;
wire _05546_ ;
wire _05547_ ;
wire _05548_ ;
wire _05549_ ;
wire _05550_ ;
wire _05551_ ;
wire _05552_ ;
wire _05553_ ;
wire _05554_ ;
wire _05555_ ;
wire _05556_ ;
wire _05557_ ;
wire _05558_ ;
wire _05559_ ;
wire _05560_ ;
wire _05561_ ;
wire _05562_ ;
wire _05563_ ;
wire _05564_ ;
wire _05565_ ;
wire _05566_ ;
wire _05567_ ;
wire _05568_ ;
wire _05569_ ;
wire _05570_ ;
wire _05571_ ;
wire _05572_ ;
wire _05573_ ;
wire _05574_ ;
wire _05575_ ;
wire _05576_ ;
wire _05577_ ;
wire _05578_ ;
wire _05579_ ;
wire _05580_ ;
wire _05581_ ;
wire _05582_ ;
wire _05583_ ;
wire _05584_ ;
wire _05585_ ;
wire _05586_ ;
wire _05587_ ;
wire _05588_ ;
wire _05589_ ;
wire _05590_ ;
wire _05591_ ;
wire _05592_ ;
wire _05593_ ;
wire _05594_ ;
wire _05595_ ;
wire _05596_ ;
wire _05597_ ;
wire _05598_ ;
wire _05599_ ;
wire _05600_ ;
wire _05601_ ;
wire _05602_ ;
wire _05603_ ;
wire _05604_ ;
wire _05605_ ;
wire _05606_ ;
wire _05607_ ;
wire _05608_ ;
wire _05609_ ;
wire _05610_ ;
wire _05611_ ;
wire _05612_ ;
wire _05613_ ;
wire _05614_ ;
wire _05615_ ;
wire _05616_ ;
wire _05617_ ;
wire _05618_ ;
wire _05619_ ;
wire _05620_ ;
wire _05621_ ;
wire _05622_ ;
wire _05623_ ;
wire _05624_ ;
wire _05625_ ;
wire _05626_ ;
wire _05627_ ;
wire _05628_ ;
wire _05629_ ;
wire _05630_ ;
wire _05631_ ;
wire _05632_ ;
wire _05633_ ;
wire _05634_ ;
wire _05635_ ;
wire _05636_ ;
wire _05637_ ;
wire _05638_ ;
wire _05639_ ;
wire _05640_ ;
wire _05641_ ;
wire _05642_ ;
wire _05643_ ;
wire _05644_ ;
wire _05645_ ;
wire _05646_ ;
wire _05647_ ;
wire _05648_ ;
wire _05649_ ;
wire _05650_ ;
wire _05651_ ;
wire _05652_ ;
wire _05653_ ;
wire _05654_ ;
wire _05655_ ;
wire _05656_ ;
wire _05657_ ;
wire _05658_ ;
wire _05659_ ;
wire _05660_ ;
wire _05661_ ;
wire _05662_ ;
wire _05663_ ;
wire _05664_ ;
wire _05665_ ;
wire _05666_ ;
wire _05667_ ;
wire _05668_ ;
wire _05669_ ;
wire _05670_ ;
wire _05671_ ;
wire _05672_ ;
wire _05673_ ;
wire _05674_ ;
wire _05675_ ;
wire _05676_ ;
wire _05677_ ;
wire _05678_ ;
wire _05679_ ;
wire _05680_ ;
wire _05681_ ;
wire _05682_ ;
wire _05683_ ;
wire _05684_ ;
wire _05685_ ;
wire _05686_ ;
wire _05687_ ;
wire _05688_ ;
wire _05689_ ;
wire _05690_ ;
wire _05691_ ;
wire _05692_ ;
wire _05693_ ;
wire _05694_ ;
wire _05695_ ;
wire _05696_ ;
wire _05697_ ;
wire _05698_ ;
wire _05699_ ;
wire _05700_ ;
wire _05701_ ;
wire _05702_ ;
wire _05703_ ;
wire _05704_ ;
wire _05705_ ;
wire _05706_ ;
wire _05707_ ;
wire _05708_ ;
wire _05709_ ;
wire _05710_ ;
wire _05711_ ;
wire _05712_ ;
wire _05713_ ;
wire _05714_ ;
wire _05715_ ;
wire _05716_ ;
wire _05717_ ;
wire _05718_ ;
wire _05719_ ;
wire _05720_ ;
wire _05721_ ;
wire _05722_ ;
wire _05723_ ;
wire _05724_ ;
wire _05725_ ;
wire _05726_ ;
wire _05727_ ;
wire _05728_ ;
wire _05729_ ;
wire _05730_ ;
wire _05731_ ;
wire _05732_ ;
wire _05733_ ;
wire _05734_ ;
wire _05735_ ;
wire _05736_ ;
wire _05737_ ;
wire _05738_ ;
wire _05739_ ;
wire _05740_ ;
wire _05741_ ;
wire _05742_ ;
wire _05743_ ;
wire _05744_ ;
wire _05745_ ;
wire _05746_ ;
wire _05747_ ;
wire _05748_ ;
wire _05749_ ;
wire _05750_ ;
wire _05751_ ;
wire _05752_ ;
wire _05753_ ;
wire _05754_ ;
wire _05755_ ;
wire _05756_ ;
wire _05757_ ;
wire _05758_ ;
wire _05759_ ;
wire _05760_ ;
wire _05761_ ;
wire _05762_ ;
wire _05763_ ;
wire _05764_ ;
wire _05765_ ;
wire _05766_ ;
wire _05767_ ;
wire _05768_ ;
wire _05769_ ;
wire _05770_ ;
wire _05771_ ;
wire _05772_ ;
wire _05773_ ;
wire _05774_ ;
wire _05775_ ;
wire _05776_ ;
wire _05777_ ;
wire _05778_ ;
wire _05779_ ;
wire _05780_ ;
wire _05781_ ;
wire _05782_ ;
wire _05783_ ;
wire _05784_ ;
wire _05785_ ;
wire _05786_ ;
wire _05787_ ;
wire _05788_ ;
wire _05789_ ;
wire _05790_ ;
wire _05791_ ;
wire _05792_ ;
wire _05793_ ;
wire _05794_ ;
wire _05795_ ;
wire _05796_ ;
wire _05797_ ;
wire _05798_ ;
wire _05799_ ;
wire _05800_ ;
wire _05801_ ;
wire _05802_ ;
wire _05803_ ;
wire _05804_ ;
wire _05805_ ;
wire _05806_ ;
wire _05807_ ;
wire _05808_ ;
wire _05809_ ;
wire _05810_ ;
wire _05811_ ;
wire _05812_ ;
wire _05813_ ;
wire _05814_ ;
wire _05815_ ;
wire _05816_ ;
wire _05817_ ;
wire _05818_ ;
wire _05819_ ;
wire _05820_ ;
wire _05821_ ;
wire _05822_ ;
wire _05823_ ;
wire _05824_ ;
wire _05825_ ;
wire _05826_ ;
wire _05827_ ;
wire _05828_ ;
wire _05829_ ;
wire _05830_ ;
wire _05831_ ;
wire _05832_ ;
wire _05833_ ;
wire _05834_ ;
wire _05835_ ;
wire _05836_ ;
wire _05837_ ;
wire _05838_ ;
wire _05839_ ;
wire _05840_ ;
wire _05841_ ;
wire _05842_ ;
wire _05843_ ;
wire _05844_ ;
wire _05845_ ;
wire _05846_ ;
wire _05847_ ;
wire _05848_ ;
wire _05849_ ;
wire _05850_ ;
wire _05851_ ;
wire _05852_ ;
wire _05853_ ;
wire _05854_ ;
wire _05855_ ;
wire _05856_ ;
wire _05857_ ;
wire _05858_ ;
wire _05859_ ;
wire _05860_ ;
wire _05861_ ;
wire _05862_ ;
wire _05863_ ;
wire _05864_ ;
wire _05865_ ;
wire _05866_ ;
wire _05867_ ;
wire _05868_ ;
wire _05869_ ;
wire _05870_ ;
wire _05871_ ;
wire _05872_ ;
wire _05873_ ;
wire _05874_ ;
wire _05875_ ;
wire _05876_ ;
wire _05877_ ;
wire _05878_ ;
wire _05879_ ;
wire _05880_ ;
wire _05881_ ;
wire _05882_ ;
wire _05883_ ;
wire _05884_ ;
wire _05885_ ;
wire _05886_ ;
wire _05887_ ;
wire _05888_ ;
wire _05889_ ;
wire _05890_ ;
wire _05891_ ;
wire _05892_ ;
wire _05893_ ;
wire _05894_ ;
wire _05895_ ;
wire _05896_ ;
wire _05897_ ;
wire _05898_ ;
wire _05899_ ;
wire _05900_ ;
wire _05901_ ;
wire _05902_ ;
wire _05903_ ;
wire _05904_ ;
wire _05905_ ;
wire _05906_ ;
wire _05907_ ;
wire _05908_ ;
wire _05909_ ;
wire _05910_ ;
wire _05911_ ;
wire _05912_ ;
wire _05913_ ;
wire _05914_ ;
wire _05915_ ;
wire _05916_ ;
wire _05917_ ;
wire _05918_ ;
wire _05919_ ;
wire _05920_ ;
wire _05921_ ;
wire _05922_ ;
wire _05923_ ;
wire _05924_ ;
wire _05925_ ;
wire _05926_ ;
wire _05927_ ;
wire _05928_ ;
wire _05929_ ;
wire _05930_ ;
wire _05931_ ;
wire _05932_ ;
wire _05933_ ;
wire _05934_ ;
wire _05935_ ;
wire _05936_ ;
wire _05937_ ;
wire _05938_ ;
wire _05939_ ;
wire _05940_ ;
wire _05941_ ;
wire _05942_ ;
wire _05943_ ;
wire _05944_ ;
wire _05945_ ;
wire _05946_ ;
wire _05947_ ;
wire _05948_ ;
wire _05949_ ;
wire _05950_ ;
wire _05951_ ;
wire _05952_ ;
wire _05953_ ;
wire _05954_ ;
wire _05955_ ;
wire _05956_ ;
wire _05957_ ;
wire _05958_ ;
wire _05959_ ;
wire _05960_ ;
wire _05961_ ;
wire _05962_ ;
wire _05963_ ;
wire _05964_ ;
wire _05965_ ;
wire _05966_ ;
wire _05967_ ;
wire _05968_ ;
wire _05969_ ;
wire _05970_ ;
wire _05971_ ;
wire _05972_ ;
wire _05973_ ;
wire _05974_ ;
wire _05975_ ;
wire _05976_ ;
wire _05977_ ;
wire _05978_ ;
wire _05979_ ;
wire _05980_ ;
wire _05981_ ;
wire _05982_ ;
wire _05983_ ;
wire _05984_ ;
wire _05985_ ;
wire _05986_ ;
wire _05987_ ;
wire _05988_ ;
wire _05989_ ;
wire _05990_ ;
wire _05991_ ;
wire _05992_ ;
wire _05993_ ;
wire _05994_ ;
wire _05995_ ;
wire _05996_ ;
wire _05997_ ;
wire _05998_ ;
wire _05999_ ;
wire _06000_ ;
wire _06001_ ;
wire _06002_ ;
wire _06003_ ;
wire _06004_ ;
wire _06005_ ;
wire _06006_ ;
wire _06007_ ;
wire _06008_ ;
wire _06009_ ;
wire _06010_ ;
wire _06011_ ;
wire _06012_ ;
wire _06013_ ;
wire _06014_ ;
wire _06015_ ;
wire _06016_ ;
wire _06017_ ;
wire _06018_ ;
wire _06019_ ;
wire _06020_ ;
wire _06021_ ;
wire _06022_ ;
wire _06023_ ;
wire _06024_ ;
wire _06025_ ;
wire _06026_ ;
wire _06027_ ;
wire _06028_ ;
wire _06029_ ;
wire _06030_ ;
wire _06031_ ;
wire _06032_ ;
wire _06033_ ;
wire _06034_ ;
wire _06035_ ;
wire _06036_ ;
wire _06037_ ;
wire _06038_ ;
wire _06039_ ;
wire _06040_ ;
wire _06041_ ;
wire _06042_ ;
wire _06043_ ;
wire _06044_ ;
wire _06045_ ;
wire _06046_ ;
wire _06047_ ;
wire _06048_ ;
wire _06049_ ;
wire _06050_ ;
wire _06051_ ;
wire _06052_ ;
wire _06053_ ;
wire _06054_ ;
wire _06055_ ;
wire _06056_ ;
wire _06057_ ;
wire _06058_ ;
wire _06059_ ;
wire _06060_ ;
wire _06061_ ;
wire _06062_ ;
wire _06063_ ;
wire _06064_ ;
wire _06065_ ;
wire _06066_ ;
wire _06067_ ;
wire _06068_ ;
wire _06069_ ;
wire _06070_ ;
wire _06071_ ;
wire _06072_ ;
wire _06073_ ;
wire _06074_ ;
wire _06075_ ;
wire _06076_ ;
wire _06077_ ;
wire _06078_ ;
wire _06079_ ;
wire _06080_ ;
wire _06081_ ;
wire _06082_ ;
wire _06083_ ;
wire _06084_ ;
wire _06085_ ;
wire _06086_ ;
wire _06087_ ;
wire _06088_ ;
wire _06089_ ;
wire _06090_ ;
wire _06091_ ;
wire _06092_ ;
wire _06093_ ;
wire _06094_ ;
wire _06095_ ;
wire _06096_ ;
wire _06097_ ;
wire _06098_ ;
wire _06099_ ;
wire _06100_ ;
wire _06101_ ;
wire _06102_ ;
wire _06103_ ;
wire _06104_ ;
wire _06105_ ;
wire _06106_ ;
wire _06107_ ;
wire _06108_ ;
wire _06109_ ;
wire _06110_ ;
wire _06111_ ;
wire _06112_ ;
wire _06113_ ;
wire _06114_ ;
wire _06115_ ;
wire _06116_ ;
wire _06117_ ;
wire _06118_ ;
wire _06119_ ;
wire _06120_ ;
wire _06121_ ;
wire _06122_ ;
wire _06123_ ;
wire _06124_ ;
wire _06125_ ;
wire _06126_ ;
wire _06127_ ;
wire _06128_ ;
wire _06129_ ;
wire _06130_ ;
wire _06131_ ;
wire _06132_ ;
wire _06133_ ;
wire _06134_ ;
wire _06135_ ;
wire _06136_ ;
wire _06137_ ;
wire _06138_ ;
wire _06139_ ;
wire _06140_ ;
wire _06141_ ;
wire _06142_ ;
wire _06143_ ;
wire _06144_ ;
wire _06145_ ;
wire _06146_ ;
wire _06147_ ;
wire _06148_ ;
wire _06149_ ;
wire _06150_ ;
wire _06151_ ;
wire _06152_ ;
wire _06153_ ;
wire _06154_ ;
wire _06155_ ;
wire _06156_ ;
wire _06157_ ;
wire _06158_ ;
wire _06159_ ;
wire _06160_ ;
wire _06161_ ;
wire _06162_ ;
wire _06163_ ;
wire _06164_ ;
wire _06165_ ;
wire _06166_ ;
wire _06167_ ;
wire _06168_ ;
wire _06169_ ;
wire _06170_ ;
wire _06171_ ;
wire _06172_ ;
wire _06173_ ;
wire _06174_ ;
wire _06175_ ;
wire _06176_ ;
wire _06177_ ;
wire _06178_ ;
wire _06179_ ;
wire _06180_ ;
wire _06181_ ;
wire _06182_ ;
wire _06183_ ;
wire _06184_ ;
wire _06185_ ;
wire _06186_ ;
wire _06187_ ;
wire _06188_ ;
wire _06189_ ;
wire _06190_ ;
wire _06191_ ;
wire _06192_ ;
wire _06193_ ;
wire _06194_ ;
wire _06195_ ;
wire _06196_ ;
wire _06197_ ;
wire _06198_ ;
wire _06199_ ;
wire _06200_ ;
wire _06201_ ;
wire _06202_ ;
wire _06203_ ;
wire _06204_ ;
wire _06205_ ;
wire _06206_ ;
wire _06207_ ;
wire _06208_ ;
wire _06209_ ;
wire _06210_ ;
wire _06211_ ;
wire _06212_ ;
wire _06213_ ;
wire _06214_ ;
wire _06215_ ;
wire _06216_ ;
wire _06217_ ;
wire _06218_ ;
wire _06219_ ;
wire _06220_ ;
wire _06221_ ;
wire _06222_ ;
wire _06223_ ;
wire _06224_ ;
wire _06225_ ;
wire _06226_ ;
wire _06227_ ;
wire _06228_ ;
wire _06229_ ;
wire _06230_ ;
wire _06231_ ;
wire _06232_ ;
wire _06233_ ;
wire _06234_ ;
wire _06235_ ;
wire _06236_ ;
wire _06237_ ;
wire _06238_ ;
wire _06239_ ;
wire _06240_ ;
wire _06241_ ;
wire _06242_ ;
wire _06243_ ;
wire _06244_ ;
wire _06245_ ;
wire _06246_ ;
wire _06247_ ;
wire _06248_ ;
wire _06249_ ;
wire _06250_ ;
wire _06251_ ;
wire _06252_ ;
wire _06253_ ;
wire _06254_ ;
wire _06255_ ;
wire _06256_ ;
wire _06257_ ;
wire _06258_ ;
wire _06259_ ;
wire _06260_ ;
wire _06261_ ;
wire _06262_ ;
wire _06263_ ;
wire _06264_ ;
wire _06265_ ;
wire _06266_ ;
wire _06267_ ;
wire _06268_ ;
wire _06269_ ;
wire _06270_ ;
wire _06271_ ;
wire _06272_ ;
wire _06273_ ;
wire _06274_ ;
wire _06275_ ;
wire _06276_ ;
wire _06277_ ;
wire _06278_ ;
wire _06279_ ;
wire _06280_ ;
wire _06281_ ;
wire _06282_ ;
wire _06283_ ;
wire _06284_ ;
wire _06285_ ;
wire _06286_ ;
wire _06287_ ;
wire _06288_ ;
wire _06289_ ;
wire _06290_ ;
wire _06291_ ;
wire _06292_ ;
wire _06293_ ;
wire _06294_ ;
wire _06295_ ;
wire _06296_ ;
wire _06297_ ;
wire _06298_ ;
wire _06299_ ;
wire _06300_ ;
wire _06301_ ;
wire _06302_ ;
wire _06303_ ;
wire _06304_ ;
wire _06305_ ;
wire _06306_ ;
wire _06307_ ;
wire _06308_ ;
wire _06309_ ;
wire _06310_ ;
wire _06311_ ;
wire _06312_ ;
wire _06313_ ;
wire _06314_ ;
wire _06315_ ;
wire _06316_ ;
wire _06317_ ;
wire _06318_ ;
wire _06319_ ;
wire _06320_ ;
wire _06321_ ;
wire _06322_ ;
wire _06323_ ;
wire _06324_ ;
wire _06325_ ;
wire _06326_ ;
wire _06327_ ;
wire _06328_ ;
wire _06329_ ;
wire _06330_ ;
wire _06331_ ;
wire _06332_ ;
wire _06333_ ;
wire _06334_ ;
wire _06335_ ;
wire _06336_ ;
wire _06337_ ;
wire _06338_ ;
wire _06339_ ;
wire _06340_ ;
wire _06341_ ;
wire _06342_ ;
wire _06343_ ;
wire _06344_ ;
wire _06345_ ;
wire _06346_ ;
wire _06347_ ;
wire _06348_ ;
wire _06349_ ;
wire _06350_ ;
wire _06351_ ;
wire _06352_ ;
wire _06353_ ;
wire _06354_ ;
wire _06355_ ;
wire _06356_ ;
wire _06357_ ;
wire _06358_ ;
wire _06359_ ;
wire _06360_ ;
wire _06361_ ;
wire _06362_ ;
wire _06363_ ;
wire _06364_ ;
wire _06365_ ;
wire _06366_ ;
wire _06367_ ;
wire _06368_ ;
wire _06369_ ;
wire _06370_ ;
wire _06371_ ;
wire _06372_ ;
wire _06373_ ;
wire _06374_ ;
wire _06375_ ;
wire _06376_ ;
wire _06377_ ;
wire _06378_ ;
wire _06379_ ;
wire _06380_ ;
wire _06381_ ;
wire _06382_ ;
wire _06383_ ;
wire _06384_ ;
wire _06385_ ;
wire _06386_ ;
wire _06387_ ;
wire _06388_ ;
wire _06389_ ;
wire _06390_ ;
wire _06391_ ;
wire _06392_ ;
wire _06393_ ;
wire _06394_ ;
wire _06395_ ;
wire _06396_ ;
wire _06397_ ;
wire _06398_ ;
wire _06399_ ;
wire _06400_ ;
wire _06401_ ;
wire _06402_ ;
wire _06403_ ;
wire _06404_ ;
wire _06405_ ;
wire _06406_ ;
wire _06407_ ;
wire _06408_ ;
wire _06409_ ;
wire _06410_ ;
wire _06411_ ;
wire _06412_ ;
wire _06413_ ;
wire _06414_ ;
wire _06415_ ;
wire _06416_ ;
wire _06417_ ;
wire _06418_ ;
wire _06419_ ;
wire _06420_ ;
wire _06421_ ;
wire _06422_ ;
wire _06423_ ;
wire _06424_ ;
wire _06425_ ;
wire _06426_ ;
wire _06427_ ;
wire _06428_ ;
wire _06429_ ;
wire _06430_ ;
wire _06431_ ;
wire _06432_ ;
wire _06433_ ;
wire _06434_ ;
wire _06435_ ;
wire _06436_ ;
wire _06437_ ;
wire _06438_ ;
wire _06439_ ;
wire _06440_ ;
wire _06441_ ;
wire _06442_ ;
wire _06443_ ;
wire _06444_ ;
wire _06445_ ;
wire _06446_ ;
wire _06447_ ;
wire _06448_ ;
wire _06449_ ;
wire _06450_ ;
wire _06451_ ;
wire _06452_ ;
wire _06453_ ;
wire _06454_ ;
wire _06455_ ;
wire _06456_ ;
wire _06457_ ;
wire _06458_ ;
wire _06459_ ;
wire _06460_ ;
wire _06461_ ;
wire _06462_ ;
wire _06463_ ;
wire _06464_ ;
wire _06465_ ;
wire _06466_ ;
wire _06467_ ;
wire _06468_ ;
wire _06469_ ;
wire _06470_ ;
wire _06471_ ;
wire _06472_ ;
wire _06473_ ;
wire _06474_ ;
wire _06475_ ;
wire _06476_ ;
wire _06477_ ;
wire _06478_ ;
wire _06479_ ;
wire _06480_ ;
wire _06481_ ;
wire _06482_ ;
wire _06483_ ;
wire _06484_ ;
wire _06485_ ;
wire _06486_ ;
wire _06487_ ;
wire _06488_ ;
wire _06489_ ;
wire _06490_ ;
wire _06491_ ;
wire _06492_ ;
wire _06493_ ;
wire _06494_ ;
wire _06495_ ;
wire _06496_ ;
wire _06497_ ;
wire _06498_ ;
wire _06499_ ;
wire _06500_ ;
wire _06501_ ;
wire _06502_ ;
wire _06503_ ;
wire _06504_ ;
wire _06505_ ;
wire _06506_ ;
wire _06507_ ;
wire _06508_ ;
wire _06509_ ;
wire _06510_ ;
wire _06511_ ;
wire _06512_ ;
wire _06513_ ;
wire _06514_ ;
wire _06515_ ;
wire _06516_ ;
wire _06517_ ;
wire _06518_ ;
wire _06519_ ;
wire _06520_ ;
wire _06521_ ;
wire _06522_ ;
wire _06523_ ;
wire _06524_ ;
wire _06525_ ;
wire _06526_ ;
wire _06527_ ;
wire _06528_ ;
wire _06529_ ;
wire _06530_ ;
wire _06531_ ;
wire _06532_ ;
wire _06533_ ;
wire _06534_ ;
wire _06535_ ;
wire _06536_ ;
wire _06537_ ;
wire _06538_ ;
wire _06539_ ;
wire _06540_ ;
wire _06541_ ;
wire _06542_ ;
wire _06543_ ;
wire _06544_ ;
wire _06545_ ;
wire _06546_ ;
wire _06547_ ;
wire _06548_ ;
wire _06549_ ;
wire _06550_ ;
wire _06551_ ;
wire _06552_ ;
wire _06553_ ;
wire _06554_ ;
wire _06555_ ;
wire _06556_ ;
wire _06557_ ;
wire _06558_ ;
wire _06559_ ;
wire _06560_ ;
wire _06561_ ;
wire _06562_ ;
wire _06563_ ;
wire _06564_ ;
wire _06565_ ;
wire _06566_ ;
wire _06567_ ;
wire _06568_ ;
wire _06569_ ;
wire _06570_ ;
wire _06571_ ;
wire _06572_ ;
wire _06573_ ;
wire _06574_ ;
wire _06575_ ;
wire _06576_ ;
wire _06577_ ;
wire _06578_ ;
wire _06579_ ;
wire _06580_ ;
wire _06581_ ;
wire _06582_ ;
wire _06583_ ;
wire _06584_ ;
wire _06585_ ;
wire _06586_ ;
wire _06587_ ;
wire _06588_ ;
wire _06589_ ;
wire _06590_ ;
wire _06591_ ;
wire _06592_ ;
wire _06593_ ;
wire _06594_ ;
wire _06595_ ;
wire _06596_ ;
wire _06597_ ;
wire _06598_ ;
wire _06599_ ;
wire _06600_ ;
wire _06601_ ;
wire _06602_ ;
wire _06603_ ;
wire _06604_ ;
wire _06605_ ;
wire _06606_ ;
wire _06607_ ;
wire _06608_ ;
wire _06609_ ;
wire _06610_ ;
wire _06611_ ;
wire _06612_ ;
wire _06613_ ;
wire _06614_ ;
wire _06615_ ;
wire _06616_ ;
wire _06617_ ;
wire _06618_ ;
wire _06619_ ;
wire _06620_ ;
wire _06621_ ;
wire _06622_ ;
wire _06623_ ;
wire _06624_ ;
wire _06625_ ;
wire _06626_ ;
wire _06627_ ;
wire _06628_ ;
wire _06629_ ;
wire _06630_ ;
wire _06631_ ;
wire _06632_ ;
wire _06633_ ;
wire _06634_ ;
wire _06635_ ;
wire _06636_ ;
wire _06637_ ;
wire _06638_ ;
wire _06639_ ;
wire _06640_ ;
wire _06641_ ;
wire _06642_ ;
wire _06643_ ;
wire _06644_ ;
wire _06645_ ;
wire _06646_ ;
wire _06647_ ;
wire _06648_ ;
wire _06649_ ;
wire _06650_ ;
wire _06651_ ;
wire _06652_ ;
wire _06653_ ;
wire _06654_ ;
wire _06655_ ;
wire _06656_ ;
wire _06657_ ;
wire _06658_ ;
wire _06659_ ;
wire _06660_ ;
wire _06661_ ;
wire _06662_ ;
wire _06663_ ;
wire _06664_ ;
wire _06665_ ;
wire _06666_ ;
wire _06667_ ;
wire _06668_ ;
wire _06669_ ;
wire _06670_ ;
wire _06671_ ;
wire _06672_ ;
wire _06673_ ;
wire _06674_ ;
wire _06675_ ;
wire _06676_ ;
wire _06677_ ;
wire _06678_ ;
wire _06679_ ;
wire _06680_ ;
wire _06681_ ;
wire _06682_ ;
wire _06683_ ;
wire _06684_ ;
wire _06685_ ;
wire _06686_ ;
wire _06687_ ;
wire _06688_ ;
wire _06689_ ;
wire _06690_ ;
wire _06691_ ;
wire _06692_ ;
wire _06693_ ;
wire _06694_ ;
wire _06695_ ;
wire _06696_ ;
wire _06697_ ;
wire _06698_ ;
wire _06699_ ;
wire _06700_ ;
wire _06701_ ;
wire _06702_ ;
wire _06703_ ;
wire _06704_ ;
wire _06705_ ;
wire _06706_ ;
wire _06707_ ;
wire _06708_ ;
wire _06709_ ;
wire _06710_ ;
wire _06711_ ;
wire _06712_ ;
wire _06713_ ;
wire _06714_ ;
wire _06715_ ;
wire _06716_ ;
wire _06717_ ;
wire _06718_ ;
wire _06719_ ;
wire _06720_ ;
wire _06721_ ;
wire _06722_ ;
wire _06723_ ;
wire _06724_ ;
wire _06725_ ;
wire _06726_ ;
wire _06727_ ;
wire _06728_ ;
wire _06729_ ;
wire _06730_ ;
wire _06731_ ;
wire _06732_ ;
wire _06733_ ;
wire _06734_ ;
wire _06735_ ;
wire _06736_ ;
wire _06737_ ;
wire _06738_ ;
wire _06739_ ;
wire _06740_ ;
wire _06741_ ;
wire _06742_ ;
wire _06743_ ;
wire _06744_ ;
wire _06745_ ;
wire _06746_ ;
wire _06747_ ;
wire _06748_ ;
wire _06749_ ;
wire _06750_ ;
wire _06751_ ;
wire _06752_ ;
wire _06753_ ;
wire _06754_ ;
wire _06755_ ;
wire _06756_ ;
wire _06757_ ;
wire _06758_ ;
wire _06759_ ;
wire _06760_ ;
wire _06761_ ;
wire _06762_ ;
wire _06763_ ;
wire _06764_ ;
wire _06765_ ;
wire _06766_ ;
wire _06767_ ;
wire _06768_ ;
wire _06769_ ;
wire _06770_ ;
wire _06771_ ;
wire _06772_ ;
wire _06773_ ;
wire _06774_ ;
wire _06775_ ;
wire _06776_ ;
wire _06777_ ;
wire _06778_ ;
wire _06779_ ;
wire _06780_ ;
wire _06781_ ;
wire _06782_ ;
wire _06783_ ;
wire _06784_ ;
wire _06785_ ;
wire _06786_ ;
wire _06787_ ;
wire _06788_ ;
wire _06789_ ;
wire _06790_ ;
wire _06791_ ;
wire _06792_ ;
wire _06793_ ;
wire _06794_ ;
wire _06795_ ;
wire _06796_ ;
wire _06797_ ;
wire _06798_ ;
wire _06799_ ;
wire _06800_ ;
wire _06801_ ;
wire _06802_ ;
wire _06803_ ;
wire _06804_ ;
wire _06805_ ;
wire _06806_ ;
wire _06807_ ;
wire _06808_ ;
wire _06809_ ;
wire _06810_ ;
wire _06811_ ;
wire _06812_ ;
wire _06813_ ;
wire _06814_ ;
wire _06815_ ;
wire _06816_ ;
wire _06817_ ;
wire _06818_ ;
wire _06819_ ;
wire _06820_ ;
wire _06821_ ;
wire _06822_ ;
wire _06823_ ;
wire _06824_ ;
wire _06825_ ;
wire _06826_ ;
wire _06827_ ;
wire _06828_ ;
wire _06829_ ;
wire _06830_ ;
wire _06831_ ;
wire _06832_ ;
wire _06833_ ;
wire _06834_ ;
wire _06835_ ;
wire _06836_ ;
wire _06837_ ;
wire _06838_ ;
wire _06839_ ;
wire _06840_ ;
wire _06841_ ;
wire _06842_ ;
wire _06843_ ;
wire _06844_ ;
wire _06845_ ;
wire _06846_ ;
wire _06847_ ;
wire _06848_ ;
wire _06849_ ;
wire _06850_ ;
wire _06851_ ;
wire _06852_ ;
wire _06853_ ;
wire _06854_ ;
wire _06855_ ;
wire _06856_ ;
wire _06857_ ;
wire _06858_ ;
wire _06859_ ;
wire _06860_ ;
wire _06861_ ;
wire _06862_ ;
wire _06863_ ;
wire _06864_ ;
wire _06865_ ;
wire _06866_ ;
wire _06867_ ;
wire _06868_ ;
wire _06869_ ;
wire _06870_ ;
wire _06871_ ;
wire _06872_ ;
wire _06873_ ;
wire _06874_ ;
wire _06875_ ;
wire _06876_ ;
wire _06877_ ;
wire _06878_ ;
wire _06879_ ;
wire _06880_ ;
wire _06881_ ;
wire _06882_ ;
wire _06883_ ;
wire _06884_ ;
wire _06885_ ;
wire _06886_ ;
wire _06887_ ;
wire _06888_ ;
wire _06889_ ;
wire _06890_ ;
wire _06891_ ;
wire _06892_ ;
wire _06893_ ;
wire _06894_ ;
wire _06895_ ;
wire _06896_ ;
wire _06897_ ;
wire _06898_ ;
wire _06899_ ;
wire _06900_ ;
wire _06901_ ;
wire _06902_ ;
wire _06903_ ;
wire _06904_ ;
wire _06905_ ;
wire _06906_ ;
wire _06907_ ;
wire _06908_ ;
wire _06909_ ;
wire _06910_ ;
wire _06911_ ;
wire _06912_ ;
wire _06913_ ;
wire _06914_ ;
wire _06915_ ;
wire _06916_ ;
wire _06917_ ;
wire _06918_ ;
wire _06919_ ;
wire _06920_ ;
wire _06921_ ;
wire _06922_ ;
wire _06923_ ;
wire _06924_ ;
wire _06925_ ;
wire _06926_ ;
wire _06927_ ;
wire _06928_ ;
wire _06929_ ;
wire _06930_ ;
wire _06931_ ;
wire _06932_ ;
wire _06933_ ;
wire _06934_ ;
wire _06935_ ;
wire _06936_ ;
wire _06937_ ;
wire _06938_ ;
wire _06939_ ;
wire _06940_ ;
wire _06941_ ;
wire _06942_ ;
wire _06943_ ;
wire _06944_ ;
wire _06945_ ;
wire _06946_ ;
wire _06947_ ;
wire _06948_ ;
wire _06949_ ;
wire _06950_ ;
wire _06951_ ;
wire _06952_ ;
wire _06953_ ;
wire _06954_ ;
wire _06955_ ;
wire _06956_ ;
wire _06957_ ;
wire _06958_ ;
wire _06959_ ;
wire _06960_ ;
wire _06961_ ;
wire _06962_ ;
wire _06963_ ;
wire _06964_ ;
wire _06965_ ;
wire _06966_ ;
wire _06967_ ;
wire _06968_ ;
wire _06969_ ;
wire _06970_ ;
wire _06971_ ;
wire _06972_ ;
wire _06973_ ;
wire _06974_ ;
wire _06975_ ;
wire _06976_ ;
wire _06977_ ;
wire _06978_ ;
wire _06979_ ;
wire _06980_ ;
wire _06981_ ;
wire _06982_ ;
wire _06983_ ;
wire _06984_ ;
wire _06985_ ;
wire _06986_ ;
wire _06987_ ;
wire _06988_ ;
wire _06989_ ;
wire _06990_ ;
wire _06991_ ;
wire _06992_ ;
wire _06993_ ;
wire _06994_ ;
wire _06995_ ;
wire _06996_ ;
wire _06997_ ;
wire _06998_ ;
wire _06999_ ;
wire _07000_ ;
wire _07001_ ;
wire _07002_ ;
wire _07003_ ;
wire _07004_ ;
wire _07005_ ;
wire _07006_ ;
wire _07007_ ;
wire _07008_ ;
wire _07009_ ;
wire _07010_ ;
wire _07011_ ;
wire _07012_ ;
wire _07013_ ;
wire _07014_ ;
wire _07015_ ;
wire _07016_ ;
wire _07017_ ;
wire _07018_ ;
wire _07019_ ;
wire _07020_ ;
wire _07021_ ;
wire _07022_ ;
wire _07023_ ;
wire _07024_ ;
wire _07025_ ;
wire _07026_ ;
wire _07027_ ;
wire _07028_ ;
wire _07029_ ;
wire _07030_ ;
wire _07031_ ;
wire _07032_ ;
wire _07033_ ;
wire _07034_ ;
wire _07035_ ;
wire _07036_ ;
wire _07037_ ;
wire _07038_ ;
wire _07039_ ;
wire _07040_ ;
wire _07041_ ;
wire _07042_ ;
wire _07043_ ;
wire _07044_ ;
wire _07045_ ;
wire _07046_ ;
wire _07047_ ;
wire _07048_ ;
wire _07049_ ;
wire _07050_ ;
wire _07051_ ;
wire _07052_ ;
wire _07053_ ;
wire _07054_ ;
wire _07055_ ;
wire _07056_ ;
wire _07057_ ;
wire _07058_ ;
wire _07059_ ;
wire _07060_ ;
wire _07061_ ;
wire _07062_ ;
wire _07063_ ;
wire _07064_ ;
wire _07065_ ;
wire _07066_ ;
wire _07067_ ;
wire _07068_ ;
wire _07069_ ;
wire _07070_ ;
wire _07071_ ;
wire _07072_ ;
wire _07073_ ;
wire _07074_ ;
wire _07075_ ;
wire _07076_ ;
wire _07077_ ;
wire _07078_ ;
wire _07079_ ;
wire _07080_ ;
wire _07081_ ;
wire _07082_ ;
wire _07083_ ;
wire _07084_ ;
wire _07085_ ;
wire _07086_ ;
wire _07087_ ;
wire _07088_ ;
wire _07089_ ;
wire _07090_ ;
wire _07091_ ;
wire _07092_ ;
wire _07093_ ;
wire _07094_ ;
wire _07095_ ;
wire _07096_ ;
wire _07097_ ;
wire _07098_ ;
wire _07099_ ;
wire _07100_ ;
wire _07101_ ;
wire _07102_ ;
wire _07103_ ;
wire _07104_ ;
wire _07105_ ;
wire _07106_ ;
wire _07107_ ;
wire _07108_ ;
wire _07109_ ;
wire _07110_ ;
wire _07111_ ;
wire _07112_ ;
wire _07113_ ;
wire _07114_ ;
wire _07115_ ;
wire _07116_ ;
wire _07117_ ;
wire _07118_ ;
wire _07119_ ;
wire _07120_ ;
wire _07121_ ;
wire _07122_ ;
wire _07123_ ;
wire _07124_ ;
wire _07125_ ;
wire _07126_ ;
wire _07127_ ;
wire _07128_ ;
wire _07129_ ;
wire _07130_ ;
wire _07131_ ;
wire _07132_ ;
wire _07133_ ;
wire _07134_ ;
wire _07135_ ;
wire _07136_ ;
wire _07137_ ;
wire _07138_ ;
wire _07139_ ;
wire _07140_ ;
wire _07141_ ;
wire _07142_ ;
wire _07143_ ;
wire _07144_ ;
wire _07145_ ;
wire _07146_ ;
wire _07147_ ;
wire _07148_ ;
wire _07149_ ;
wire _07150_ ;
wire _07151_ ;
wire _07152_ ;
wire _07153_ ;
wire _07154_ ;
wire _07155_ ;
wire _07156_ ;
wire _07157_ ;
wire _07158_ ;
wire _07159_ ;
wire _07160_ ;
wire _07161_ ;
wire _07162_ ;
wire _07163_ ;
wire _07164_ ;
wire _07165_ ;
wire _07166_ ;
wire _07167_ ;
wire _07168_ ;
wire _07169_ ;
wire _07170_ ;
wire _07171_ ;
wire _07172_ ;
wire _07173_ ;
wire _07174_ ;
wire _07175_ ;
wire _07176_ ;
wire _07177_ ;
wire _07178_ ;
wire _07179_ ;
wire _07180_ ;
wire _07181_ ;
wire _07182_ ;
wire _07183_ ;
wire _07184_ ;
wire _07185_ ;
wire _07186_ ;
wire _07187_ ;
wire _07188_ ;
wire _07189_ ;
wire _07190_ ;
wire _07191_ ;
wire _07192_ ;
wire _07193_ ;
wire _07194_ ;
wire _07195_ ;
wire _07196_ ;
wire _07197_ ;
wire _07198_ ;
wire _07199_ ;
wire _07200_ ;
wire _07201_ ;
wire _07202_ ;
wire _07203_ ;
wire _07204_ ;
wire _07205_ ;
wire _07206_ ;
wire _07207_ ;
wire _07208_ ;
wire _07209_ ;
wire _07210_ ;
wire _07211_ ;
wire _07212_ ;
wire _07213_ ;
wire _07214_ ;
wire _07215_ ;
wire _07216_ ;
wire _07217_ ;
wire _07218_ ;
wire _07219_ ;
wire _07220_ ;
wire _07221_ ;
wire _07222_ ;
wire _07223_ ;
wire _07224_ ;
wire _07225_ ;
wire _07226_ ;
wire _07227_ ;
wire _07228_ ;
wire _07229_ ;
wire _07230_ ;
wire _07231_ ;
wire _07232_ ;
wire _07233_ ;
wire _07234_ ;
wire _07235_ ;
wire _07236_ ;
wire _07237_ ;
wire _07238_ ;
wire _07239_ ;
wire _07240_ ;
wire _07241_ ;
wire _07242_ ;
wire _07243_ ;
wire _07244_ ;
wire _07245_ ;
wire _07246_ ;
wire _07247_ ;
wire _07248_ ;
wire _07249_ ;
wire _07250_ ;
wire _07251_ ;
wire _07252_ ;
wire _07253_ ;
wire _07254_ ;
wire _07255_ ;
wire _07256_ ;
wire _07257_ ;
wire _07258_ ;
wire _07259_ ;
wire _07260_ ;
wire _07261_ ;
wire _07262_ ;
wire _07263_ ;
wire _07264_ ;
wire _07265_ ;
wire _07266_ ;
wire _07267_ ;
wire _07268_ ;
wire _07269_ ;
wire _07270_ ;
wire _07271_ ;
wire _07272_ ;
wire _07273_ ;
wire _07274_ ;
wire _07275_ ;
wire _07276_ ;
wire _07277_ ;
wire _07278_ ;
wire _07279_ ;
wire _07280_ ;
wire _07281_ ;
wire _07282_ ;
wire _07283_ ;
wire _07284_ ;
wire _07285_ ;
wire _07286_ ;
wire _07287_ ;
wire _07288_ ;
wire _07289_ ;
wire _07290_ ;
wire _07291_ ;
wire _07292_ ;
wire _07293_ ;
wire _07294_ ;
wire _07295_ ;
wire _07296_ ;
wire _07297_ ;
wire _07298_ ;
wire _07299_ ;
wire _07300_ ;
wire _07301_ ;
wire _07302_ ;
wire _07303_ ;
wire _07304_ ;
wire _07305_ ;
wire _07306_ ;
wire _07307_ ;
wire _07308_ ;
wire _07309_ ;
wire _07310_ ;
wire _07311_ ;
wire _07312_ ;
wire _07313_ ;
wire _07314_ ;
wire _07315_ ;
wire _07316_ ;
wire _07317_ ;
wire _07318_ ;
wire _07319_ ;
wire _07320_ ;
wire _07321_ ;
wire _07322_ ;
wire _07323_ ;
wire _07324_ ;
wire _07325_ ;
wire _07326_ ;
wire _07327_ ;
wire _07328_ ;
wire _07329_ ;
wire _07330_ ;
wire _07331_ ;
wire _07332_ ;
wire _07333_ ;
wire _07334_ ;
wire _07335_ ;
wire _07336_ ;
wire _07337_ ;
wire _07338_ ;
wire _07339_ ;
wire _07340_ ;
wire _07341_ ;
wire _07342_ ;
wire _07343_ ;
wire _07344_ ;
wire _07345_ ;
wire _07346_ ;
wire _07347_ ;
wire _07348_ ;
wire _07349_ ;
wire _07350_ ;
wire _07351_ ;
wire _07352_ ;
wire _07353_ ;
wire _07354_ ;
wire _07355_ ;
wire _07356_ ;
wire _07357_ ;
wire _07358_ ;
wire _07359_ ;
wire _07360_ ;
wire _07361_ ;
wire _07362_ ;
wire _07363_ ;
wire _07364_ ;
wire _07365_ ;
wire _07366_ ;
wire _07367_ ;
wire _07368_ ;
wire _07369_ ;
wire _07370_ ;
wire _07371_ ;
wire _07372_ ;
wire _07373_ ;
wire _07374_ ;
wire _07375_ ;
wire _07376_ ;
wire _07377_ ;
wire _07378_ ;
wire _07379_ ;
wire _07380_ ;
wire _07381_ ;
wire _07382_ ;
wire _07383_ ;
wire _07384_ ;
wire _07385_ ;
wire _07386_ ;
wire _07387_ ;
wire _07388_ ;
wire _07389_ ;
wire _07390_ ;
wire _07391_ ;
wire _07392_ ;
wire _07393_ ;
wire _07394_ ;
wire _07395_ ;
wire _07396_ ;
wire _07397_ ;
wire _07398_ ;
wire _07399_ ;
wire _07400_ ;
wire _07401_ ;
wire _07402_ ;
wire _07403_ ;
wire _07404_ ;
wire _07405_ ;
wire _07406_ ;
wire _07407_ ;
wire _07408_ ;
wire _07409_ ;
wire _07410_ ;
wire _07411_ ;
wire _07412_ ;
wire _07413_ ;
wire _07414_ ;
wire _07415_ ;
wire _07416_ ;
wire _07417_ ;
wire _07418_ ;
wire _07419_ ;
wire _07420_ ;
wire _07421_ ;
wire _07422_ ;
wire _07423_ ;
wire _07424_ ;
wire _07425_ ;
wire _07426_ ;
wire _07427_ ;
wire _07428_ ;
wire _07429_ ;
wire _07430_ ;
wire _07431_ ;
wire _07432_ ;
wire _07433_ ;
wire _07434_ ;
wire _07435_ ;
wire _07436_ ;
wire _07437_ ;
wire _07438_ ;
wire _07439_ ;
wire _07440_ ;
wire _07441_ ;
wire _07442_ ;
wire _07443_ ;
wire _07444_ ;
wire _07445_ ;
wire _07446_ ;
wire _07447_ ;
wire _07448_ ;
wire _07449_ ;
wire _07450_ ;
wire _07451_ ;
wire _07452_ ;
wire _07453_ ;
wire _07454_ ;
wire _07455_ ;
wire _07456_ ;
wire _07457_ ;
wire _07458_ ;
wire _07459_ ;
wire _07460_ ;
wire _07461_ ;
wire _07462_ ;
wire _07463_ ;
wire _07464_ ;
wire _07465_ ;
wire _07466_ ;
wire _07467_ ;
wire _07468_ ;
wire _07469_ ;
wire _07470_ ;
wire _07471_ ;
wire _07472_ ;
wire _07473_ ;
wire _07474_ ;
wire _07475_ ;
wire _07476_ ;
wire _07477_ ;
wire _07478_ ;
wire _07479_ ;
wire _07480_ ;
wire _07481_ ;
wire _07482_ ;
wire _07483_ ;
wire _07484_ ;
wire _07485_ ;
wire _07486_ ;
wire _07487_ ;
wire _07488_ ;
wire _07489_ ;
wire _07490_ ;
wire _07491_ ;
wire _07492_ ;
wire _07493_ ;
wire _07494_ ;
wire _07495_ ;
wire _07496_ ;
wire _07497_ ;
wire _07498_ ;
wire _07499_ ;
wire _07500_ ;
wire _07501_ ;
wire _07502_ ;
wire _07503_ ;
wire _07504_ ;
wire _07505_ ;
wire _07506_ ;
wire _07507_ ;
wire _07508_ ;
wire _07509_ ;
wire _07510_ ;
wire _07511_ ;
wire _07512_ ;
wire _07513_ ;
wire _07514_ ;
wire _07515_ ;
wire _07516_ ;
wire _07517_ ;
wire _07518_ ;
wire _07519_ ;
wire _07520_ ;
wire _07521_ ;
wire _07522_ ;
wire _07523_ ;
wire _07524_ ;
wire _07525_ ;
wire _07526_ ;
wire _07527_ ;
wire _07528_ ;
wire _07529_ ;
wire _07530_ ;
wire _07531_ ;
wire _07532_ ;
wire _07533_ ;
wire _07534_ ;
wire _07535_ ;
wire _07536_ ;
wire _07537_ ;
wire _07538_ ;
wire _07539_ ;
wire _07540_ ;
wire _07541_ ;
wire _07542_ ;
wire _07543_ ;
wire _07544_ ;
wire _07545_ ;
wire _07546_ ;
wire _07547_ ;
wire _07548_ ;
wire _07549_ ;
wire _07550_ ;
wire _07551_ ;
wire _07552_ ;
wire _07553_ ;
wire _07554_ ;
wire _07555_ ;
wire _07556_ ;
wire _07557_ ;
wire _07558_ ;
wire _07559_ ;
wire _07560_ ;
wire _07561_ ;
wire _07562_ ;
wire _07563_ ;
wire _07564_ ;
wire _07565_ ;
wire _07566_ ;
wire _07567_ ;
wire _07568_ ;
wire _07569_ ;
wire _07570_ ;
wire _07571_ ;
wire _07572_ ;
wire _07573_ ;
wire _07574_ ;
wire _07575_ ;
wire _07576_ ;
wire _07577_ ;
wire _07578_ ;
wire _07579_ ;
wire _07580_ ;
wire _07581_ ;
wire _07582_ ;
wire _07583_ ;
wire _07584_ ;
wire _07585_ ;
wire _07586_ ;
wire _07587_ ;
wire _07588_ ;
wire _07589_ ;
wire _07590_ ;
wire _07591_ ;
wire _07592_ ;
wire _07593_ ;
wire _07594_ ;
wire _07595_ ;
wire _07596_ ;
wire _07597_ ;
wire _07598_ ;
wire _07599_ ;
wire _07600_ ;
wire _07601_ ;
wire _07602_ ;
wire _07603_ ;
wire _07604_ ;
wire _07605_ ;
wire _07606_ ;
wire _07607_ ;
wire _07608_ ;
wire _07609_ ;
wire _07610_ ;
wire _07611_ ;
wire _07612_ ;
wire _07613_ ;
wire _07614_ ;
wire _07615_ ;
wire _07616_ ;
wire _07617_ ;
wire _07618_ ;
wire _07619_ ;
wire _07620_ ;
wire _07621_ ;
wire _07622_ ;
wire _07623_ ;
wire _07624_ ;
wire _07625_ ;
wire _07626_ ;
wire _07627_ ;
wire _07628_ ;
wire _07629_ ;
wire _07630_ ;
wire _07631_ ;
wire _07632_ ;
wire _07633_ ;
wire _07634_ ;
wire _07635_ ;
wire _07636_ ;
wire _07637_ ;
wire _07638_ ;
wire _07639_ ;
wire _07640_ ;
wire _07641_ ;
wire _07642_ ;
wire _07643_ ;
wire _07644_ ;
wire _07645_ ;
wire _07646_ ;
wire _07647_ ;
wire _07648_ ;
wire _07649_ ;
wire _07650_ ;
wire _07651_ ;
wire _07652_ ;
wire _07653_ ;
wire _07654_ ;
wire _07655_ ;
wire _07656_ ;
wire _07657_ ;
wire _07658_ ;
wire _07659_ ;
wire _07660_ ;
wire _07661_ ;
wire _07662_ ;
wire _07663_ ;
wire _07664_ ;
wire _07665_ ;
wire _07666_ ;
wire _07667_ ;
wire _07668_ ;
wire _07669_ ;
wire _07670_ ;
wire _07671_ ;
wire _07672_ ;
wire _07673_ ;
wire _07674_ ;
wire _07675_ ;
wire _07676_ ;
wire _07677_ ;
wire _07678_ ;
wire _07679_ ;
wire _07680_ ;
wire _07681_ ;
wire _07682_ ;
wire _07683_ ;
wire _07684_ ;
wire _07685_ ;
wire _07686_ ;
wire _07687_ ;
wire _07688_ ;
wire _07689_ ;
wire _07690_ ;
wire _07691_ ;
wire _07692_ ;
wire _07693_ ;
wire _07694_ ;
wire _07695_ ;
wire _07696_ ;
wire _07697_ ;
wire _07698_ ;
wire _07699_ ;
wire _07700_ ;
wire _07701_ ;
wire _07702_ ;
wire _07703_ ;
wire _07704_ ;
wire _07705_ ;
wire _07706_ ;
wire _07707_ ;
wire _07708_ ;
wire _07709_ ;
wire _07710_ ;
wire _07711_ ;
wire _07712_ ;
wire _07713_ ;
wire _07714_ ;
wire _07715_ ;
wire _07716_ ;
wire _07717_ ;
wire _07718_ ;
wire _07719_ ;
wire _07720_ ;
wire _07721_ ;
wire _07722_ ;
wire _07723_ ;
wire _07724_ ;
wire _07725_ ;
wire _07726_ ;
wire _07727_ ;
wire _07728_ ;
wire _07729_ ;
wire _07730_ ;
wire _07731_ ;
wire _07732_ ;
wire _07733_ ;
wire _07734_ ;
wire _07735_ ;
wire _07736_ ;
wire _07737_ ;
wire _07738_ ;
wire _07739_ ;
wire _07740_ ;
wire _07741_ ;
wire _07742_ ;
wire _07743_ ;
wire _07744_ ;
wire _07745_ ;
wire _07746_ ;
wire _07747_ ;
wire _07748_ ;
wire _07749_ ;
wire _07750_ ;
wire _07751_ ;
wire _07752_ ;
wire _07753_ ;
wire _07754_ ;
wire _07755_ ;
wire _07756_ ;
wire _07757_ ;
wire _07758_ ;
wire _07759_ ;
wire _07760_ ;
wire _07761_ ;
wire _07762_ ;
wire _07763_ ;
wire _07764_ ;
wire _07765_ ;
wire _07766_ ;
wire _07767_ ;
wire _07768_ ;
wire _07769_ ;
wire _07770_ ;
wire _07771_ ;
wire _07772_ ;
wire _07773_ ;
wire _07774_ ;
wire _07775_ ;
wire _07776_ ;
wire _07777_ ;
wire _07778_ ;
wire _07779_ ;
wire _07780_ ;
wire _07781_ ;
wire _07782_ ;
wire _07783_ ;
wire _07784_ ;
wire _07785_ ;
wire _07786_ ;
wire _07787_ ;
wire _07788_ ;
wire _07789_ ;
wire _07790_ ;
wire _07791_ ;
wire _07792_ ;
wire _07793_ ;
wire _07794_ ;
wire _07795_ ;
wire _07796_ ;
wire _07797_ ;
wire _07798_ ;
wire _07799_ ;
wire _07800_ ;
wire _07801_ ;
wire _07802_ ;
wire _07803_ ;
wire _07804_ ;
wire _07805_ ;
wire _07806_ ;
wire _07807_ ;
wire _07808_ ;
wire _07809_ ;
wire _07810_ ;
wire _07811_ ;
wire _07812_ ;
wire _07813_ ;
wire _07814_ ;
wire _07815_ ;
wire _07816_ ;
wire _07817_ ;
wire _07818_ ;
wire _07819_ ;
wire _07820_ ;
wire _07821_ ;
wire _07822_ ;
wire _07823_ ;
wire _07824_ ;
wire _07825_ ;
wire _07826_ ;
wire _07827_ ;
wire _07828_ ;
wire _07829_ ;
wire _07830_ ;
wire _07831_ ;
wire _07832_ ;
wire _07833_ ;
wire _07834_ ;
wire _07835_ ;
wire _07836_ ;
wire _07837_ ;
wire _07838_ ;
wire _07839_ ;
wire _07840_ ;
wire _07841_ ;
wire _07842_ ;
wire _07843_ ;
wire _07844_ ;
wire _07845_ ;
wire _07846_ ;
wire _07847_ ;
wire _07848_ ;
wire _07849_ ;
wire _07850_ ;
wire _07851_ ;
wire _07852_ ;
wire _07853_ ;
wire _07854_ ;
wire _07855_ ;
wire _07856_ ;
wire _07857_ ;
wire _07858_ ;
wire _07859_ ;
wire _07860_ ;
wire _07861_ ;
wire _07862_ ;
wire _07863_ ;
wire _07864_ ;
wire _07865_ ;
wire _07866_ ;
wire _07867_ ;
wire _07868_ ;
wire _07869_ ;
wire _07870_ ;
wire _07871_ ;
wire _07872_ ;
wire _07873_ ;
wire _07874_ ;
wire _07875_ ;
wire _07876_ ;
wire _07877_ ;
wire _07878_ ;
wire _07879_ ;
wire _07880_ ;
wire _07881_ ;
wire _07882_ ;
wire _07883_ ;
wire _07884_ ;
wire _07885_ ;
wire _07886_ ;
wire _07887_ ;
wire _07888_ ;
wire _07889_ ;
wire _07890_ ;
wire _07891_ ;
wire _07892_ ;
wire _07893_ ;
wire _07894_ ;
wire _07895_ ;
wire _07896_ ;
wire _07897_ ;
wire _07898_ ;
wire _07899_ ;
wire _07900_ ;
wire _07901_ ;
wire _07902_ ;
wire _07903_ ;
wire _07904_ ;
wire _07905_ ;
wire _07906_ ;
wire _07907_ ;
wire _07908_ ;
wire _07909_ ;
wire _07910_ ;
wire _07911_ ;
wire _07912_ ;
wire _07913_ ;
wire _07914_ ;
wire _07915_ ;
wire _07916_ ;
wire _07917_ ;
wire _07918_ ;
wire _07919_ ;
wire _07920_ ;
wire _07921_ ;
wire _07922_ ;
wire _07923_ ;
wire _07924_ ;
wire _07925_ ;
wire _07926_ ;
wire _07927_ ;
wire _07928_ ;
wire _07929_ ;
wire _07930_ ;
wire _07931_ ;
wire _07932_ ;
wire _07933_ ;
wire _07934_ ;
wire _07935_ ;
wire _07936_ ;
wire _07937_ ;
wire _07938_ ;
wire _07939_ ;
wire _07940_ ;
wire _07941_ ;
wire _07942_ ;
wire _07943_ ;
wire _07944_ ;
wire _07945_ ;
wire _07946_ ;
wire _07947_ ;
wire _07948_ ;
wire _07949_ ;
wire _07950_ ;
wire _07951_ ;
wire _07952_ ;
wire _07953_ ;
wire _07954_ ;
wire _07955_ ;
wire _07956_ ;
wire _07957_ ;
wire _07958_ ;
wire _07959_ ;
wire _07960_ ;
wire _07961_ ;
wire _07962_ ;
wire _07963_ ;
wire _07964_ ;
wire _07965_ ;
wire _07966_ ;
wire _07967_ ;
wire _07968_ ;
wire _07969_ ;
wire _07970_ ;
wire _07971_ ;
wire _07972_ ;
wire _07973_ ;
wire _07974_ ;
wire _07975_ ;
wire _07976_ ;
wire _07977_ ;
wire _07978_ ;
wire _07979_ ;
wire _07980_ ;
wire _07981_ ;
wire _07982_ ;
wire _07983_ ;
wire _07984_ ;
wire _07985_ ;
wire _07986_ ;
wire _07987_ ;
wire _07988_ ;
wire _07989_ ;
wire _07990_ ;
wire _07991_ ;
wire _07992_ ;
wire _07993_ ;
wire _07994_ ;
wire _07995_ ;
wire _07996_ ;
wire _07997_ ;
wire _07998_ ;
wire _07999_ ;
wire _08000_ ;
wire _08001_ ;
wire _08002_ ;
wire _08003_ ;
wire _08004_ ;
wire _08005_ ;
wire _08006_ ;
wire _08007_ ;
wire _08008_ ;
wire _08009_ ;
wire _08010_ ;
wire _08011_ ;
wire _08012_ ;
wire _08013_ ;
wire _08014_ ;
wire _08015_ ;
wire _08016_ ;
wire _08017_ ;
wire _08018_ ;
wire _08019_ ;
wire _08020_ ;
wire _08021_ ;
wire _08022_ ;
wire _08023_ ;
wire _08024_ ;
wire _08025_ ;
wire _08026_ ;
wire _08027_ ;
wire _08028_ ;
wire _08029_ ;
wire _08030_ ;
wire _08031_ ;
wire _08032_ ;
wire _08033_ ;
wire _08034_ ;
wire _08035_ ;
wire _08036_ ;
wire _08037_ ;
wire _08038_ ;
wire _08039_ ;
wire _08040_ ;
wire _08041_ ;
wire _08042_ ;
wire _08043_ ;
wire _08044_ ;
wire _08045_ ;
wire _08046_ ;
wire _08047_ ;
wire _08048_ ;
wire _08049_ ;
wire _08050_ ;
wire _08051_ ;
wire _08052_ ;
wire _08053_ ;
wire _08054_ ;
wire _08055_ ;
wire _08056_ ;
wire _08057_ ;
wire _08058_ ;
wire _08059_ ;
wire _08060_ ;
wire _08061_ ;
wire _08062_ ;
wire _08063_ ;
wire _08064_ ;
wire _08065_ ;
wire _08066_ ;
wire _08067_ ;
wire _08068_ ;
wire _08069_ ;
wire _08070_ ;
wire _08071_ ;
wire _08072_ ;
wire _08073_ ;
wire _08074_ ;
wire _08075_ ;
wire _08076_ ;
wire _08077_ ;
wire _08078_ ;
wire _08079_ ;
wire _08080_ ;
wire _08081_ ;
wire _08082_ ;
wire _08083_ ;
wire _08084_ ;
wire _08085_ ;
wire _08086_ ;
wire _08087_ ;
wire _08088_ ;
wire _08089_ ;
wire _08090_ ;
wire _08091_ ;
wire _08092_ ;
wire _08093_ ;
wire _08094_ ;
wire _08095_ ;
wire _08096_ ;
wire _08097_ ;
wire _08098_ ;
wire _08099_ ;
wire _08100_ ;
wire _08101_ ;
wire _08102_ ;
wire _08103_ ;
wire _08104_ ;
wire _08105_ ;
wire _08106_ ;
wire _08107_ ;
wire _08108_ ;
wire _08109_ ;
wire _08110_ ;
wire _08111_ ;
wire _08112_ ;
wire _08113_ ;
wire _08114_ ;
wire _08115_ ;
wire _08116_ ;
wire _08117_ ;
wire _08118_ ;
wire _08119_ ;
wire _08120_ ;
wire _08121_ ;
wire _08122_ ;
wire _08123_ ;
wire _08124_ ;
wire _08125_ ;
wire _08126_ ;
wire _08127_ ;
wire _08128_ ;
wire _08129_ ;
wire _08130_ ;
wire _08131_ ;
wire _08132_ ;
wire _08133_ ;
wire _08134_ ;
wire _08135_ ;
wire _08136_ ;
wire _08137_ ;
wire _08138_ ;
wire _08139_ ;
wire _08140_ ;
wire _08141_ ;
wire _08142_ ;
wire _08143_ ;
wire _08144_ ;
wire _08145_ ;
wire _08146_ ;
wire _08147_ ;
wire _08148_ ;
wire _08149_ ;
wire _08150_ ;
wire _08151_ ;
wire _08152_ ;
wire _08153_ ;
wire _08154_ ;
wire _08155_ ;
wire _08156_ ;
wire _08157_ ;
wire _08158_ ;
wire _08159_ ;
wire _08160_ ;
wire _08161_ ;
wire _08162_ ;
wire _08163_ ;
wire _08164_ ;
wire _08165_ ;
wire _08166_ ;
wire _08167_ ;
wire _08168_ ;
wire _08169_ ;
wire _08170_ ;
wire _08171_ ;
wire _08172_ ;
wire _08173_ ;
wire _08174_ ;
wire _08175_ ;
wire _08176_ ;
wire _08177_ ;
wire _08178_ ;
wire _08179_ ;
wire _08180_ ;
wire _08181_ ;
wire _08182_ ;
wire _08183_ ;
wire _08184_ ;
wire _08185_ ;
wire _08186_ ;
wire _08187_ ;
wire _08188_ ;
wire _08189_ ;
wire _08190_ ;
wire _08191_ ;
wire _08192_ ;
wire _08193_ ;
wire _08194_ ;
wire _08195_ ;
wire _08196_ ;
wire _08197_ ;
wire _08198_ ;
wire _08199_ ;
wire _08200_ ;
wire _08201_ ;
wire _08202_ ;
wire _08203_ ;
wire _08204_ ;
wire _08205_ ;
wire _08206_ ;
wire _08207_ ;
wire _08208_ ;
wire _08209_ ;
wire _08210_ ;
wire _08211_ ;
wire _08212_ ;
wire _08213_ ;
wire _08214_ ;
wire _08215_ ;
wire _08216_ ;
wire _08217_ ;
wire _08218_ ;
wire _08219_ ;
wire _08220_ ;
wire _08221_ ;
wire _08222_ ;
wire _08223_ ;
wire _08224_ ;
wire _08225_ ;
wire _08226_ ;
wire _08227_ ;
wire _08228_ ;
wire _08229_ ;
wire _08230_ ;
wire _08231_ ;
wire _08232_ ;
wire _08233_ ;
wire _08234_ ;
wire _08235_ ;
wire _08236_ ;
wire _08237_ ;
wire _08238_ ;
wire _08239_ ;
wire _08240_ ;
wire _08241_ ;
wire _08242_ ;
wire _08243_ ;
wire _08244_ ;
wire _08245_ ;
wire _08246_ ;
wire _08247_ ;
wire _08248_ ;
wire _08249_ ;
wire _08250_ ;
wire _08251_ ;
wire _08252_ ;
wire _08253_ ;
wire _08254_ ;
wire _08255_ ;
wire _08256_ ;
wire _08257_ ;
wire _08258_ ;
wire _08259_ ;
wire _08260_ ;
wire _08261_ ;
wire _08262_ ;
wire _08263_ ;
wire _08264_ ;
wire _08265_ ;
wire _08266_ ;
wire _08267_ ;
wire _08268_ ;
wire _08269_ ;
wire _08270_ ;
wire _08271_ ;
wire _08272_ ;
wire _08273_ ;
wire _08274_ ;
wire _08275_ ;
wire _08276_ ;
wire _08277_ ;
wire _08278_ ;
wire _08279_ ;
wire _08280_ ;
wire _08281_ ;
wire _08282_ ;
wire _08283_ ;
wire _08284_ ;
wire _08285_ ;
wire _08286_ ;
wire _08287_ ;
wire _08288_ ;
wire _08289_ ;
wire _08290_ ;
wire _08291_ ;
wire _08292_ ;
wire _08293_ ;
wire _08294_ ;
wire _08295_ ;
wire _08296_ ;
wire _08297_ ;
wire _08298_ ;
wire _08299_ ;
wire _08300_ ;
wire _08301_ ;
wire _08302_ ;
wire _08303_ ;
wire _08304_ ;
wire _08305_ ;
wire _08306_ ;
wire _08307_ ;
wire _08308_ ;
wire _08309_ ;
wire _08310_ ;
wire _08311_ ;
wire _08312_ ;
wire _08313_ ;
wire _08314_ ;
wire _08315_ ;
wire _08316_ ;
wire _08317_ ;
wire _08318_ ;
wire _08319_ ;
wire _08320_ ;
wire _08321_ ;
wire _08322_ ;
wire _08323_ ;
wire _08324_ ;
wire _08325_ ;
wire _08326_ ;
wire _08327_ ;
wire _08328_ ;
wire _08329_ ;
wire _08330_ ;
wire _08331_ ;
wire _08332_ ;
wire _08333_ ;
wire _08334_ ;
wire _08335_ ;
wire _08336_ ;
wire _08337_ ;
wire _08338_ ;
wire _08339_ ;
wire _08340_ ;
wire _08341_ ;
wire _08342_ ;
wire _08343_ ;
wire _08344_ ;
wire _08345_ ;
wire _08346_ ;
wire _08347_ ;
wire _08348_ ;
wire _08349_ ;
wire _08350_ ;
wire _08351_ ;
wire _08352_ ;
wire _08353_ ;
wire _08354_ ;
wire _08355_ ;
wire _08356_ ;
wire _08357_ ;
wire _08358_ ;
wire _08359_ ;
wire _08360_ ;
wire _08361_ ;
wire _08362_ ;
wire _08363_ ;
wire _08364_ ;
wire _08365_ ;
wire _08366_ ;
wire _08367_ ;
wire _08368_ ;
wire _08369_ ;
wire _08370_ ;
wire _08371_ ;
wire _08372_ ;
wire _08373_ ;
wire _08374_ ;
wire _08375_ ;
wire _08376_ ;
wire _08377_ ;
wire _08378_ ;
wire _08379_ ;
wire _08380_ ;
wire _08381_ ;
wire _08382_ ;
wire _08383_ ;
wire _08384_ ;
wire _08385_ ;
wire _08386_ ;
wire _08387_ ;
wire _08388_ ;
wire _08389_ ;
wire _08390_ ;
wire _08391_ ;
wire _08392_ ;
wire _08393_ ;
wire _08394_ ;
wire _08395_ ;
wire _08396_ ;
wire _08397_ ;
wire _08398_ ;
wire _08399_ ;
wire _08400_ ;
wire _08401_ ;
wire _08402_ ;
wire _08403_ ;
wire _08404_ ;
wire _08405_ ;
wire _08406_ ;
wire _08407_ ;
wire _08408_ ;
wire _08409_ ;
wire _08410_ ;
wire _08411_ ;
wire _08412_ ;
wire _08413_ ;
wire _08414_ ;
wire _08415_ ;
wire _08416_ ;
wire _08417_ ;
wire _08418_ ;
wire _08419_ ;
wire _08420_ ;
wire _08421_ ;
wire _08422_ ;
wire _08423_ ;
wire _08424_ ;
wire _08425_ ;
wire _08426_ ;
wire _08427_ ;
wire _08428_ ;
wire _08429_ ;
wire _08430_ ;
wire _08431_ ;
wire _08432_ ;
wire _08433_ ;
wire _08434_ ;
wire _08435_ ;
wire _08436_ ;
wire _08437_ ;
wire _08438_ ;
wire _08439_ ;
wire _08440_ ;
wire _08441_ ;
wire _08442_ ;
wire _08443_ ;
wire _08444_ ;
wire _08445_ ;
wire _08446_ ;
wire _08447_ ;
wire _08448_ ;
wire _08449_ ;
wire _08450_ ;
wire _08451_ ;
wire _08452_ ;
wire _08453_ ;
wire _08454_ ;
wire _08455_ ;
wire _08456_ ;
wire _08457_ ;
wire _08458_ ;
wire _08459_ ;
wire _08460_ ;
wire _08461_ ;
wire _08462_ ;
wire _08463_ ;
wire _08464_ ;
wire _08465_ ;
wire _08466_ ;
wire _08467_ ;
wire _08468_ ;
wire _08469_ ;
wire _08470_ ;
wire _08471_ ;
wire _08472_ ;
wire _08473_ ;
wire _08474_ ;
wire _08475_ ;
wire _08476_ ;
wire _08477_ ;
wire _08478_ ;
wire _08479_ ;
wire _08480_ ;
wire _08481_ ;
wire _08482_ ;
wire _08483_ ;
wire _08484_ ;
wire _08485_ ;
wire _08486_ ;
wire _08487_ ;
wire _08488_ ;
wire _08489_ ;
wire _08490_ ;
wire _08491_ ;
wire _08492_ ;
wire _08493_ ;
wire _08494_ ;
wire _08495_ ;
wire _08496_ ;
wire _08497_ ;
wire _08498_ ;
wire _08499_ ;
wire _08500_ ;
wire _08501_ ;
wire _08502_ ;
wire _08503_ ;
wire _08504_ ;
wire _08505_ ;
wire _08506_ ;
wire _08507_ ;
wire _08508_ ;
wire _08509_ ;
wire _08510_ ;
wire _08511_ ;
wire _08512_ ;
wire _08513_ ;
wire _08514_ ;
wire _08515_ ;
wire _08516_ ;
wire _08517_ ;
wire _08518_ ;
wire _08519_ ;
wire _08520_ ;
wire _08521_ ;
wire _08522_ ;
wire _08523_ ;
wire _08524_ ;
wire _08525_ ;
wire _08526_ ;
wire _08527_ ;
wire _08528_ ;
wire _08529_ ;
wire _08530_ ;
wire _08531_ ;
wire _08532_ ;
wire _08533_ ;
wire _08534_ ;
wire _08535_ ;
wire _08536_ ;
wire _08537_ ;
wire _08538_ ;
wire _08539_ ;
wire _08540_ ;
wire _08541_ ;
wire _08542_ ;
wire _08543_ ;
wire _08544_ ;
wire _08545_ ;
wire _08546_ ;
wire _08547_ ;
wire _08548_ ;
wire _08549_ ;
wire _08550_ ;
wire _08551_ ;
wire _08552_ ;
wire _08553_ ;
wire _08554_ ;
wire _08555_ ;
wire _08556_ ;
wire _08557_ ;
wire _08558_ ;
wire _08559_ ;
wire _08560_ ;
wire _08561_ ;
wire _08562_ ;
wire _08563_ ;
wire _08564_ ;
wire _08565_ ;
wire _08566_ ;
wire _08567_ ;
wire _08568_ ;
wire _08569_ ;
wire _08570_ ;
wire _08571_ ;
wire _08572_ ;
wire _08573_ ;
wire _08574_ ;
wire _08575_ ;
wire _08576_ ;
wire _08577_ ;
wire _08578_ ;
wire _08579_ ;
wire _08580_ ;
wire _08581_ ;
wire _08582_ ;
wire _08583_ ;
wire _08584_ ;
wire _08585_ ;
wire _08586_ ;
wire _08587_ ;
wire _08588_ ;
wire _08589_ ;
wire _08590_ ;
wire _08591_ ;
wire _08592_ ;
wire _08593_ ;
wire _08594_ ;
wire _08595_ ;
wire _08596_ ;
wire _08597_ ;
wire _08598_ ;
wire _08599_ ;
wire _08600_ ;
wire _08601_ ;
wire _08602_ ;
wire _08603_ ;
wire _08604_ ;
wire _08605_ ;
wire _08606_ ;
wire _08607_ ;
wire _08608_ ;
wire _08609_ ;
wire _08610_ ;
wire _08611_ ;
wire _08612_ ;
wire _08613_ ;
wire _08614_ ;
wire _08615_ ;
wire _08616_ ;
wire _08617_ ;
wire _08618_ ;
wire _08619_ ;
wire _08620_ ;
wire _08621_ ;
wire _08622_ ;
wire _08623_ ;
wire _08624_ ;
wire _08625_ ;
wire _08626_ ;
wire _08627_ ;
wire _08628_ ;
wire _08629_ ;
wire _08630_ ;
wire _08631_ ;
wire _08632_ ;
wire _08633_ ;
wire _08634_ ;
wire _08635_ ;
wire _08636_ ;
wire _08637_ ;
wire _08638_ ;
wire _08639_ ;
wire _08640_ ;
wire _08641_ ;
wire _08642_ ;
wire _08643_ ;
wire _08644_ ;
wire _08645_ ;
wire _08646_ ;
wire _08647_ ;
wire _08648_ ;
wire _08649_ ;
wire _08650_ ;
wire _08651_ ;
wire _08652_ ;
wire _08653_ ;
wire _08654_ ;
wire _08655_ ;
wire _08656_ ;
wire _08657_ ;
wire _08658_ ;
wire _08659_ ;
wire _08660_ ;
wire _08661_ ;
wire _08662_ ;
wire _08663_ ;
wire _08664_ ;
wire _08665_ ;
wire _08666_ ;
wire _08667_ ;
wire _08668_ ;
wire _08669_ ;
wire _08670_ ;
wire _08671_ ;
wire _08672_ ;
wire _08673_ ;
wire _08674_ ;
wire _08675_ ;
wire _08676_ ;
wire _08677_ ;
wire _08678_ ;
wire _08679_ ;
wire _08680_ ;
wire _08681_ ;
wire _08682_ ;
wire _08683_ ;
wire _08684_ ;
wire _08685_ ;
wire _08686_ ;
wire _08687_ ;
wire _08688_ ;
wire _08689_ ;
wire _08690_ ;
wire _08691_ ;
wire _08692_ ;
wire _08693_ ;
wire _08694_ ;
wire _08695_ ;
wire _08696_ ;
wire _08697_ ;
wire _08698_ ;
wire _08699_ ;
wire _08700_ ;
wire _08701_ ;
wire _08702_ ;
wire _08703_ ;
wire _08704_ ;
wire _08705_ ;
wire _08706_ ;
wire _08707_ ;
wire _08708_ ;
wire _08709_ ;
wire _08710_ ;
wire _08711_ ;
wire _08712_ ;
wire _08713_ ;
wire _08714_ ;
wire _08715_ ;
wire _08716_ ;
wire _08717_ ;
wire _08718_ ;
wire _08719_ ;
wire _08720_ ;
wire _08721_ ;
wire _08722_ ;
wire _08723_ ;
wire _08724_ ;
wire _08725_ ;
wire _08726_ ;
wire _08727_ ;
wire _08728_ ;
wire _08729_ ;
wire _08730_ ;
wire _08731_ ;
wire _08732_ ;
wire _08733_ ;
wire _08734_ ;
wire _08735_ ;
wire _08736_ ;
wire _08737_ ;
wire _08738_ ;
wire _08739_ ;
wire _08740_ ;
wire _08741_ ;
wire _08742_ ;
wire _08743_ ;
wire _08744_ ;
wire _08745_ ;
wire _08746_ ;
wire _08747_ ;
wire _08748_ ;
wire _08749_ ;
wire _08750_ ;
wire _08751_ ;
wire _08752_ ;
wire _08753_ ;
wire _08754_ ;
wire _08755_ ;
wire _08756_ ;
wire _08757_ ;
wire _08758_ ;
wire _08759_ ;
wire _08760_ ;
wire _08761_ ;
wire _08762_ ;
wire _08763_ ;
wire _08764_ ;
wire _08765_ ;
wire _08766_ ;
wire _08767_ ;
wire _08768_ ;
wire _08769_ ;
wire _08770_ ;
wire _08771_ ;
wire _08772_ ;
wire _08773_ ;
wire _08774_ ;
wire _08775_ ;
wire _08776_ ;
wire _08777_ ;
wire _08778_ ;
wire _08779_ ;
wire _08780_ ;
wire _08781_ ;
wire _08782_ ;
wire _08783_ ;
wire _08784_ ;
wire _08785_ ;
wire _08786_ ;
wire _08787_ ;
wire _08788_ ;
wire _08789_ ;
wire _08790_ ;
wire _08791_ ;
wire _08792_ ;
wire _08793_ ;
wire _08794_ ;
wire _08795_ ;
wire _08796_ ;
wire _08797_ ;
wire _08798_ ;
wire _08799_ ;
wire _08800_ ;
wire _08801_ ;
wire _08802_ ;
wire _08803_ ;
wire _08804_ ;
wire _08805_ ;
wire _08806_ ;
wire _08807_ ;
wire _08808_ ;
wire _08809_ ;
wire _08810_ ;
wire _08811_ ;
wire _08812_ ;
wire _08813_ ;
wire _08814_ ;
wire _08815_ ;
wire _08816_ ;
wire _08817_ ;
wire _08818_ ;
wire _08819_ ;
wire _08820_ ;
wire _08821_ ;
wire _08822_ ;
wire _08823_ ;
wire _08824_ ;
wire _08825_ ;
wire _08826_ ;
wire _08827_ ;
wire _08828_ ;
wire _08829_ ;
wire _08830_ ;
wire _08831_ ;
wire _08832_ ;
wire _08833_ ;
wire _08834_ ;
wire _08835_ ;
wire _08836_ ;
wire _08837_ ;
wire _08838_ ;
wire _08839_ ;
wire _08840_ ;
wire _08841_ ;
wire _08842_ ;
wire _08843_ ;
wire _08844_ ;
wire _08845_ ;
wire _08846_ ;
wire _08847_ ;
wire _08848_ ;
wire _08849_ ;
wire _08850_ ;
wire _08851_ ;
wire _08852_ ;
wire _08853_ ;
wire _08854_ ;
wire _08855_ ;
wire _08856_ ;
wire _08857_ ;
wire _08858_ ;
wire _08859_ ;
wire _08860_ ;
wire _08861_ ;
wire _08862_ ;
wire _08863_ ;
wire _08864_ ;
wire _08865_ ;
wire _08866_ ;
wire _08867_ ;
wire _08868_ ;
wire _08869_ ;
wire _08870_ ;
wire _08871_ ;
wire _08872_ ;
wire _08873_ ;
wire _08874_ ;
wire _08875_ ;
wire _08876_ ;
wire _08877_ ;
wire _08878_ ;
wire _08879_ ;
wire _08880_ ;
wire _08881_ ;
wire _08882_ ;
wire _08883_ ;
wire _08884_ ;
wire _08885_ ;
wire _08886_ ;
wire _08887_ ;
wire _08888_ ;
wire _08889_ ;
wire _08890_ ;
wire _08891_ ;
wire _08892_ ;
wire _08893_ ;
wire _08894_ ;
wire _08895_ ;
wire _08896_ ;
wire _08897_ ;
wire _08898_ ;
wire _08899_ ;
wire _08900_ ;
wire _08901_ ;
wire _08902_ ;
wire _08903_ ;
wire _08904_ ;
wire _08905_ ;
wire _08906_ ;
wire _08907_ ;
wire _08908_ ;
wire _08909_ ;
wire _08910_ ;
wire _08911_ ;
wire _08912_ ;
wire _08913_ ;
wire _08914_ ;
wire _08915_ ;
wire _08916_ ;
wire _08917_ ;
wire _08918_ ;
wire _08919_ ;
wire _08920_ ;
wire _08921_ ;
wire _08922_ ;
wire _08923_ ;
wire _08924_ ;
wire _08925_ ;
wire _08926_ ;
wire _08927_ ;
wire _08928_ ;
wire _08929_ ;
wire _08930_ ;
wire _08931_ ;
wire _08932_ ;
wire _08933_ ;
wire _08934_ ;
wire _08935_ ;
wire _08936_ ;
wire _08937_ ;
wire _08938_ ;
wire _08939_ ;
wire _08940_ ;
wire _08941_ ;
wire _08942_ ;
wire _08943_ ;
wire EXU_valid_LSU ;
wire IDU_ready_IFU ;
wire IDU_valid_EXU ;
wire LS_WB_pc ;
wire LS_WB_wen_reg ;
wire check_assert ;
wire check_quest ;
wire exception_quest_IDU ;
wire excp_written ;
wire fc_disenable ;
wire io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ;
wire io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ;
wire io_master_wready_$_NOR__B_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ;
wire io_master_wready_$_NOR__B_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ;
wire loaduse_clear ;
wire \myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ;
wire \myclint.rvalid ;
wire \myclint.state_r_$_NOT__A_Y ;
wire \mycsreg.CSReg[0][0] ;
wire \mycsreg.CSReg[0][10] ;
wire \mycsreg.CSReg[0][11] ;
wire \mycsreg.CSReg[0][12] ;
wire \mycsreg.CSReg[0][13] ;
wire \mycsreg.CSReg[0][14] ;
wire \mycsreg.CSReg[0][15] ;
wire \mycsreg.CSReg[0][16] ;
wire \mycsreg.CSReg[0][17] ;
wire \mycsreg.CSReg[0][18] ;
wire \mycsreg.CSReg[0][19] ;
wire \mycsreg.CSReg[0][1] ;
wire \mycsreg.CSReg[0][20] ;
wire \mycsreg.CSReg[0][21] ;
wire \mycsreg.CSReg[0][22] ;
wire \mycsreg.CSReg[0][23] ;
wire \mycsreg.CSReg[0][24] ;
wire \mycsreg.CSReg[0][25] ;
wire \mycsreg.CSReg[0][26] ;
wire \mycsreg.CSReg[0][27] ;
wire \mycsreg.CSReg[0][28] ;
wire \mycsreg.CSReg[0][29] ;
wire \mycsreg.CSReg[0][2] ;
wire \mycsreg.CSReg[0][30] ;
wire \mycsreg.CSReg[0][31] ;
wire \mycsreg.CSReg[0][3] ;
wire \mycsreg.CSReg[0][4] ;
wire \mycsreg.CSReg[0][5] ;
wire \mycsreg.CSReg[0][6] ;
wire \mycsreg.CSReg[0][7] ;
wire \mycsreg.CSReg[0][8] ;
wire \mycsreg.CSReg[0][9] ;
wire \mycsreg.CSReg[3][0] ;
wire \mycsreg.CSReg[3][10] ;
wire \mycsreg.CSReg[3][11] ;
wire \mycsreg.CSReg[3][12] ;
wire \mycsreg.CSReg[3][13] ;
wire \mycsreg.CSReg[3][14] ;
wire \mycsreg.CSReg[3][15] ;
wire \mycsreg.CSReg[3][16] ;
wire \mycsreg.CSReg[3][17] ;
wire \mycsreg.CSReg[3][18] ;
wire \mycsreg.CSReg[3][19] ;
wire \mycsreg.CSReg[3][1] ;
wire \mycsreg.CSReg[3][20] ;
wire \mycsreg.CSReg[3][21] ;
wire \mycsreg.CSReg[3][22] ;
wire \mycsreg.CSReg[3][23] ;
wire \mycsreg.CSReg[3][24] ;
wire \mycsreg.CSReg[3][25] ;
wire \mycsreg.CSReg[3][26] ;
wire \mycsreg.CSReg[3][27] ;
wire \mycsreg.CSReg[3][28] ;
wire \mycsreg.CSReg[3][29] ;
wire \mycsreg.CSReg[3][2] ;
wire \mycsreg.CSReg[3][30] ;
wire \mycsreg.CSReg[3][31] ;
wire \mycsreg.CSReg[3][3] ;
wire \mycsreg.CSReg[3][4] ;
wire \mycsreg.CSReg[3][5] ;
wire \mycsreg.CSReg[3][6] ;
wire \mycsreg.CSReg[3][7] ;
wire \mycsreg.CSReg[3][8] ;
wire \mycsreg.CSReg[3][9] ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ;
wire \mycsreg.CSReg[3]_$_DFFE_PP__Q_D ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_OR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_10_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_11_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_12_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_13_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_14_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_15_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_16_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_17_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_18_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_19_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_1_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_20_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_21_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_22_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_23_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_24_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_25_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_26_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_27_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_28_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_29_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_2_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_30_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_31_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_3_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_4_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_5_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_6_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_7_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_8_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_9_D ;
wire \myec.mepc_tmp_$_DFFE_PP__Q_D ;
wire \myec.state_$_SDFFE_PP0P__Q_E ;
wire \myexu.check_quest_$_DFF_PP0__Q_D ;
wire \myexu.check_quest_$_DFF_PP0__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.dest_reg_$_DFFE_PP0P__Q_1_D ;
wire \myexu.dest_reg_$_DFFE_PP0P__Q_2_D ;
wire \myexu.dest_reg_$_DFFE_PP0P__Q_3_D ;
wire \myexu.dest_reg_$_DFFE_PP0P__Q_4_D ;
wire \myexu.dest_reg_$_DFFE_PP0P__Q_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_10_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_11_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_12_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_13_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_14_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_15_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_16_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_17_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_18_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_19_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_1_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_20_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_21_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_22_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_23_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_24_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_25_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_26_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_27_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_28_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_29_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_29_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_2_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_30_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_30_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_3_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_4_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_5_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_6_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_7_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_8_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_9_D ;
wire \myexu.pc_jump_$_DFFE_PP0P__Q_D ;
wire \myexu.pc_jump_$_DFFE_PP1P__Q_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_10_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_11_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_12_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_13_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_14_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_15_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_16_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_17_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_18_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_19_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_1_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_20_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_21_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_22_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_23_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_24_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_25_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_26_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_27_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_28_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_29_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_2_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_30_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_31_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_3_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_4_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_5_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_6_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_7_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_8_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_9_D ;
wire \myexu.pc_out_$_DFFE_PP0P__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_10_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_12_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_13_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_14_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_15_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_16_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_17_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_18_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_19_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_20_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_21_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_22_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_23_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_24_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_26_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_27_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_28_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_2_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_30_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ;
wire \myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__B_A_$_OR__A_Y_$_OR__A_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_4_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_6_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_7_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_8_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D ;
wire \myexu.result_reg_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ;
wire \myexu.result_reg_$_DFFE_PP__Q_D ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_1_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_3_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ;
wire \myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_B ;
wire \myexu.state_$_DFF_PP0__Q_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_1_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_2_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_3_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_4_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_5_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_6_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_7_D ;
wire \myexu.typ_out_$_DFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ;
wire \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y ;
wire \myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E ;
wire \myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ;
wire \myidu.stall_quest_fencei ;
wire \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ;
wire \myidu.stall_quest_loaduse ;
wire \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ;
wire \myidu.state_$_DFF_P__Q_1_D ;
wire \myidu.state_$_DFF_P__Q_2_D ;
wire \myidu.state_$_DFF_P__Q_D ;
wire \myidu.typ_$_SDFFE_PP0P__Q_E ;
wire \myifu.check_assert_$_DFFE_PP__Q_E ;
wire \myifu.check_assert_$_ORNOT__A_Y_$_MUX__A_S_$_OR__A_Y_$_ANDNOT__A_B_$_NOR__B_Y ;
wire \myifu.check_assert_$_ORNOT__A_Y_$_MUX__A_S_$_OR__A_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.myicache.data[0][0] ;
wire \myifu.myicache.data[0][10] ;
wire \myifu.myicache.data[0][11] ;
wire \myifu.myicache.data[0][12] ;
wire \myifu.myicache.data[0][13] ;
wire \myifu.myicache.data[0][14] ;
wire \myifu.myicache.data[0][15] ;
wire \myifu.myicache.data[0][16] ;
wire \myifu.myicache.data[0][17] ;
wire \myifu.myicache.data[0][18] ;
wire \myifu.myicache.data[0][19] ;
wire \myifu.myicache.data[0][1] ;
wire \myifu.myicache.data[0][20] ;
wire \myifu.myicache.data[0][21] ;
wire \myifu.myicache.data[0][22] ;
wire \myifu.myicache.data[0][23] ;
wire \myifu.myicache.data[0][24] ;
wire \myifu.myicache.data[0][25] ;
wire \myifu.myicache.data[0][26] ;
wire \myifu.myicache.data[0][27] ;
wire \myifu.myicache.data[0][28] ;
wire \myifu.myicache.data[0][29] ;
wire \myifu.myicache.data[0][2] ;
wire \myifu.myicache.data[0][30] ;
wire \myifu.myicache.data[0][31] ;
wire \myifu.myicache.data[0][3] ;
wire \myifu.myicache.data[0][4] ;
wire \myifu.myicache.data[0][5] ;
wire \myifu.myicache.data[0][6] ;
wire \myifu.myicache.data[0][7] ;
wire \myifu.myicache.data[0][8] ;
wire \myifu.myicache.data[0][9] ;
wire \myifu.myicache.data[1][0] ;
wire \myifu.myicache.data[1][10] ;
wire \myifu.myicache.data[1][11] ;
wire \myifu.myicache.data[1][12] ;
wire \myifu.myicache.data[1][13] ;
wire \myifu.myicache.data[1][14] ;
wire \myifu.myicache.data[1][15] ;
wire \myifu.myicache.data[1][16] ;
wire \myifu.myicache.data[1][17] ;
wire \myifu.myicache.data[1][18] ;
wire \myifu.myicache.data[1][19] ;
wire \myifu.myicache.data[1][1] ;
wire \myifu.myicache.data[1][20] ;
wire \myifu.myicache.data[1][21] ;
wire \myifu.myicache.data[1][22] ;
wire \myifu.myicache.data[1][23] ;
wire \myifu.myicache.data[1][24] ;
wire \myifu.myicache.data[1][25] ;
wire \myifu.myicache.data[1][26] ;
wire \myifu.myicache.data[1][27] ;
wire \myifu.myicache.data[1][28] ;
wire \myifu.myicache.data[1][29] ;
wire \myifu.myicache.data[1][2] ;
wire \myifu.myicache.data[1][30] ;
wire \myifu.myicache.data[1][31] ;
wire \myifu.myicache.data[1][3] ;
wire \myifu.myicache.data[1][4] ;
wire \myifu.myicache.data[1][5] ;
wire \myifu.myicache.data[1][6] ;
wire \myifu.myicache.data[1][7] ;
wire \myifu.myicache.data[1][8] ;
wire \myifu.myicache.data[1][9] ;
wire \myifu.myicache.data[2][0] ;
wire \myifu.myicache.data[2][10] ;
wire \myifu.myicache.data[2][11] ;
wire \myifu.myicache.data[2][12] ;
wire \myifu.myicache.data[2][13] ;
wire \myifu.myicache.data[2][14] ;
wire \myifu.myicache.data[2][15] ;
wire \myifu.myicache.data[2][16] ;
wire \myifu.myicache.data[2][17] ;
wire \myifu.myicache.data[2][18] ;
wire \myifu.myicache.data[2][19] ;
wire \myifu.myicache.data[2][1] ;
wire \myifu.myicache.data[2][20] ;
wire \myifu.myicache.data[2][21] ;
wire \myifu.myicache.data[2][22] ;
wire \myifu.myicache.data[2][23] ;
wire \myifu.myicache.data[2][24] ;
wire \myifu.myicache.data[2][25] ;
wire \myifu.myicache.data[2][26] ;
wire \myifu.myicache.data[2][27] ;
wire \myifu.myicache.data[2][28] ;
wire \myifu.myicache.data[2][29] ;
wire \myifu.myicache.data[2][2] ;
wire \myifu.myicache.data[2][30] ;
wire \myifu.myicache.data[2][31] ;
wire \myifu.myicache.data[2][3] ;
wire \myifu.myicache.data[2][4] ;
wire \myifu.myicache.data[2][5] ;
wire \myifu.myicache.data[2][6] ;
wire \myifu.myicache.data[2][7] ;
wire \myifu.myicache.data[2][8] ;
wire \myifu.myicache.data[2][9] ;
wire \myifu.myicache.data[3][0] ;
wire \myifu.myicache.data[3][10] ;
wire \myifu.myicache.data[3][11] ;
wire \myifu.myicache.data[3][12] ;
wire \myifu.myicache.data[3][13] ;
wire \myifu.myicache.data[3][14] ;
wire \myifu.myicache.data[3][15] ;
wire \myifu.myicache.data[3][16] ;
wire \myifu.myicache.data[3][17] ;
wire \myifu.myicache.data[3][18] ;
wire \myifu.myicache.data[3][19] ;
wire \myifu.myicache.data[3][1] ;
wire \myifu.myicache.data[3][20] ;
wire \myifu.myicache.data[3][21] ;
wire \myifu.myicache.data[3][22] ;
wire \myifu.myicache.data[3][23] ;
wire \myifu.myicache.data[3][24] ;
wire \myifu.myicache.data[3][25] ;
wire \myifu.myicache.data[3][26] ;
wire \myifu.myicache.data[3][27] ;
wire \myifu.myicache.data[3][28] ;
wire \myifu.myicache.data[3][29] ;
wire \myifu.myicache.data[3][2] ;
wire \myifu.myicache.data[3][30] ;
wire \myifu.myicache.data[3][31] ;
wire \myifu.myicache.data[3][3] ;
wire \myifu.myicache.data[3][4] ;
wire \myifu.myicache.data[3][5] ;
wire \myifu.myicache.data[3][6] ;
wire \myifu.myicache.data[3][7] ;
wire \myifu.myicache.data[3][8] ;
wire \myifu.myicache.data[3][9] ;
wire \myifu.myicache.data[4][0] ;
wire \myifu.myicache.data[4][10] ;
wire \myifu.myicache.data[4][11] ;
wire \myifu.myicache.data[4][12] ;
wire \myifu.myicache.data[4][13] ;
wire \myifu.myicache.data[4][14] ;
wire \myifu.myicache.data[4][15] ;
wire \myifu.myicache.data[4][16] ;
wire \myifu.myicache.data[4][17] ;
wire \myifu.myicache.data[4][18] ;
wire \myifu.myicache.data[4][19] ;
wire \myifu.myicache.data[4][1] ;
wire \myifu.myicache.data[4][20] ;
wire \myifu.myicache.data[4][21] ;
wire \myifu.myicache.data[4][22] ;
wire \myifu.myicache.data[4][23] ;
wire \myifu.myicache.data[4][24] ;
wire \myifu.myicache.data[4][25] ;
wire \myifu.myicache.data[4][26] ;
wire \myifu.myicache.data[4][27] ;
wire \myifu.myicache.data[4][28] ;
wire \myifu.myicache.data[4][29] ;
wire \myifu.myicache.data[4][2] ;
wire \myifu.myicache.data[4][30] ;
wire \myifu.myicache.data[4][31] ;
wire \myifu.myicache.data[4][3] ;
wire \myifu.myicache.data[4][4] ;
wire \myifu.myicache.data[4][5] ;
wire \myifu.myicache.data[4][6] ;
wire \myifu.myicache.data[4][7] ;
wire \myifu.myicache.data[4][8] ;
wire \myifu.myicache.data[4][9] ;
wire \myifu.myicache.data[5][0] ;
wire \myifu.myicache.data[5][10] ;
wire \myifu.myicache.data[5][11] ;
wire \myifu.myicache.data[5][12] ;
wire \myifu.myicache.data[5][13] ;
wire \myifu.myicache.data[5][14] ;
wire \myifu.myicache.data[5][15] ;
wire \myifu.myicache.data[5][16] ;
wire \myifu.myicache.data[5][17] ;
wire \myifu.myicache.data[5][18] ;
wire \myifu.myicache.data[5][19] ;
wire \myifu.myicache.data[5][1] ;
wire \myifu.myicache.data[5][20] ;
wire \myifu.myicache.data[5][21] ;
wire \myifu.myicache.data[5][22] ;
wire \myifu.myicache.data[5][23] ;
wire \myifu.myicache.data[5][24] ;
wire \myifu.myicache.data[5][25] ;
wire \myifu.myicache.data[5][26] ;
wire \myifu.myicache.data[5][27] ;
wire \myifu.myicache.data[5][28] ;
wire \myifu.myicache.data[5][29] ;
wire \myifu.myicache.data[5][2] ;
wire \myifu.myicache.data[5][30] ;
wire \myifu.myicache.data[5][31] ;
wire \myifu.myicache.data[5][3] ;
wire \myifu.myicache.data[5][4] ;
wire \myifu.myicache.data[5][5] ;
wire \myifu.myicache.data[5][6] ;
wire \myifu.myicache.data[5][7] ;
wire \myifu.myicache.data[5][8] ;
wire \myifu.myicache.data[5][9] ;
wire \myifu.myicache.data[6][0] ;
wire \myifu.myicache.data[6][10] ;
wire \myifu.myicache.data[6][11] ;
wire \myifu.myicache.data[6][12] ;
wire \myifu.myicache.data[6][13] ;
wire \myifu.myicache.data[6][14] ;
wire \myifu.myicache.data[6][15] ;
wire \myifu.myicache.data[6][16] ;
wire \myifu.myicache.data[6][17] ;
wire \myifu.myicache.data[6][18] ;
wire \myifu.myicache.data[6][19] ;
wire \myifu.myicache.data[6][1] ;
wire \myifu.myicache.data[6][20] ;
wire \myifu.myicache.data[6][21] ;
wire \myifu.myicache.data[6][22] ;
wire \myifu.myicache.data[6][23] ;
wire \myifu.myicache.data[6][24] ;
wire \myifu.myicache.data[6][25] ;
wire \myifu.myicache.data[6][26] ;
wire \myifu.myicache.data[6][27] ;
wire \myifu.myicache.data[6][28] ;
wire \myifu.myicache.data[6][29] ;
wire \myifu.myicache.data[6][2] ;
wire \myifu.myicache.data[6][30] ;
wire \myifu.myicache.data[6][31] ;
wire \myifu.myicache.data[6][3] ;
wire \myifu.myicache.data[6][4] ;
wire \myifu.myicache.data[6][5] ;
wire \myifu.myicache.data[6][6] ;
wire \myifu.myicache.data[6][7] ;
wire \myifu.myicache.data[6][8] ;
wire \myifu.myicache.data[6][9] ;
wire \myifu.myicache.data[7][0] ;
wire \myifu.myicache.data[7][10] ;
wire \myifu.myicache.data[7][11] ;
wire \myifu.myicache.data[7][12] ;
wire \myifu.myicache.data[7][13] ;
wire \myifu.myicache.data[7][14] ;
wire \myifu.myicache.data[7][15] ;
wire \myifu.myicache.data[7][16] ;
wire \myifu.myicache.data[7][17] ;
wire \myifu.myicache.data[7][18] ;
wire \myifu.myicache.data[7][19] ;
wire \myifu.myicache.data[7][1] ;
wire \myifu.myicache.data[7][20] ;
wire \myifu.myicache.data[7][21] ;
wire \myifu.myicache.data[7][22] ;
wire \myifu.myicache.data[7][23] ;
wire \myifu.myicache.data[7][24] ;
wire \myifu.myicache.data[7][25] ;
wire \myifu.myicache.data[7][26] ;
wire \myifu.myicache.data[7][27] ;
wire \myifu.myicache.data[7][28] ;
wire \myifu.myicache.data[7][29] ;
wire \myifu.myicache.data[7][2] ;
wire \myifu.myicache.data[7][30] ;
wire \myifu.myicache.data[7][31] ;
wire \myifu.myicache.data[7][3] ;
wire \myifu.myicache.data[7][4] ;
wire \myifu.myicache.data[7][5] ;
wire \myifu.myicache.data[7][6] ;
wire \myifu.myicache.data[7][7] ;
wire \myifu.myicache.data[7][8] ;
wire \myifu.myicache.data[7][9] ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ;
wire \myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ;
wire \myifu.myicache.tag[0][0] ;
wire \myifu.myicache.tag[0][10] ;
wire \myifu.myicache.tag[0][11] ;
wire \myifu.myicache.tag[0][12] ;
wire \myifu.myicache.tag[0][13] ;
wire \myifu.myicache.tag[0][14] ;
wire \myifu.myicache.tag[0][15] ;
wire \myifu.myicache.tag[0][16] ;
wire \myifu.myicache.tag[0][17] ;
wire \myifu.myicache.tag[0][18] ;
wire \myifu.myicache.tag[0][19] ;
wire \myifu.myicache.tag[0][1] ;
wire \myifu.myicache.tag[0][20] ;
wire \myifu.myicache.tag[0][21] ;
wire \myifu.myicache.tag[0][22] ;
wire \myifu.myicache.tag[0][23] ;
wire \myifu.myicache.tag[0][24] ;
wire \myifu.myicache.tag[0][25] ;
wire \myifu.myicache.tag[0][26] ;
wire \myifu.myicache.tag[0][2] ;
wire \myifu.myicache.tag[0][3] ;
wire \myifu.myicache.tag[0][4] ;
wire \myifu.myicache.tag[0][5] ;
wire \myifu.myicache.tag[0][6] ;
wire \myifu.myicache.tag[0][7] ;
wire \myifu.myicache.tag[0][8] ;
wire \myifu.myicache.tag[0][9] ;
wire \myifu.myicache.tag[1][0] ;
wire \myifu.myicache.tag[1][10] ;
wire \myifu.myicache.tag[1][11] ;
wire \myifu.myicache.tag[1][12] ;
wire \myifu.myicache.tag[1][13] ;
wire \myifu.myicache.tag[1][14] ;
wire \myifu.myicache.tag[1][15] ;
wire \myifu.myicache.tag[1][16] ;
wire \myifu.myicache.tag[1][17] ;
wire \myifu.myicache.tag[1][18] ;
wire \myifu.myicache.tag[1][19] ;
wire \myifu.myicache.tag[1][1] ;
wire \myifu.myicache.tag[1][20] ;
wire \myifu.myicache.tag[1][21] ;
wire \myifu.myicache.tag[1][22] ;
wire \myifu.myicache.tag[1][23] ;
wire \myifu.myicache.tag[1][24] ;
wire \myifu.myicache.tag[1][25] ;
wire \myifu.myicache.tag[1][26] ;
wire \myifu.myicache.tag[1][2] ;
wire \myifu.myicache.tag[1][3] ;
wire \myifu.myicache.tag[1][4] ;
wire \myifu.myicache.tag[1][5] ;
wire \myifu.myicache.tag[1][6] ;
wire \myifu.myicache.tag[1][7] ;
wire \myifu.myicache.tag[1][8] ;
wire \myifu.myicache.tag[1][9] ;
wire \myifu.myicache.tag[2][0] ;
wire \myifu.myicache.tag[2][10] ;
wire \myifu.myicache.tag[2][11] ;
wire \myifu.myicache.tag[2][12] ;
wire \myifu.myicache.tag[2][13] ;
wire \myifu.myicache.tag[2][14] ;
wire \myifu.myicache.tag[2][15] ;
wire \myifu.myicache.tag[2][16] ;
wire \myifu.myicache.tag[2][17] ;
wire \myifu.myicache.tag[2][18] ;
wire \myifu.myicache.tag[2][19] ;
wire \myifu.myicache.tag[2][1] ;
wire \myifu.myicache.tag[2][20] ;
wire \myifu.myicache.tag[2][21] ;
wire \myifu.myicache.tag[2][22] ;
wire \myifu.myicache.tag[2][23] ;
wire \myifu.myicache.tag[2][24] ;
wire \myifu.myicache.tag[2][25] ;
wire \myifu.myicache.tag[2][26] ;
wire \myifu.myicache.tag[2][2] ;
wire \myifu.myicache.tag[2][3] ;
wire \myifu.myicache.tag[2][4] ;
wire \myifu.myicache.tag[2][5] ;
wire \myifu.myicache.tag[2][6] ;
wire \myifu.myicache.tag[2][7] ;
wire \myifu.myicache.tag[2][8] ;
wire \myifu.myicache.tag[2][9] ;
wire \myifu.myicache.tag[3][0] ;
wire \myifu.myicache.tag[3][10] ;
wire \myifu.myicache.tag[3][11] ;
wire \myifu.myicache.tag[3][12] ;
wire \myifu.myicache.tag[3][13] ;
wire \myifu.myicache.tag[3][14] ;
wire \myifu.myicache.tag[3][15] ;
wire \myifu.myicache.tag[3][16] ;
wire \myifu.myicache.tag[3][17] ;
wire \myifu.myicache.tag[3][18] ;
wire \myifu.myicache.tag[3][19] ;
wire \myifu.myicache.tag[3][1] ;
wire \myifu.myicache.tag[3][20] ;
wire \myifu.myicache.tag[3][21] ;
wire \myifu.myicache.tag[3][22] ;
wire \myifu.myicache.tag[3][23] ;
wire \myifu.myicache.tag[3][24] ;
wire \myifu.myicache.tag[3][25] ;
wire \myifu.myicache.tag[3][26] ;
wire \myifu.myicache.tag[3][2] ;
wire \myifu.myicache.tag[3][3] ;
wire \myifu.myicache.tag[3][4] ;
wire \myifu.myicache.tag[3][5] ;
wire \myifu.myicache.tag[3][6] ;
wire \myifu.myicache.tag[3][7] ;
wire \myifu.myicache.tag[3][8] ;
wire \myifu.myicache.tag[3][9] ;
wire \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ;
wire \myifu.myicache.valid[3]_$_DFFE_PP__Q_E ;
wire \myifu.myicache.valid_data_in ;
wire \myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ;
wire \myifu.pc_$_SDFFE_PP0P__Q_E ;
wire \myifu.pc_$_SDFFE_PP1P__Q_E ;
wire \myifu.state_$_DFF_P__Q_1_D ;
wire \myifu.state_$_DFF_P__Q_2_D ;
wire \myifu.state_$_DFF_P__Q_D ;
wire \myifu.tmp_offset_$_SDFFE_PP0P__Q_E ;
wire \myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ;
wire \myifu.to_reset ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ;
wire \myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_B_$_MUX__Y_A_$_NOR__B_Y ;
wire \myifu.wen_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ;
wire \myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ;
wire \myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.pc_out_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ;
wire \mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ;
wire \mylsu.state_$_DFF_P__Q_1_D ;
wire \mylsu.state_$_DFF_P__Q_2_D ;
wire \mylsu.state_$_DFF_P__Q_3_D ;
wire \mylsu.state_$_DFF_P__Q_4_D ;
wire \mylsu.state_$_DFF_P__Q_D ;
wire \mylsu.typ_tmp_$_NOT__A_Y ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_csreg_$_DFFE_PP__Q_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_10_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_11_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_12_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_13_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_14_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_15_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_16_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_17_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_18_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_19_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_1_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_20_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_21_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_22_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_23_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_24_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_25_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_26_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_27_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_28_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_29_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_2_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_30_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_31_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_3_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_4_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_5_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_6_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_7_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_8_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_9_D ;
wire \mylsu.wdata_reg_$_DFFE_PP__Q_D ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ;
wire \mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ;
wire \myminixbar.state_$_DFF_P__Q_1_D ;
wire \myminixbar.state_$_DFF_P__Q_D ;
wire \myreg.Reg[0][0] ;
wire \myreg.Reg[0][10] ;
wire \myreg.Reg[0][11] ;
wire \myreg.Reg[0][12] ;
wire \myreg.Reg[0][13] ;
wire \myreg.Reg[0][14] ;
wire \myreg.Reg[0][15] ;
wire \myreg.Reg[0][16] ;
wire \myreg.Reg[0][17] ;
wire \myreg.Reg[0][18] ;
wire \myreg.Reg[0][19] ;
wire \myreg.Reg[0][1] ;
wire \myreg.Reg[0][20] ;
wire \myreg.Reg[0][21] ;
wire \myreg.Reg[0][22] ;
wire \myreg.Reg[0][23] ;
wire \myreg.Reg[0][24] ;
wire \myreg.Reg[0][25] ;
wire \myreg.Reg[0][26] ;
wire \myreg.Reg[0][27] ;
wire \myreg.Reg[0][28] ;
wire \myreg.Reg[0][29] ;
wire \myreg.Reg[0][2] ;
wire \myreg.Reg[0][30] ;
wire \myreg.Reg[0][31] ;
wire \myreg.Reg[0][3] ;
wire \myreg.Reg[0][4] ;
wire \myreg.Reg[0][5] ;
wire \myreg.Reg[0][6] ;
wire \myreg.Reg[0][7] ;
wire \myreg.Reg[0][8] ;
wire \myreg.Reg[0][9] ;
wire \myreg.Reg[10][0] ;
wire \myreg.Reg[10][10] ;
wire \myreg.Reg[10][11] ;
wire \myreg.Reg[10][12] ;
wire \myreg.Reg[10][13] ;
wire \myreg.Reg[10][14] ;
wire \myreg.Reg[10][15] ;
wire \myreg.Reg[10][16] ;
wire \myreg.Reg[10][17] ;
wire \myreg.Reg[10][18] ;
wire \myreg.Reg[10][19] ;
wire \myreg.Reg[10][1] ;
wire \myreg.Reg[10][20] ;
wire \myreg.Reg[10][21] ;
wire \myreg.Reg[10][22] ;
wire \myreg.Reg[10][23] ;
wire \myreg.Reg[10][24] ;
wire \myreg.Reg[10][25] ;
wire \myreg.Reg[10][26] ;
wire \myreg.Reg[10][27] ;
wire \myreg.Reg[10][28] ;
wire \myreg.Reg[10][29] ;
wire \myreg.Reg[10][2] ;
wire \myreg.Reg[10][30] ;
wire \myreg.Reg[10][31] ;
wire \myreg.Reg[10][3] ;
wire \myreg.Reg[10][4] ;
wire \myreg.Reg[10][5] ;
wire \myreg.Reg[10][6] ;
wire \myreg.Reg[10][7] ;
wire \myreg.Reg[10][8] ;
wire \myreg.Reg[10][9] ;
wire \myreg.Reg[11][0] ;
wire \myreg.Reg[11][10] ;
wire \myreg.Reg[11][11] ;
wire \myreg.Reg[11][12] ;
wire \myreg.Reg[11][13] ;
wire \myreg.Reg[11][14] ;
wire \myreg.Reg[11][15] ;
wire \myreg.Reg[11][16] ;
wire \myreg.Reg[11][17] ;
wire \myreg.Reg[11][18] ;
wire \myreg.Reg[11][19] ;
wire \myreg.Reg[11][1] ;
wire \myreg.Reg[11][20] ;
wire \myreg.Reg[11][21] ;
wire \myreg.Reg[11][22] ;
wire \myreg.Reg[11][23] ;
wire \myreg.Reg[11][24] ;
wire \myreg.Reg[11][25] ;
wire \myreg.Reg[11][26] ;
wire \myreg.Reg[11][27] ;
wire \myreg.Reg[11][28] ;
wire \myreg.Reg[11][29] ;
wire \myreg.Reg[11][2] ;
wire \myreg.Reg[11][30] ;
wire \myreg.Reg[11][31] ;
wire \myreg.Reg[11][3] ;
wire \myreg.Reg[11][4] ;
wire \myreg.Reg[11][5] ;
wire \myreg.Reg[11][6] ;
wire \myreg.Reg[11][7] ;
wire \myreg.Reg[11][8] ;
wire \myreg.Reg[11][9] ;
wire \myreg.Reg[12][0] ;
wire \myreg.Reg[12][10] ;
wire \myreg.Reg[12][11] ;
wire \myreg.Reg[12][12] ;
wire \myreg.Reg[12][13] ;
wire \myreg.Reg[12][14] ;
wire \myreg.Reg[12][15] ;
wire \myreg.Reg[12][16] ;
wire \myreg.Reg[12][17] ;
wire \myreg.Reg[12][18] ;
wire \myreg.Reg[12][19] ;
wire \myreg.Reg[12][1] ;
wire \myreg.Reg[12][20] ;
wire \myreg.Reg[12][21] ;
wire \myreg.Reg[12][22] ;
wire \myreg.Reg[12][23] ;
wire \myreg.Reg[12][24] ;
wire \myreg.Reg[12][25] ;
wire \myreg.Reg[12][26] ;
wire \myreg.Reg[12][27] ;
wire \myreg.Reg[12][28] ;
wire \myreg.Reg[12][29] ;
wire \myreg.Reg[12][2] ;
wire \myreg.Reg[12][30] ;
wire \myreg.Reg[12][31] ;
wire \myreg.Reg[12][3] ;
wire \myreg.Reg[12][4] ;
wire \myreg.Reg[12][5] ;
wire \myreg.Reg[12][6] ;
wire \myreg.Reg[12][7] ;
wire \myreg.Reg[12][8] ;
wire \myreg.Reg[12][9] ;
wire \myreg.Reg[13][0] ;
wire \myreg.Reg[13][10] ;
wire \myreg.Reg[13][11] ;
wire \myreg.Reg[13][12] ;
wire \myreg.Reg[13][13] ;
wire \myreg.Reg[13][14] ;
wire \myreg.Reg[13][15] ;
wire \myreg.Reg[13][16] ;
wire \myreg.Reg[13][17] ;
wire \myreg.Reg[13][18] ;
wire \myreg.Reg[13][19] ;
wire \myreg.Reg[13][1] ;
wire \myreg.Reg[13][20] ;
wire \myreg.Reg[13][21] ;
wire \myreg.Reg[13][22] ;
wire \myreg.Reg[13][23] ;
wire \myreg.Reg[13][24] ;
wire \myreg.Reg[13][25] ;
wire \myreg.Reg[13][26] ;
wire \myreg.Reg[13][27] ;
wire \myreg.Reg[13][28] ;
wire \myreg.Reg[13][29] ;
wire \myreg.Reg[13][2] ;
wire \myreg.Reg[13][30] ;
wire \myreg.Reg[13][31] ;
wire \myreg.Reg[13][3] ;
wire \myreg.Reg[13][4] ;
wire \myreg.Reg[13][5] ;
wire \myreg.Reg[13][6] ;
wire \myreg.Reg[13][7] ;
wire \myreg.Reg[13][8] ;
wire \myreg.Reg[13][9] ;
wire \myreg.Reg[14][0] ;
wire \myreg.Reg[14][10] ;
wire \myreg.Reg[14][11] ;
wire \myreg.Reg[14][12] ;
wire \myreg.Reg[14][13] ;
wire \myreg.Reg[14][14] ;
wire \myreg.Reg[14][15] ;
wire \myreg.Reg[14][16] ;
wire \myreg.Reg[14][17] ;
wire \myreg.Reg[14][18] ;
wire \myreg.Reg[14][19] ;
wire \myreg.Reg[14][1] ;
wire \myreg.Reg[14][20] ;
wire \myreg.Reg[14][21] ;
wire \myreg.Reg[14][22] ;
wire \myreg.Reg[14][23] ;
wire \myreg.Reg[14][24] ;
wire \myreg.Reg[14][25] ;
wire \myreg.Reg[14][26] ;
wire \myreg.Reg[14][27] ;
wire \myreg.Reg[14][28] ;
wire \myreg.Reg[14][29] ;
wire \myreg.Reg[14][2] ;
wire \myreg.Reg[14][30] ;
wire \myreg.Reg[14][31] ;
wire \myreg.Reg[14][3] ;
wire \myreg.Reg[14][4] ;
wire \myreg.Reg[14][5] ;
wire \myreg.Reg[14][6] ;
wire \myreg.Reg[14][7] ;
wire \myreg.Reg[14][8] ;
wire \myreg.Reg[14][9] ;
wire \myreg.Reg[15][0] ;
wire \myreg.Reg[15][10] ;
wire \myreg.Reg[15][11] ;
wire \myreg.Reg[15][12] ;
wire \myreg.Reg[15][13] ;
wire \myreg.Reg[15][14] ;
wire \myreg.Reg[15][15] ;
wire \myreg.Reg[15][16] ;
wire \myreg.Reg[15][17] ;
wire \myreg.Reg[15][18] ;
wire \myreg.Reg[15][19] ;
wire \myreg.Reg[15][1] ;
wire \myreg.Reg[15][20] ;
wire \myreg.Reg[15][21] ;
wire \myreg.Reg[15][22] ;
wire \myreg.Reg[15][23] ;
wire \myreg.Reg[15][24] ;
wire \myreg.Reg[15][25] ;
wire \myreg.Reg[15][26] ;
wire \myreg.Reg[15][27] ;
wire \myreg.Reg[15][28] ;
wire \myreg.Reg[15][29] ;
wire \myreg.Reg[15][2] ;
wire \myreg.Reg[15][30] ;
wire \myreg.Reg[15][31] ;
wire \myreg.Reg[15][3] ;
wire \myreg.Reg[15][4] ;
wire \myreg.Reg[15][5] ;
wire \myreg.Reg[15][6] ;
wire \myreg.Reg[15][7] ;
wire \myreg.Reg[15][8] ;
wire \myreg.Reg[15][9] ;
wire \myreg.Reg[1][0] ;
wire \myreg.Reg[1][10] ;
wire \myreg.Reg[1][11] ;
wire \myreg.Reg[1][12] ;
wire \myreg.Reg[1][13] ;
wire \myreg.Reg[1][14] ;
wire \myreg.Reg[1][15] ;
wire \myreg.Reg[1][16] ;
wire \myreg.Reg[1][17] ;
wire \myreg.Reg[1][18] ;
wire \myreg.Reg[1][19] ;
wire \myreg.Reg[1][1] ;
wire \myreg.Reg[1][20] ;
wire \myreg.Reg[1][21] ;
wire \myreg.Reg[1][22] ;
wire \myreg.Reg[1][23] ;
wire \myreg.Reg[1][24] ;
wire \myreg.Reg[1][25] ;
wire \myreg.Reg[1][26] ;
wire \myreg.Reg[1][27] ;
wire \myreg.Reg[1][28] ;
wire \myreg.Reg[1][29] ;
wire \myreg.Reg[1][2] ;
wire \myreg.Reg[1][30] ;
wire \myreg.Reg[1][31] ;
wire \myreg.Reg[1][3] ;
wire \myreg.Reg[1][4] ;
wire \myreg.Reg[1][5] ;
wire \myreg.Reg[1][6] ;
wire \myreg.Reg[1][7] ;
wire \myreg.Reg[1][8] ;
wire \myreg.Reg[1][9] ;
wire \myreg.Reg[2][0] ;
wire \myreg.Reg[2][10] ;
wire \myreg.Reg[2][11] ;
wire \myreg.Reg[2][12] ;
wire \myreg.Reg[2][13] ;
wire \myreg.Reg[2][14] ;
wire \myreg.Reg[2][15] ;
wire \myreg.Reg[2][16] ;
wire \myreg.Reg[2][17] ;
wire \myreg.Reg[2][18] ;
wire \myreg.Reg[2][19] ;
wire \myreg.Reg[2][1] ;
wire \myreg.Reg[2][20] ;
wire \myreg.Reg[2][21] ;
wire \myreg.Reg[2][22] ;
wire \myreg.Reg[2][23] ;
wire \myreg.Reg[2][24] ;
wire \myreg.Reg[2][25] ;
wire \myreg.Reg[2][26] ;
wire \myreg.Reg[2][27] ;
wire \myreg.Reg[2][28] ;
wire \myreg.Reg[2][29] ;
wire \myreg.Reg[2][2] ;
wire \myreg.Reg[2][30] ;
wire \myreg.Reg[2][31] ;
wire \myreg.Reg[2][3] ;
wire \myreg.Reg[2][4] ;
wire \myreg.Reg[2][5] ;
wire \myreg.Reg[2][6] ;
wire \myreg.Reg[2][7] ;
wire \myreg.Reg[2][8] ;
wire \myreg.Reg[2][9] ;
wire \myreg.Reg[3][0] ;
wire \myreg.Reg[3][10] ;
wire \myreg.Reg[3][11] ;
wire \myreg.Reg[3][12] ;
wire \myreg.Reg[3][13] ;
wire \myreg.Reg[3][14] ;
wire \myreg.Reg[3][15] ;
wire \myreg.Reg[3][16] ;
wire \myreg.Reg[3][17] ;
wire \myreg.Reg[3][18] ;
wire \myreg.Reg[3][19] ;
wire \myreg.Reg[3][1] ;
wire \myreg.Reg[3][20] ;
wire \myreg.Reg[3][21] ;
wire \myreg.Reg[3][22] ;
wire \myreg.Reg[3][23] ;
wire \myreg.Reg[3][24] ;
wire \myreg.Reg[3][25] ;
wire \myreg.Reg[3][26] ;
wire \myreg.Reg[3][27] ;
wire \myreg.Reg[3][28] ;
wire \myreg.Reg[3][29] ;
wire \myreg.Reg[3][2] ;
wire \myreg.Reg[3][30] ;
wire \myreg.Reg[3][31] ;
wire \myreg.Reg[3][3] ;
wire \myreg.Reg[3][4] ;
wire \myreg.Reg[3][5] ;
wire \myreg.Reg[3][6] ;
wire \myreg.Reg[3][7] ;
wire \myreg.Reg[3][8] ;
wire \myreg.Reg[3][9] ;
wire \myreg.Reg[4][0] ;
wire \myreg.Reg[4][10] ;
wire \myreg.Reg[4][11] ;
wire \myreg.Reg[4][12] ;
wire \myreg.Reg[4][13] ;
wire \myreg.Reg[4][14] ;
wire \myreg.Reg[4][15] ;
wire \myreg.Reg[4][16] ;
wire \myreg.Reg[4][17] ;
wire \myreg.Reg[4][18] ;
wire \myreg.Reg[4][19] ;
wire \myreg.Reg[4][1] ;
wire \myreg.Reg[4][20] ;
wire \myreg.Reg[4][21] ;
wire \myreg.Reg[4][22] ;
wire \myreg.Reg[4][23] ;
wire \myreg.Reg[4][24] ;
wire \myreg.Reg[4][25] ;
wire \myreg.Reg[4][26] ;
wire \myreg.Reg[4][27] ;
wire \myreg.Reg[4][28] ;
wire \myreg.Reg[4][29] ;
wire \myreg.Reg[4][2] ;
wire \myreg.Reg[4][30] ;
wire \myreg.Reg[4][31] ;
wire \myreg.Reg[4][3] ;
wire \myreg.Reg[4][4] ;
wire \myreg.Reg[4][5] ;
wire \myreg.Reg[4][6] ;
wire \myreg.Reg[4][7] ;
wire \myreg.Reg[4][8] ;
wire \myreg.Reg[4][9] ;
wire \myreg.Reg[5][0] ;
wire \myreg.Reg[5][10] ;
wire \myreg.Reg[5][11] ;
wire \myreg.Reg[5][12] ;
wire \myreg.Reg[5][13] ;
wire \myreg.Reg[5][14] ;
wire \myreg.Reg[5][15] ;
wire \myreg.Reg[5][16] ;
wire \myreg.Reg[5][17] ;
wire \myreg.Reg[5][18] ;
wire \myreg.Reg[5][19] ;
wire \myreg.Reg[5][1] ;
wire \myreg.Reg[5][20] ;
wire \myreg.Reg[5][21] ;
wire \myreg.Reg[5][22] ;
wire \myreg.Reg[5][23] ;
wire \myreg.Reg[5][24] ;
wire \myreg.Reg[5][25] ;
wire \myreg.Reg[5][26] ;
wire \myreg.Reg[5][27] ;
wire \myreg.Reg[5][28] ;
wire \myreg.Reg[5][29] ;
wire \myreg.Reg[5][2] ;
wire \myreg.Reg[5][30] ;
wire \myreg.Reg[5][31] ;
wire \myreg.Reg[5][3] ;
wire \myreg.Reg[5][4] ;
wire \myreg.Reg[5][5] ;
wire \myreg.Reg[5][6] ;
wire \myreg.Reg[5][7] ;
wire \myreg.Reg[5][8] ;
wire \myreg.Reg[5][9] ;
wire \myreg.Reg[6][0] ;
wire \myreg.Reg[6][10] ;
wire \myreg.Reg[6][11] ;
wire \myreg.Reg[6][12] ;
wire \myreg.Reg[6][13] ;
wire \myreg.Reg[6][14] ;
wire \myreg.Reg[6][15] ;
wire \myreg.Reg[6][16] ;
wire \myreg.Reg[6][17] ;
wire \myreg.Reg[6][18] ;
wire \myreg.Reg[6][19] ;
wire \myreg.Reg[6][1] ;
wire \myreg.Reg[6][20] ;
wire \myreg.Reg[6][21] ;
wire \myreg.Reg[6][22] ;
wire \myreg.Reg[6][23] ;
wire \myreg.Reg[6][24] ;
wire \myreg.Reg[6][25] ;
wire \myreg.Reg[6][26] ;
wire \myreg.Reg[6][27] ;
wire \myreg.Reg[6][28] ;
wire \myreg.Reg[6][29] ;
wire \myreg.Reg[6][2] ;
wire \myreg.Reg[6][30] ;
wire \myreg.Reg[6][31] ;
wire \myreg.Reg[6][3] ;
wire \myreg.Reg[6][4] ;
wire \myreg.Reg[6][5] ;
wire \myreg.Reg[6][6] ;
wire \myreg.Reg[6][7] ;
wire \myreg.Reg[6][8] ;
wire \myreg.Reg[6][9] ;
wire \myreg.Reg[7][0] ;
wire \myreg.Reg[7][10] ;
wire \myreg.Reg[7][11] ;
wire \myreg.Reg[7][12] ;
wire \myreg.Reg[7][13] ;
wire \myreg.Reg[7][14] ;
wire \myreg.Reg[7][15] ;
wire \myreg.Reg[7][16] ;
wire \myreg.Reg[7][17] ;
wire \myreg.Reg[7][18] ;
wire \myreg.Reg[7][19] ;
wire \myreg.Reg[7][1] ;
wire \myreg.Reg[7][20] ;
wire \myreg.Reg[7][21] ;
wire \myreg.Reg[7][22] ;
wire \myreg.Reg[7][23] ;
wire \myreg.Reg[7][24] ;
wire \myreg.Reg[7][25] ;
wire \myreg.Reg[7][26] ;
wire \myreg.Reg[7][27] ;
wire \myreg.Reg[7][28] ;
wire \myreg.Reg[7][29] ;
wire \myreg.Reg[7][2] ;
wire \myreg.Reg[7][30] ;
wire \myreg.Reg[7][31] ;
wire \myreg.Reg[7][3] ;
wire \myreg.Reg[7][4] ;
wire \myreg.Reg[7][5] ;
wire \myreg.Reg[7][6] ;
wire \myreg.Reg[7][7] ;
wire \myreg.Reg[7][8] ;
wire \myreg.Reg[7][9] ;
wire \myreg.Reg[8][0] ;
wire \myreg.Reg[8][10] ;
wire \myreg.Reg[8][11] ;
wire \myreg.Reg[8][12] ;
wire \myreg.Reg[8][13] ;
wire \myreg.Reg[8][14] ;
wire \myreg.Reg[8][15] ;
wire \myreg.Reg[8][16] ;
wire \myreg.Reg[8][17] ;
wire \myreg.Reg[8][18] ;
wire \myreg.Reg[8][19] ;
wire \myreg.Reg[8][1] ;
wire \myreg.Reg[8][20] ;
wire \myreg.Reg[8][21] ;
wire \myreg.Reg[8][22] ;
wire \myreg.Reg[8][23] ;
wire \myreg.Reg[8][24] ;
wire \myreg.Reg[8][25] ;
wire \myreg.Reg[8][26] ;
wire \myreg.Reg[8][27] ;
wire \myreg.Reg[8][28] ;
wire \myreg.Reg[8][29] ;
wire \myreg.Reg[8][2] ;
wire \myreg.Reg[8][30] ;
wire \myreg.Reg[8][31] ;
wire \myreg.Reg[8][3] ;
wire \myreg.Reg[8][4] ;
wire \myreg.Reg[8][5] ;
wire \myreg.Reg[8][6] ;
wire \myreg.Reg[8][7] ;
wire \myreg.Reg[8][8] ;
wire \myreg.Reg[8][9] ;
wire \myreg.Reg[9][0] ;
wire \myreg.Reg[9][10] ;
wire \myreg.Reg[9][11] ;
wire \myreg.Reg[9][12] ;
wire \myreg.Reg[9][13] ;
wire \myreg.Reg[9][14] ;
wire \myreg.Reg[9][15] ;
wire \myreg.Reg[9][16] ;
wire \myreg.Reg[9][17] ;
wire \myreg.Reg[9][18] ;
wire \myreg.Reg[9][19] ;
wire \myreg.Reg[9][1] ;
wire \myreg.Reg[9][20] ;
wire \myreg.Reg[9][21] ;
wire \myreg.Reg[9][22] ;
wire \myreg.Reg[9][23] ;
wire \myreg.Reg[9][24] ;
wire \myreg.Reg[9][25] ;
wire \myreg.Reg[9][26] ;
wire \myreg.Reg[9][27] ;
wire \myreg.Reg[9][28] ;
wire \myreg.Reg[9][29] ;
wire \myreg.Reg[9][2] ;
wire \myreg.Reg[9][30] ;
wire \myreg.Reg[9][31] ;
wire \myreg.Reg[9][3] ;
wire \myreg.Reg[9][4] ;
wire \myreg.Reg[9][5] ;
wire \myreg.Reg[9][6] ;
wire \myreg.Reg[9][7] ;
wire \myreg.Reg[9][8] ;
wire \myreg.Reg[9][9] ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_10_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_11_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_12_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_13_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_14_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_15_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_16_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_17_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_18_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_19_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_1_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_20_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_21_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_22_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_23_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_24_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_25_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_26_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_27_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_28_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_29_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_2_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_30_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_31_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_3_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_4_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_5_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_6_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_7_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_8_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_9_D ;
wire \myreg.Reg[9]_$_DFFE_PP__Q_D ;
wire \mysc.state_$_DFF_P__Q_1_D ;
wire \mysc.state_$_DFF_P__Q_2_D ;
wire \mysc.state_$_DFF_P__Q_D ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire fanout_net_21 ;
wire fanout_net_22 ;
wire fanout_net_23 ;
wire fanout_net_24 ;
wire fanout_net_25 ;
wire fanout_net_26 ;
wire fanout_net_27 ;
wire fanout_net_28 ;
wire fanout_net_29 ;
wire fanout_net_30 ;
wire fanout_net_31 ;
wire fanout_net_32 ;
wire fanout_net_33 ;
wire fanout_net_34 ;
wire fanout_net_35 ;
wire fanout_net_36 ;
wire fanout_net_37 ;
wire fanout_net_38 ;
wire fanout_net_39 ;
wire fanout_net_40 ;
wire fanout_net_41 ;
wire fanout_net_42 ;
wire fanout_net_43 ;
wire fanout_net_44 ;
wire fanout_net_45 ;
wire fanout_net_46 ;
wire fanout_net_47 ;
wire fanout_net_48 ;
wire fanout_net_49 ;
wire [31:0] io_master_awaddr ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [1:0] io_master_awburst ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [1:0] io_master_bresp ;
wire [3:0] io_master_bid ;
wire [31:0] io_master_araddr ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [1:0] io_master_arburst ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [31:0] io_slave_awaddr ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [1:0] io_slave_awburst ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] io_slave_bresp ;
wire [3:0] io_slave_bid ;
wire [31:0] io_slave_araddr ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [1:0] io_slave_arburst ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [31:0] EX_LS_dest_csreg_mem ;
wire [4:0] EX_LS_dest_reg ;
wire [2:0] EX_LS_flag ;
wire [31:0] EX_LS_pc ;
wire [31:0] EX_LS_result_csreg_mem ;
wire [31:0] EX_LS_result_reg ;
wire [4:0] EX_LS_typ ;
wire [11:0] ID_EX_csr ;
wire [31:0] ID_EX_imm ;
wire [31:0] ID_EX_pc ;
wire [4:0] ID_EX_rd ;
wire [4:0] ID_EX_rs1 ;
wire [4:0] ID_EX_rs2 ;
wire [7:0] ID_EX_typ ;
wire [31:0] IF_ID_inst ;
wire [31:0] IF_ID_pc ;
wire [11:0] LS_WB_waddr_csreg ;
wire [3:0] LS_WB_waddr_reg ;
wire [31:0] LS_WB_wdata_csreg ;
wire [31:0] LS_WB_wdata_reg ;
wire [7:0] LS_WB_wen_csreg ;
wire [31:0] mepc ;
wire [31:0] mtvec ;
wire [63:0] \myclint.mtime ;
wire [0:0] \myclint.mtime_$_SDFF_PP0__Q_63_D ;
wire [31:0] \myec.mepc_tmp ;
wire [1:0] \myec.state ;
wire [31:0] \myexu.pc_jump ;
wire [3:0] \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [3:0] \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [2:0] \myidu.state ;
wire [31:0] \myifu.data_in ;
wire [3:0] \myifu.myicache.valid ;
wire [1:0] \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y ;
wire [31:0] \myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y ;
wire [2:0] \myifu.state ;
wire [2:0] \myifu.tmp_offset ;
wire [31:0] \mylsu.araddr_tmp ;
wire [31:0] \mylsu.awaddr_tmp ;
wire [4:0] \mylsu.state ;
wire [2:0] \mylsu.typ_tmp ;
wire [2:0] \myminixbar.state ;
wire [2:0] \mysc.state ;

assign \io_master_awid [1] = \io_master_awid [0] ;
assign \io_master_awid [2] = \io_master_arburst [1] ;
assign \io_master_awid [3] = \io_master_arburst [1] ;
assign \io_master_awlen [0] = \io_master_arburst [1] ;
assign \io_master_awlen [1] = \io_master_arburst [1] ;
assign \io_master_awlen [2] = \io_master_arburst [1] ;
assign \io_master_awlen [3] = \io_master_arburst [1] ;
assign \io_master_awlen [4] = \io_master_arburst [1] ;
assign \io_master_awlen [5] = \io_master_arburst [1] ;
assign \io_master_awlen [6] = \io_master_arburst [1] ;
assign \io_master_awlen [7] = \io_master_arburst [1] ;
assign \io_master_awsize [2] = \io_master_arburst [1] ;
assign \io_master_awburst [0] = \io_master_arburst [1] ;
assign \io_master_awburst [1] = \io_master_arburst [1] ;
assign io_master_wlast = \io_master_awid [0] ;
assign \io_master_arid [0] = \io_master_arburst [0] ;
assign \io_master_arid [2] = \io_master_arburst [1] ;
assign \io_master_arid [3] = \io_master_arburst [1] ;
assign \io_master_arlen [0] = \io_master_arburst [0] ;
assign \io_master_arlen [1] = \io_master_arburst [1] ;
assign \io_master_arlen [2] = \io_master_arburst [1] ;
assign \io_master_arlen [3] = \io_master_arburst [1] ;
assign \io_master_arlen [4] = \io_master_arburst [1] ;
assign \io_master_arlen [5] = \io_master_arburst [1] ;
assign \io_master_arlen [6] = \io_master_arburst [1] ;
assign \io_master_arlen [7] = \io_master_arburst [1] ;
assign io_slave_awready = \io_master_arburst [1] ;
assign io_slave_wready = \io_master_arburst [1] ;
assign io_slave_bvalid = \io_master_arburst [1] ;
assign \io_slave_bresp [0] = \io_master_arburst [1] ;
assign \io_slave_bresp [1] = \io_master_arburst [1] ;
assign \io_slave_bid [0] = \io_master_arburst [1] ;
assign \io_slave_bid [1] = \io_master_arburst [1] ;
assign \io_slave_bid [2] = \io_master_arburst [1] ;
assign \io_slave_bid [3] = \io_master_arburst [1] ;
assign io_slave_arready = \io_master_arburst [1] ;
assign io_slave_rvalid = \io_master_arburst [1] ;
assign \io_slave_rresp [0] = \io_master_arburst [1] ;
assign \io_slave_rresp [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [0] = \io_master_arburst [1] ;
assign \io_slave_rdata [1] = \io_master_arburst [1] ;
assign \io_slave_rdata [2] = \io_master_arburst [1] ;
assign \io_slave_rdata [3] = \io_master_arburst [1] ;
assign \io_slave_rdata [4] = \io_master_arburst [1] ;
assign \io_slave_rdata [5] = \io_master_arburst [1] ;
assign \io_slave_rdata [6] = \io_master_arburst [1] ;
assign \io_slave_rdata [7] = \io_master_arburst [1] ;
assign \io_slave_rdata [8] = \io_master_arburst [1] ;
assign \io_slave_rdata [9] = \io_master_arburst [1] ;
assign \io_slave_rdata [10] = \io_master_arburst [1] ;
assign \io_slave_rdata [11] = \io_master_arburst [1] ;
assign \io_slave_rdata [12] = \io_master_arburst [1] ;
assign \io_slave_rdata [13] = \io_master_arburst [1] ;
assign \io_slave_rdata [14] = \io_master_arburst [1] ;
assign \io_slave_rdata [15] = \io_master_arburst [1] ;
assign \io_slave_rdata [16] = \io_master_arburst [1] ;
assign \io_slave_rdata [17] = \io_master_arburst [1] ;
assign \io_slave_rdata [18] = \io_master_arburst [1] ;
assign \io_slave_rdata [19] = \io_master_arburst [1] ;
assign \io_slave_rdata [20] = \io_master_arburst [1] ;
assign \io_slave_rdata [21] = \io_master_arburst [1] ;
assign \io_slave_rdata [22] = \io_master_arburst [1] ;
assign \io_slave_rdata [23] = \io_master_arburst [1] ;
assign \io_slave_rdata [24] = \io_master_arburst [1] ;
assign \io_slave_rdata [25] = \io_master_arburst [1] ;
assign \io_slave_rdata [26] = \io_master_arburst [1] ;
assign \io_slave_rdata [27] = \io_master_arburst [1] ;
assign \io_slave_rdata [28] = \io_master_arburst [1] ;
assign \io_slave_rdata [29] = \io_master_arburst [1] ;
assign \io_slave_rdata [30] = \io_master_arburst [1] ;
assign \io_slave_rdata [31] = \io_master_arburst [1] ;
assign io_slave_rlast = \io_master_arburst [1] ;
assign \io_slave_rid [0] = \io_master_arburst [1] ;
assign \io_slave_rid [1] = \io_master_arburst [1] ;
assign \io_slave_rid [2] = \io_master_arburst [1] ;
assign \io_slave_rid [3] = \io_master_arburst [1] ;

INV_X1 _08944_ ( .A(\myec.state [1] ), .ZN(_01455_ ) );
AOI21_X1 _08945_ ( .A(excp_written ), .B1(_01455_ ), .B2(\myec.state [0] ), .ZN(_00000_ ) );
INV_X1 _08946_ ( .A(fanout_net_1 ), .ZN(_01456_ ) );
BUF_X4 _08947_ ( .A(_01456_ ), .Z(_01457_ ) );
BUF_X4 _08948_ ( .A(_01457_ ), .Z(_01458_ ) );
AND3_X4 _08949_ ( .A1(\myclint.mtime [2] ), .A2(\myclint.mtime [1] ), .A3(\myclint.mtime [0] ), .ZN(_01459_ ) );
AND3_X4 _08950_ ( .A1(_01459_ ), .A2(\myclint.mtime [4] ), .A3(\myclint.mtime [3] ), .ZN(_01460_ ) );
AND3_X4 _08951_ ( .A1(_01460_ ), .A2(\myclint.mtime [6] ), .A3(\myclint.mtime [5] ), .ZN(_01461_ ) );
AND3_X4 _08952_ ( .A1(_01461_ ), .A2(\myclint.mtime [8] ), .A3(\myclint.mtime [7] ), .ZN(_01462_ ) );
AND3_X4 _08953_ ( .A1(_01462_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [9] ), .ZN(_01463_ ) );
AND3_X4 _08954_ ( .A1(_01463_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [11] ), .ZN(_01464_ ) );
AND3_X4 _08955_ ( .A1(_01464_ ), .A2(\myclint.mtime [14] ), .A3(\myclint.mtime [13] ), .ZN(_01465_ ) );
AND3_X4 _08956_ ( .A1(_01465_ ), .A2(\myclint.mtime [16] ), .A3(\myclint.mtime [15] ), .ZN(_01466_ ) );
AND3_X4 _08957_ ( .A1(_01466_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [17] ), .ZN(_01467_ ) );
AND3_X4 _08958_ ( .A1(_01467_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [19] ), .ZN(_01468_ ) );
AND3_X4 _08959_ ( .A1(_01468_ ), .A2(\myclint.mtime [22] ), .A3(\myclint.mtime [21] ), .ZN(_01469_ ) );
AND3_X4 _08960_ ( .A1(_01469_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [23] ), .ZN(_01470_ ) );
AND3_X4 _08961_ ( .A1(_01470_ ), .A2(\myclint.mtime [26] ), .A3(\myclint.mtime [25] ), .ZN(_01471_ ) );
AND2_X4 _08962_ ( .A1(_01471_ ), .A2(\myclint.mtime [27] ), .ZN(_01472_ ) );
AND2_X1 _08963_ ( .A1(\myclint.mtime [30] ), .A2(\myclint.mtime [31] ), .ZN(_01473_ ) );
AND2_X1 _08964_ ( .A1(\myclint.mtime [28] ), .A2(\myclint.mtime [29] ), .ZN(_01474_ ) );
AND4_X2 _08965_ ( .A1(\myclint.mtime [33] ), .A2(_01472_ ), .A3(_01473_ ), .A4(_01474_ ), .ZN(_01475_ ) );
AND3_X4 _08966_ ( .A1(_01475_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [32] ), .ZN(_01476_ ) );
AND3_X4 _08967_ ( .A1(_01476_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [35] ), .ZN(_01477_ ) );
NAND3_X4 _08968_ ( .A1(_01477_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [37] ), .ZN(_01478_ ) );
INV_X1 _08969_ ( .A(\myclint.mtime [40] ), .ZN(_01479_ ) );
INV_X1 _08970_ ( .A(\myclint.mtime [39] ), .ZN(_01480_ ) );
NOR3_X2 _08971_ ( .A1(_01478_ ), .A2(_01479_ ), .A3(_01480_ ), .ZN(_01481_ ) );
AND2_X2 _08972_ ( .A1(_01481_ ), .A2(\myclint.mtime [41] ), .ZN(_01482_ ) );
AND2_X2 _08973_ ( .A1(\myclint.mtime [42] ), .A2(\myclint.mtime [43] ), .ZN(_01483_ ) );
AND2_X2 _08974_ ( .A1(_01482_ ), .A2(_01483_ ), .ZN(_01484_ ) );
AND2_X1 _08975_ ( .A1(\myclint.mtime [44] ), .A2(\myclint.mtime [45] ), .ZN(_01485_ ) );
AND3_X1 _08976_ ( .A1(_01485_ ), .A2(\myclint.mtime [46] ), .A3(\myclint.mtime [47] ), .ZN(_01486_ ) );
NAND2_X1 _08977_ ( .A1(_01484_ ), .A2(_01486_ ), .ZN(_01487_ ) );
AND2_X1 _08978_ ( .A1(\myclint.mtime [48] ), .A2(\myclint.mtime [49] ), .ZN(_01488_ ) );
INV_X1 _08979_ ( .A(_01488_ ), .ZN(_01489_ ) );
NOR2_X1 _08980_ ( .A1(_01487_ ), .A2(_01489_ ), .ZN(_01490_ ) );
AND2_X1 _08981_ ( .A1(\myclint.mtime [50] ), .A2(\myclint.mtime [51] ), .ZN(_01491_ ) );
AND2_X1 _08982_ ( .A1(_01490_ ), .A2(_01491_ ), .ZN(_01492_ ) );
AND2_X1 _08983_ ( .A1(\myclint.mtime [52] ), .A2(\myclint.mtime [53] ), .ZN(_01493_ ) );
AND2_X2 _08984_ ( .A1(_01492_ ), .A2(_01493_ ), .ZN(_01494_ ) );
AND2_X1 _08985_ ( .A1(\myclint.mtime [54] ), .A2(\myclint.mtime [55] ), .ZN(_01495_ ) );
NAND2_X1 _08986_ ( .A1(_01494_ ), .A2(_01495_ ), .ZN(_01496_ ) );
AND2_X1 _08987_ ( .A1(\myclint.mtime [56] ), .A2(\myclint.mtime [57] ), .ZN(_01497_ ) );
INV_X1 _08988_ ( .A(_01497_ ), .ZN(_01498_ ) );
NOR2_X2 _08989_ ( .A1(_01496_ ), .A2(_01498_ ), .ZN(_01499_ ) );
AND2_X1 _08990_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [59] ), .ZN(_01500_ ) );
AND2_X2 _08991_ ( .A1(_01499_ ), .A2(_01500_ ), .ZN(_01501_ ) );
NAND3_X2 _08992_ ( .A1(_01501_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01502_ ) );
NOR2_X2 _08993_ ( .A1(_01502_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01503_ ) );
OAI21_X1 _08994_ ( .A(_01458_ ), .B1(_01503_ ), .B2(\myclint.mtime [63] ), .ZN(_01504_ ) );
AND2_X2 _08995_ ( .A1(_01472_ ), .A2(_01474_ ), .ZN(_01505_ ) );
AND2_X1 _08996_ ( .A1(\myclint.mtime [33] ), .A2(\myclint.mtime [32] ), .ZN(_01506_ ) );
AND3_X2 _08997_ ( .A1(_01505_ ), .A2(_01506_ ), .A3(_01473_ ), .ZN(_01507_ ) );
AND3_X2 _08998_ ( .A1(_01507_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01508_ ) );
AND3_X2 _08999_ ( .A1(_01508_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .ZN(_01509_ ) );
NAND2_X1 _09000_ ( .A1(_01509_ ), .A2(\myclint.mtime [38] ), .ZN(_01510_ ) );
NOR3_X2 _09001_ ( .A1(_01510_ ), .A2(_01479_ ), .A3(_01480_ ), .ZN(_01511_ ) );
AND2_X2 _09002_ ( .A1(_01511_ ), .A2(\myclint.mtime [41] ), .ZN(_01512_ ) );
AND2_X2 _09003_ ( .A1(_01512_ ), .A2(_01483_ ), .ZN(_01513_ ) );
AND2_X2 _09004_ ( .A1(_01513_ ), .A2(_01486_ ), .ZN(_01514_ ) );
AND2_X2 _09005_ ( .A1(_01514_ ), .A2(_01488_ ), .ZN(_01515_ ) );
AND2_X1 _09006_ ( .A1(_01515_ ), .A2(_01491_ ), .ZN(_01516_ ) );
AND2_X2 _09007_ ( .A1(_01516_ ), .A2(_01493_ ), .ZN(_01517_ ) );
AND2_X2 _09008_ ( .A1(_01517_ ), .A2(_01495_ ), .ZN(_01518_ ) );
AND2_X2 _09009_ ( .A1(_01518_ ), .A2(_01497_ ), .ZN(_01519_ ) );
AND2_X1 _09010_ ( .A1(_01519_ ), .A2(_01500_ ), .ZN(_01520_ ) );
NAND3_X1 _09011_ ( .A1(_01520_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01521_ ) );
NOR2_X1 _09012_ ( .A1(_01521_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01522_ ) );
AOI21_X1 _09013_ ( .A(_01504_ ), .B1(_01522_ ), .B2(\myclint.mtime [63] ), .ZN(_00001_ ) );
AND2_X2 _09014_ ( .A1(_01461_ ), .A2(\myclint.mtime [7] ), .ZN(_01523_ ) );
AND4_X1 _09015_ ( .A1(\myclint.mtime [14] ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .A4(\myclint.mtime [15] ), .ZN(_01524_ ) );
AND2_X1 _09016_ ( .A1(\myclint.mtime [8] ), .A2(\myclint.mtime [9] ), .ZN(_01525_ ) );
AND4_X1 _09017_ ( .A1(\myclint.mtime [10] ), .A2(_01524_ ), .A3(\myclint.mtime [11] ), .A4(_01525_ ), .ZN(_01526_ ) );
NAND2_X1 _09018_ ( .A1(_01523_ ), .A2(_01526_ ), .ZN(_01527_ ) );
AND2_X1 _09019_ ( .A1(\myclint.mtime [16] ), .A2(\myclint.mtime [17] ), .ZN(_01528_ ) );
AND3_X1 _09020_ ( .A1(_01528_ ), .A2(\myclint.mtime [18] ), .A3(\myclint.mtime [19] ), .ZN(_01529_ ) );
AND4_X1 _09021_ ( .A1(\myclint.mtime [22] ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .A4(\myclint.mtime [23] ), .ZN(_01530_ ) );
AND2_X1 _09022_ ( .A1(_01529_ ), .A2(_01530_ ), .ZN(_01531_ ) );
AND2_X1 _09023_ ( .A1(\myclint.mtime [26] ), .A2(\myclint.mtime [27] ), .ZN(_01532_ ) );
AND3_X1 _09024_ ( .A1(_01532_ ), .A2(\myclint.mtime [24] ), .A3(\myclint.mtime [25] ), .ZN(_01533_ ) );
NAND4_X1 _09025_ ( .A1(_01531_ ), .A2(_01473_ ), .A3(_01474_ ), .A4(_01533_ ), .ZN(_01534_ ) );
NOR2_X1 _09026_ ( .A1(_01527_ ), .A2(_01534_ ), .ZN(_01535_ ) );
AND3_X1 _09027_ ( .A1(_01483_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01536_ ) );
AND3_X1 _09028_ ( .A1(_01506_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01537_ ) );
AND4_X1 _09029_ ( .A1(\myclint.mtime [38] ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .A4(\myclint.mtime [39] ), .ZN(_01538_ ) );
AND4_X1 _09030_ ( .A1(_01486_ ), .A2(_01536_ ), .A3(_01537_ ), .A4(_01538_ ), .ZN(_01539_ ) );
AND2_X1 _09031_ ( .A1(_01535_ ), .A2(_01539_ ), .ZN(_01540_ ) );
AND4_X1 _09032_ ( .A1(_01495_ ), .A2(_01493_ ), .A3(_01491_ ), .A4(_01488_ ), .ZN(_01541_ ) );
AND2_X1 _09033_ ( .A1(_01540_ ), .A2(_01541_ ), .ZN(_01542_ ) );
AND4_X1 _09034_ ( .A1(\myclint.mtime [58] ), .A2(\myclint.mtime [56] ), .A3(\myclint.mtime [57] ), .A4(\myclint.mtime [59] ), .ZN(_01543_ ) );
AND2_X1 _09035_ ( .A1(_01542_ ), .A2(_01543_ ), .ZN(_01544_ ) );
AND3_X1 _09036_ ( .A1(_01544_ ), .A2(\myclint.mtime [60] ), .A3(\myclint.mtime [61] ), .ZN(_01545_ ) );
XNOR2_X1 _09037_ ( .A(_01545_ ), .B(\myclint.mtime [62] ), .ZN(_01546_ ) );
NOR2_X1 _09038_ ( .A1(_01546_ ), .A2(fanout_net_1 ), .ZN(_00002_ ) );
INV_X1 _09039_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01547_ ) );
AND3_X1 _09040_ ( .A1(_01490_ ), .A2(_01547_ ), .A3(_01491_ ), .ZN(_01548_ ) );
OAI21_X1 _09041_ ( .A(_01458_ ), .B1(_01548_ ), .B2(\myclint.mtime [53] ), .ZN(_01549_ ) );
AND3_X1 _09042_ ( .A1(_01515_ ), .A2(_01547_ ), .A3(_01491_ ), .ZN(_01550_ ) );
AOI21_X1 _09043_ ( .A(_01549_ ), .B1(_01550_ ), .B2(\myclint.mtime [53] ), .ZN(_00003_ ) );
AND2_X1 _09044_ ( .A1(_01491_ ), .A2(_01488_ ), .ZN(_01551_ ) );
AND2_X1 _09045_ ( .A1(_01540_ ), .A2(_01551_ ), .ZN(_01552_ ) );
XNOR2_X1 _09046_ ( .A(_01552_ ), .B(\myclint.mtime [52] ), .ZN(_01553_ ) );
NOR2_X1 _09047_ ( .A1(_01553_ ), .A2(fanout_net_1 ), .ZN(_00004_ ) );
NOR3_X1 _09048_ ( .A1(_01487_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01489_ ), .ZN(_01554_ ) );
OAI21_X1 _09049_ ( .A(_01458_ ), .B1(_01554_ ), .B2(\myclint.mtime [51] ), .ZN(_01555_ ) );
INV_X1 _09050_ ( .A(_01514_ ), .ZN(_01556_ ) );
NOR3_X1 _09051_ ( .A1(_01556_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01489_ ), .ZN(_01557_ ) );
AOI21_X1 _09052_ ( .A(_01555_ ), .B1(_01557_ ), .B2(\myclint.mtime [51] ), .ZN(_00005_ ) );
INV_X1 _09053_ ( .A(_01535_ ), .ZN(_01558_ ) );
INV_X1 _09054_ ( .A(_01539_ ), .ZN(_01559_ ) );
OR4_X1 _09055_ ( .A1(\myclint.mtime [50] ), .A2(_01558_ ), .A3(_01489_ ), .A4(_01559_ ), .ZN(_01560_ ) );
AND3_X1 _09056_ ( .A1(_01535_ ), .A2(_01488_ ), .A3(_01539_ ), .ZN(_01561_ ) );
INV_X1 _09057_ ( .A(_01561_ ), .ZN(_01562_ ) );
NAND2_X1 _09058_ ( .A1(_01562_ ), .A2(\myclint.mtime [50] ), .ZN(_01563_ ) );
AOI21_X1 _09059_ ( .A(fanout_net_1 ), .B1(_01560_ ), .B2(_01563_ ), .ZN(_00006_ ) );
CLKBUF_X2 _09060_ ( .A(_01457_ ), .Z(_01564_ ) );
INV_X1 _09061_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01565_ ) );
AND3_X1 _09062_ ( .A1(_01484_ ), .A2(_01565_ ), .A3(_01486_ ), .ZN(_01566_ ) );
OAI21_X1 _09063_ ( .A(_01564_ ), .B1(_01566_ ), .B2(\myclint.mtime [49] ), .ZN(_01567_ ) );
AND4_X1 _09064_ ( .A1(\myclint.mtime [49] ), .A2(_01513_ ), .A3(_01565_ ), .A4(_01486_ ), .ZN(_01568_ ) );
NOR2_X1 _09065_ ( .A1(_01567_ ), .A2(_01568_ ), .ZN(_00007_ ) );
OAI21_X1 _09066_ ( .A(\myclint.mtime [48] ), .B1(_01558_ ), .B2(_01559_ ), .ZN(_01569_ ) );
OR4_X1 _09067_ ( .A1(\myclint.mtime [48] ), .A2(_01527_ ), .A3(_01534_ ), .A4(_01559_ ), .ZN(_01570_ ) );
AOI21_X1 _09068_ ( .A(fanout_net_1 ), .B1(_01569_ ), .B2(_01570_ ), .ZN(_00008_ ) );
NAND3_X1 _09069_ ( .A1(_01482_ ), .A2(_01485_ ), .A3(_01483_ ), .ZN(_01571_ ) );
NOR2_X1 _09070_ ( .A1(_01571_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01572_ ) );
OAI21_X1 _09071_ ( .A(_01458_ ), .B1(_01572_ ), .B2(\myclint.mtime [47] ), .ZN(_01573_ ) );
NAND3_X1 _09072_ ( .A1(_01512_ ), .A2(\myclint.mtime [44] ), .A3(_01483_ ), .ZN(_01574_ ) );
INV_X1 _09073_ ( .A(\myclint.mtime [45] ), .ZN(_01575_ ) );
NOR3_X1 _09074_ ( .A1(_01574_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01575_ ), .ZN(_01576_ ) );
AOI21_X1 _09075_ ( .A(_01573_ ), .B1(\myclint.mtime [47] ), .B2(_01576_ ), .ZN(_00009_ ) );
AND2_X1 _09076_ ( .A1(_01537_ ), .A2(_01538_ ), .ZN(_01577_ ) );
AND2_X1 _09077_ ( .A1(_01535_ ), .A2(_01577_ ), .ZN(_01578_ ) );
AND3_X1 _09078_ ( .A1(_01578_ ), .A2(_01485_ ), .A3(_01536_ ), .ZN(_01579_ ) );
XNOR2_X1 _09079_ ( .A(_01579_ ), .B(\myclint.mtime [46] ), .ZN(_01580_ ) );
NOR2_X1 _09080_ ( .A1(_01580_ ), .A2(fanout_net_1 ), .ZN(_00010_ ) );
INV_X1 _09081_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01581_ ) );
NAND3_X1 _09082_ ( .A1(_01482_ ), .A2(_01581_ ), .A3(_01483_ ), .ZN(_01582_ ) );
AOI21_X1 _09083_ ( .A(fanout_net_1 ), .B1(_01582_ ), .B2(_01575_ ), .ZN(_01583_ ) );
NAND4_X1 _09084_ ( .A1(_01512_ ), .A2(\myclint.mtime [45] ), .A3(_01581_ ), .A4(_01483_ ), .ZN(_01584_ ) );
AND2_X1 _09085_ ( .A1(_01583_ ), .A2(_01584_ ), .ZN(_00011_ ) );
AND2_X1 _09086_ ( .A1(_01578_ ), .A2(_01536_ ), .ZN(_01585_ ) );
XNOR2_X1 _09087_ ( .A(_01585_ ), .B(\myclint.mtime [44] ), .ZN(_01586_ ) );
NOR2_X1 _09088_ ( .A1(_01586_ ), .A2(fanout_net_1 ), .ZN(_00012_ ) );
INV_X1 _09089_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01587_ ) );
AND3_X1 _09090_ ( .A1(_01499_ ), .A2(_01587_ ), .A3(_01500_ ), .ZN(_01588_ ) );
OAI21_X1 _09091_ ( .A(_01458_ ), .B1(_01588_ ), .B2(\myclint.mtime [61] ), .ZN(_01589_ ) );
AND3_X1 _09092_ ( .A1(_01519_ ), .A2(_01587_ ), .A3(_01500_ ), .ZN(_01590_ ) );
AOI21_X1 _09093_ ( .A(_01589_ ), .B1(_01590_ ), .B2(\myclint.mtime [61] ), .ZN(_00013_ ) );
INV_X1 _09094_ ( .A(_01481_ ), .ZN(_01591_ ) );
INV_X1 _09095_ ( .A(\myclint.mtime [41] ), .ZN(_01592_ ) );
NOR3_X1 _09096_ ( .A1(_01591_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01592_ ), .ZN(_01593_ ) );
OAI21_X1 _09097_ ( .A(_01458_ ), .B1(_01593_ ), .B2(\myclint.mtime [43] ), .ZN(_01594_ ) );
INV_X1 _09098_ ( .A(_01511_ ), .ZN(_01595_ ) );
NOR3_X1 _09099_ ( .A1(_01595_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01592_ ), .ZN(_01596_ ) );
AOI21_X1 _09100_ ( .A(_01594_ ), .B1(\myclint.mtime [43] ), .B2(_01596_ ), .ZN(_00014_ ) );
INV_X1 _09101_ ( .A(_01578_ ), .ZN(_01597_ ) );
OR4_X1 _09102_ ( .A1(\myclint.mtime [42] ), .A2(_01597_ ), .A3(_01479_ ), .A4(_01592_ ), .ZN(_01598_ ) );
AND3_X1 _09103_ ( .A1(_01578_ ), .A2(\myclint.mtime [40] ), .A3(\myclint.mtime [41] ), .ZN(_01599_ ) );
INV_X1 _09104_ ( .A(_01599_ ), .ZN(_01600_ ) );
NAND2_X1 _09105_ ( .A1(_01600_ ), .A2(\myclint.mtime [42] ), .ZN(_01601_ ) );
AOI21_X1 _09106_ ( .A(fanout_net_1 ), .B1(_01598_ ), .B2(_01601_ ), .ZN(_00015_ ) );
BUF_X4 _09107_ ( .A(_01457_ ), .Z(_01602_ ) );
NOR3_X1 _09108_ ( .A1(_01478_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01480_ ), .ZN(_01603_ ) );
OAI21_X1 _09109_ ( .A(_01602_ ), .B1(_01603_ ), .B2(\myclint.mtime [41] ), .ZN(_01604_ ) );
NOR4_X1 _09110_ ( .A1(_01510_ ), .A2(_01592_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A4(_01480_ ), .ZN(_01605_ ) );
NOR2_X1 _09111_ ( .A1(_01604_ ), .A2(_01605_ ), .ZN(_00016_ ) );
NAND4_X1 _09112_ ( .A1(_01472_ ), .A2(\myclint.mtime [33] ), .A3(_01473_ ), .A4(_01474_ ), .ZN(_01606_ ) );
INV_X1 _09113_ ( .A(\myclint.mtime [32] ), .ZN(_01607_ ) );
NOR2_X1 _09114_ ( .A1(_01606_ ), .A2(_01607_ ), .ZN(_01608_ ) );
AND3_X1 _09115_ ( .A1(_01608_ ), .A2(\myclint.mtime [34] ), .A3(\myclint.mtime [35] ), .ZN(_01609_ ) );
AND3_X1 _09116_ ( .A1(_01609_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .ZN(_01610_ ) );
AND3_X1 _09117_ ( .A1(_01610_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [39] ), .ZN(_01611_ ) );
OAI21_X1 _09118_ ( .A(_01602_ ), .B1(_01611_ ), .B2(\myclint.mtime [40] ), .ZN(_01612_ ) );
NOR2_X1 _09119_ ( .A1(_01612_ ), .A2(_01481_ ), .ZN(_00017_ ) );
AND2_X1 _09120_ ( .A1(_01535_ ), .A2(_01537_ ), .ZN(_01613_ ) );
NAND3_X1 _09121_ ( .A1(_01613_ ), .A2(\myclint.mtime [36] ), .A3(\myclint.mtime [37] ), .ZN(_01614_ ) );
NOR2_X1 _09122_ ( .A1(_01614_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01615_ ) );
XNOR2_X1 _09123_ ( .A(_01615_ ), .B(\myclint.mtime [39] ), .ZN(_01616_ ) );
NOR2_X1 _09124_ ( .A1(_01616_ ), .A2(fanout_net_1 ), .ZN(_00018_ ) );
OAI21_X1 _09125_ ( .A(_01602_ ), .B1(_01610_ ), .B2(\myclint.mtime [38] ), .ZN(_01617_ ) );
AND3_X1 _09126_ ( .A1(_01477_ ), .A2(\myclint.mtime [38] ), .A3(\myclint.mtime [37] ), .ZN(_01618_ ) );
NOR2_X1 _09127_ ( .A1(_01617_ ), .A2(_01618_ ), .ZN(_00019_ ) );
INV_X1 _09128_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01619_ ) );
AND3_X1 _09129_ ( .A1(_01476_ ), .A2(_01619_ ), .A3(\myclint.mtime [35] ), .ZN(_01620_ ) );
OAI21_X1 _09130_ ( .A(_01602_ ), .B1(_01620_ ), .B2(\myclint.mtime [37] ), .ZN(_01621_ ) );
AND3_X1 _09131_ ( .A1(_01508_ ), .A2(\myclint.mtime [37] ), .A3(_01619_ ), .ZN(_01622_ ) );
NOR2_X1 _09132_ ( .A1(_01621_ ), .A2(_01622_ ), .ZN(_00020_ ) );
OAI21_X1 _09133_ ( .A(_01602_ ), .B1(_01609_ ), .B2(\myclint.mtime [36] ), .ZN(_01623_ ) );
NOR2_X1 _09134_ ( .A1(_01623_ ), .A2(_01477_ ), .ZN(_00021_ ) );
INV_X1 _09135_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01624_ ) );
AND3_X1 _09136_ ( .A1(_01507_ ), .A2(_01624_ ), .A3(\myclint.mtime [35] ), .ZN(_01625_ ) );
BUF_X4 _09137_ ( .A(_01457_ ), .Z(_01626_ ) );
NOR3_X1 _09138_ ( .A1(_01606_ ), .A2(_01607_ ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01627_ ) );
OAI21_X1 _09139_ ( .A(_01626_ ), .B1(_01627_ ), .B2(\myclint.mtime [35] ), .ZN(_01628_ ) );
NOR2_X1 _09140_ ( .A1(_01625_ ), .A2(_01628_ ), .ZN(_00022_ ) );
OAI21_X1 _09141_ ( .A(_01602_ ), .B1(_01608_ ), .B2(\myclint.mtime [34] ), .ZN(_01629_ ) );
NOR2_X1 _09142_ ( .A1(_01629_ ), .A2(_01476_ ), .ZN(_00023_ ) );
XNOR2_X1 _09143_ ( .A(_01544_ ), .B(\myclint.mtime [60] ), .ZN(_01630_ ) );
NOR2_X1 _09144_ ( .A1(_01630_ ), .A2(fanout_net_1 ), .ZN(_00024_ ) );
OR3_X1 _09145_ ( .A1(_01527_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_01534_ ), .ZN(_01631_ ) );
NAND2_X1 _09146_ ( .A1(_01631_ ), .A2(\myclint.mtime [33] ), .ZN(_01632_ ) );
OR4_X1 _09147_ ( .A1(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A2(_01527_ ), .A3(\myclint.mtime [33] ), .A4(_01534_ ), .ZN(_01633_ ) );
AOI21_X1 _09148_ ( .A(fanout_net_1 ), .B1(_01632_ ), .B2(_01633_ ), .ZN(_00025_ ) );
OAI21_X1 _09149_ ( .A(\myclint.mtime [32] ), .B1(_01527_ ), .B2(_01534_ ), .ZN(_01634_ ) );
AND4_X1 _09150_ ( .A1(_01473_ ), .A2(_01531_ ), .A3(_01474_ ), .A4(_01533_ ), .ZN(_01635_ ) );
NAND4_X1 _09151_ ( .A1(_01635_ ), .A2(_01523_ ), .A3(_01607_ ), .A4(_01526_ ), .ZN(_01636_ ) );
AOI21_X1 _09152_ ( .A(fanout_net_1 ), .B1(_01634_ ), .B2(_01636_ ), .ZN(_00026_ ) );
AND2_X1 _09153_ ( .A1(_01523_ ), .A2(_01526_ ), .ZN(_01637_ ) );
AND2_X1 _09154_ ( .A1(_01637_ ), .A2(_01531_ ), .ZN(_01638_ ) );
NAND3_X1 _09155_ ( .A1(_01638_ ), .A2(_01474_ ), .A3(_01533_ ), .ZN(_01639_ ) );
OR3_X1 _09156_ ( .A1(_01639_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [31] ), .ZN(_01640_ ) );
OAI21_X1 _09157_ ( .A(\myclint.mtime [31] ), .B1(_01639_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01641_ ) );
AOI21_X1 _09158_ ( .A(fanout_net_1 ), .B1(_01640_ ), .B2(_01641_ ), .ZN(_00027_ ) );
OR2_X1 _09159_ ( .A1(_01639_ ), .A2(\myclint.mtime [30] ), .ZN(_01642_ ) );
NAND2_X1 _09160_ ( .A1(_01639_ ), .A2(\myclint.mtime [30] ), .ZN(_01643_ ) );
AOI21_X1 _09161_ ( .A(fanout_net_1 ), .B1(_01642_ ), .B2(_01643_ ), .ZN(_00028_ ) );
INV_X1 _09162_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01644_ ) );
AND3_X1 _09163_ ( .A1(_01471_ ), .A2(_01644_ ), .A3(\myclint.mtime [27] ), .ZN(_01645_ ) );
AND2_X1 _09164_ ( .A1(_01645_ ), .A2(\myclint.mtime [29] ), .ZN(_01646_ ) );
OAI21_X1 _09165_ ( .A(_01626_ ), .B1(_01645_ ), .B2(\myclint.mtime [29] ), .ZN(_01647_ ) );
NOR2_X1 _09166_ ( .A1(_01646_ ), .A2(_01647_ ), .ZN(_00029_ ) );
NAND2_X1 _09167_ ( .A1(_01638_ ), .A2(_01533_ ), .ZN(_01648_ ) );
OR2_X1 _09168_ ( .A1(_01648_ ), .A2(\myclint.mtime [28] ), .ZN(_01649_ ) );
NAND2_X1 _09169_ ( .A1(_01648_ ), .A2(\myclint.mtime [28] ), .ZN(_01650_ ) );
AOI21_X1 _09170_ ( .A(fanout_net_1 ), .B1(_01649_ ), .B2(_01650_ ), .ZN(_00030_ ) );
INV_X1 _09171_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01651_ ) );
AND3_X1 _09172_ ( .A1(_01470_ ), .A2(_01651_ ), .A3(\myclint.mtime [25] ), .ZN(_01652_ ) );
AND2_X1 _09173_ ( .A1(_01652_ ), .A2(\myclint.mtime [27] ), .ZN(_01653_ ) );
OAI21_X1 _09174_ ( .A(_01626_ ), .B1(_01652_ ), .B2(\myclint.mtime [27] ), .ZN(_01654_ ) );
NOR2_X1 _09175_ ( .A1(_01653_ ), .A2(_01654_ ), .ZN(_00031_ ) );
AND2_X1 _09176_ ( .A1(_01470_ ), .A2(\myclint.mtime [25] ), .ZN(_01655_ ) );
OAI21_X1 _09177_ ( .A(_01602_ ), .B1(_01655_ ), .B2(\myclint.mtime [26] ), .ZN(_01656_ ) );
NOR2_X1 _09178_ ( .A1(_01656_ ), .A2(_01471_ ), .ZN(_00032_ ) );
INV_X1 _09179_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01657_ ) );
AND3_X1 _09180_ ( .A1(_01469_ ), .A2(_01657_ ), .A3(\myclint.mtime [23] ), .ZN(_01658_ ) );
AND2_X1 _09181_ ( .A1(_01658_ ), .A2(\myclint.mtime [25] ), .ZN(_01659_ ) );
OAI21_X1 _09182_ ( .A(_01626_ ), .B1(_01658_ ), .B2(\myclint.mtime [25] ), .ZN(_01660_ ) );
NOR2_X1 _09183_ ( .A1(_01659_ ), .A2(_01660_ ), .ZN(_00033_ ) );
AND2_X1 _09184_ ( .A1(_01469_ ), .A2(\myclint.mtime [23] ), .ZN(_01661_ ) );
OAI21_X1 _09185_ ( .A(_01602_ ), .B1(_01661_ ), .B2(\myclint.mtime [24] ), .ZN(_01662_ ) );
NOR2_X1 _09186_ ( .A1(_01662_ ), .A2(_01470_ ), .ZN(_00034_ ) );
NOR3_X1 _09187_ ( .A1(_01496_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_01498_ ), .ZN(_01663_ ) );
OAI21_X1 _09188_ ( .A(_01458_ ), .B1(_01663_ ), .B2(\myclint.mtime [59] ), .ZN(_01664_ ) );
INV_X1 _09189_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01665_ ) );
AND3_X1 _09190_ ( .A1(_01518_ ), .A2(_01665_ ), .A3(_01497_ ), .ZN(_01666_ ) );
AOI21_X1 _09191_ ( .A(_01664_ ), .B1(_01666_ ), .B2(\myclint.mtime [59] ), .ZN(_00035_ ) );
AND2_X1 _09192_ ( .A1(_01637_ ), .A2(_01529_ ), .ZN(_01667_ ) );
NAND3_X1 _09193_ ( .A1(_01667_ ), .A2(\myclint.mtime [20] ), .A3(\myclint.mtime [21] ), .ZN(_01668_ ) );
OR3_X1 _09194_ ( .A1(_01668_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [23] ), .ZN(_01669_ ) );
OAI21_X1 _09195_ ( .A(\myclint.mtime [23] ), .B1(_01668_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01670_ ) );
AOI21_X1 _09196_ ( .A(fanout_net_1 ), .B1(_01669_ ), .B2(_01670_ ), .ZN(_00036_ ) );
AND2_X1 _09197_ ( .A1(_01468_ ), .A2(\myclint.mtime [21] ), .ZN(_01671_ ) );
OAI21_X1 _09198_ ( .A(_01602_ ), .B1(_01671_ ), .B2(\myclint.mtime [22] ), .ZN(_01672_ ) );
NOR2_X1 _09199_ ( .A1(_01672_ ), .A2(_01469_ ), .ZN(_00037_ ) );
INV_X1 _09200_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01673_ ) );
AND3_X1 _09201_ ( .A1(_01467_ ), .A2(_01673_ ), .A3(\myclint.mtime [19] ), .ZN(_01674_ ) );
AND2_X1 _09202_ ( .A1(_01674_ ), .A2(\myclint.mtime [21] ), .ZN(_01675_ ) );
OAI21_X1 _09203_ ( .A(_01626_ ), .B1(_01674_ ), .B2(\myclint.mtime [21] ), .ZN(_01676_ ) );
NOR2_X1 _09204_ ( .A1(_01675_ ), .A2(_01676_ ), .ZN(_00038_ ) );
AND2_X1 _09205_ ( .A1(_01467_ ), .A2(\myclint.mtime [19] ), .ZN(_01677_ ) );
OAI21_X1 _09206_ ( .A(_01602_ ), .B1(_01677_ ), .B2(\myclint.mtime [20] ), .ZN(_01678_ ) );
NOR2_X1 _09207_ ( .A1(_01678_ ), .A2(_01468_ ), .ZN(_00039_ ) );
NAND3_X1 _09208_ ( .A1(_01523_ ), .A2(_01526_ ), .A3(_01528_ ), .ZN(_01679_ ) );
OR3_X1 _09209_ ( .A1(_01679_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [19] ), .ZN(_01680_ ) );
OAI21_X1 _09210_ ( .A(\myclint.mtime [19] ), .B1(_01679_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01681_ ) );
AOI21_X1 _09211_ ( .A(fanout_net_1 ), .B1(_01680_ ), .B2(_01681_ ), .ZN(_00040_ ) );
BUF_X2 _09212_ ( .A(_01457_ ), .Z(_01682_ ) );
AND2_X1 _09213_ ( .A1(_01466_ ), .A2(\myclint.mtime [17] ), .ZN(_01683_ ) );
OAI21_X1 _09214_ ( .A(_01682_ ), .B1(_01683_ ), .B2(\myclint.mtime [18] ), .ZN(_01684_ ) );
NOR2_X1 _09215_ ( .A1(_01684_ ), .A2(_01467_ ), .ZN(_00041_ ) );
INV_X1 _09216_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01685_ ) );
AND3_X1 _09217_ ( .A1(_01465_ ), .A2(_01685_ ), .A3(\myclint.mtime [15] ), .ZN(_01686_ ) );
AND2_X1 _09218_ ( .A1(_01686_ ), .A2(\myclint.mtime [17] ), .ZN(_01687_ ) );
OAI21_X1 _09219_ ( .A(_01626_ ), .B1(_01686_ ), .B2(\myclint.mtime [17] ), .ZN(_01688_ ) );
NOR2_X1 _09220_ ( .A1(_01687_ ), .A2(_01688_ ), .ZN(_00042_ ) );
AND2_X1 _09221_ ( .A1(_01465_ ), .A2(\myclint.mtime [15] ), .ZN(_01689_ ) );
OAI21_X1 _09222_ ( .A(_01682_ ), .B1(_01689_ ), .B2(\myclint.mtime [16] ), .ZN(_01690_ ) );
NOR2_X1 _09223_ ( .A1(_01690_ ), .A2(_01466_ ), .ZN(_00043_ ) );
AND3_X1 _09224_ ( .A1(_01525_ ), .A2(\myclint.mtime [10] ), .A3(\myclint.mtime [11] ), .ZN(_01691_ ) );
AND2_X1 _09225_ ( .A1(_01523_ ), .A2(_01691_ ), .ZN(_01692_ ) );
NAND3_X1 _09226_ ( .A1(_01692_ ), .A2(\myclint.mtime [12] ), .A3(\myclint.mtime [13] ), .ZN(_01693_ ) );
OR3_X1 _09227_ ( .A1(_01693_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [15] ), .ZN(_01694_ ) );
OAI21_X1 _09228_ ( .A(\myclint.mtime [15] ), .B1(_01693_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01695_ ) );
AOI21_X1 _09229_ ( .A(fanout_net_1 ), .B1(_01694_ ), .B2(_01695_ ), .ZN(_00044_ ) );
AND2_X1 _09230_ ( .A1(_01464_ ), .A2(\myclint.mtime [13] ), .ZN(_01696_ ) );
OAI21_X1 _09231_ ( .A(_01682_ ), .B1(_01696_ ), .B2(\myclint.mtime [14] ), .ZN(_01697_ ) );
NOR2_X1 _09232_ ( .A1(_01697_ ), .A2(_01465_ ), .ZN(_00045_ ) );
NAND3_X1 _09233_ ( .A1(_01540_ ), .A2(_01497_ ), .A3(_01541_ ), .ZN(_01698_ ) );
OR2_X1 _09234_ ( .A1(_01698_ ), .A2(\myclint.mtime [58] ), .ZN(_01699_ ) );
NAND2_X1 _09235_ ( .A1(_01698_ ), .A2(\myclint.mtime [58] ), .ZN(_01700_ ) );
AOI21_X1 _09236_ ( .A(fanout_net_1 ), .B1(_01699_ ), .B2(_01700_ ), .ZN(_00046_ ) );
INV_X1 _09237_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01701_ ) );
AND3_X1 _09238_ ( .A1(_01463_ ), .A2(_01701_ ), .A3(\myclint.mtime [11] ), .ZN(_01702_ ) );
AND2_X1 _09239_ ( .A1(_01702_ ), .A2(\myclint.mtime [13] ), .ZN(_01703_ ) );
OAI21_X1 _09240_ ( .A(_01626_ ), .B1(_01702_ ), .B2(\myclint.mtime [13] ), .ZN(_01704_ ) );
NOR2_X1 _09241_ ( .A1(_01703_ ), .A2(_01704_ ), .ZN(_00047_ ) );
AND2_X1 _09242_ ( .A1(_01463_ ), .A2(\myclint.mtime [11] ), .ZN(_01705_ ) );
OAI21_X1 _09243_ ( .A(_01682_ ), .B1(_01705_ ), .B2(\myclint.mtime [12] ), .ZN(_01706_ ) );
NOR2_X1 _09244_ ( .A1(_01706_ ), .A2(_01464_ ), .ZN(_00048_ ) );
NAND3_X1 _09245_ ( .A1(_01461_ ), .A2(\myclint.mtime [7] ), .A3(_01525_ ), .ZN(_01707_ ) );
OR3_X1 _09246_ ( .A1(_01707_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [11] ), .ZN(_01708_ ) );
OAI21_X1 _09247_ ( .A(\myclint.mtime [11] ), .B1(_01707_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01709_ ) );
AOI21_X1 _09248_ ( .A(fanout_net_1 ), .B1(_01708_ ), .B2(_01709_ ), .ZN(_00049_ ) );
AOI21_X1 _09249_ ( .A(\myclint.mtime [10] ), .B1(_01462_ ), .B2(\myclint.mtime [9] ), .ZN(_01710_ ) );
NOR3_X1 _09250_ ( .A1(_01463_ ), .A2(_01710_ ), .A3(fanout_net_1 ), .ZN(_00050_ ) );
INV_X1 _09251_ ( .A(_01523_ ), .ZN(_01711_ ) );
OR3_X1 _09252_ ( .A1(_01711_ ), .A2(\myclint.mtime [9] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01712_ ) );
OAI21_X1 _09253_ ( .A(\myclint.mtime [9] ), .B1(_01711_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01713_ ) );
AOI21_X1 _09254_ ( .A(fanout_net_1 ), .B1(_01712_ ), .B2(_01713_ ), .ZN(_00051_ ) );
OAI21_X1 _09255_ ( .A(_01682_ ), .B1(_01523_ ), .B2(\myclint.mtime [8] ), .ZN(_01714_ ) );
NOR2_X1 _09256_ ( .A1(_01714_ ), .A2(_01462_ ), .ZN(_00052_ ) );
AND2_X1 _09257_ ( .A1(_01460_ ), .A2(\myclint.mtime [5] ), .ZN(_01715_ ) );
INV_X1 _09258_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01716_ ) );
AND3_X1 _09259_ ( .A1(_01715_ ), .A2(_01716_ ), .A3(\myclint.mtime [7] ), .ZN(_01717_ ) );
AOI21_X1 _09260_ ( .A(\myclint.mtime [7] ), .B1(_01715_ ), .B2(_01716_ ), .ZN(_01718_ ) );
NOR3_X1 _09261_ ( .A1(_01717_ ), .A2(_01718_ ), .A3(fanout_net_1 ), .ZN(_00053_ ) );
OAI21_X1 _09262_ ( .A(_01682_ ), .B1(_01715_ ), .B2(\myclint.mtime [6] ), .ZN(_01719_ ) );
NOR2_X1 _09263_ ( .A1(_01719_ ), .A2(_01461_ ), .ZN(_00054_ ) );
AND2_X1 _09264_ ( .A1(_01459_ ), .A2(\myclint.mtime [3] ), .ZN(_01720_ ) );
INV_X1 _09265_ ( .A(_01720_ ), .ZN(_01721_ ) );
OR3_X1 _09266_ ( .A1(_01721_ ), .A2(\myclint.mtime [5] ), .A3(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01722_ ) );
OAI21_X1 _09267_ ( .A(\myclint.mtime [5] ), .B1(_01721_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01723_ ) );
AOI21_X1 _09268_ ( .A(fanout_net_1 ), .B1(_01722_ ), .B2(_01723_ ), .ZN(_00055_ ) );
OAI21_X1 _09269_ ( .A(_01682_ ), .B1(_01720_ ), .B2(\myclint.mtime [4] ), .ZN(_01724_ ) );
NOR2_X1 _09270_ ( .A1(_01724_ ), .A2(_01460_ ), .ZN(_00056_ ) );
INV_X1 _09271_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01725_ ) );
AND3_X1 _09272_ ( .A1(_01494_ ), .A2(_01725_ ), .A3(_01495_ ), .ZN(_01726_ ) );
OAI21_X1 _09273_ ( .A(_01458_ ), .B1(_01726_ ), .B2(\myclint.mtime [57] ), .ZN(_01727_ ) );
AND3_X1 _09274_ ( .A1(_01517_ ), .A2(_01725_ ), .A3(_01495_ ), .ZN(_01728_ ) );
AOI21_X1 _09275_ ( .A(_01727_ ), .B1(_01728_ ), .B2(\myclint.mtime [57] ), .ZN(_00057_ ) );
AND2_X1 _09276_ ( .A1(\myclint.mtime [1] ), .A2(\myclint.mtime [0] ), .ZN(_01729_ ) );
INV_X1 _09277_ ( .A(_01729_ ), .ZN(_01730_ ) );
OR3_X1 _09278_ ( .A1(_01730_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .A3(\myclint.mtime [3] ), .ZN(_01731_ ) );
OAI21_X1 _09279_ ( .A(\myclint.mtime [3] ), .B1(_01730_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_01732_ ) );
AOI21_X1 _09280_ ( .A(fanout_net_1 ), .B1(_01731_ ), .B2(_01732_ ), .ZN(_00058_ ) );
AOI21_X1 _09281_ ( .A(\myclint.mtime [2] ), .B1(\myclint.mtime [1] ), .B2(\myclint.mtime [0] ), .ZN(_01733_ ) );
NOR3_X1 _09282_ ( .A1(_01459_ ), .A2(_01733_ ), .A3(fanout_net_1 ), .ZN(_00059_ ) );
NOR2_X1 _09283_ ( .A1(\myclint.mtime [1] ), .A2(\myclint.mtime [0] ), .ZN(_01734_ ) );
NOR3_X1 _09284_ ( .A1(_01729_ ), .A2(_01734_ ), .A3(fanout_net_1 ), .ZN(_00060_ ) );
CLKBUF_X2 _09285_ ( .A(_01457_ ), .Z(_01735_ ) );
AND2_X1 _09286_ ( .A1(_01735_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .ZN(_00061_ ) );
XNOR2_X1 _09287_ ( .A(_01542_ ), .B(\myclint.mtime [56] ), .ZN(_01736_ ) );
NOR2_X1 _09288_ ( .A1(_01736_ ), .A2(fanout_net_1 ), .ZN(_00062_ ) );
NAND3_X1 _09289_ ( .A1(_01540_ ), .A2(_01493_ ), .A3(_01551_ ), .ZN(_01737_ ) );
OR3_X1 _09290_ ( .A1(_01737_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(\myclint.mtime [55] ), .ZN(_01738_ ) );
OAI21_X1 _09291_ ( .A(\myclint.mtime [55] ), .B1(_01737_ ), .B2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_01739_ ) );
AOI21_X1 _09292_ ( .A(fanout_net_1 ), .B1(_01738_ ), .B2(_01739_ ), .ZN(_00063_ ) );
OR2_X1 _09293_ ( .A1(_01737_ ), .A2(\myclint.mtime [54] ), .ZN(_01740_ ) );
NAND2_X1 _09294_ ( .A1(_01737_ ), .A2(\myclint.mtime [54] ), .ZN(_01741_ ) );
AOI21_X1 _09295_ ( .A(fanout_net_2 ), .B1(_01740_ ), .B2(_01741_ ), .ZN(_00064_ ) );
INV_X32 _09296_ ( .A(fanout_net_48 ), .ZN(_01742_ ) );
BUF_X32 _09297_ ( .A(_01742_ ), .Z(_01743_ ) );
OR2_X1 _09298_ ( .A1(_01743_ ), .A2(\myifu.myicache.tag[3][1] ), .ZN(_01744_ ) );
OAI211_X1 _09299_ ( .A(_01744_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_48 ), .C2(\myifu.myicache.tag[2][1] ), .ZN(_01745_ ) );
OR2_X1 _09300_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][1] ), .ZN(_01746_ ) );
INV_X32 _09301_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01747_ ) );
BUF_X2 _09302_ ( .A(_01747_ ), .Z(_01748_ ) );
BUF_X8 _09303_ ( .A(_01743_ ), .Z(_01749_ ) );
OAI211_X1 _09304_ ( .A(_01746_ ), .B(_01748_ ), .C1(_01749_ ), .C2(\myifu.myicache.tag[1][1] ), .ZN(_01750_ ) );
AND3_X1 _09305_ ( .A1(_01745_ ), .A2(\IF_ID_pc [6] ), .A3(_01750_ ), .ZN(_01751_ ) );
OR2_X1 _09306_ ( .A1(_01742_ ), .A2(\myifu.myicache.tag[3][12] ), .ZN(_01752_ ) );
OAI211_X1 _09307_ ( .A(_01752_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_48 ), .C2(\myifu.myicache.tag[2][12] ), .ZN(_01753_ ) );
OR2_X1 _09308_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][12] ), .ZN(_01754_ ) );
BUF_X32 _09309_ ( .A(_01747_ ), .Z(_01755_ ) );
BUF_X16 _09310_ ( .A(_01742_ ), .Z(_01756_ ) );
OAI211_X1 _09311_ ( .A(_01754_ ), .B(_01755_ ), .C1(_01756_ ), .C2(\myifu.myicache.tag[1][12] ), .ZN(_01757_ ) );
NAND2_X1 _09312_ ( .A1(_01753_ ), .A2(_01757_ ), .ZN(_01758_ ) );
INV_X1 _09313_ ( .A(\IF_ID_pc [17] ), .ZN(_01759_ ) );
XNOR2_X1 _09314_ ( .A(_01758_ ), .B(_01759_ ), .ZN(_01760_ ) );
OR2_X4 _09315_ ( .A1(_01742_ ), .A2(\myifu.myicache.tag[1][26] ), .ZN(_01761_ ) );
OAI211_X1 _09316_ ( .A(_01761_ ), .B(_01755_ ), .C1(fanout_net_48 ), .C2(\myifu.myicache.tag[0][26] ), .ZN(_01762_ ) );
OR2_X1 _09317_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][26] ), .ZN(_01763_ ) );
OAI211_X1 _09318_ ( .A(_01763_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01743_ ), .C2(\myifu.myicache.tag[3][26] ), .ZN(_01764_ ) );
INV_X1 _09319_ ( .A(\IF_ID_pc [31] ), .ZN(_01765_ ) );
AND3_X1 _09320_ ( .A1(_01762_ ), .A2(_01764_ ), .A3(_01765_ ), .ZN(_01766_ ) );
AOI21_X1 _09321_ ( .A(_01765_ ), .B1(_01762_ ), .B2(_01764_ ), .ZN(_01767_ ) );
OR2_X1 _09322_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][0] ), .ZN(_01768_ ) );
OAI211_X1 _09323_ ( .A(_01768_ ), .B(_01755_ ), .C1(_01743_ ), .C2(\myifu.myicache.tag[1][0] ), .ZN(_01769_ ) );
OR2_X2 _09324_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][0] ), .ZN(_01770_ ) );
OAI211_X1 _09325_ ( .A(_01770_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01743_ ), .C2(\myifu.myicache.tag[3][0] ), .ZN(_01771_ ) );
AND3_X2 _09326_ ( .A1(_01769_ ), .A2(_01771_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_01772_ ) );
AOI21_X1 _09327_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B1(_01769_ ), .B2(_01771_ ), .ZN(_01773_ ) );
OAI22_X1 _09328_ ( .A1(_01766_ ), .A2(_01767_ ), .B1(_01772_ ), .B2(_01773_ ), .ZN(_01774_ ) );
AOI21_X1 _09329_ ( .A(\IF_ID_pc [6] ), .B1(_01745_ ), .B2(_01750_ ), .ZN(_01775_ ) );
OR4_X1 _09330_ ( .A1(_01751_ ), .A2(_01760_ ), .A3(_01774_ ), .A4(_01775_ ), .ZN(_01776_ ) );
OR2_X1 _09331_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][10] ), .ZN(_01777_ ) );
OAI211_X1 _09332_ ( .A(_01777_ ), .B(_01755_ ), .C1(_01756_ ), .C2(\myifu.myicache.tag[1][10] ), .ZN(_01778_ ) );
OR2_X1 _09333_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][10] ), .ZN(_01779_ ) );
OAI211_X1 _09334_ ( .A(_01779_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01743_ ), .C2(\myifu.myicache.tag[3][10] ), .ZN(_01780_ ) );
NAND2_X1 _09335_ ( .A1(_01778_ ), .A2(_01780_ ), .ZN(_01781_ ) );
XOR2_X1 _09336_ ( .A(_01781_ ), .B(\IF_ID_pc [15] ), .Z(_01782_ ) );
OR2_X1 _09337_ ( .A1(_01742_ ), .A2(\myifu.myicache.tag[3][17] ), .ZN(_01783_ ) );
OAI211_X1 _09338_ ( .A(_01783_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(fanout_net_48 ), .C2(\myifu.myicache.tag[2][17] ), .ZN(_01784_ ) );
INV_X1 _09339_ ( .A(\IF_ID_pc [22] ), .ZN(_01785_ ) );
OR2_X1 _09340_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][17] ), .ZN(_01786_ ) );
OAI211_X1 _09341_ ( .A(_01786_ ), .B(_01755_ ), .C1(_01743_ ), .C2(\myifu.myicache.tag[1][17] ), .ZN(_01787_ ) );
AND3_X1 _09342_ ( .A1(_01784_ ), .A2(_01785_ ), .A3(_01787_ ), .ZN(_01788_ ) );
AOI21_X1 _09343_ ( .A(_01785_ ), .B1(_01784_ ), .B2(_01787_ ), .ZN(_01789_ ) );
OR2_X1 _09344_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][4] ), .ZN(_01790_ ) );
OAI211_X1 _09345_ ( .A(_01790_ ), .B(_01755_ ), .C1(_01743_ ), .C2(\myifu.myicache.tag[1][4] ), .ZN(_01791_ ) );
OR2_X2 _09346_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][4] ), .ZN(_01792_ ) );
OAI211_X1 _09347_ ( .A(_01792_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01742_ ), .C2(\myifu.myicache.tag[3][4] ), .ZN(_01793_ ) );
INV_X1 _09348_ ( .A(\IF_ID_pc [9] ), .ZN(_01794_ ) );
AND3_X2 _09349_ ( .A1(_01791_ ), .A2(_01793_ ), .A3(_01794_ ), .ZN(_01795_ ) );
AOI21_X1 _09350_ ( .A(_01794_ ), .B1(_01791_ ), .B2(_01793_ ), .ZN(_01796_ ) );
OAI22_X1 _09351_ ( .A1(_01788_ ), .A2(_01789_ ), .B1(_01795_ ), .B2(_01796_ ), .ZN(_01797_ ) );
OR2_X1 _09352_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][8] ), .ZN(_01798_ ) );
OAI211_X1 _09353_ ( .A(_01798_ ), .B(_01755_ ), .C1(_01756_ ), .C2(\myifu.myicache.tag[1][8] ), .ZN(_01799_ ) );
OR2_X1 _09354_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][8] ), .ZN(_01800_ ) );
OAI211_X1 _09355_ ( .A(_01800_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01756_ ), .C2(\myifu.myicache.tag[3][8] ), .ZN(_01801_ ) );
AND3_X1 _09356_ ( .A1(_01799_ ), .A2(_01801_ ), .A3(\IF_ID_pc [13] ), .ZN(_01802_ ) );
AOI21_X1 _09357_ ( .A(\IF_ID_pc [13] ), .B1(_01799_ ), .B2(_01801_ ), .ZN(_01803_ ) );
OR4_X2 _09358_ ( .A1(_01782_ ), .A2(_01797_ ), .A3(_01802_ ), .A4(_01803_ ), .ZN(_01804_ ) );
OR2_X1 _09359_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][6] ), .ZN(_01805_ ) );
OAI211_X1 _09360_ ( .A(_01805_ ), .B(_01748_ ), .C1(_01749_ ), .C2(\myifu.myicache.tag[1][6] ), .ZN(_01806_ ) );
OR2_X1 _09361_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][6] ), .ZN(_01807_ ) );
OAI211_X1 _09362_ ( .A(_01807_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01749_ ), .C2(\myifu.myicache.tag[3][6] ), .ZN(_01808_ ) );
AND3_X1 _09363_ ( .A1(_01806_ ), .A2(_01808_ ), .A3(\IF_ID_pc [11] ), .ZN(_01809_ ) );
OR2_X4 _09364_ ( .A1(_01743_ ), .A2(\myifu.myicache.tag[1][14] ), .ZN(_01810_ ) );
OAI211_X1 _09365_ ( .A(_01810_ ), .B(_01748_ ), .C1(fanout_net_48 ), .C2(\myifu.myicache.tag[0][14] ), .ZN(_01811_ ) );
OR2_X1 _09366_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][14] ), .ZN(_01812_ ) );
OAI211_X1 _09367_ ( .A(_01812_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01749_ ), .C2(\myifu.myicache.tag[3][14] ), .ZN(_01813_ ) );
AOI21_X1 _09368_ ( .A(\IF_ID_pc [19] ), .B1(_01811_ ), .B2(_01813_ ), .ZN(_01814_ ) );
OR2_X1 _09369_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][23] ), .ZN(_01815_ ) );
OAI211_X1 _09370_ ( .A(_01815_ ), .B(_01755_ ), .C1(_01756_ ), .C2(\myifu.myicache.tag[1][23] ), .ZN(_01816_ ) );
OR2_X1 _09371_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][23] ), .ZN(_01817_ ) );
OAI211_X1 _09372_ ( .A(_01817_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01756_ ), .C2(\myifu.myicache.tag[3][23] ), .ZN(_01818_ ) );
AND3_X1 _09373_ ( .A1(_01816_ ), .A2(_01818_ ), .A3(\IF_ID_pc [28] ), .ZN(_01819_ ) );
AOI21_X1 _09374_ ( .A(\IF_ID_pc [11] ), .B1(_01806_ ), .B2(_01808_ ), .ZN(_01820_ ) );
OR4_X2 _09375_ ( .A1(_01809_ ), .A2(_01814_ ), .A3(_01819_ ), .A4(_01820_ ), .ZN(_01821_ ) );
MUX2_X1 _09376_ ( .A(\myifu.myicache.valid [0] ), .B(\myifu.myicache.valid [1] ), .S(fanout_net_48 ), .Z(_01822_ ) );
MUX2_X1 _09377_ ( .A(\myifu.myicache.valid [2] ), .B(\myifu.myicache.valid [3] ), .S(fanout_net_48 ), .Z(_01823_ ) );
MUX2_X1 _09378_ ( .A(_01822_ ), .B(_01823_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01824_ ) );
NAND3_X1 _09379_ ( .A1(_01811_ ), .A2(_01813_ ), .A3(\IF_ID_pc [19] ), .ZN(_01825_ ) );
OR2_X1 _09380_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[0][21] ), .ZN(_01826_ ) );
OAI211_X1 _09381_ ( .A(_01826_ ), .B(_01748_ ), .C1(_01749_ ), .C2(\myifu.myicache.tag[1][21] ), .ZN(_01827_ ) );
OR2_X1 _09382_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][21] ), .ZN(_01828_ ) );
OAI211_X1 _09383_ ( .A(_01828_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01749_ ), .C2(\myifu.myicache.tag[3][21] ), .ZN(_01829_ ) );
INV_X1 _09384_ ( .A(\IF_ID_pc [26] ), .ZN(_01830_ ) );
AND3_X1 _09385_ ( .A1(_01827_ ), .A2(_01829_ ), .A3(_01830_ ), .ZN(_01831_ ) );
AOI21_X1 _09386_ ( .A(_01830_ ), .B1(_01827_ ), .B2(_01829_ ), .ZN(_01832_ ) );
OAI211_X1 _09387_ ( .A(_01824_ ), .B(_01825_ ), .C1(_01831_ ), .C2(_01832_ ), .ZN(_01833_ ) );
NOR4_X4 _09388_ ( .A1(_01776_ ), .A2(_01804_ ), .A3(_01821_ ), .A4(_01833_ ), .ZN(_01834_ ) );
OR2_X1 _09389_ ( .A1(_01756_ ), .A2(\myifu.myicache.tag[1][5] ), .ZN(_01835_ ) );
OAI211_X1 _09390_ ( .A(_01835_ ), .B(_01748_ ), .C1(fanout_net_48 ), .C2(\myifu.myicache.tag[0][5] ), .ZN(_01836_ ) );
OR2_X1 _09391_ ( .A1(fanout_net_48 ), .A2(\myifu.myicache.tag[2][5] ), .ZN(_01837_ ) );
OAI211_X1 _09392_ ( .A(_01837_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01749_ ), .C2(\myifu.myicache.tag[3][5] ), .ZN(_01838_ ) );
AOI21_X1 _09393_ ( .A(\IF_ID_pc [10] ), .B1(_01836_ ), .B2(_01838_ ), .ZN(_01839_ ) );
MUX2_X1 _09394_ ( .A(\myifu.myicache.tag[0][9] ), .B(\myifu.myicache.tag[1][9] ), .S(fanout_net_48 ), .Z(_01840_ ) );
MUX2_X1 _09395_ ( .A(\myifu.myicache.tag[2][9] ), .B(\myifu.myicache.tag[3][9] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01841_ ) );
MUX2_X1 _09396_ ( .A(_01840_ ), .B(_01841_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01842_ ) );
INV_X1 _09397_ ( .A(_01842_ ), .ZN(_01843_ ) );
AOI21_X1 _09398_ ( .A(_01839_ ), .B1(_01843_ ), .B2(\IF_ID_pc [14] ), .ZN(_01844_ ) );
MUX2_X1 _09399_ ( .A(\myifu.myicache.tag[0][11] ), .B(\myifu.myicache.tag[1][11] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01845_ ) );
MUX2_X1 _09400_ ( .A(\myifu.myicache.tag[2][11] ), .B(\myifu.myicache.tag[3][11] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01846_ ) );
MUX2_X1 _09401_ ( .A(_01845_ ), .B(_01846_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01847_ ) );
INV_X1 _09402_ ( .A(_01847_ ), .ZN(_01848_ ) );
INV_X1 _09403_ ( .A(\IF_ID_pc [12] ), .ZN(_01849_ ) );
OR2_X1 _09404_ ( .A1(_01756_ ), .A2(\myifu.myicache.tag[1][7] ), .ZN(_01850_ ) );
OAI211_X1 _09405_ ( .A(_01850_ ), .B(_01748_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][7] ), .ZN(_01851_ ) );
OR2_X1 _09406_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][7] ), .ZN(_01852_ ) );
OAI211_X1 _09407_ ( .A(_01852_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01749_ ), .C2(\myifu.myicache.tag[3][7] ), .ZN(_01853_ ) );
NAND2_X1 _09408_ ( .A1(_01851_ ), .A2(_01853_ ), .ZN(_01854_ ) );
OAI221_X1 _09409_ ( .A(_01844_ ), .B1(\IF_ID_pc [16] ), .B2(_01848_ ), .C1(_01849_ ), .C2(_01854_ ), .ZN(_01855_ ) );
INV_X1 _09410_ ( .A(\IF_ID_pc [29] ), .ZN(_01856_ ) );
MUX2_X1 _09411_ ( .A(\myifu.myicache.tag[0][24] ), .B(\myifu.myicache.tag[1][24] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01857_ ) );
MUX2_X1 _09412_ ( .A(\myifu.myicache.tag[2][24] ), .B(\myifu.myicache.tag[3][24] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01858_ ) );
MUX2_X1 _09413_ ( .A(_01857_ ), .B(_01858_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01859_ ) );
MUX2_X1 _09414_ ( .A(\myifu.myicache.tag[0][15] ), .B(\myifu.myicache.tag[1][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01860_ ) );
MUX2_X1 _09415_ ( .A(\myifu.myicache.tag[2][15] ), .B(\myifu.myicache.tag[3][15] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01861_ ) );
MUX2_X1 _09416_ ( .A(_01860_ ), .B(_01861_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01862_ ) );
INV_X1 _09417_ ( .A(\IF_ID_pc [20] ), .ZN(_01863_ ) );
AOI22_X1 _09418_ ( .A1(_01856_ ), .A2(_01859_ ), .B1(_01862_ ), .B2(_01863_ ), .ZN(_01864_ ) );
MUX2_X1 _09419_ ( .A(\myifu.myicache.tag[2][2] ), .B(\myifu.myicache.tag[3][2] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01865_ ) );
OR2_X1 _09420_ ( .A1(_01865_ ), .A2(_01748_ ), .ZN(_01866_ ) );
MUX2_X1 _09421_ ( .A(\myifu.myicache.tag[0][2] ), .B(\myifu.myicache.tag[1][2] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01867_ ) );
OR2_X1 _09422_ ( .A1(_01867_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01868_ ) );
INV_X1 _09423_ ( .A(\IF_ID_pc [7] ), .ZN(_01869_ ) );
NAND3_X1 _09424_ ( .A1(_01866_ ), .A2(_01868_ ), .A3(_01869_ ), .ZN(_01870_ ) );
OAI211_X1 _09425_ ( .A(_01864_ ), .B(_01870_ ), .C1(\IF_ID_pc [14] ), .C2(_01843_ ), .ZN(_01871_ ) );
OR2_X1 _09426_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][20] ), .ZN(_01872_ ) );
OAI211_X1 _09427_ ( .A(_01872_ ), .B(_01755_ ), .C1(_01743_ ), .C2(\myifu.myicache.tag[1][20] ), .ZN(_01873_ ) );
OR2_X1 _09428_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][20] ), .ZN(_01874_ ) );
OAI211_X1 _09429_ ( .A(_01874_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01742_ ), .C2(\myifu.myicache.tag[3][20] ), .ZN(_01875_ ) );
NAND3_X1 _09430_ ( .A1(_01873_ ), .A2(_01875_ ), .A3(\IF_ID_pc [25] ), .ZN(_01876_ ) );
OR2_X1 _09431_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[0][3] ), .ZN(_01877_ ) );
OAI211_X1 _09432_ ( .A(_01877_ ), .B(_01755_ ), .C1(_01742_ ), .C2(\myifu.myicache.tag[1][3] ), .ZN(_01878_ ) );
OR2_X1 _09433_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][3] ), .ZN(_01879_ ) );
OAI211_X1 _09434_ ( .A(_01879_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01742_ ), .C2(\myifu.myicache.tag[3][3] ), .ZN(_01880_ ) );
NAND3_X1 _09435_ ( .A1(_01878_ ), .A2(_01880_ ), .A3(\IF_ID_pc [8] ), .ZN(_01881_ ) );
AND2_X1 _09436_ ( .A1(_01876_ ), .A2(_01881_ ), .ZN(_01882_ ) );
INV_X1 _09437_ ( .A(\IF_ID_pc [21] ), .ZN(_01883_ ) );
MUX2_X1 _09438_ ( .A(\myifu.myicache.tag[0][16] ), .B(\myifu.myicache.tag[1][16] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01884_ ) );
MUX2_X1 _09439_ ( .A(\myifu.myicache.tag[2][16] ), .B(\myifu.myicache.tag[3][16] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01885_ ) );
MUX2_X1 _09440_ ( .A(_01884_ ), .B(_01885_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01886_ ) );
OAI221_X1 _09441_ ( .A(_01882_ ), .B1(_01856_ ), .B2(_01859_ ), .C1(_01883_ ), .C2(_01886_ ), .ZN(_01887_ ) );
AOI22_X1 _09442_ ( .A1(_01886_ ), .A2(_01883_ ), .B1(_01854_ ), .B2(_01849_ ), .ZN(_01888_ ) );
INV_X1 _09443_ ( .A(\IF_ID_pc [27] ), .ZN(_01889_ ) );
MUX2_X1 _09444_ ( .A(\myifu.myicache.tag[0][22] ), .B(\myifu.myicache.tag[1][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01890_ ) );
MUX2_X1 _09445_ ( .A(\myifu.myicache.tag[2][22] ), .B(\myifu.myicache.tag[3][22] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01891_ ) );
MUX2_X1 _09446_ ( .A(_01890_ ), .B(_01891_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01892_ ) );
OAI21_X1 _09447_ ( .A(_01888_ ), .B1(_01889_ ), .B2(_01892_ ), .ZN(_01893_ ) );
NOR4_X1 _09448_ ( .A1(_01855_ ), .A2(_01871_ ), .A3(_01887_ ), .A4(_01893_ ), .ZN(_01894_ ) );
AOI21_X1 _09449_ ( .A(\IF_ID_pc [25] ), .B1(_01873_ ), .B2(_01875_ ), .ZN(_01895_ ) );
AOI21_X1 _09450_ ( .A(\IF_ID_pc [8] ), .B1(_01878_ ), .B2(_01880_ ), .ZN(_01896_ ) );
OR2_X2 _09451_ ( .A1(_01895_ ), .A2(_01896_ ), .ZN(_01897_ ) );
INV_X1 _09452_ ( .A(\IF_ID_pc [23] ), .ZN(_01898_ ) );
MUX2_X1 _09453_ ( .A(\myifu.myicache.tag[0][18] ), .B(\myifu.myicache.tag[1][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01899_ ) );
MUX2_X1 _09454_ ( .A(\myifu.myicache.tag[2][18] ), .B(\myifu.myicache.tag[3][18] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01900_ ) );
MUX2_X1 _09455_ ( .A(_01899_ ), .B(_01900_ ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_01901_ ) );
MUX2_X1 _09456_ ( .A(\myifu.myicache.tag[0][13] ), .B(\myifu.myicache.tag[1][13] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01902_ ) );
OR2_X1 _09457_ ( .A1(_01902_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .ZN(_01903_ ) );
MUX2_X1 _09458_ ( .A(\myifu.myicache.tag[2][13] ), .B(\myifu.myicache.tag[3][13] ), .S(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_01904_ ) );
OAI21_X1 _09459_ ( .A(_01903_ ), .B1(_01748_ ), .B2(_01904_ ), .ZN(_01905_ ) );
AOI221_X4 _09460_ ( .A(_01897_ ), .B1(_01898_ ), .B2(_01901_ ), .C1(\IF_ID_pc [18] ), .C2(_01905_ ), .ZN(_01906_ ) );
NOR2_X1 _09461_ ( .A1(_01905_ ), .A2(\IF_ID_pc [18] ), .ZN(_01907_ ) );
OAI22_X1 _09462_ ( .A1(_01898_ ), .A2(_01901_ ), .B1(_01862_ ), .B2(_01863_ ), .ZN(_01908_ ) );
AOI211_X1 _09463_ ( .A(_01907_ ), .B(_01908_ ), .C1(\IF_ID_pc [16] ), .C2(_01848_ ), .ZN(_01909_ ) );
AND2_X1 _09464_ ( .A1(_01892_ ), .A2(_01889_ ), .ZN(_01910_ ) );
AOI21_X1 _09465_ ( .A(\IF_ID_pc [28] ), .B1(_01816_ ), .B2(_01818_ ), .ZN(_01911_ ) );
OR2_X1 _09466_ ( .A1(_01756_ ), .A2(\myifu.myicache.tag[1][19] ), .ZN(_01912_ ) );
OAI211_X1 _09467_ ( .A(_01912_ ), .B(_01748_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][19] ), .ZN(_01913_ ) );
OR2_X1 _09468_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][19] ), .ZN(_01914_ ) );
OAI211_X1 _09469_ ( .A(_01914_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01749_ ), .C2(\myifu.myicache.tag[3][19] ), .ZN(_01915_ ) );
AND3_X1 _09470_ ( .A1(_01913_ ), .A2(_01915_ ), .A3(\IF_ID_pc [24] ), .ZN(_01916_ ) );
AND3_X1 _09471_ ( .A1(_01836_ ), .A2(\IF_ID_pc [10] ), .A3(_01838_ ), .ZN(_01917_ ) );
NOR4_X1 _09472_ ( .A1(_01910_ ), .A2(_01911_ ), .A3(_01916_ ), .A4(_01917_ ), .ZN(_01918_ ) );
AOI21_X1 _09473_ ( .A(_01869_ ), .B1(_01866_ ), .B2(_01868_ ), .ZN(_01919_ ) );
OR2_X1 _09474_ ( .A1(_01756_ ), .A2(\myifu.myicache.tag[1][25] ), .ZN(_01920_ ) );
OAI211_X1 _09475_ ( .A(_01920_ ), .B(_01748_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myifu.myicache.tag[0][25] ), .ZN(_01921_ ) );
OR2_X1 _09476_ ( .A1(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myifu.myicache.tag[2][25] ), .ZN(_01922_ ) );
OAI211_X1 _09477_ ( .A(_01922_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(_01749_ ), .C2(\myifu.myicache.tag[3][25] ), .ZN(_01923_ ) );
AND3_X1 _09478_ ( .A1(_01921_ ), .A2(\IF_ID_pc [30] ), .A3(_01923_ ), .ZN(_01924_ ) );
AOI21_X1 _09479_ ( .A(\IF_ID_pc [24] ), .B1(_01913_ ), .B2(_01915_ ), .ZN(_01925_ ) );
AOI21_X1 _09480_ ( .A(\IF_ID_pc [30] ), .B1(_01921_ ), .B2(_01923_ ), .ZN(_01926_ ) );
NOR4_X1 _09481_ ( .A1(_01919_ ), .A2(_01924_ ), .A3(_01925_ ), .A4(_01926_ ), .ZN(_01927_ ) );
AND4_X4 _09482_ ( .A1(_01906_ ), .A2(_01909_ ), .A3(_01918_ ), .A4(_01927_ ), .ZN(_01928_ ) );
NAND3_X2 _09483_ ( .A1(_01834_ ), .A2(_01894_ ), .A3(_01928_ ), .ZN(_01929_ ) );
AND2_X4 _09484_ ( .A1(_01929_ ), .A2(\myifu.state [0] ), .ZN(_01930_ ) );
INV_X1 _09485_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01931_ ) );
NOR2_X4 _09486_ ( .A1(_01930_ ), .A2(_01931_ ), .ZN(_01932_ ) );
NOR2_X1 _09487_ ( .A1(\myminixbar.state [2] ), .A2(\myminixbar.state [0] ), .ZN(_01933_ ) );
NOR2_X4 _09488_ ( .A1(_01932_ ), .A2(_01933_ ), .ZN(_01934_ ) );
INV_X1 _09489_ ( .A(\EX_LS_flag [2] ), .ZN(_01935_ ) );
NAND4_X1 _09490_ ( .A1(_01935_ ), .A2(\EX_LS_flag [1] ), .A3(\EX_LS_flag [0] ), .A4(EXU_valid_LSU ), .ZN(_01936_ ) );
NOR2_X1 _09491_ ( .A1(_01936_ ), .A2(fanout_net_20 ), .ZN(_01937_ ) );
INV_X1 _09492_ ( .A(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ), .ZN(_01938_ ) );
NOR2_X1 _09493_ ( .A1(_01937_ ), .A2(_01938_ ), .ZN(_01939_ ) );
NOR2_X4 _09494_ ( .A1(_01934_ ), .A2(_01939_ ), .ZN(_01940_ ) );
INV_X1 _09495_ ( .A(EXU_valid_LSU ), .ZN(_01941_ ) );
NOR2_X1 _09496_ ( .A1(_01941_ ), .A2(fanout_net_20 ), .ZN(_01942_ ) );
INV_X1 _09497_ ( .A(\EX_LS_dest_csreg_mem [25] ), .ZN(_01943_ ) );
AND2_X4 _09498_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_01944_ ) );
BUF_X4 _09499_ ( .A(_01935_ ), .Z(_01945_ ) );
NAND4_X1 _09500_ ( .A1(_01942_ ), .A2(_01943_ ), .A3(_01944_ ), .A4(_01945_ ), .ZN(_01946_ ) );
BUF_X4 _09501_ ( .A(_01937_ ), .Z(_01947_ ) );
OAI211_X1 _09502_ ( .A(_01940_ ), .B(_01946_ ), .C1(\mylsu.araddr_tmp [25] ), .C2(_01947_ ), .ZN(_01948_ ) );
INV_X1 _09503_ ( .A(\IF_ID_pc [25] ), .ZN(_01949_ ) );
INV_X2 _09504_ ( .A(_01934_ ), .ZN(_01950_ ) );
OAI21_X1 _09505_ ( .A(_01948_ ), .B1(_01949_ ), .B2(_01950_ ), .ZN(\io_master_araddr [25] ) );
BUF_X4 _09506_ ( .A(_01940_ ), .Z(_01951_ ) );
INV_X1 _09507_ ( .A(\EX_LS_dest_csreg_mem [24] ), .ZN(_01952_ ) );
NAND4_X1 _09508_ ( .A1(_01942_ ), .A2(_01952_ ), .A3(_01944_ ), .A4(_01945_ ), .ZN(_01953_ ) );
OAI211_X1 _09509_ ( .A(_01951_ ), .B(_01953_ ), .C1(\mylsu.araddr_tmp [24] ), .C2(_01947_ ), .ZN(_01954_ ) );
INV_X1 _09510_ ( .A(\IF_ID_pc [24] ), .ZN(_01955_ ) );
BUF_X4 _09511_ ( .A(_01950_ ), .Z(_01956_ ) );
OAI211_X1 _09512_ ( .A(\io_master_araddr [25] ), .B(_01954_ ), .C1(_01955_ ), .C2(_01956_ ), .ZN(_01957_ ) );
CLKBUF_X2 _09513_ ( .A(_01936_ ), .Z(_01958_ ) );
OR3_X1 _09514_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [26] ), .A3(fanout_net_20 ), .ZN(_01959_ ) );
OAI211_X1 _09515_ ( .A(_01951_ ), .B(_01959_ ), .C1(\mylsu.araddr_tmp [26] ), .C2(_01947_ ), .ZN(_01960_ ) );
OAI21_X1 _09516_ ( .A(_01960_ ), .B1(_01830_ ), .B2(_01950_ ), .ZN(\io_master_araddr [26] ) );
INV_X1 _09517_ ( .A(_01939_ ), .ZN(_01961_ ) );
OR3_X1 _09518_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(fanout_net_20 ), .ZN(_01962_ ) );
OAI211_X1 _09519_ ( .A(_01961_ ), .B(_01962_ ), .C1(\mylsu.araddr_tmp [27] ), .C2(_01937_ ), .ZN(_01963_ ) );
CLKBUF_X2 _09520_ ( .A(_01934_ ), .Z(_01964_ ) );
MUX2_X1 _09521_ ( .A(_01963_ ), .B(_01889_ ), .S(_01964_ ), .Z(_01965_ ) );
INV_X1 _09522_ ( .A(_01965_ ), .ZN(\io_master_araddr [27] ) );
OR3_X2 _09523_ ( .A1(_01957_ ), .A2(\io_master_araddr [26] ), .A3(\io_master_araddr [27] ), .ZN(_01966_ ) );
OR3_X1 _09524_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [31] ), .A3(fanout_net_20 ), .ZN(_01967_ ) );
OAI211_X1 _09525_ ( .A(_01951_ ), .B(_01967_ ), .C1(\mylsu.araddr_tmp [31] ), .C2(_01947_ ), .ZN(_01968_ ) );
OAI221_X1 _09526_ ( .A(\IF_ID_pc [31] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01930_ ), .C2(_01931_ ), .ZN(_01969_ ) );
AND2_X1 _09527_ ( .A1(_01968_ ), .A2(_01969_ ), .ZN(_01970_ ) );
INV_X1 _09528_ ( .A(_01970_ ), .ZN(\io_master_araddr [31] ) );
CLKBUF_X2 _09529_ ( .A(_01958_ ), .Z(_01971_ ) );
OR3_X1 _09530_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .A3(fanout_net_20 ), .ZN(_01972_ ) );
BUF_X4 _09531_ ( .A(_01947_ ), .Z(_01973_ ) );
OAI211_X1 _09532_ ( .A(_01951_ ), .B(_01972_ ), .C1(\mylsu.araddr_tmp [28] ), .C2(_01973_ ), .ZN(_01974_ ) );
INV_X1 _09533_ ( .A(\IF_ID_pc [28] ), .ZN(_01975_ ) );
OAI21_X1 _09534_ ( .A(_01974_ ), .B1(_01975_ ), .B2(_01956_ ), .ZN(\io_master_araddr [28] ) );
OR3_X4 _09535_ ( .A1(_01966_ ), .A2(\io_master_araddr [31] ), .A3(\io_master_araddr [28] ), .ZN(_01976_ ) );
OR3_X1 _09536_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [29] ), .A3(fanout_net_20 ), .ZN(_01977_ ) );
OAI211_X1 _09537_ ( .A(_01951_ ), .B(_01977_ ), .C1(\mylsu.araddr_tmp [29] ), .C2(_01947_ ), .ZN(_01978_ ) );
OAI21_X1 _09538_ ( .A(_01978_ ), .B1(_01856_ ), .B2(_01956_ ), .ZN(\io_master_araddr [29] ) );
BUF_X2 _09539_ ( .A(_01951_ ), .Z(_01979_ ) );
OR3_X1 _09540_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [30] ), .A3(fanout_net_20 ), .ZN(_01980_ ) );
OAI211_X1 _09541_ ( .A(_01979_ ), .B(_01980_ ), .C1(\mylsu.araddr_tmp [30] ), .C2(_01973_ ), .ZN(_01981_ ) );
INV_X1 _09542_ ( .A(\IF_ID_pc [30] ), .ZN(_01982_ ) );
OAI21_X1 _09543_ ( .A(_01981_ ), .B1(_01982_ ), .B2(_01956_ ), .ZN(\io_master_araddr [30] ) );
OR3_X4 _09544_ ( .A1(_01976_ ), .A2(\io_master_araddr [29] ), .A3(\io_master_araddr [30] ), .ZN(_01983_ ) );
OR3_X1 _09545_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [18] ), .A3(fanout_net_20 ), .ZN(_01984_ ) );
OAI211_X1 _09546_ ( .A(_01951_ ), .B(_01984_ ), .C1(\mylsu.araddr_tmp [18] ), .C2(_01947_ ), .ZN(_01985_ ) );
INV_X1 _09547_ ( .A(\IF_ID_pc [18] ), .ZN(_01986_ ) );
OAI21_X1 _09548_ ( .A(_01985_ ), .B1(_01986_ ), .B2(_01950_ ), .ZN(\io_master_araddr [18] ) );
OR3_X1 _09549_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [20] ), .A3(fanout_net_20 ), .ZN(_01987_ ) );
OAI211_X1 _09550_ ( .A(_01940_ ), .B(_01987_ ), .C1(\mylsu.araddr_tmp [20] ), .C2(_01947_ ), .ZN(_01988_ ) );
OAI21_X1 _09551_ ( .A(_01988_ ), .B1(_01863_ ), .B2(_01950_ ), .ZN(\io_master_araddr [20] ) );
OR3_X1 _09552_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [17] ), .A3(fanout_net_20 ), .ZN(_01989_ ) );
OAI211_X1 _09553_ ( .A(_01940_ ), .B(_01989_ ), .C1(\mylsu.araddr_tmp [17] ), .C2(_01937_ ), .ZN(_01990_ ) );
OAI21_X1 _09554_ ( .A(_01990_ ), .B1(_01759_ ), .B2(_01950_ ), .ZN(\io_master_araddr [17] ) );
OR3_X1 _09555_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [23] ), .A3(fanout_net_20 ), .ZN(_01991_ ) );
OAI211_X1 _09556_ ( .A(_01940_ ), .B(_01991_ ), .C1(\mylsu.araddr_tmp [23] ), .C2(_01937_ ), .ZN(_01992_ ) );
OAI21_X1 _09557_ ( .A(_01992_ ), .B1(_01898_ ), .B2(_01950_ ), .ZN(\io_master_araddr [23] ) );
OR4_X2 _09558_ ( .A1(\io_master_araddr [18] ), .A2(\io_master_araddr [20] ), .A3(\io_master_araddr [17] ), .A4(\io_master_araddr [23] ), .ZN(_01993_ ) );
OR3_X1 _09559_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [21] ), .A3(fanout_net_20 ), .ZN(_01994_ ) );
OAI211_X1 _09560_ ( .A(_01951_ ), .B(_01994_ ), .C1(\mylsu.araddr_tmp [21] ), .C2(_01947_ ), .ZN(_01995_ ) );
OAI21_X1 _09561_ ( .A(_01995_ ), .B1(_01883_ ), .B2(_01956_ ), .ZN(\io_master_araddr [21] ) );
OR3_X1 _09562_ ( .A1(_01958_ ), .A2(\EX_LS_dest_csreg_mem [22] ), .A3(fanout_net_20 ), .ZN(_01996_ ) );
OAI211_X1 _09563_ ( .A(_01951_ ), .B(_01996_ ), .C1(\mylsu.araddr_tmp [22] ), .C2(_01947_ ), .ZN(_01997_ ) );
OAI21_X1 _09564_ ( .A(_01997_ ), .B1(_01785_ ), .B2(_01956_ ), .ZN(\io_master_araddr [22] ) );
OR3_X1 _09565_ ( .A1(_01993_ ), .A2(\io_master_araddr [21] ), .A3(\io_master_araddr [22] ), .ZN(_01998_ ) );
OR3_X1 _09566_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [19] ), .A3(fanout_net_20 ), .ZN(_01999_ ) );
OAI211_X1 _09567_ ( .A(_01979_ ), .B(_01999_ ), .C1(\mylsu.araddr_tmp [19] ), .C2(_01973_ ), .ZN(_02000_ ) );
INV_X1 _09568_ ( .A(\IF_ID_pc [19] ), .ZN(_02001_ ) );
OAI21_X1 _09569_ ( .A(_02000_ ), .B1(_02001_ ), .B2(_01956_ ), .ZN(\io_master_araddr [19] ) );
OR3_X1 _09570_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [16] ), .A3(fanout_net_20 ), .ZN(_02002_ ) );
OAI211_X1 _09571_ ( .A(_01951_ ), .B(_02002_ ), .C1(\mylsu.araddr_tmp [16] ), .C2(_01973_ ), .ZN(_02003_ ) );
INV_X1 _09572_ ( .A(\IF_ID_pc [16] ), .ZN(_02004_ ) );
OAI21_X1 _09573_ ( .A(_02003_ ), .B1(_02004_ ), .B2(_01956_ ), .ZN(\io_master_araddr [16] ) );
OR3_X4 _09574_ ( .A1(_01998_ ), .A2(\io_master_araddr [19] ), .A3(\io_master_araddr [16] ), .ZN(_02005_ ) );
NOR2_X4 _09575_ ( .A1(_01983_ ), .A2(_02005_ ), .ZN(_02006_ ) );
BUF_X4 _09576_ ( .A(_02006_ ), .Z(_02007_ ) );
BUF_X2 _09577_ ( .A(_02007_ ), .Z(_02008_ ) );
BUF_X2 _09578_ ( .A(_02008_ ), .Z(_02009_ ) );
CLKBUF_X2 _09579_ ( .A(_01964_ ), .Z(_02010_ ) );
CLKBUF_X2 _09580_ ( .A(_02010_ ), .Z(_02011_ ) );
CLKBUF_X2 _09581_ ( .A(_02011_ ), .Z(_02012_ ) );
NAND2_X1 _09582_ ( .A1(_01952_ ), .A2(_01943_ ), .ZN(_02013_ ) );
OR3_X1 _09583_ ( .A1(_02013_ ), .A2(\EX_LS_dest_csreg_mem [27] ), .A3(\EX_LS_dest_csreg_mem [26] ), .ZN(_02014_ ) );
OR4_X1 _09584_ ( .A1(\EX_LS_dest_csreg_mem [31] ), .A2(_02014_ ), .A3(\EX_LS_dest_csreg_mem [30] ), .A4(\EX_LS_dest_csreg_mem [29] ), .ZN(_02015_ ) );
OR2_X1 _09585_ ( .A1(_02015_ ), .A2(\EX_LS_dest_csreg_mem [28] ), .ZN(_02016_ ) );
AND2_X2 _09586_ ( .A1(_01944_ ), .A2(_01945_ ), .ZN(_02017_ ) );
INV_X1 _09587_ ( .A(_02017_ ), .ZN(_02018_ ) );
NOR2_X1 _09588_ ( .A1(_02016_ ), .A2(_02018_ ), .ZN(_02019_ ) );
INV_X1 _09589_ ( .A(\EX_LS_typ [0] ), .ZN(_02020_ ) );
NOR2_X1 _09590_ ( .A1(fanout_net_7 ), .A2(\EX_LS_dest_csreg_mem [1] ), .ZN(_02021_ ) );
INV_X1 _09591_ ( .A(\EX_LS_typ [2] ), .ZN(_02022_ ) );
NOR4_X1 _09592_ ( .A1(_02021_ ), .A2(_02022_ ), .A3(\EX_LS_typ [1] ), .A4(\EX_LS_typ [3] ), .ZN(_02023_ ) );
AND2_X1 _09593_ ( .A1(fanout_net_7 ), .A2(\EX_LS_typ [1] ), .ZN(_02024_ ) );
NOR2_X1 _09594_ ( .A1(\EX_LS_typ [3] ), .A2(\EX_LS_typ [2] ), .ZN(_02025_ ) );
AND2_X1 _09595_ ( .A1(_02024_ ), .A2(_02025_ ), .ZN(_02026_ ) );
OAI21_X1 _09596_ ( .A(_02020_ ), .B1(_02023_ ), .B2(_02026_ ), .ZN(_02027_ ) );
NAND3_X1 _09597_ ( .A1(_02024_ ), .A2(_02025_ ), .A3(\EX_LS_typ [0] ), .ZN(_02028_ ) );
NAND2_X1 _09598_ ( .A1(_02027_ ), .A2(_02028_ ), .ZN(_02029_ ) );
INV_X1 _09599_ ( .A(\EX_LS_typ [4] ), .ZN(_02030_ ) );
AND2_X1 _09600_ ( .A1(_02017_ ), .A2(_02030_ ), .ZN(_02031_ ) );
AND2_X1 _09601_ ( .A1(_02029_ ), .A2(_02031_ ), .ZN(_02032_ ) );
NOR2_X1 _09602_ ( .A1(_02019_ ), .A2(_02032_ ), .ZN(_02033_ ) );
INV_X1 _09603_ ( .A(\EX_LS_flag [1] ), .ZN(_02034_ ) );
NOR2_X1 _09604_ ( .A1(_02034_ ), .A2(\EX_LS_flag [0] ), .ZN(_02035_ ) );
AND2_X2 _09605_ ( .A1(_02035_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02036_ ) );
INV_X1 _09606_ ( .A(_02036_ ), .ZN(_02037_ ) );
NOR2_X1 _09607_ ( .A1(_02016_ ), .A2(_02037_ ), .ZN(_02038_ ) );
NAND3_X1 _09608_ ( .A1(_01945_ ), .A2(_02030_ ), .A3(\EX_LS_typ [0] ), .ZN(_02039_ ) );
NOR3_X1 _09609_ ( .A1(_02039_ ), .A2(_02034_ ), .A3(\EX_LS_flag [0] ), .ZN(_02040_ ) );
INV_X1 _09610_ ( .A(_02040_ ), .ZN(_02041_ ) );
INV_X1 _09611_ ( .A(_02021_ ), .ZN(_02042_ ) );
AND3_X1 _09612_ ( .A1(\EX_LS_typ [1] ), .A2(\EX_LS_typ [3] ), .A3(\EX_LS_typ [2] ), .ZN(_02043_ ) );
AOI22_X1 _09613_ ( .A1(_02042_ ), .A2(_02043_ ), .B1(_02024_ ), .B2(_02025_ ), .ZN(_02044_ ) );
NOR2_X1 _09614_ ( .A1(_02041_ ), .A2(_02044_ ), .ZN(_02045_ ) );
NOR2_X1 _09615_ ( .A1(_02038_ ), .A2(_02045_ ), .ZN(_02046_ ) );
AND2_X1 _09616_ ( .A1(_02033_ ), .A2(_02046_ ), .ZN(_02047_ ) );
AOI211_X1 _09617_ ( .A(_01938_ ), .B(_02012_ ), .C1(_01973_ ), .C2(_02047_ ), .ZN(_02048_ ) );
NOR2_X1 _09618_ ( .A1(fanout_net_2 ), .A2(\myidu.stall_quest_fencei ), .ZN(_02049_ ) );
AND3_X1 _09619_ ( .A1(_01929_ ), .A2(\myifu.state [0] ), .A3(_02049_ ), .ZN(_02050_ ) );
NOR4_X1 _09620_ ( .A1(_01932_ ), .A2(_01931_ ), .A3(_01933_ ), .A4(_02050_ ), .ZN(_02051_ ) );
NOR2_X1 _09621_ ( .A1(_02048_ ), .A2(_02051_ ), .ZN(_02052_ ) );
AND3_X1 _09622_ ( .A1(_02009_ ), .A2(\myclint.rvalid ), .A3(_02052_ ), .ZN(_02053_ ) );
OR4_X1 _09623_ ( .A1(\io_master_araddr [29] ), .A2(\io_master_araddr [26] ), .A3(\io_master_araddr [18] ), .A4(\io_master_araddr [20] ), .ZN(_02054_ ) );
NAND2_X1 _09624_ ( .A1(_01970_ ), .A2(\io_master_araddr [25] ), .ZN(_02055_ ) );
NOR4_X2 _09625_ ( .A1(_02054_ ), .A2(_02055_ ), .A3(\io_master_araddr [27] ), .A4(\io_master_araddr [28] ), .ZN(_02056_ ) );
NOR4_X1 _09626_ ( .A1(\io_master_araddr [17] ), .A2(\io_master_araddr [23] ), .A3(\io_master_araddr [19] ), .A4(\io_master_araddr [21] ), .ZN(_02057_ ) );
OAI21_X1 _09627_ ( .A(_01954_ ), .B1(_01955_ ), .B2(_01956_ ), .ZN(\io_master_araddr [24] ) );
NOR4_X1 _09628_ ( .A1(\io_master_araddr [30] ), .A2(\io_master_araddr [24] ), .A3(\io_master_araddr [16] ), .A4(\io_master_araddr [22] ), .ZN(_02058_ ) );
AND2_X1 _09629_ ( .A1(_02057_ ), .A2(_02058_ ), .ZN(_02059_ ) );
AND2_X2 _09630_ ( .A1(_02056_ ), .A2(_02059_ ), .ZN(_02060_ ) );
INV_X1 _09631_ ( .A(_02060_ ), .ZN(_02061_ ) );
BUF_X2 _09632_ ( .A(_02061_ ), .Z(_02062_ ) );
AOI21_X1 _09633_ ( .A(_02012_ ), .B1(_01973_ ), .B2(_02047_ ), .ZN(_02063_ ) );
AOI211_X1 _09634_ ( .A(_01933_ ), .B(_01932_ ), .C1(\myifu.state [0] ), .C2(_02049_ ), .ZN(_02064_ ) );
NOR3_X1 _09635_ ( .A1(_02062_ ), .A2(_02063_ ), .A3(_02064_ ), .ZN(_02065_ ) );
OAI21_X1 _09636_ ( .A(_01626_ ), .B1(_02065_ ), .B2(\myclint.rvalid ), .ZN(_02066_ ) );
NOR2_X1 _09637_ ( .A1(_02053_ ), .A2(_02066_ ), .ZN(_00065_ ) );
INV_X1 _09638_ ( .A(\LS_WB_wen_csreg [6] ), .ZN(_02067_ ) );
CLKBUF_X2 _09639_ ( .A(_02067_ ), .Z(_02068_ ) );
AND2_X1 _09640_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [5] ), .ZN(_00066_ ) );
INV_X1 _09641_ ( .A(\LS_WB_wdata_csreg [4] ), .ZN(_02069_ ) );
NOR2_X1 _09642_ ( .A1(_02069_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00067_ ) );
AND2_X1 _09643_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [23] ), .ZN(_00068_ ) );
AND2_X1 _09644_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [22] ), .ZN(_00069_ ) );
INV_X1 _09645_ ( .A(\LS_WB_wdata_csreg [21] ), .ZN(_02070_ ) );
NOR2_X1 _09646_ ( .A1(_02070_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00070_ ) );
AND2_X1 _09647_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [20] ), .ZN(_00071_ ) );
AND2_X1 _09648_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [19] ), .ZN(_00072_ ) );
AND2_X1 _09649_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [18] ), .ZN(_00073_ ) );
AND2_X1 _09650_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [17] ), .ZN(_00074_ ) );
AND2_X1 _09651_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [16] ), .ZN(_00075_ ) );
AND2_X1 _09652_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [15] ), .ZN(_00076_ ) );
AND2_X1 _09653_ ( .A1(_02068_ ), .A2(\LS_WB_wdata_csreg [14] ), .ZN(_00077_ ) );
CLKBUF_X2 _09654_ ( .A(_02067_ ), .Z(_02071_ ) );
AND2_X1 _09655_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [31] ), .ZN(_00078_ ) );
AND2_X1 _09656_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [13] ), .ZN(_00079_ ) );
AND2_X1 _09657_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [12] ), .ZN(_00080_ ) );
AND2_X1 _09658_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [11] ), .ZN(_00081_ ) );
AND2_X1 _09659_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [10] ), .ZN(_00082_ ) );
INV_X1 _09660_ ( .A(\LS_WB_wdata_csreg [9] ), .ZN(_02072_ ) );
NOR2_X1 _09661_ ( .A1(_02072_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00083_ ) );
AND2_X1 _09662_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [8] ), .ZN(_00084_ ) );
AND2_X1 _09663_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [7] ), .ZN(_00085_ ) );
INV_X1 _09664_ ( .A(\LS_WB_wdata_csreg [6] ), .ZN(_02073_ ) );
NOR2_X1 _09665_ ( .A1(_02073_ ), .A2(\LS_WB_wen_csreg [6] ), .ZN(_00086_ ) );
AND2_X1 _09666_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [30] ), .ZN(_00087_ ) );
AND2_X1 _09667_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [29] ), .ZN(_00088_ ) );
AND2_X1 _09668_ ( .A1(_02071_ ), .A2(\LS_WB_wdata_csreg [28] ), .ZN(_00089_ ) );
AND2_X1 _09669_ ( .A1(_02067_ ), .A2(\LS_WB_wdata_csreg [27] ), .ZN(_00090_ ) );
AND2_X1 _09670_ ( .A1(_02067_ ), .A2(\LS_WB_wdata_csreg [26] ), .ZN(_00091_ ) );
AND2_X1 _09671_ ( .A1(_02067_ ), .A2(\LS_WB_wdata_csreg [25] ), .ZN(_00092_ ) );
AND2_X1 _09672_ ( .A1(_02067_ ), .A2(\LS_WB_wdata_csreg [24] ), .ZN(_00093_ ) );
INV_X1 _09673_ ( .A(_02033_ ), .ZN(_02074_ ) );
INV_X1 _09674_ ( .A(_02046_ ), .ZN(_02075_ ) );
NOR2_X1 _09675_ ( .A1(\myec.state [0] ), .A2(\myec.state [1] ), .ZN(_02076_ ) );
AND2_X1 _09676_ ( .A1(_02076_ ), .A2(_01456_ ), .ZN(_02077_ ) );
INV_X1 _09677_ ( .A(_02077_ ), .ZN(_02078_ ) );
OR2_X1 _09678_ ( .A1(\myexu.pc_jump [25] ), .A2(\myexu.pc_jump [24] ), .ZN(_02079_ ) );
OR3_X1 _09679_ ( .A1(_02079_ ), .A2(\myexu.pc_jump [27] ), .A3(\myexu.pc_jump [26] ), .ZN(_02080_ ) );
OR4_X1 _09680_ ( .A1(\myexu.pc_jump [31] ), .A2(\myexu.pc_jump [30] ), .A3(\myexu.pc_jump [29] ), .A4(\myexu.pc_jump [28] ), .ZN(_02081_ ) );
NOR2_X1 _09681_ ( .A1(_02080_ ), .A2(_02081_ ), .ZN(_02082_ ) );
NOR2_X1 _09682_ ( .A1(\myexu.pc_jump [0] ), .A2(\myexu.pc_jump [1] ), .ZN(_02083_ ) );
INV_X1 _09683_ ( .A(_02083_ ), .ZN(_02084_ ) );
NOR3_X1 _09684_ ( .A1(_02082_ ), .A2(exception_quest_IDU ), .A3(_02084_ ), .ZN(_02085_ ) );
NOR4_X1 _09685_ ( .A1(_02074_ ), .A2(_02075_ ), .A3(_02078_ ), .A4(_02085_ ), .ZN(_00095_ ) );
AOI21_X1 _09686_ ( .A(_02078_ ), .B1(_02047_ ), .B2(exception_quest_IDU ), .ZN(_00096_ ) );
INV_X1 _09687_ ( .A(fanout_net_34 ), .ZN(_02086_ ) );
BUF_X4 _09688_ ( .A(_02086_ ), .Z(_02087_ ) );
BUF_X4 _09689_ ( .A(_02087_ ), .Z(_02088_ ) );
BUF_X4 _09690_ ( .A(_02088_ ), .Z(_02089_ ) );
INV_X32 _09691_ ( .A(fanout_net_21 ), .ZN(_02090_ ) );
BUF_X2 _09692_ ( .A(_02090_ ), .Z(_02091_ ) );
BUF_X4 _09693_ ( .A(_02091_ ), .Z(_02092_ ) );
CLKBUF_X2 _09694_ ( .A(_02092_ ), .Z(_02093_ ) );
BUF_X4 _09695_ ( .A(_02093_ ), .Z(_02094_ ) );
CLKBUF_X2 _09696_ ( .A(_02094_ ), .Z(_02095_ ) );
CLKBUF_X2 _09697_ ( .A(_02095_ ), .Z(_02096_ ) );
OR2_X1 _09698_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02097_ ) );
INV_X2 _09699_ ( .A(fanout_net_29 ), .ZN(_02098_ ) );
BUF_X4 _09700_ ( .A(_02098_ ), .Z(_02099_ ) );
BUF_X4 _09701_ ( .A(_02099_ ), .Z(_02100_ ) );
BUF_X4 _09702_ ( .A(_02100_ ), .Z(_02101_ ) );
BUF_X4 _09703_ ( .A(_02101_ ), .Z(_02102_ ) );
BUF_X4 _09704_ ( .A(_02102_ ), .Z(_02103_ ) );
BUF_X4 _09705_ ( .A(_02103_ ), .Z(_02104_ ) );
OAI211_X1 _09706_ ( .A(_02097_ ), .B(_02104_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02105_ ) );
OR2_X1 _09707_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02106_ ) );
OAI211_X1 _09708_ ( .A(_02106_ ), .B(fanout_net_29 ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02107_ ) );
NAND3_X1 _09709_ ( .A1(_02105_ ), .A2(_02107_ ), .A3(fanout_net_32 ), .ZN(_02108_ ) );
MUX2_X1 _09710_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02109_ ) );
MUX2_X1 _09711_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02110_ ) );
MUX2_X1 _09712_ ( .A(_02109_ ), .B(_02110_ ), .S(_02104_ ), .Z(_02111_ ) );
OAI211_X1 _09713_ ( .A(_02089_ ), .B(_02108_ ), .C1(_02111_ ), .C2(fanout_net_32 ), .ZN(_02112_ ) );
INV_X1 _09714_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02113_ ) );
AOI21_X1 _09715_ ( .A(fanout_net_29 ), .B1(_02113_ ), .B2(fanout_net_21 ), .ZN(_02114_ ) );
OR2_X1 _09716_ ( .A1(fanout_net_21 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02115_ ) );
MUX2_X1 _09717_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02116_ ) );
AOI221_X4 _09718_ ( .A(fanout_net_32 ), .B1(_02114_ ), .B2(_02115_ ), .C1(_02116_ ), .C2(fanout_net_29 ), .ZN(_02117_ ) );
MUX2_X1 _09719_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02118_ ) );
MUX2_X1 _09720_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02119_ ) );
MUX2_X1 _09721_ ( .A(_02118_ ), .B(_02119_ ), .S(fanout_net_29 ), .Z(_02120_ ) );
INV_X1 _09722_ ( .A(fanout_net_32 ), .ZN(_02121_ ) );
BUF_X4 _09723_ ( .A(_02121_ ), .Z(_02122_ ) );
BUF_X4 _09724_ ( .A(_02122_ ), .Z(_02123_ ) );
BUF_X4 _09725_ ( .A(_02123_ ), .Z(_02124_ ) );
BUF_X4 _09726_ ( .A(_02124_ ), .Z(_02125_ ) );
BUF_X4 _09727_ ( .A(_02125_ ), .Z(_02126_ ) );
OAI21_X1 _09728_ ( .A(fanout_net_34 ), .B1(_02120_ ), .B2(_02126_ ), .ZN(_02127_ ) );
INV_X32 _09729_ ( .A(\ID_EX_rs1 [3] ), .ZN(_02128_ ) );
NAND2_X4 _09730_ ( .A1(_02128_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_02129_ ) );
INV_X16 _09731_ ( .A(\EX_LS_dest_reg [1] ), .ZN(_02130_ ) );
OAI21_X2 _09732_ ( .A(_02129_ ), .B1(\ID_EX_rs1 [1] ), .B2(_02130_ ), .ZN(_02131_ ) );
OR4_X4 _09733_ ( .A1(\EX_LS_dest_reg [3] ), .A2(\EX_LS_dest_reg [2] ), .A3(\EX_LS_dest_reg [1] ), .A4(\EX_LS_dest_reg [0] ), .ZN(_02132_ ) );
NOR2_X4 _09734_ ( .A1(_02132_ ), .A2(\EX_LS_dest_reg [4] ), .ZN(_02133_ ) );
AOI211_X2 _09735_ ( .A(_02131_ ), .B(_02133_ ), .C1(\ID_EX_rs1 [1] ), .C2(_02130_ ), .ZN(_02134_ ) );
INV_X16 _09736_ ( .A(\ID_EX_rs1 [2] ), .ZN(_02135_ ) );
NAND2_X1 _09737_ ( .A1(_02135_ ), .A2(\EX_LS_dest_reg [2] ), .ZN(_02136_ ) );
INV_X16 _09738_ ( .A(\ID_EX_rs1 [4] ), .ZN(_02137_ ) );
OAI21_X1 _09739_ ( .A(_02136_ ), .B1(_02137_ ), .B2(\EX_LS_dest_reg [4] ), .ZN(_02138_ ) );
XOR2_X2 _09740_ ( .A(\ID_EX_rs1 [0] ), .B(\EX_LS_dest_reg [0] ), .Z(_02139_ ) );
NAND2_X1 _09741_ ( .A1(_02137_ ), .A2(\EX_LS_dest_reg [4] ), .ZN(_02140_ ) );
OAI21_X1 _09742_ ( .A(_02140_ ), .B1(_02128_ ), .B2(\EX_LS_dest_reg [3] ), .ZN(_02141_ ) );
OAI21_X1 _09743_ ( .A(\myidu.fc_disenable_$_NOT__A_Y ), .B1(_02135_ ), .B2(\EX_LS_dest_reg [2] ), .ZN(_02142_ ) );
NOR4_X4 _09744_ ( .A1(_02138_ ), .A2(_02139_ ), .A3(_02141_ ), .A4(_02142_ ), .ZN(_02143_ ) );
NAND2_X4 _09745_ ( .A1(_02134_ ), .A2(_02143_ ), .ZN(_02144_ ) );
BUF_X8 _09746_ ( .A(_02144_ ), .Z(_02145_ ) );
BUF_X2 _09747_ ( .A(_02145_ ), .Z(_02146_ ) );
BUF_X2 _09748_ ( .A(_02146_ ), .Z(_02147_ ) );
BUF_X2 _09749_ ( .A(_02147_ ), .Z(_02148_ ) );
NAND3_X1 _09750_ ( .A1(_02034_ ), .A2(\EX_LS_flag [0] ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_02149_ ) );
INV_X2 _09751_ ( .A(_01944_ ), .ZN(_02150_ ) );
OAI21_X1 _09752_ ( .A(_02149_ ), .B1(_02150_ ), .B2(\EX_LS_flag [2] ), .ZN(_02151_ ) );
NOR2_X2 _09753_ ( .A1(\EX_LS_flag [1] ), .A2(\EX_LS_flag [0] ), .ZN(_02152_ ) );
NOR3_X1 _09754_ ( .A1(_01944_ ), .A2(_02152_ ), .A3(_01935_ ), .ZN(_02153_ ) );
NOR2_X2 _09755_ ( .A1(_02151_ ), .A2(_02153_ ), .ZN(_02154_ ) );
BUF_X4 _09756_ ( .A(_02154_ ), .Z(_02155_ ) );
BUF_X2 _09757_ ( .A(_02155_ ), .Z(_02156_ ) );
BUF_X4 _09758_ ( .A(_02156_ ), .Z(_02157_ ) );
BUF_X2 _09759_ ( .A(_02157_ ), .Z(_02158_ ) );
BUF_X2 _09760_ ( .A(_02158_ ), .Z(_02159_ ) );
OAI221_X1 _09761_ ( .A(_02112_ ), .B1(_02117_ ), .B2(_02127_ ), .C1(_02148_ ), .C2(_02159_ ), .ZN(_02160_ ) );
OR3_X1 _09762_ ( .A1(_02147_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02158_ ), .ZN(_02161_ ) );
NAND2_X1 _09763_ ( .A1(_02160_ ), .A2(_02161_ ), .ZN(_02162_ ) );
INV_X1 _09764_ ( .A(\ID_EX_imm [24] ), .ZN(_02163_ ) );
XNOR2_X1 _09765_ ( .A(_02162_ ), .B(_02163_ ), .ZN(_02164_ ) );
OR3_X4 _09766_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02155_ ), .ZN(_02165_ ) );
INV_X1 _09767_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02166_ ) );
NAND2_X1 _09768_ ( .A1(_02166_ ), .A2(fanout_net_21 ), .ZN(_02167_ ) );
OAI211_X1 _09769_ ( .A(_02167_ ), .B(_02099_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02168_ ) );
INV_X1 _09770_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02169_ ) );
NAND2_X1 _09771_ ( .A1(_02169_ ), .A2(fanout_net_21 ), .ZN(_02170_ ) );
OAI211_X1 _09772_ ( .A(_02170_ ), .B(fanout_net_29 ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02171_ ) );
NAND3_X1 _09773_ ( .A1(_02168_ ), .A2(_02171_ ), .A3(fanout_net_32 ), .ZN(_02172_ ) );
MUX2_X1 _09774_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02173_ ) );
MUX2_X1 _09775_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02174_ ) );
MUX2_X1 _09776_ ( .A(_02173_ ), .B(_02174_ ), .S(_02099_ ), .Z(_02175_ ) );
OAI211_X1 _09777_ ( .A(_02087_ ), .B(_02172_ ), .C1(_02175_ ), .C2(fanout_net_32 ), .ZN(_02176_ ) );
NOR2_X1 _09778_ ( .A1(_02092_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02177_ ) );
OAI21_X1 _09779_ ( .A(fanout_net_29 ), .B1(fanout_net_21 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02178_ ) );
INV_X1 _09780_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02179_ ) );
INV_X1 _09781_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02180_ ) );
MUX2_X1 _09782_ ( .A(_02179_ ), .B(_02180_ ), .S(fanout_net_21 ), .Z(_02181_ ) );
OAI221_X1 _09783_ ( .A(_02122_ ), .B1(_02177_ ), .B2(_02178_ ), .C1(_02181_ ), .C2(fanout_net_29 ), .ZN(_02182_ ) );
MUX2_X1 _09784_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02183_ ) );
MUX2_X1 _09785_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02184_ ) );
MUX2_X1 _09786_ ( .A(_02183_ ), .B(_02184_ ), .S(fanout_net_29 ), .Z(_02185_ ) );
OAI211_X1 _09787_ ( .A(fanout_net_34 ), .B(_02182_ ), .C1(_02185_ ), .C2(_02122_ ), .ZN(_02186_ ) );
OAI211_X4 _09788_ ( .A(_02176_ ), .B(_02186_ ), .C1(_02145_ ), .C2(_02155_ ), .ZN(_02187_ ) );
NAND2_X4 _09789_ ( .A1(_02165_ ), .A2(_02187_ ), .ZN(_02188_ ) );
XNOR2_X2 _09790_ ( .A(_02188_ ), .B(\ID_EX_imm [5] ), .ZN(_02189_ ) );
OR3_X4 _09791_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02155_ ), .ZN(_02190_ ) );
OR2_X1 _09792_ ( .A1(_02092_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02191_ ) );
OAI211_X1 _09793_ ( .A(_02191_ ), .B(_02100_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02192_ ) );
OR2_X1 _09794_ ( .A1(_02092_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02193_ ) );
OAI211_X1 _09795_ ( .A(_02193_ ), .B(fanout_net_29 ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02194_ ) );
NAND3_X1 _09796_ ( .A1(_02192_ ), .A2(_02194_ ), .A3(_02122_ ), .ZN(_02195_ ) );
MUX2_X1 _09797_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02196_ ) );
MUX2_X1 _09798_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02197_ ) );
MUX2_X1 _09799_ ( .A(_02196_ ), .B(_02197_ ), .S(_02099_ ), .Z(_02198_ ) );
OAI211_X1 _09800_ ( .A(_02087_ ), .B(_02195_ ), .C1(_02198_ ), .C2(_02122_ ), .ZN(_02199_ ) );
OR2_X1 _09801_ ( .A1(_02092_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02200_ ) );
OAI211_X1 _09802_ ( .A(_02200_ ), .B(fanout_net_29 ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02201_ ) );
OR2_X1 _09803_ ( .A1(_02091_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02202_ ) );
OAI211_X1 _09804_ ( .A(_02202_ ), .B(_02099_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02203_ ) );
NAND3_X1 _09805_ ( .A1(_02201_ ), .A2(_02203_ ), .A3(fanout_net_32 ), .ZN(_02204_ ) );
MUX2_X1 _09806_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02205_ ) );
MUX2_X1 _09807_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_21 ), .Z(_02206_ ) );
MUX2_X1 _09808_ ( .A(_02205_ ), .B(_02206_ ), .S(fanout_net_29 ), .Z(_02207_ ) );
OAI211_X1 _09809_ ( .A(fanout_net_34 ), .B(_02204_ ), .C1(_02207_ ), .C2(fanout_net_32 ), .ZN(_02208_ ) );
OAI211_X1 _09810_ ( .A(_02199_ ), .B(_02208_ ), .C1(_02145_ ), .C2(_02155_ ), .ZN(_02209_ ) );
NAND2_X1 _09811_ ( .A1(_02190_ ), .A2(_02209_ ), .ZN(_02210_ ) );
NAND2_X1 _09812_ ( .A1(_02210_ ), .A2(\ID_EX_imm [4] ), .ZN(_02211_ ) );
OR2_X1 _09813_ ( .A1(_02189_ ), .A2(_02211_ ), .ZN(_02212_ ) );
INV_X1 _09814_ ( .A(_02188_ ), .ZN(_02213_ ) );
OAI21_X4 _09815_ ( .A(_02212_ ), .B1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .B2(_02213_ ), .ZN(_02214_ ) );
OR3_X4 _09816_ ( .A1(_02144_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02154_ ), .ZN(_02215_ ) );
OR2_X1 _09817_ ( .A1(_02090_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02216_ ) );
OAI211_X1 _09818_ ( .A(_02216_ ), .B(_02098_ ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02217_ ) );
OR2_X1 _09819_ ( .A1(_02090_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02218_ ) );
OAI211_X1 _09820_ ( .A(_02218_ ), .B(fanout_net_29 ), .C1(fanout_net_21 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02219_ ) );
NAND3_X1 _09821_ ( .A1(_02217_ ), .A2(_02219_ ), .A3(_02121_ ), .ZN(_02220_ ) );
MUX2_X1 _09822_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02221_ ) );
MUX2_X1 _09823_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02222_ ) );
MUX2_X1 _09824_ ( .A(_02221_ ), .B(_02222_ ), .S(_02098_ ), .Z(_02223_ ) );
OAI211_X1 _09825_ ( .A(_02086_ ), .B(_02220_ ), .C1(_02223_ ), .C2(_02121_ ), .ZN(_02224_ ) );
OR2_X1 _09826_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02225_ ) );
OAI211_X1 _09827_ ( .A(_02225_ ), .B(fanout_net_29 ), .C1(_02091_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02226_ ) );
OR2_X1 _09828_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02227_ ) );
OAI211_X1 _09829_ ( .A(_02227_ ), .B(_02098_ ), .C1(_02091_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02228_ ) );
NAND3_X1 _09830_ ( .A1(_02226_ ), .A2(_02228_ ), .A3(fanout_net_32 ), .ZN(_02229_ ) );
MUX2_X1 _09831_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02230_ ) );
MUX2_X1 _09832_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02231_ ) );
MUX2_X1 _09833_ ( .A(_02230_ ), .B(_02231_ ), .S(fanout_net_29 ), .Z(_02232_ ) );
OAI211_X1 _09834_ ( .A(fanout_net_34 ), .B(_02229_ ), .C1(_02232_ ), .C2(fanout_net_32 ), .ZN(_02233_ ) );
OAI211_X2 _09835_ ( .A(_02224_ ), .B(_02233_ ), .C1(_02144_ ), .C2(_02154_ ), .ZN(_02234_ ) );
NAND2_X4 _09836_ ( .A1(_02215_ ), .A2(_02234_ ), .ZN(_02235_ ) );
INV_X1 _09837_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_02236_ ) );
XNOR2_X2 _09838_ ( .A(_02235_ ), .B(_02236_ ), .ZN(_02237_ ) );
OR3_X4 _09839_ ( .A1(_02144_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02154_ ), .ZN(_02238_ ) );
OR2_X1 _09840_ ( .A1(_02090_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02239_ ) );
OAI211_X1 _09841_ ( .A(_02239_ ), .B(_02098_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02240_ ) );
OR2_X1 _09842_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02241_ ) );
OAI211_X1 _09843_ ( .A(_02241_ ), .B(fanout_net_29 ), .C1(_02091_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02242_ ) );
NAND3_X1 _09844_ ( .A1(_02240_ ), .A2(_02121_ ), .A3(_02242_ ), .ZN(_02243_ ) );
MUX2_X1 _09845_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02244_ ) );
MUX2_X1 _09846_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02245_ ) );
MUX2_X1 _09847_ ( .A(_02244_ ), .B(_02245_ ), .S(_02098_ ), .Z(_02246_ ) );
OAI211_X1 _09848_ ( .A(_02086_ ), .B(_02243_ ), .C1(_02246_ ), .C2(_02121_ ), .ZN(_02247_ ) );
OR2_X1 _09849_ ( .A1(_02090_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02248_ ) );
OAI211_X1 _09850_ ( .A(_02248_ ), .B(_02098_ ), .C1(fanout_net_22 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02249_ ) );
OR2_X1 _09851_ ( .A1(fanout_net_22 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02250_ ) );
OAI211_X1 _09852_ ( .A(_02250_ ), .B(fanout_net_29 ), .C1(_02090_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02251_ ) );
NAND3_X1 _09853_ ( .A1(_02249_ ), .A2(fanout_net_32 ), .A3(_02251_ ), .ZN(_02252_ ) );
MUX2_X1 _09854_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02253_ ) );
MUX2_X1 _09855_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02254_ ) );
MUX2_X1 _09856_ ( .A(_02253_ ), .B(_02254_ ), .S(fanout_net_29 ), .Z(_02255_ ) );
OAI211_X1 _09857_ ( .A(fanout_net_34 ), .B(_02252_ ), .C1(_02255_ ), .C2(fanout_net_32 ), .ZN(_02256_ ) );
OAI211_X2 _09858_ ( .A(_02247_ ), .B(_02256_ ), .C1(_02144_ ), .C2(_02154_ ), .ZN(_02257_ ) );
NAND2_X4 _09859_ ( .A1(_02238_ ), .A2(_02257_ ), .ZN(_02258_ ) );
INV_X1 _09860_ ( .A(\ID_EX_imm [2] ), .ZN(_02259_ ) );
XNOR2_X1 _09861_ ( .A(_02258_ ), .B(_02259_ ), .ZN(_02260_ ) );
INV_X4 _09862_ ( .A(_02260_ ), .ZN(_02261_ ) );
OR3_X2 _09863_ ( .A1(_02144_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02154_ ), .ZN(_02262_ ) );
OR2_X1 _09864_ ( .A1(_02090_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02263_ ) );
OAI211_X1 _09865_ ( .A(_02263_ ), .B(_02099_ ), .C1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .C2(fanout_net_22 ), .ZN(_02264_ ) );
OR2_X1 _09866_ ( .A1(_02090_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02265_ ) );
OAI211_X1 _09867_ ( .A(_02265_ ), .B(fanout_net_29 ), .C1(fanout_net_22 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02266_ ) );
NAND3_X1 _09868_ ( .A1(_02264_ ), .A2(_02266_ ), .A3(_02121_ ), .ZN(_02267_ ) );
MUX2_X1 _09869_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02268_ ) );
MUX2_X1 _09870_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02269_ ) );
MUX2_X1 _09871_ ( .A(_02268_ ), .B(_02269_ ), .S(_02098_ ), .Z(_02270_ ) );
OAI211_X1 _09872_ ( .A(_02086_ ), .B(_02267_ ), .C1(_02270_ ), .C2(_02122_ ), .ZN(_02271_ ) );
OR2_X1 _09873_ ( .A1(_02090_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02272_ ) );
OAI211_X1 _09874_ ( .A(_02272_ ), .B(fanout_net_29 ), .C1(fanout_net_22 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02273_ ) );
OR2_X1 _09875_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02274_ ) );
OAI211_X1 _09876_ ( .A(_02274_ ), .B(_02099_ ), .C1(_02091_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02275_ ) );
NAND3_X1 _09877_ ( .A1(_02273_ ), .A2(fanout_net_32 ), .A3(_02275_ ), .ZN(_02276_ ) );
MUX2_X1 _09878_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02277_ ) );
MUX2_X1 _09879_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02278_ ) );
MUX2_X1 _09880_ ( .A(_02277_ ), .B(_02278_ ), .S(fanout_net_29 ), .Z(_02279_ ) );
OAI211_X1 _09881_ ( .A(fanout_net_34 ), .B(_02276_ ), .C1(_02279_ ), .C2(fanout_net_32 ), .ZN(_02280_ ) );
OAI211_X2 _09882_ ( .A(_02271_ ), .B(_02280_ ), .C1(_02144_ ), .C2(_02154_ ), .ZN(_02281_ ) );
NAND2_X4 _09883_ ( .A1(_02262_ ), .A2(_02281_ ), .ZN(_02282_ ) );
INV_X1 _09884_ ( .A(_02282_ ), .ZN(_02283_ ) );
OR2_X4 _09885_ ( .A1(_02283_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02284_ ) );
INV_X1 _09886_ ( .A(\ID_EX_imm [1] ), .ZN(_02285_ ) );
XNOR2_X2 _09887_ ( .A(_02282_ ), .B(_02285_ ), .ZN(_02286_ ) );
OR2_X1 _09888_ ( .A1(_02091_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02287_ ) );
OAI211_X1 _09889_ ( .A(_02287_ ), .B(_02099_ ), .C1(fanout_net_22 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02288_ ) );
OR2_X1 _09890_ ( .A1(_02091_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02289_ ) );
OAI211_X1 _09891_ ( .A(_02289_ ), .B(fanout_net_29 ), .C1(fanout_net_22 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02290_ ) );
NAND3_X1 _09892_ ( .A1(_02288_ ), .A2(_02290_ ), .A3(_02122_ ), .ZN(_02291_ ) );
MUX2_X1 _09893_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02292_ ) );
MUX2_X1 _09894_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02293_ ) );
MUX2_X1 _09895_ ( .A(_02292_ ), .B(_02293_ ), .S(_02099_ ), .Z(_02294_ ) );
OAI211_X1 _09896_ ( .A(_02086_ ), .B(_02291_ ), .C1(_02294_ ), .C2(_02122_ ), .ZN(_02295_ ) );
OR2_X1 _09897_ ( .A1(_02091_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02296_ ) );
OAI211_X1 _09898_ ( .A(_02296_ ), .B(_02099_ ), .C1(fanout_net_22 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02297_ ) );
OR2_X1 _09899_ ( .A1(fanout_net_22 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02298_ ) );
OAI211_X1 _09900_ ( .A(_02298_ ), .B(fanout_net_29 ), .C1(_02091_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02299_ ) );
NAND3_X1 _09901_ ( .A1(_02297_ ), .A2(fanout_net_32 ), .A3(_02299_ ), .ZN(_02300_ ) );
MUX2_X1 _09902_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02301_ ) );
MUX2_X1 _09903_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_22 ), .Z(_02302_ ) );
MUX2_X1 _09904_ ( .A(_02301_ ), .B(_02302_ ), .S(fanout_net_29 ), .Z(_02303_ ) );
OAI211_X1 _09905_ ( .A(fanout_net_34 ), .B(_02300_ ), .C1(_02303_ ), .C2(fanout_net_32 ), .ZN(_02304_ ) );
NAND2_X1 _09906_ ( .A1(_02295_ ), .A2(_02304_ ), .ZN(_02305_ ) );
OAI21_X4 _09907_ ( .A(_02305_ ), .B1(_02145_ ), .B2(_02155_ ), .ZN(_02306_ ) );
INV_X1 _09908_ ( .A(_02154_ ), .ZN(_02307_ ) );
NAND4_X1 _09909_ ( .A1(_02134_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .A3(_02307_ ), .A4(_02143_ ), .ZN(_02308_ ) );
AND3_X1 _09910_ ( .A1(_02306_ ), .A2(\ID_EX_imm [0] ), .A3(_02308_ ), .ZN(_02309_ ) );
NAND2_X2 _09911_ ( .A1(_02286_ ), .A2(_02309_ ), .ZN(_02310_ ) );
AOI211_X2 _09912_ ( .A(_02237_ ), .B(_02261_ ), .C1(_02284_ ), .C2(_02310_ ), .ZN(_02311_ ) );
AOI21_X1 _09913_ ( .A(_02259_ ), .B1(_02238_ ), .B2(_02257_ ), .ZN(_02312_ ) );
INV_X1 _09914_ ( .A(_02312_ ), .ZN(_02313_ ) );
OR2_X1 _09915_ ( .A1(_02237_ ), .A2(_02313_ ), .ZN(_02314_ ) );
INV_X1 _09916_ ( .A(_02235_ ), .ZN(_02315_ ) );
OAI21_X2 _09917_ ( .A(_02314_ ), .B1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ), .B2(_02315_ ), .ZN(_02316_ ) );
NOR2_X2 _09918_ ( .A1(_02311_ ), .A2(_02316_ ), .ZN(_02317_ ) );
INV_X2 _09919_ ( .A(_02317_ ), .ZN(_02318_ ) );
BUF_X4 _09920_ ( .A(_02210_ ), .Z(_02319_ ) );
INV_X1 _09921_ ( .A(\ID_EX_imm [4] ), .ZN(_02320_ ) );
XNOR2_X1 _09922_ ( .A(_02319_ ), .B(_02320_ ), .ZN(_02321_ ) );
AND2_X4 _09923_ ( .A1(_02318_ ), .A2(_02321_ ), .ZN(_02322_ ) );
INV_X1 _09924_ ( .A(_02189_ ), .ZN(_02323_ ) );
AOI21_X4 _09925_ ( .A(_02214_ ), .B1(_02322_ ), .B2(_02323_ ), .ZN(_02324_ ) );
OR3_X1 _09926_ ( .A1(_02145_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .A3(_02155_ ), .ZN(_02325_ ) );
OR2_X1 _09927_ ( .A1(_02092_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02326_ ) );
OAI211_X1 _09928_ ( .A(_02326_ ), .B(_02100_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02327_ ) );
OR2_X1 _09929_ ( .A1(_02092_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02328_ ) );
OAI211_X1 _09930_ ( .A(_02328_ ), .B(fanout_net_29 ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02329_ ) );
NAND3_X1 _09931_ ( .A1(_02327_ ), .A2(_02329_ ), .A3(_02122_ ), .ZN(_02330_ ) );
MUX2_X1 _09932_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02331_ ) );
MUX2_X1 _09933_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02332_ ) );
MUX2_X1 _09934_ ( .A(_02331_ ), .B(_02332_ ), .S(_02100_ ), .Z(_02333_ ) );
OAI211_X1 _09935_ ( .A(_02087_ ), .B(_02330_ ), .C1(_02333_ ), .C2(_02123_ ), .ZN(_02334_ ) );
OR2_X1 _09936_ ( .A1(_02092_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02335_ ) );
OAI211_X1 _09937_ ( .A(_02335_ ), .B(_02100_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02336_ ) );
OR2_X1 _09938_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02337_ ) );
OAI211_X1 _09939_ ( .A(_02337_ ), .B(fanout_net_29 ), .C1(_02093_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02338_ ) );
NAND3_X1 _09940_ ( .A1(_02336_ ), .A2(fanout_net_32 ), .A3(_02338_ ), .ZN(_02339_ ) );
MUX2_X1 _09941_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02340_ ) );
MUX2_X1 _09942_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02341_ ) );
MUX2_X1 _09943_ ( .A(_02340_ ), .B(_02341_ ), .S(fanout_net_29 ), .Z(_02342_ ) );
OAI211_X1 _09944_ ( .A(fanout_net_34 ), .B(_02339_ ), .C1(_02342_ ), .C2(fanout_net_32 ), .ZN(_02343_ ) );
OAI211_X1 _09945_ ( .A(_02334_ ), .B(_02343_ ), .C1(_02145_ ), .C2(_02155_ ), .ZN(_02344_ ) );
NAND2_X2 _09946_ ( .A1(_02325_ ), .A2(_02344_ ), .ZN(_02345_ ) );
XOR2_X1 _09947_ ( .A(_02345_ ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .Z(_02346_ ) );
BUF_X8 _09948_ ( .A(_02145_ ), .Z(_02347_ ) );
OR3_X4 _09949_ ( .A1(_02347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02156_ ), .ZN(_02348_ ) );
CLKBUF_X3 _09950_ ( .A(_02092_ ), .Z(_02349_ ) );
OR2_X1 _09951_ ( .A1(_02349_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02350_ ) );
OAI211_X1 _09952_ ( .A(_02350_ ), .B(fanout_net_29 ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02351_ ) );
OR2_X1 _09953_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02352_ ) );
BUF_X4 _09954_ ( .A(_02100_ ), .Z(_02353_ ) );
OAI211_X1 _09955_ ( .A(_02352_ ), .B(_02353_ ), .C1(_02094_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02354_ ) );
NAND3_X1 _09956_ ( .A1(_02351_ ), .A2(_02123_ ), .A3(_02354_ ), .ZN(_02355_ ) );
MUX2_X1 _09957_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02356_ ) );
MUX2_X1 _09958_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02357_ ) );
MUX2_X1 _09959_ ( .A(_02356_ ), .B(_02357_ ), .S(_02353_ ), .Z(_02358_ ) );
BUF_X4 _09960_ ( .A(_02123_ ), .Z(_02359_ ) );
OAI211_X1 _09961_ ( .A(fanout_net_34 ), .B(_02355_ ), .C1(_02358_ ), .C2(_02359_ ), .ZN(_02360_ ) );
OR2_X1 _09962_ ( .A1(_02349_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02361_ ) );
OAI211_X1 _09963_ ( .A(_02361_ ), .B(_02101_ ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02362_ ) );
OR2_X1 _09964_ ( .A1(_02093_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02363_ ) );
OAI211_X1 _09965_ ( .A(_02363_ ), .B(fanout_net_29 ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02364_ ) );
NAND3_X1 _09966_ ( .A1(_02362_ ), .A2(_02364_ ), .A3(_02123_ ), .ZN(_02365_ ) );
MUX2_X1 _09967_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02366_ ) );
MUX2_X1 _09968_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02367_ ) );
MUX2_X1 _09969_ ( .A(_02366_ ), .B(_02367_ ), .S(_02353_ ), .Z(_02368_ ) );
OAI211_X1 _09970_ ( .A(_02087_ ), .B(_02365_ ), .C1(_02368_ ), .C2(_02359_ ), .ZN(_02369_ ) );
OAI211_X1 _09971_ ( .A(_02360_ ), .B(_02369_ ), .C1(_02347_ ), .C2(_02156_ ), .ZN(_02370_ ) );
NAND2_X2 _09972_ ( .A1(_02348_ ), .A2(_02370_ ), .ZN(_02371_ ) );
XNOR2_X1 _09973_ ( .A(_02371_ ), .B(\ID_EX_imm [6] ), .ZN(_02372_ ) );
NOR3_X4 _09974_ ( .A1(_02324_ ), .A2(_02346_ ), .A3(_02372_ ), .ZN(_02373_ ) );
NAND2_X1 _09975_ ( .A1(_02371_ ), .A2(\ID_EX_imm [6] ), .ZN(_02374_ ) );
OR2_X1 _09976_ ( .A1(_02346_ ), .A2(_02374_ ), .ZN(_02375_ ) );
INV_X1 _09977_ ( .A(_02345_ ), .ZN(_02376_ ) );
OAI21_X1 _09978_ ( .A(_02375_ ), .B1(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .B2(_02376_ ), .ZN(_02377_ ) );
OR2_X4 _09979_ ( .A1(_02373_ ), .A2(_02377_ ), .ZN(_02378_ ) );
OR3_X1 _09980_ ( .A1(_02145_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02155_ ), .ZN(_02379_ ) );
OR2_X1 _09981_ ( .A1(_02092_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02380_ ) );
OAI211_X1 _09982_ ( .A(_02380_ ), .B(fanout_net_29 ), .C1(fanout_net_23 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02381_ ) );
OR2_X1 _09983_ ( .A1(fanout_net_23 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02382_ ) );
OAI211_X1 _09984_ ( .A(_02382_ ), .B(_02100_ ), .C1(_02349_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02383_ ) );
NAND3_X1 _09985_ ( .A1(_02381_ ), .A2(fanout_net_32 ), .A3(_02383_ ), .ZN(_02384_ ) );
MUX2_X1 _09986_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02385_ ) );
MUX2_X1 _09987_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02386_ ) );
MUX2_X1 _09988_ ( .A(_02385_ ), .B(_02386_ ), .S(_02100_ ), .Z(_02387_ ) );
OAI211_X1 _09989_ ( .A(_02087_ ), .B(_02384_ ), .C1(_02387_ ), .C2(fanout_net_32 ), .ZN(_02388_ ) );
NOR2_X1 _09990_ ( .A1(_02349_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02389_ ) );
OAI21_X1 _09991_ ( .A(fanout_net_30 ), .B1(fanout_net_23 ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02390_ ) );
NOR2_X1 _09992_ ( .A1(fanout_net_23 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02391_ ) );
OAI21_X1 _09993_ ( .A(_02100_ ), .B1(_02349_ ), .B2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02392_ ) );
OAI221_X1 _09994_ ( .A(_02122_ ), .B1(_02389_ ), .B2(_02390_ ), .C1(_02391_ ), .C2(_02392_ ), .ZN(_02393_ ) );
MUX2_X1 _09995_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02394_ ) );
MUX2_X1 _09996_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02395_ ) );
MUX2_X1 _09997_ ( .A(_02394_ ), .B(_02395_ ), .S(fanout_net_30 ), .Z(_02396_ ) );
OAI211_X1 _09998_ ( .A(fanout_net_34 ), .B(_02393_ ), .C1(_02396_ ), .C2(_02123_ ), .ZN(_02397_ ) );
OAI211_X2 _09999_ ( .A(_02388_ ), .B(_02397_ ), .C1(_02347_ ), .C2(_02156_ ), .ZN(_02398_ ) );
NAND2_X4 _10000_ ( .A1(_02379_ ), .A2(_02398_ ), .ZN(_02399_ ) );
XNOR2_X2 _10001_ ( .A(_02399_ ), .B(\ID_EX_imm [11] ), .ZN(_02400_ ) );
OR3_X4 _10002_ ( .A1(_02347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02156_ ), .ZN(_02401_ ) );
OR2_X1 _10003_ ( .A1(_02349_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02402_ ) );
OAI211_X1 _10004_ ( .A(_02402_ ), .B(fanout_net_30 ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02403_ ) );
OR2_X1 _10005_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02404_ ) );
CLKBUF_X2 _10006_ ( .A(_02093_ ), .Z(_02405_ ) );
OAI211_X1 _10007_ ( .A(_02404_ ), .B(_02101_ ), .C1(_02405_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02406_ ) );
NAND3_X1 _10008_ ( .A1(_02403_ ), .A2(_02123_ ), .A3(_02406_ ), .ZN(_02407_ ) );
MUX2_X1 _10009_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02408_ ) );
MUX2_X1 _10010_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_23 ), .Z(_02409_ ) );
MUX2_X1 _10011_ ( .A(_02408_ ), .B(_02409_ ), .S(_02353_ ), .Z(_02410_ ) );
OAI211_X1 _10012_ ( .A(_02087_ ), .B(_02407_ ), .C1(_02410_ ), .C2(_02359_ ), .ZN(_02411_ ) );
OR2_X1 _10013_ ( .A1(_02349_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02412_ ) );
OAI211_X1 _10014_ ( .A(_02412_ ), .B(fanout_net_30 ), .C1(fanout_net_23 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02413_ ) );
OR2_X1 _10015_ ( .A1(fanout_net_23 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02414_ ) );
OAI211_X1 _10016_ ( .A(_02414_ ), .B(_02101_ ), .C1(_02405_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02415_ ) );
NAND3_X1 _10017_ ( .A1(_02413_ ), .A2(fanout_net_32 ), .A3(_02415_ ), .ZN(_02416_ ) );
MUX2_X1 _10018_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02417_ ) );
MUX2_X1 _10019_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02418_ ) );
MUX2_X1 _10020_ ( .A(_02417_ ), .B(_02418_ ), .S(fanout_net_30 ), .Z(_02419_ ) );
OAI211_X1 _10021_ ( .A(fanout_net_34 ), .B(_02416_ ), .C1(_02419_ ), .C2(fanout_net_32 ), .ZN(_02420_ ) );
OAI211_X1 _10022_ ( .A(_02411_ ), .B(_02420_ ), .C1(_02347_ ), .C2(_02156_ ), .ZN(_02421_ ) );
NAND2_X2 _10023_ ( .A1(_02401_ ), .A2(_02421_ ), .ZN(_02422_ ) );
XNOR2_X1 _10024_ ( .A(_02422_ ), .B(\ID_EX_imm [10] ), .ZN(_02423_ ) );
NOR2_X2 _10025_ ( .A1(_02400_ ), .A2(_02423_ ), .ZN(_02424_ ) );
OR3_X1 _10026_ ( .A1(_02146_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02156_ ), .ZN(_02425_ ) );
OR2_X1 _10027_ ( .A1(_02094_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02426_ ) );
BUF_X4 _10028_ ( .A(_02353_ ), .Z(_02427_ ) );
OAI211_X1 _10029_ ( .A(_02426_ ), .B(_02427_ ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02428_ ) );
OR2_X1 _10030_ ( .A1(fanout_net_24 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02429_ ) );
CLKBUF_X2 _10031_ ( .A(_02349_ ), .Z(_02430_ ) );
OAI211_X1 _10032_ ( .A(_02429_ ), .B(fanout_net_30 ), .C1(_02430_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02431_ ) );
NAND3_X1 _10033_ ( .A1(_02428_ ), .A2(_02359_ ), .A3(_02431_ ), .ZN(_02432_ ) );
MUX2_X1 _10034_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02433_ ) );
MUX2_X1 _10035_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02434_ ) );
MUX2_X1 _10036_ ( .A(_02433_ ), .B(_02434_ ), .S(_02101_ ), .Z(_02435_ ) );
OAI211_X1 _10037_ ( .A(_02088_ ), .B(_02432_ ), .C1(_02435_ ), .C2(_02124_ ), .ZN(_02436_ ) );
OR2_X1 _10038_ ( .A1(_02094_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02437_ ) );
OAI211_X1 _10039_ ( .A(_02437_ ), .B(_02427_ ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02438_ ) );
OR2_X1 _10040_ ( .A1(fanout_net_24 ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02439_ ) );
BUF_X2 _10041_ ( .A(_02349_ ), .Z(_02440_ ) );
OAI211_X1 _10042_ ( .A(_02439_ ), .B(fanout_net_30 ), .C1(_02440_ ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02441_ ) );
NAND3_X1 _10043_ ( .A1(_02438_ ), .A2(fanout_net_32 ), .A3(_02441_ ), .ZN(_02442_ ) );
MUX2_X1 _10044_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02443_ ) );
MUX2_X1 _10045_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02444_ ) );
MUX2_X1 _10046_ ( .A(_02443_ ), .B(_02444_ ), .S(fanout_net_30 ), .Z(_02445_ ) );
OAI211_X1 _10047_ ( .A(fanout_net_34 ), .B(_02442_ ), .C1(_02445_ ), .C2(fanout_net_32 ), .ZN(_02446_ ) );
OAI211_X1 _10048_ ( .A(_02436_ ), .B(_02446_ ), .C1(_02146_ ), .C2(_02157_ ), .ZN(_02447_ ) );
NAND2_X2 _10049_ ( .A1(_02425_ ), .A2(_02447_ ), .ZN(_02448_ ) );
INV_X1 _10050_ ( .A(\ID_EX_imm [8] ), .ZN(_02449_ ) );
XNOR2_X1 _10051_ ( .A(_02448_ ), .B(_02449_ ), .ZN(_02450_ ) );
INV_X1 _10052_ ( .A(_02450_ ), .ZN(_02451_ ) );
OR3_X4 _10053_ ( .A1(_02347_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02155_ ), .ZN(_02452_ ) );
OR2_X1 _10054_ ( .A1(_02093_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02453_ ) );
OAI211_X1 _10055_ ( .A(_02453_ ), .B(_02353_ ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02454_ ) );
OR2_X1 _10056_ ( .A1(_02093_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02455_ ) );
OAI211_X1 _10057_ ( .A(_02455_ ), .B(fanout_net_30 ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02456_ ) );
NAND3_X1 _10058_ ( .A1(_02454_ ), .A2(_02456_ ), .A3(_02123_ ), .ZN(_02457_ ) );
MUX2_X1 _10059_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02458_ ) );
MUX2_X1 _10060_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02459_ ) );
MUX2_X1 _10061_ ( .A(_02458_ ), .B(_02459_ ), .S(_02353_ ), .Z(_02460_ ) );
OAI211_X1 _10062_ ( .A(_02087_ ), .B(_02457_ ), .C1(_02460_ ), .C2(_02359_ ), .ZN(_02461_ ) );
OR2_X1 _10063_ ( .A1(_02093_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02462_ ) );
OAI211_X1 _10064_ ( .A(_02462_ ), .B(fanout_net_30 ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02463_ ) );
OR2_X1 _10065_ ( .A1(_02093_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02464_ ) );
OAI211_X1 _10066_ ( .A(_02464_ ), .B(_02353_ ), .C1(fanout_net_24 ), .C2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02465_ ) );
NAND3_X1 _10067_ ( .A1(_02463_ ), .A2(_02465_ ), .A3(fanout_net_32 ), .ZN(_02466_ ) );
MUX2_X1 _10068_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02467_ ) );
MUX2_X1 _10069_ ( .A(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02468_ ) );
MUX2_X1 _10070_ ( .A(_02467_ ), .B(_02468_ ), .S(fanout_net_30 ), .Z(_02469_ ) );
OAI211_X1 _10071_ ( .A(fanout_net_34 ), .B(_02466_ ), .C1(_02469_ ), .C2(fanout_net_32 ), .ZN(_02470_ ) );
OAI211_X1 _10072_ ( .A(_02461_ ), .B(_02470_ ), .C1(_02347_ ), .C2(_02156_ ), .ZN(_02471_ ) );
NAND2_X2 _10073_ ( .A1(_02452_ ), .A2(_02471_ ), .ZN(_02472_ ) );
XNOR2_X2 _10074_ ( .A(_02472_ ), .B(\ID_EX_imm [9] ), .ZN(_02473_ ) );
NOR2_X1 _10075_ ( .A1(_02451_ ), .A2(_02473_ ), .ZN(_02474_ ) );
NAND3_X4 _10076_ ( .A1(_02378_ ), .A2(_02424_ ), .A3(_02474_ ), .ZN(_02475_ ) );
OR3_X1 _10077_ ( .A1(_02146_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02157_ ), .ZN(_02476_ ) );
OR2_X1 _10078_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02477_ ) );
OAI211_X1 _10079_ ( .A(_02477_ ), .B(_02427_ ), .C1(_02430_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02478_ ) );
OR2_X1 _10080_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02479_ ) );
OAI211_X1 _10081_ ( .A(_02479_ ), .B(fanout_net_30 ), .C1(_02430_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02480_ ) );
NAND3_X1 _10082_ ( .A1(_02478_ ), .A2(_02480_ ), .A3(fanout_net_32 ), .ZN(_02481_ ) );
MUX2_X1 _10083_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02482_ ) );
MUX2_X1 _10084_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02483_ ) );
MUX2_X1 _10085_ ( .A(_02482_ ), .B(_02483_ ), .S(_02427_ ), .Z(_02484_ ) );
OAI211_X1 _10086_ ( .A(_02088_ ), .B(_02481_ ), .C1(_02484_ ), .C2(fanout_net_32 ), .ZN(_02485_ ) );
NOR2_X1 _10087_ ( .A1(_02440_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02486_ ) );
OAI21_X1 _10088_ ( .A(fanout_net_30 ), .B1(fanout_net_24 ), .B2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02487_ ) );
NOR2_X1 _10089_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02488_ ) );
OAI21_X1 _10090_ ( .A(_02101_ ), .B1(_02440_ ), .B2(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02489_ ) );
OAI221_X1 _10091_ ( .A(_02359_ ), .B1(_02486_ ), .B2(_02487_ ), .C1(_02488_ ), .C2(_02489_ ), .ZN(_02490_ ) );
MUX2_X1 _10092_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02491_ ) );
MUX2_X1 _10093_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02492_ ) );
MUX2_X1 _10094_ ( .A(_02491_ ), .B(_02492_ ), .S(fanout_net_30 ), .Z(_02493_ ) );
OAI211_X1 _10095_ ( .A(fanout_net_34 ), .B(_02490_ ), .C1(_02493_ ), .C2(_02124_ ), .ZN(_02494_ ) );
OAI211_X1 _10096_ ( .A(_02485_ ), .B(_02494_ ), .C1(_02146_ ), .C2(_02157_ ), .ZN(_02495_ ) );
NAND2_X1 _10097_ ( .A1(_02476_ ), .A2(_02495_ ), .ZN(_02496_ ) );
XNOR2_X1 _10098_ ( .A(_02496_ ), .B(\ID_EX_imm [14] ), .ZN(_02497_ ) );
OR3_X1 _10099_ ( .A1(_02347_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02156_ ), .ZN(_02498_ ) );
OR2_X1 _10100_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02499_ ) );
OAI211_X1 _10101_ ( .A(_02499_ ), .B(_02101_ ), .C1(_02440_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02500_ ) );
OR2_X1 _10102_ ( .A1(fanout_net_24 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02501_ ) );
OAI211_X1 _10103_ ( .A(_02501_ ), .B(fanout_net_30 ), .C1(_02440_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02502_ ) );
NAND3_X1 _10104_ ( .A1(_02500_ ), .A2(_02502_ ), .A3(_02359_ ), .ZN(_02503_ ) );
MUX2_X1 _10105_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02504_ ) );
MUX2_X1 _10106_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_24 ), .Z(_02505_ ) );
MUX2_X1 _10107_ ( .A(_02504_ ), .B(_02505_ ), .S(_02101_ ), .Z(_02506_ ) );
OAI211_X1 _10108_ ( .A(_02087_ ), .B(_02503_ ), .C1(_02506_ ), .C2(_02359_ ), .ZN(_02507_ ) );
OR2_X1 _10109_ ( .A1(_02349_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02508_ ) );
OAI211_X1 _10110_ ( .A(_02508_ ), .B(fanout_net_30 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02509_ ) );
OR2_X1 _10111_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02510_ ) );
OAI211_X1 _10112_ ( .A(_02510_ ), .B(_02101_ ), .C1(_02440_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02511_ ) );
NAND3_X1 _10113_ ( .A1(_02509_ ), .A2(fanout_net_32 ), .A3(_02511_ ), .ZN(_02512_ ) );
MUX2_X1 _10114_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02513_ ) );
MUX2_X1 _10115_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02514_ ) );
MUX2_X1 _10116_ ( .A(_02513_ ), .B(_02514_ ), .S(fanout_net_30 ), .Z(_02515_ ) );
OAI211_X1 _10117_ ( .A(fanout_net_34 ), .B(_02512_ ), .C1(_02515_ ), .C2(fanout_net_32 ), .ZN(_02516_ ) );
OAI211_X1 _10118_ ( .A(_02507_ ), .B(_02516_ ), .C1(_02146_ ), .C2(_02157_ ), .ZN(_02517_ ) );
NAND2_X2 _10119_ ( .A1(_02498_ ), .A2(_02517_ ), .ZN(_02518_ ) );
XNOR2_X1 _10120_ ( .A(_02518_ ), .B(\ID_EX_imm [15] ), .ZN(_02519_ ) );
NOR2_X1 _10121_ ( .A1(_02497_ ), .A2(_02519_ ), .ZN(_02520_ ) );
OR3_X1 _10122_ ( .A1(_02146_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02157_ ), .ZN(_02521_ ) );
OR2_X1 _10123_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02522_ ) );
OAI211_X1 _10124_ ( .A(_02522_ ), .B(_02102_ ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02523_ ) );
OR2_X1 _10125_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02524_ ) );
OAI211_X1 _10126_ ( .A(_02524_ ), .B(fanout_net_30 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02525_ ) );
NAND3_X1 _10127_ ( .A1(_02523_ ), .A2(_02525_ ), .A3(_02124_ ), .ZN(_02526_ ) );
MUX2_X1 _10128_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02527_ ) );
MUX2_X1 _10129_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02528_ ) );
MUX2_X1 _10130_ ( .A(_02527_ ), .B(_02528_ ), .S(_02427_ ), .Z(_02529_ ) );
OAI211_X1 _10131_ ( .A(_02088_ ), .B(_02526_ ), .C1(_02529_ ), .C2(_02124_ ), .ZN(_02530_ ) );
OR2_X1 _10132_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02531_ ) );
OAI211_X1 _10133_ ( .A(_02531_ ), .B(_02427_ ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02532_ ) );
OR2_X1 _10134_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02533_ ) );
OAI211_X1 _10135_ ( .A(_02533_ ), .B(fanout_net_30 ), .C1(_02430_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02534_ ) );
NAND3_X1 _10136_ ( .A1(_02532_ ), .A2(fanout_net_33 ), .A3(_02534_ ), .ZN(_02535_ ) );
MUX2_X1 _10137_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02536_ ) );
MUX2_X1 _10138_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02537_ ) );
MUX2_X1 _10139_ ( .A(_02536_ ), .B(_02537_ ), .S(fanout_net_30 ), .Z(_02538_ ) );
OAI211_X1 _10140_ ( .A(fanout_net_34 ), .B(_02535_ ), .C1(_02538_ ), .C2(fanout_net_33 ), .ZN(_02539_ ) );
BUF_X4 _10141_ ( .A(_02347_ ), .Z(_02540_ ) );
BUF_X2 _10142_ ( .A(_02156_ ), .Z(_02541_ ) );
OAI211_X1 _10143_ ( .A(_02530_ ), .B(_02539_ ), .C1(_02540_ ), .C2(_02541_ ), .ZN(_02542_ ) );
NAND2_X1 _10144_ ( .A1(_02521_ ), .A2(_02542_ ), .ZN(_02543_ ) );
XNOR2_X1 _10145_ ( .A(_02543_ ), .B(\ID_EX_imm [12] ), .ZN(_02544_ ) );
OR3_X1 _10146_ ( .A1(_02146_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02157_ ), .ZN(_02545_ ) );
OR2_X1 _10147_ ( .A1(_02094_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02546_ ) );
OAI211_X1 _10148_ ( .A(_02546_ ), .B(_02427_ ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02547_ ) );
OR2_X1 _10149_ ( .A1(_02094_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02548_ ) );
OAI211_X1 _10150_ ( .A(_02548_ ), .B(fanout_net_30 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02549_ ) );
NAND3_X1 _10151_ ( .A1(_02547_ ), .A2(_02549_ ), .A3(_02359_ ), .ZN(_02550_ ) );
MUX2_X1 _10152_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02551_ ) );
MUX2_X1 _10153_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02552_ ) );
MUX2_X1 _10154_ ( .A(_02551_ ), .B(_02552_ ), .S(_02427_ ), .Z(_02553_ ) );
OAI211_X1 _10155_ ( .A(_02088_ ), .B(_02550_ ), .C1(_02553_ ), .C2(_02124_ ), .ZN(_02554_ ) );
OR2_X1 _10156_ ( .A1(_02094_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02555_ ) );
OAI211_X1 _10157_ ( .A(_02555_ ), .B(fanout_net_30 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02556_ ) );
OR2_X1 _10158_ ( .A1(_02094_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02557_ ) );
OAI211_X1 _10159_ ( .A(_02557_ ), .B(_02427_ ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02558_ ) );
NAND3_X1 _10160_ ( .A1(_02556_ ), .A2(_02558_ ), .A3(fanout_net_33 ), .ZN(_02559_ ) );
MUX2_X1 _10161_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02560_ ) );
MUX2_X1 _10162_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02561_ ) );
MUX2_X1 _10163_ ( .A(_02560_ ), .B(_02561_ ), .S(fanout_net_30 ), .Z(_02562_ ) );
OAI211_X1 _10164_ ( .A(fanout_net_34 ), .B(_02559_ ), .C1(_02562_ ), .C2(fanout_net_33 ), .ZN(_02563_ ) );
OAI211_X1 _10165_ ( .A(_02554_ ), .B(_02563_ ), .C1(_02146_ ), .C2(_02541_ ), .ZN(_02564_ ) );
NAND2_X1 _10166_ ( .A1(_02545_ ), .A2(_02564_ ), .ZN(_02565_ ) );
NAND2_X1 _10167_ ( .A1(_02565_ ), .A2(\ID_EX_imm [13] ), .ZN(_02566_ ) );
INV_X1 _10168_ ( .A(\ID_EX_imm [13] ), .ZN(_02567_ ) );
NAND3_X1 _10169_ ( .A1(_02545_ ), .A2(_02564_ ), .A3(_02567_ ), .ZN(_02568_ ) );
NAND2_X1 _10170_ ( .A1(_02566_ ), .A2(_02568_ ), .ZN(_02569_ ) );
NOR2_X1 _10171_ ( .A1(_02544_ ), .A2(_02569_ ), .ZN(_02570_ ) );
NAND2_X1 _10172_ ( .A1(_02520_ ), .A2(_02570_ ), .ZN(_02571_ ) );
OR2_X4 _10173_ ( .A1(_02475_ ), .A2(_02571_ ), .ZN(_02572_ ) );
INV_X1 _10174_ ( .A(\ID_EX_imm [10] ), .ZN(_02573_ ) );
INV_X1 _10175_ ( .A(_02422_ ), .ZN(_02574_ ) );
OR3_X2 _10176_ ( .A1(_02400_ ), .A2(_02573_ ), .A3(_02574_ ), .ZN(_02575_ ) );
INV_X1 _10177_ ( .A(\ID_EX_imm [11] ), .ZN(_02576_ ) );
INV_X1 _10178_ ( .A(_02399_ ), .ZN(_02577_ ) );
OAI21_X1 _10179_ ( .A(_02575_ ), .B1(_02576_ ), .B2(_02577_ ), .ZN(_02578_ ) );
NAND2_X1 _10180_ ( .A1(_02448_ ), .A2(\ID_EX_imm [8] ), .ZN(_02579_ ) );
OR2_X4 _10181_ ( .A1(_02473_ ), .A2(_02579_ ), .ZN(_02580_ ) );
INV_X1 _10182_ ( .A(\ID_EX_imm [9] ), .ZN(_02581_ ) );
INV_X1 _10183_ ( .A(_02472_ ), .ZN(_02582_ ) );
OAI21_X1 _10184_ ( .A(_02580_ ), .B1(_02581_ ), .B2(_02582_ ), .ZN(_02583_ ) );
AOI21_X1 _10185_ ( .A(_02578_ ), .B1(_02583_ ), .B2(_02424_ ), .ZN(_02584_ ) );
NOR2_X1 _10186_ ( .A1(_02584_ ), .A2(_02571_ ), .ZN(_02585_ ) );
INV_X1 _10187_ ( .A(\ID_EX_imm [15] ), .ZN(_02586_ ) );
AOI21_X1 _10188_ ( .A(_02586_ ), .B1(_02498_ ), .B2(_02517_ ), .ZN(_02587_ ) );
BUF_X4 _10189_ ( .A(_02543_ ), .Z(_02588_ ) );
NAND2_X1 _10190_ ( .A1(_02588_ ), .A2(\ID_EX_imm [12] ), .ZN(_02589_ ) );
NAND2_X1 _10191_ ( .A1(_02589_ ), .A2(_02566_ ), .ZN(_02590_ ) );
AND3_X1 _10192_ ( .A1(_02520_ ), .A2(_02568_ ), .A3(_02590_ ), .ZN(_02591_ ) );
BUF_X4 _10193_ ( .A(_02496_ ), .Z(_02592_ ) );
NAND2_X1 _10194_ ( .A1(_02592_ ), .A2(\ID_EX_imm [14] ), .ZN(_02593_ ) );
NOR2_X1 _10195_ ( .A1(_02519_ ), .A2(_02593_ ), .ZN(_02594_ ) );
NOR4_X4 _10196_ ( .A1(_02585_ ), .A2(_02587_ ), .A3(_02591_ ), .A4(_02594_ ), .ZN(_02595_ ) );
NAND2_X4 _10197_ ( .A1(_02572_ ), .A2(_02595_ ), .ZN(_02596_ ) );
OR3_X1 _10198_ ( .A1(_02540_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02157_ ), .ZN(_02597_ ) );
OR2_X1 _10199_ ( .A1(_02440_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02598_ ) );
OAI211_X1 _10200_ ( .A(_02598_ ), .B(_02102_ ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02599_ ) );
OR2_X1 _10201_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02600_ ) );
OAI211_X1 _10202_ ( .A(_02600_ ), .B(fanout_net_30 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02601_ ) );
NAND3_X1 _10203_ ( .A1(_02599_ ), .A2(_02601_ ), .A3(_02124_ ), .ZN(_02602_ ) );
MUX2_X1 _10204_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02603_ ) );
MUX2_X1 _10205_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02604_ ) );
MUX2_X1 _10206_ ( .A(_02603_ ), .B(_02604_ ), .S(_02102_ ), .Z(_02605_ ) );
BUF_X4 _10207_ ( .A(_02359_ ), .Z(_02606_ ) );
OAI211_X1 _10208_ ( .A(_02088_ ), .B(_02602_ ), .C1(_02605_ ), .C2(_02606_ ), .ZN(_02607_ ) );
OR2_X1 _10209_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02608_ ) );
OAI211_X1 _10210_ ( .A(_02608_ ), .B(fanout_net_30 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02609_ ) );
OR2_X1 _10211_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02610_ ) );
OAI211_X1 _10212_ ( .A(_02610_ ), .B(_02102_ ), .C1(_02095_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02611_ ) );
NAND3_X1 _10213_ ( .A1(_02609_ ), .A2(fanout_net_33 ), .A3(_02611_ ), .ZN(_02612_ ) );
MUX2_X1 _10214_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02613_ ) );
MUX2_X1 _10215_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_25 ), .Z(_02614_ ) );
MUX2_X1 _10216_ ( .A(_02613_ ), .B(_02614_ ), .S(fanout_net_30 ), .Z(_02615_ ) );
OAI211_X1 _10217_ ( .A(fanout_net_34 ), .B(_02612_ ), .C1(_02615_ ), .C2(fanout_net_33 ), .ZN(_02616_ ) );
OAI211_X1 _10218_ ( .A(_02607_ ), .B(_02616_ ), .C1(_02540_ ), .C2(_02541_ ), .ZN(_02617_ ) );
NAND2_X4 _10219_ ( .A1(_02597_ ), .A2(_02617_ ), .ZN(_02618_ ) );
INV_X1 _10220_ ( .A(\ID_EX_imm [19] ), .ZN(_02619_ ) );
XNOR2_X1 _10221_ ( .A(_02618_ ), .B(_02619_ ), .ZN(_02620_ ) );
OR2_X1 _10222_ ( .A1(_02430_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02621_ ) );
OAI211_X1 _10223_ ( .A(_02621_ ), .B(fanout_net_30 ), .C1(fanout_net_25 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02622_ ) );
OR2_X1 _10224_ ( .A1(fanout_net_25 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02623_ ) );
BUF_X4 _10225_ ( .A(_02101_ ), .Z(_02624_ ) );
CLKBUF_X2 _10226_ ( .A(_02440_ ), .Z(_02625_ ) );
OAI211_X1 _10227_ ( .A(_02623_ ), .B(_02624_ ), .C1(_02625_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02626_ ) );
NAND3_X1 _10228_ ( .A1(_02622_ ), .A2(_02606_ ), .A3(_02626_ ), .ZN(_02627_ ) );
MUX2_X1 _10229_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02628_ ) );
MUX2_X1 _10230_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02629_ ) );
MUX2_X1 _10231_ ( .A(_02628_ ), .B(_02629_ ), .S(_02624_ ), .Z(_02630_ ) );
OAI211_X1 _10232_ ( .A(fanout_net_34 ), .B(_02627_ ), .C1(_02630_ ), .C2(_02125_ ), .ZN(_02631_ ) );
MUX2_X1 _10233_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02632_ ) );
AND2_X1 _10234_ ( .A1(_02632_ ), .A2(fanout_net_30 ), .ZN(_02633_ ) );
MUX2_X1 _10235_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02634_ ) );
AOI211_X1 _10236_ ( .A(fanout_net_33 ), .B(_02633_ ), .C1(_02103_ ), .C2(_02634_ ), .ZN(_02635_ ) );
MUX2_X1 _10237_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02636_ ) );
MUX2_X1 _10238_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02637_ ) );
MUX2_X1 _10239_ ( .A(_02636_ ), .B(_02637_ ), .S(_02102_ ), .Z(_02638_ ) );
OAI21_X1 _10240_ ( .A(_02088_ ), .B1(_02638_ ), .B2(_02606_ ), .ZN(_02639_ ) );
OAI221_X1 _10241_ ( .A(_02631_ ), .B1(_02635_ ), .B2(_02639_ ), .C1(_02540_ ), .C2(_02158_ ), .ZN(_02640_ ) );
OR3_X1 _10242_ ( .A1(_02540_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02541_ ), .ZN(_02641_ ) );
NAND2_X2 _10243_ ( .A1(_02640_ ), .A2(_02641_ ), .ZN(_02642_ ) );
INV_X1 _10244_ ( .A(\ID_EX_imm [18] ), .ZN(_02643_ ) );
XNOR2_X1 _10245_ ( .A(_02642_ ), .B(_02643_ ), .ZN(_02644_ ) );
OR3_X1 _10246_ ( .A1(_02147_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02541_ ), .ZN(_02645_ ) );
OR2_X1 _10247_ ( .A1(_02095_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02646_ ) );
OAI211_X1 _10248_ ( .A(_02646_ ), .B(fanout_net_30 ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02647_ ) );
OR2_X1 _10249_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02648_ ) );
OAI211_X1 _10250_ ( .A(_02648_ ), .B(_02103_ ), .C1(_02625_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02649_ ) );
NAND3_X1 _10251_ ( .A1(_02647_ ), .A2(_02606_ ), .A3(_02649_ ), .ZN(_02650_ ) );
MUX2_X1 _10252_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02651_ ) );
MUX2_X1 _10253_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02652_ ) );
MUX2_X1 _10254_ ( .A(_02651_ ), .B(_02652_ ), .S(_02103_ ), .Z(_02653_ ) );
OAI211_X1 _10255_ ( .A(fanout_net_34 ), .B(_02650_ ), .C1(_02653_ ), .C2(_02125_ ), .ZN(_02654_ ) );
OR2_X1 _10256_ ( .A1(_02095_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02655_ ) );
OAI211_X1 _10257_ ( .A(_02655_ ), .B(_02103_ ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02656_ ) );
OR2_X1 _10258_ ( .A1(_02095_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02657_ ) );
OAI211_X1 _10259_ ( .A(_02657_ ), .B(fanout_net_30 ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02658_ ) );
NAND3_X1 _10260_ ( .A1(_02656_ ), .A2(_02658_ ), .A3(_02606_ ), .ZN(_02659_ ) );
MUX2_X1 _10261_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02660_ ) );
MUX2_X1 _10262_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02661_ ) );
MUX2_X1 _10263_ ( .A(_02660_ ), .B(_02661_ ), .S(_02103_ ), .Z(_02662_ ) );
OAI211_X1 _10264_ ( .A(_02089_ ), .B(_02659_ ), .C1(_02662_ ), .C2(_02125_ ), .ZN(_02663_ ) );
OAI211_X1 _10265_ ( .A(_02654_ ), .B(_02663_ ), .C1(_02147_ ), .C2(_02158_ ), .ZN(_02664_ ) );
NAND2_X1 _10266_ ( .A1(_02645_ ), .A2(_02664_ ), .ZN(_02665_ ) );
BUF_X4 _10267_ ( .A(_02665_ ), .Z(_02666_ ) );
XOR2_X1 _10268_ ( .A(_02666_ ), .B(\ID_EX_imm [16] ), .Z(_02667_ ) );
OR3_X1 _10269_ ( .A1(_02146_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02157_ ), .ZN(_02668_ ) );
OR2_X1 _10270_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02669_ ) );
OAI211_X1 _10271_ ( .A(_02669_ ), .B(_02102_ ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02670_ ) );
OR2_X1 _10272_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02671_ ) );
OAI211_X1 _10273_ ( .A(_02671_ ), .B(fanout_net_31 ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02672_ ) );
NAND3_X1 _10274_ ( .A1(_02670_ ), .A2(_02672_ ), .A3(_02124_ ), .ZN(_02673_ ) );
MUX2_X1 _10275_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02674_ ) );
MUX2_X1 _10276_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02675_ ) );
MUX2_X1 _10277_ ( .A(_02674_ ), .B(_02675_ ), .S(_02102_ ), .Z(_02676_ ) );
OAI211_X1 _10278_ ( .A(fanout_net_34 ), .B(_02673_ ), .C1(_02676_ ), .C2(_02606_ ), .ZN(_02677_ ) );
OR2_X1 _10279_ ( .A1(_02405_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02678_ ) );
OAI211_X1 _10280_ ( .A(_02678_ ), .B(_02102_ ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02679_ ) );
OR2_X1 _10281_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02680_ ) );
OAI211_X1 _10282_ ( .A(_02680_ ), .B(fanout_net_31 ), .C1(_02095_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02681_ ) );
NAND3_X1 _10283_ ( .A1(_02679_ ), .A2(_02124_ ), .A3(_02681_ ), .ZN(_02682_ ) );
MUX2_X1 _10284_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02683_ ) );
MUX2_X1 _10285_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02684_ ) );
MUX2_X1 _10286_ ( .A(_02683_ ), .B(_02684_ ), .S(_02427_ ), .Z(_02685_ ) );
OAI211_X1 _10287_ ( .A(_02088_ ), .B(_02682_ ), .C1(_02685_ ), .C2(_02606_ ), .ZN(_02686_ ) );
OAI211_X1 _10288_ ( .A(_02677_ ), .B(_02686_ ), .C1(_02540_ ), .C2(_02541_ ), .ZN(_02687_ ) );
NAND2_X2 _10289_ ( .A1(_02668_ ), .A2(_02687_ ), .ZN(_02688_ ) );
AND2_X1 _10290_ ( .A1(_02688_ ), .A2(\ID_EX_imm [17] ), .ZN(_02689_ ) );
INV_X1 _10291_ ( .A(_02689_ ), .ZN(_02690_ ) );
INV_X1 _10292_ ( .A(\ID_EX_imm [17] ), .ZN(_02691_ ) );
AND3_X1 _10293_ ( .A1(_02668_ ), .A2(_02691_ ), .A3(_02687_ ), .ZN(_02692_ ) );
INV_X1 _10294_ ( .A(_02692_ ), .ZN(_02693_ ) );
AND3_X1 _10295_ ( .A1(_02667_ ), .A2(_02690_ ), .A3(_02693_ ), .ZN(_02694_ ) );
NAND4_X4 _10296_ ( .A1(_02596_ ), .A2(_02620_ ), .A3(_02644_ ), .A4(_02694_ ), .ZN(_02695_ ) );
NAND2_X1 _10297_ ( .A1(_02666_ ), .A2(\ID_EX_imm [16] ), .ZN(_02696_ ) );
OAI21_X1 _10298_ ( .A(_02690_ ), .B1(_02692_ ), .B2(_02696_ ), .ZN(_02697_ ) );
AND3_X1 _10299_ ( .A1(_02697_ ), .A2(_02620_ ), .A3(_02644_ ), .ZN(_02698_ ) );
AOI21_X1 _10300_ ( .A(_02619_ ), .B1(_02597_ ), .B2(_02617_ ), .ZN(_02699_ ) );
AND2_X1 _10301_ ( .A1(_02642_ ), .A2(\ID_EX_imm [18] ), .ZN(_02700_ ) );
AND2_X1 _10302_ ( .A1(_02620_ ), .A2(_02700_ ), .ZN(_02701_ ) );
NOR3_X1 _10303_ ( .A1(_02698_ ), .A2(_02699_ ), .A3(_02701_ ), .ZN(_02702_ ) );
AND2_X4 _10304_ ( .A1(_02695_ ), .A2(_02702_ ), .ZN(_02703_ ) );
OR2_X1 _10305_ ( .A1(_02093_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02704_ ) );
OAI211_X1 _10306_ ( .A(_02704_ ), .B(fanout_net_31 ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02705_ ) );
OR2_X1 _10307_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02706_ ) );
OAI211_X1 _10308_ ( .A(_02706_ ), .B(_02353_ ), .C1(_02094_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02707_ ) );
NAND3_X1 _10309_ ( .A1(_02705_ ), .A2(_02123_ ), .A3(_02707_ ), .ZN(_02708_ ) );
MUX2_X1 _10310_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02709_ ) );
MUX2_X1 _10311_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02710_ ) );
MUX2_X1 _10312_ ( .A(_02709_ ), .B(_02710_ ), .S(_02100_ ), .Z(_02711_ ) );
OAI211_X1 _10313_ ( .A(_02087_ ), .B(_02708_ ), .C1(_02711_ ), .C2(_02123_ ), .ZN(_02712_ ) );
OR2_X1 _10314_ ( .A1(_02093_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02713_ ) );
OAI211_X1 _10315_ ( .A(_02713_ ), .B(_02353_ ), .C1(fanout_net_26 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02714_ ) );
OR2_X1 _10316_ ( .A1(fanout_net_26 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02715_ ) );
OAI211_X1 _10317_ ( .A(_02715_ ), .B(fanout_net_31 ), .C1(_02094_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02716_ ) );
NAND3_X1 _10318_ ( .A1(_02714_ ), .A2(fanout_net_33 ), .A3(_02716_ ), .ZN(_02717_ ) );
MUX2_X1 _10319_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02718_ ) );
MUX2_X1 _10320_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_26 ), .Z(_02719_ ) );
MUX2_X1 _10321_ ( .A(_02718_ ), .B(_02719_ ), .S(fanout_net_31 ), .Z(_02720_ ) );
OAI211_X1 _10322_ ( .A(fanout_net_34 ), .B(_02717_ ), .C1(_02720_ ), .C2(fanout_net_33 ), .ZN(_02721_ ) );
NAND2_X1 _10323_ ( .A1(_02712_ ), .A2(_02721_ ), .ZN(_02722_ ) );
OAI21_X1 _10324_ ( .A(_02722_ ), .B1(_02347_ ), .B2(_02157_ ), .ZN(_02723_ ) );
NAND4_X1 _10325_ ( .A1(_02134_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02307_ ), .A4(_02143_ ), .ZN(_02724_ ) );
AND2_X1 _10326_ ( .A1(_02723_ ), .A2(_02724_ ), .ZN(_02725_ ) );
BUF_X4 _10327_ ( .A(_02725_ ), .Z(_02726_ ) );
XNOR2_X1 _10328_ ( .A(_02726_ ), .B(\ID_EX_imm [23] ), .ZN(_02727_ ) );
OR3_X1 _10329_ ( .A1(_02540_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02541_ ), .ZN(_02728_ ) );
OR2_X1 _10330_ ( .A1(_02440_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02729_ ) );
OAI211_X1 _10331_ ( .A(_02729_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02730_ ) );
OR2_X1 _10332_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02731_ ) );
OAI211_X1 _10333_ ( .A(_02731_ ), .B(_02624_ ), .C1(_02095_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02732_ ) );
NAND3_X1 _10334_ ( .A1(_02730_ ), .A2(_02124_ ), .A3(_02732_ ), .ZN(_02733_ ) );
MUX2_X1 _10335_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02734_ ) );
MUX2_X1 _10336_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02735_ ) );
MUX2_X1 _10337_ ( .A(_02734_ ), .B(_02735_ ), .S(_02102_ ), .Z(_02736_ ) );
OAI211_X1 _10338_ ( .A(_02088_ ), .B(_02733_ ), .C1(_02736_ ), .C2(_02606_ ), .ZN(_02737_ ) );
OR2_X1 _10339_ ( .A1(_02440_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02738_ ) );
OAI211_X1 _10340_ ( .A(_02738_ ), .B(_02624_ ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02739_ ) );
OR2_X1 _10341_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02740_ ) );
OAI211_X1 _10342_ ( .A(_02740_ ), .B(fanout_net_31 ), .C1(_02095_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02741_ ) );
NAND3_X1 _10343_ ( .A1(_02739_ ), .A2(fanout_net_33 ), .A3(_02741_ ), .ZN(_02742_ ) );
MUX2_X1 _10344_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02743_ ) );
MUX2_X1 _10345_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02744_ ) );
MUX2_X1 _10346_ ( .A(_02743_ ), .B(_02744_ ), .S(fanout_net_31 ), .Z(_02745_ ) );
OAI211_X1 _10347_ ( .A(fanout_net_34 ), .B(_02742_ ), .C1(_02745_ ), .C2(fanout_net_33 ), .ZN(_02746_ ) );
OAI211_X1 _10348_ ( .A(_02737_ ), .B(_02746_ ), .C1(_02540_ ), .C2(_02541_ ), .ZN(_02747_ ) );
NAND2_X2 _10349_ ( .A1(_02728_ ), .A2(_02747_ ), .ZN(_02748_ ) );
XNOR2_X1 _10350_ ( .A(_02748_ ), .B(\ID_EX_imm [22] ), .ZN(_02749_ ) );
OR3_X1 _10351_ ( .A1(_02540_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02541_ ), .ZN(_02750_ ) );
OR2_X1 _10352_ ( .A1(_02095_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02751_ ) );
OAI211_X1 _10353_ ( .A(_02751_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02752_ ) );
OR2_X1 _10354_ ( .A1(fanout_net_27 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02753_ ) );
OAI211_X1 _10355_ ( .A(_02753_ ), .B(_02624_ ), .C1(_02625_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02754_ ) );
NAND3_X1 _10356_ ( .A1(_02752_ ), .A2(_02606_ ), .A3(_02754_ ), .ZN(_02755_ ) );
MUX2_X1 _10357_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02756_ ) );
MUX2_X1 _10358_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02757_ ) );
MUX2_X1 _10359_ ( .A(_02756_ ), .B(_02757_ ), .S(_02624_ ), .Z(_02758_ ) );
OAI211_X1 _10360_ ( .A(_02089_ ), .B(_02755_ ), .C1(_02758_ ), .C2(_02125_ ), .ZN(_02759_ ) );
OR2_X1 _10361_ ( .A1(_02095_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02760_ ) );
OAI211_X1 _10362_ ( .A(_02760_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02761_ ) );
OR2_X1 _10363_ ( .A1(_02430_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02762_ ) );
OAI211_X1 _10364_ ( .A(_02762_ ), .B(_02624_ ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02763_ ) );
NAND3_X1 _10365_ ( .A1(_02761_ ), .A2(_02763_ ), .A3(fanout_net_33 ), .ZN(_02764_ ) );
MUX2_X1 _10366_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02765_ ) );
MUX2_X1 _10367_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02766_ ) );
MUX2_X1 _10368_ ( .A(_02765_ ), .B(_02766_ ), .S(fanout_net_31 ), .Z(_02767_ ) );
OAI211_X1 _10369_ ( .A(fanout_net_34 ), .B(_02764_ ), .C1(_02767_ ), .C2(fanout_net_33 ), .ZN(_02768_ ) );
OAI211_X1 _10370_ ( .A(_02759_ ), .B(_02768_ ), .C1(_02147_ ), .C2(_02158_ ), .ZN(_02769_ ) );
NAND2_X2 _10371_ ( .A1(_02750_ ), .A2(_02769_ ), .ZN(_02770_ ) );
INV_X1 _10372_ ( .A(\ID_EX_imm [20] ), .ZN(_02771_ ) );
XNOR2_X1 _10373_ ( .A(_02770_ ), .B(_02771_ ), .ZN(_02772_ ) );
OR3_X1 _10374_ ( .A1(_02540_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ), .A3(_02541_ ), .ZN(_02773_ ) );
OR2_X1 _10375_ ( .A1(_02430_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02774_ ) );
OAI211_X1 _10376_ ( .A(_02774_ ), .B(_02624_ ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02775_ ) );
OR2_X1 _10377_ ( .A1(_02430_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02776_ ) );
OAI211_X1 _10378_ ( .A(_02776_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02777_ ) );
NAND3_X1 _10379_ ( .A1(_02775_ ), .A2(_02777_ ), .A3(_02606_ ), .ZN(_02778_ ) );
MUX2_X1 _10380_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02779_ ) );
MUX2_X1 _10381_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02780_ ) );
MUX2_X1 _10382_ ( .A(_02779_ ), .B(_02780_ ), .S(_02624_ ), .Z(_02781_ ) );
OAI211_X1 _10383_ ( .A(_02088_ ), .B(_02778_ ), .C1(_02781_ ), .C2(_02125_ ), .ZN(_02782_ ) );
OR2_X1 _10384_ ( .A1(_02430_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02783_ ) );
OAI211_X1 _10385_ ( .A(_02783_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02784_ ) );
OR2_X1 _10386_ ( .A1(_02430_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02785_ ) );
OAI211_X1 _10387_ ( .A(_02785_ ), .B(_02624_ ), .C1(fanout_net_27 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02786_ ) );
NAND3_X1 _10388_ ( .A1(_02784_ ), .A2(_02786_ ), .A3(fanout_net_33 ), .ZN(_02787_ ) );
MUX2_X1 _10389_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02788_ ) );
MUX2_X1 _10390_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02789_ ) );
MUX2_X1 _10391_ ( .A(_02788_ ), .B(_02789_ ), .S(fanout_net_31 ), .Z(_02790_ ) );
OAI211_X1 _10392_ ( .A(fanout_net_34 ), .B(_02787_ ), .C1(_02790_ ), .C2(fanout_net_33 ), .ZN(_02791_ ) );
OAI211_X1 _10393_ ( .A(_02782_ ), .B(_02791_ ), .C1(_02147_ ), .C2(_02158_ ), .ZN(_02792_ ) );
NAND2_X2 _10394_ ( .A1(_02773_ ), .A2(_02792_ ), .ZN(_02793_ ) );
OR2_X1 _10395_ ( .A1(_02793_ ), .A2(\ID_EX_imm [21] ), .ZN(_02794_ ) );
NAND2_X1 _10396_ ( .A1(_02793_ ), .A2(\ID_EX_imm [21] ), .ZN(_02795_ ) );
NAND3_X1 _10397_ ( .A1(_02772_ ), .A2(_02794_ ), .A3(_02795_ ), .ZN(_02796_ ) );
NOR4_X4 _10398_ ( .A1(_02703_ ), .A2(_02727_ ), .A3(_02749_ ), .A4(_02796_ ), .ZN(_02797_ ) );
NOR2_X1 _10399_ ( .A1(_02749_ ), .A2(_02727_ ), .ZN(_02798_ ) );
INV_X1 _10400_ ( .A(_02770_ ), .ZN(_02799_ ) );
OAI21_X1 _10401_ ( .A(_02795_ ), .B1(_02799_ ), .B2(_02771_ ), .ZN(_02800_ ) );
NAND3_X1 _10402_ ( .A1(_02798_ ), .A2(_02794_ ), .A3(_02800_ ), .ZN(_02801_ ) );
INV_X1 _10403_ ( .A(_02727_ ), .ZN(_02802_ ) );
INV_X1 _10404_ ( .A(\ID_EX_imm [22] ), .ZN(_02803_ ) );
AOI21_X1 _10405_ ( .A(_02803_ ), .B1(_02728_ ), .B2(_02747_ ), .ZN(_02804_ ) );
NAND2_X1 _10406_ ( .A1(_02802_ ), .A2(_02804_ ), .ZN(_02805_ ) );
INV_X1 _10407_ ( .A(_02726_ ), .ZN(_02806_ ) );
OR2_X1 _10408_ ( .A1(_02806_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_02807_ ) );
NAND3_X1 _10409_ ( .A1(_02801_ ), .A2(_02805_ ), .A3(_02807_ ), .ZN(_02808_ ) );
OAI21_X4 _10410_ ( .A(_02164_ ), .B1(_02797_ ), .B2(_02808_ ), .ZN(_02809_ ) );
NAND2_X1 _10411_ ( .A1(_02162_ ), .A2(\ID_EX_imm [24] ), .ZN(_02810_ ) );
INV_X1 _10412_ ( .A(\ID_EX_imm [25] ), .ZN(_02811_ ) );
OR3_X1 _10413_ ( .A1(_02148_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02159_ ), .ZN(_02812_ ) );
OR2_X1 _10414_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02813_ ) );
OAI211_X1 _10415_ ( .A(_02813_ ), .B(fanout_net_31 ), .C1(fanout_net_27 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02814_ ) );
OR2_X1 _10416_ ( .A1(fanout_net_27 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02815_ ) );
BUF_X4 _10417_ ( .A(_02103_ ), .Z(_02816_ ) );
BUF_X2 _10418_ ( .A(_02625_ ), .Z(_02817_ ) );
OAI211_X1 _10419_ ( .A(_02815_ ), .B(_02816_ ), .C1(_02817_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02818_ ) );
NAND3_X1 _10420_ ( .A1(_02814_ ), .A2(_02126_ ), .A3(_02818_ ), .ZN(_02819_ ) );
MUX2_X1 _10421_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02820_ ) );
MUX2_X1 _10422_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_27 ), .Z(_02821_ ) );
MUX2_X1 _10423_ ( .A(_02820_ ), .B(_02821_ ), .S(_02816_ ), .Z(_02822_ ) );
OAI211_X1 _10424_ ( .A(_02089_ ), .B(_02819_ ), .C1(_02822_ ), .C2(_02126_ ), .ZN(_02823_ ) );
OR2_X1 _10425_ ( .A1(fanout_net_27 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02824_ ) );
OAI211_X1 _10426_ ( .A(_02824_ ), .B(_02816_ ), .C1(_02817_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02825_ ) );
NOR2_X1 _10427_ ( .A1(_02817_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02826_ ) );
OAI21_X1 _10428_ ( .A(fanout_net_31 ), .B1(fanout_net_27 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02827_ ) );
OAI211_X1 _10429_ ( .A(_02825_ ), .B(fanout_net_33 ), .C1(_02826_ ), .C2(_02827_ ), .ZN(_02828_ ) );
MUX2_X1 _10430_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02829_ ) );
MUX2_X1 _10431_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02830_ ) );
MUX2_X1 _10432_ ( .A(_02829_ ), .B(_02830_ ), .S(fanout_net_31 ), .Z(_02831_ ) );
OAI211_X1 _10433_ ( .A(fanout_net_34 ), .B(_02828_ ), .C1(_02831_ ), .C2(fanout_net_33 ), .ZN(_02832_ ) );
OAI211_X1 _10434_ ( .A(_02823_ ), .B(_02832_ ), .C1(_02148_ ), .C2(_02159_ ), .ZN(_02833_ ) );
NAND2_X2 _10435_ ( .A1(_02812_ ), .A2(_02833_ ), .ZN(_02834_ ) );
INV_X1 _10436_ ( .A(_02834_ ), .ZN(_02835_ ) );
OAI211_X2 _10437_ ( .A(_02809_ ), .B(_02810_ ), .C1(_02811_ ), .C2(_02835_ ), .ZN(_02836_ ) );
OAI21_X2 _10438_ ( .A(_02836_ ), .B1(\ID_EX_imm [25] ), .B2(_02834_ ), .ZN(_02837_ ) );
OR3_X1 _10439_ ( .A1(_02147_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02158_ ), .ZN(_02838_ ) );
OR2_X1 _10440_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02839_ ) );
OAI211_X1 _10441_ ( .A(_02839_ ), .B(_02104_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02840_ ) );
OR2_X1 _10442_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02841_ ) );
OAI211_X1 _10443_ ( .A(_02841_ ), .B(fanout_net_31 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02842_ ) );
NAND3_X1 _10444_ ( .A1(_02840_ ), .A2(_02842_ ), .A3(_02125_ ), .ZN(_02843_ ) );
MUX2_X1 _10445_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02844_ ) );
MUX2_X1 _10446_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02845_ ) );
MUX2_X1 _10447_ ( .A(_02844_ ), .B(_02845_ ), .S(_02104_ ), .Z(_02846_ ) );
OAI211_X1 _10448_ ( .A(_02089_ ), .B(_02843_ ), .C1(_02846_ ), .C2(_02126_ ), .ZN(_02847_ ) );
OR2_X1 _10449_ ( .A1(_02625_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02848_ ) );
OAI211_X1 _10450_ ( .A(_02848_ ), .B(_02104_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02849_ ) );
NOR2_X1 _10451_ ( .A1(_02817_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02850_ ) );
OAI21_X1 _10452_ ( .A(fanout_net_31 ), .B1(fanout_net_28 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02851_ ) );
OAI211_X1 _10453_ ( .A(_02849_ ), .B(fanout_net_33 ), .C1(_02850_ ), .C2(_02851_ ), .ZN(_02852_ ) );
MUX2_X1 _10454_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02853_ ) );
MUX2_X1 _10455_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02854_ ) );
MUX2_X1 _10456_ ( .A(_02853_ ), .B(_02854_ ), .S(fanout_net_31 ), .Z(_02855_ ) );
OAI211_X1 _10457_ ( .A(_02852_ ), .B(fanout_net_34 ), .C1(_02855_ ), .C2(fanout_net_33 ), .ZN(_02856_ ) );
OAI211_X1 _10458_ ( .A(_02847_ ), .B(_02856_ ), .C1(_02148_ ), .C2(_02159_ ), .ZN(_02857_ ) );
NAND2_X1 _10459_ ( .A1(_02838_ ), .A2(_02857_ ), .ZN(_02858_ ) );
XNOR2_X1 _10460_ ( .A(_02858_ ), .B(\ID_EX_imm [27] ), .ZN(_02859_ ) );
OR3_X1 _10461_ ( .A1(_02147_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ), .A3(_02158_ ), .ZN(_02860_ ) );
OR2_X1 _10462_ ( .A1(_02625_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02861_ ) );
OAI211_X1 _10463_ ( .A(_02861_ ), .B(_02104_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02862_ ) );
OR2_X1 _10464_ ( .A1(_02625_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02863_ ) );
OAI211_X1 _10465_ ( .A(_02863_ ), .B(fanout_net_31 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02864_ ) );
NAND3_X1 _10466_ ( .A1(_02862_ ), .A2(_02864_ ), .A3(_02125_ ), .ZN(_02865_ ) );
MUX2_X1 _10467_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02866_ ) );
MUX2_X1 _10468_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02867_ ) );
MUX2_X1 _10469_ ( .A(_02866_ ), .B(_02867_ ), .S(_02103_ ), .Z(_02868_ ) );
OAI211_X1 _10470_ ( .A(_02089_ ), .B(_02865_ ), .C1(_02868_ ), .C2(_02126_ ), .ZN(_02869_ ) );
OR2_X1 _10471_ ( .A1(_02625_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02870_ ) );
OAI211_X1 _10472_ ( .A(_02870_ ), .B(_02104_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02871_ ) );
NOR2_X1 _10473_ ( .A1(_02817_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02872_ ) );
OAI21_X1 _10474_ ( .A(fanout_net_31 ), .B1(fanout_net_28 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02873_ ) );
OAI211_X1 _10475_ ( .A(_02871_ ), .B(fanout_net_33 ), .C1(_02872_ ), .C2(_02873_ ), .ZN(_02874_ ) );
MUX2_X1 _10476_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02875_ ) );
MUX2_X1 _10477_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02876_ ) );
MUX2_X1 _10478_ ( .A(_02875_ ), .B(_02876_ ), .S(fanout_net_31 ), .Z(_02877_ ) );
OAI211_X1 _10479_ ( .A(_02874_ ), .B(fanout_net_34 ), .C1(_02877_ ), .C2(fanout_net_33 ), .ZN(_02878_ ) );
OAI211_X1 _10480_ ( .A(_02869_ ), .B(_02878_ ), .C1(_02148_ ), .C2(_02159_ ), .ZN(_02879_ ) );
NAND2_X1 _10481_ ( .A1(_02860_ ), .A2(_02879_ ), .ZN(_02880_ ) );
XNOR2_X1 _10482_ ( .A(_02880_ ), .B(\ID_EX_imm [26] ), .ZN(_02881_ ) );
NOR3_X4 _10483_ ( .A1(_02837_ ), .A2(_02859_ ), .A3(_02881_ ), .ZN(_02882_ ) );
INV_X1 _10484_ ( .A(\ID_EX_imm [27] ), .ZN(_02883_ ) );
AOI21_X1 _10485_ ( .A(_02883_ ), .B1(_02838_ ), .B2(_02857_ ), .ZN(_02884_ ) );
INV_X1 _10486_ ( .A(_02880_ ), .ZN(_02885_ ) );
OR2_X1 _10487_ ( .A1(_02885_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_3_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02886_ ) );
NOR2_X1 _10488_ ( .A1(_02859_ ), .A2(_02886_ ), .ZN(_02887_ ) );
NOR3_X4 _10489_ ( .A1(_02882_ ), .A2(_02884_ ), .A3(_02887_ ), .ZN(_02888_ ) );
OR3_X1 _10490_ ( .A1(_02147_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02158_ ), .ZN(_02889_ ) );
OR2_X1 _10491_ ( .A1(_02625_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02890_ ) );
OAI211_X1 _10492_ ( .A(_02890_ ), .B(_02104_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02891_ ) );
OR2_X1 _10493_ ( .A1(_02625_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02892_ ) );
OAI211_X1 _10494_ ( .A(_02892_ ), .B(fanout_net_31 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02893_ ) );
NAND3_X1 _10495_ ( .A1(_02891_ ), .A2(_02893_ ), .A3(fanout_net_33 ), .ZN(_02894_ ) );
MUX2_X1 _10496_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02895_ ) );
MUX2_X1 _10497_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02896_ ) );
MUX2_X1 _10498_ ( .A(_02895_ ), .B(_02896_ ), .S(_02103_ ), .Z(_02897_ ) );
OAI211_X1 _10499_ ( .A(_02089_ ), .B(_02894_ ), .C1(_02897_ ), .C2(fanout_net_33 ), .ZN(_02898_ ) );
NOR2_X1 _10500_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02899_ ) );
OAI21_X1 _10501_ ( .A(fanout_net_31 ), .B1(fanout_net_28 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02900_ ) );
NOR2_X1 _10502_ ( .A1(fanout_net_28 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02901_ ) );
OAI21_X1 _10503_ ( .A(_02103_ ), .B1(_02096_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02902_ ) );
OAI221_X1 _10504_ ( .A(_02125_ ), .B1(_02899_ ), .B2(_02900_ ), .C1(_02901_ ), .C2(_02902_ ), .ZN(_02903_ ) );
MUX2_X1 _10505_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02904_ ) );
MUX2_X1 _10506_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02905_ ) );
MUX2_X1 _10507_ ( .A(_02904_ ), .B(_02905_ ), .S(fanout_net_31 ), .Z(_02906_ ) );
OAI211_X1 _10508_ ( .A(fanout_net_34 ), .B(_02903_ ), .C1(_02906_ ), .C2(_02125_ ), .ZN(_02907_ ) );
OAI211_X1 _10509_ ( .A(_02898_ ), .B(_02907_ ), .C1(_02147_ ), .C2(_02158_ ), .ZN(_02908_ ) );
NAND2_X1 _10510_ ( .A1(_02889_ ), .A2(_02908_ ), .ZN(_02909_ ) );
XNOR2_X1 _10511_ ( .A(_02909_ ), .B(\ID_EX_imm [29] ), .ZN(_02910_ ) );
OR2_X1 _10512_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02911_ ) );
OAI211_X1 _10513_ ( .A(_02911_ ), .B(_02816_ ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02912_ ) );
OR2_X1 _10514_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02913_ ) );
OAI211_X1 _10515_ ( .A(_02913_ ), .B(fanout_net_31 ), .C1(fanout_net_28 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02914_ ) );
NAND3_X1 _10516_ ( .A1(_02912_ ), .A2(_02914_ ), .A3(_02126_ ), .ZN(_02915_ ) );
MUX2_X1 _10517_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02916_ ) );
MUX2_X1 _10518_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_28 ), .Z(_02917_ ) );
MUX2_X1 _10519_ ( .A(_02916_ ), .B(_02917_ ), .S(_02104_ ), .Z(_02918_ ) );
OAI211_X1 _10520_ ( .A(_02089_ ), .B(_02915_ ), .C1(_02918_ ), .C2(_02126_ ), .ZN(_02919_ ) );
OR2_X1 _10521_ ( .A1(_02096_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02920_ ) );
OAI211_X1 _10522_ ( .A(_02920_ ), .B(fanout_net_31 ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02921_ ) );
INV_X1 _10523_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02922_ ) );
NAND2_X1 _10524_ ( .A1(_02922_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .ZN(_02923_ ) );
OAI211_X1 _10525_ ( .A(_02923_ ), .B(_02104_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02924_ ) );
NAND3_X1 _10526_ ( .A1(_02921_ ), .A2(_02924_ ), .A3(fanout_net_33 ), .ZN(_02925_ ) );
MUX2_X1 _10527_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02926_ ) );
MUX2_X1 _10528_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02927_ ) );
MUX2_X1 _10529_ ( .A(_02926_ ), .B(_02927_ ), .S(fanout_net_31 ), .Z(_02928_ ) );
OAI211_X1 _10530_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02925_ ), .C1(_02928_ ), .C2(fanout_net_33 ), .ZN(_02929_ ) );
NAND2_X1 _10531_ ( .A1(_02919_ ), .A2(_02929_ ), .ZN(_02930_ ) );
OAI21_X1 _10532_ ( .A(_02930_ ), .B1(_02148_ ), .B2(_02159_ ), .ZN(_02931_ ) );
NAND4_X1 _10533_ ( .A1(_02134_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02307_ ), .A4(_02143_ ), .ZN(_02932_ ) );
AND2_X2 _10534_ ( .A1(_02931_ ), .A2(_02932_ ), .ZN(_02933_ ) );
XNOR2_X1 _10535_ ( .A(_02933_ ), .B(\ID_EX_imm [28] ), .ZN(_02934_ ) );
OR3_X4 _10536_ ( .A1(_02888_ ), .A2(_02910_ ), .A3(_02934_ ), .ZN(_02935_ ) );
INV_X1 _10537_ ( .A(_02910_ ), .ZN(_02936_ ) );
INV_X1 _10538_ ( .A(_02933_ ), .ZN(_02937_ ) );
NOR2_X1 _10539_ ( .A1(_02937_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_1_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02938_ ) );
INV_X1 _10540_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_02939_ ) );
AOI22_X1 _10541_ ( .A1(_02936_ ), .A2(_02938_ ), .B1(_02939_ ), .B2(_02909_ ), .ZN(_02940_ ) );
AND2_X4 _10542_ ( .A1(_02935_ ), .A2(_02940_ ), .ZN(_02941_ ) );
NOR2_X1 _10543_ ( .A1(_02817_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02942_ ) );
OAI21_X1 _10544_ ( .A(fanout_net_31 ), .B1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02943_ ) );
NOR2_X1 _10545_ ( .A1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02944_ ) );
OAI21_X1 _10546_ ( .A(_02816_ ), .B1(_02817_ ), .B2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02945_ ) );
OAI221_X1 _10547_ ( .A(fanout_net_33 ), .B1(_02942_ ), .B2(_02943_ ), .C1(_02944_ ), .C2(_02945_ ), .ZN(_02946_ ) );
MUX2_X1 _10548_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02947_ ) );
MUX2_X1 _10549_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02948_ ) );
MUX2_X1 _10550_ ( .A(_02947_ ), .B(_02948_ ), .S(_02816_ ), .Z(_02949_ ) );
OAI211_X1 _10551_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02946_ ), .C1(_02949_ ), .C2(fanout_net_33 ), .ZN(_02950_ ) );
MUX2_X1 _10552_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02951_ ) );
AND2_X1 _10553_ ( .A1(_02951_ ), .A2(_02816_ ), .ZN(_02952_ ) );
MUX2_X1 _10554_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02953_ ) );
AOI211_X1 _10555_ ( .A(fanout_net_33 ), .B(_02952_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C2(_02953_ ), .ZN(_02954_ ) );
MUX2_X1 _10556_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02955_ ) );
MUX2_X1 _10557_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02956_ ) );
MUX2_X1 _10558_ ( .A(_02955_ ), .B(_02956_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02957_ ) );
OAI21_X1 _10559_ ( .A(_02089_ ), .B1(_02957_ ), .B2(_02126_ ), .ZN(_02958_ ) );
OAI221_X1 _10560_ ( .A(_02950_ ), .B1(_02954_ ), .B2(_02958_ ), .C1(_02148_ ), .C2(_02159_ ), .ZN(_02959_ ) );
OR3_X1 _10561_ ( .A1(_02148_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_02159_ ), .ZN(_02960_ ) );
AND2_X1 _10562_ ( .A1(_02959_ ), .A2(_02960_ ), .ZN(_02961_ ) );
BUF_X4 _10563_ ( .A(_02961_ ), .Z(_02962_ ) );
XNOR2_X1 _10564_ ( .A(_02962_ ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_02963_ ) );
OR2_X4 _10565_ ( .A1(_02941_ ), .A2(_02963_ ), .ZN(_02964_ ) );
OAI21_X4 _10566_ ( .A(_02964_ ), .B1(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B ), .B2(_02962_ ), .ZN(_02965_ ) );
OR3_X1 _10567_ ( .A1(_02148_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_02159_ ), .ZN(_02966_ ) );
OR2_X1 _10568_ ( .A1(_02817_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02967_ ) );
OAI211_X1 _10569_ ( .A(_02967_ ), .B(_02816_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02968_ ) );
INV_X1 _10570_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02969_ ) );
NAND2_X1 _10571_ ( .A1(_02969_ ), .A2(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .ZN(_02970_ ) );
OAI211_X1 _10572_ ( .A(_02970_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02971_ ) );
NAND3_X1 _10573_ ( .A1(_02968_ ), .A2(_02971_ ), .A3(_02126_ ), .ZN(_02972_ ) );
MUX2_X1 _10574_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02973_ ) );
MUX2_X1 _10575_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02974_ ) );
MUX2_X1 _10576_ ( .A(_02973_ ), .B(_02974_ ), .S(_02816_ ), .Z(_02975_ ) );
OAI211_X1 _10577_ ( .A(_02089_ ), .B(_02972_ ), .C1(_02975_ ), .C2(_02126_ ), .ZN(_02976_ ) );
OR2_X1 _10578_ ( .A1(_02817_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_02977_ ) );
OAI211_X1 _10579_ ( .A(_02977_ ), .B(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_02978_ ) );
OR2_X1 _10580_ ( .A1(_02817_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_02979_ ) );
OAI211_X1 _10581_ ( .A(_02979_ ), .B(_02816_ ), .C1(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_02980_ ) );
NAND3_X1 _10582_ ( .A1(_02978_ ), .A2(_02980_ ), .A3(fanout_net_33 ), .ZN(_02981_ ) );
MUX2_X1 _10583_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02982_ ) );
MUX2_X1 _10584_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_02983_ ) );
MUX2_X1 _10585_ ( .A(_02982_ ), .B(_02983_ ), .S(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_02984_ ) );
OAI211_X1 _10586_ ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_02981_ ), .C1(_02984_ ), .C2(fanout_net_33 ), .ZN(_02985_ ) );
OAI211_X1 _10587_ ( .A(_02976_ ), .B(_02985_ ), .C1(_02148_ ), .C2(_02159_ ), .ZN(_02986_ ) );
NAND2_X1 _10588_ ( .A1(_02966_ ), .A2(_02986_ ), .ZN(_02987_ ) );
BUF_X2 _10589_ ( .A(_02987_ ), .Z(_02988_ ) );
XNOR2_X1 _10590_ ( .A(_02988_ ), .B(\ID_EX_imm [31] ), .ZN(_02989_ ) );
XOR2_X2 _10591_ ( .A(_02965_ ), .B(_02989_ ), .Z(_02990_ ) );
AND2_X1 _10592_ ( .A1(\ID_EX_typ [7] ), .A2(\ID_EX_typ [6] ), .ZN(_02991_ ) );
BUF_X4 _10593_ ( .A(_02991_ ), .Z(_02992_ ) );
BUF_X4 _10594_ ( .A(_02992_ ), .Z(_02993_ ) );
NOR2_X1 _10595_ ( .A1(_02990_ ), .A2(_02993_ ), .ZN(_00097_ ) );
XNOR2_X1 _10596_ ( .A(_02941_ ), .B(_02963_ ), .ZN(_02994_ ) );
NOR2_X1 _10597_ ( .A1(_02994_ ), .A2(_02993_ ), .ZN(_00098_ ) );
INV_X1 _10598_ ( .A(_02772_ ), .ZN(_02995_ ) );
AOI21_X1 _10599_ ( .A(_02995_ ), .B1(_02695_ ), .B2(_02702_ ), .ZN(_02996_ ) );
AND2_X1 _10600_ ( .A1(_02770_ ), .A2(\ID_EX_imm [20] ), .ZN(_02997_ ) );
NOR2_X1 _10601_ ( .A1(_02996_ ), .A2(_02997_ ), .ZN(_02998_ ) );
XNOR2_X1 _10602_ ( .A(_02793_ ), .B(\ID_EX_imm [21] ), .ZN(_02999_ ) );
XNOR2_X1 _10603_ ( .A(_02998_ ), .B(_02999_ ), .ZN(_03000_ ) );
NOR2_X1 _10604_ ( .A1(_03000_ ), .A2(_02993_ ), .ZN(_00099_ ) );
XNOR2_X1 _10605_ ( .A(_02703_ ), .B(_02995_ ), .ZN(_03001_ ) );
NOR2_X1 _10606_ ( .A1(_03001_ ), .A2(_02993_ ), .ZN(_00100_ ) );
AOI21_X1 _10607_ ( .A(_02697_ ), .B1(_02596_ ), .B2(_02694_ ), .ZN(_03002_ ) );
INV_X1 _10608_ ( .A(_02644_ ), .ZN(_03003_ ) );
NOR2_X1 _10609_ ( .A1(_03002_ ), .A2(_03003_ ), .ZN(_03004_ ) );
NOR2_X1 _10610_ ( .A1(_03004_ ), .A2(_02700_ ), .ZN(_03005_ ) );
XNOR2_X1 _10611_ ( .A(_03005_ ), .B(_02620_ ), .ZN(_03006_ ) );
INV_X1 _10612_ ( .A(_02991_ ), .ZN(_03007_ ) );
CLKBUF_X2 _10613_ ( .A(_03007_ ), .Z(_03008_ ) );
AND2_X1 _10614_ ( .A1(_03006_ ), .A2(_03008_ ), .ZN(_00101_ ) );
XNOR2_X1 _10615_ ( .A(_03002_ ), .B(_03003_ ), .ZN(_03009_ ) );
NOR2_X1 _10616_ ( .A1(_03009_ ), .A2(_02993_ ), .ZN(_00102_ ) );
NAND2_X1 _10617_ ( .A1(_02596_ ), .A2(_02667_ ), .ZN(_03010_ ) );
AND4_X1 _10618_ ( .A1(_02690_ ), .A2(_03010_ ), .A3(_02693_ ), .A4(_02696_ ), .ZN(_03011_ ) );
AOI22_X1 _10619_ ( .A1(_03010_ ), .A2(_02696_ ), .B1(_02690_ ), .B2(_02693_ ), .ZN(_03012_ ) );
NOR2_X1 _10620_ ( .A1(_03011_ ), .A2(_03012_ ), .ZN(_03013_ ) );
NOR2_X1 _10621_ ( .A1(_03013_ ), .A2(_02993_ ), .ZN(_00103_ ) );
XNOR2_X1 _10622_ ( .A(_02596_ ), .B(_02667_ ), .ZN(_03014_ ) );
NOR2_X1 _10623_ ( .A1(_03014_ ), .A2(_02993_ ), .ZN(_00104_ ) );
AOI21_X1 _10624_ ( .A(_02544_ ), .B1(_02475_ ), .B2(_02584_ ), .ZN(_03015_ ) );
OAI21_X1 _10625_ ( .A(_02568_ ), .B1(_03015_ ), .B2(_02590_ ), .ZN(_03016_ ) );
OR2_X1 _10626_ ( .A1(_03016_ ), .A2(_02497_ ), .ZN(_03017_ ) );
NAND2_X1 _10627_ ( .A1(_03017_ ), .A2(_02593_ ), .ZN(_03018_ ) );
XNOR2_X1 _10628_ ( .A(_03018_ ), .B(_02519_ ), .ZN(_03019_ ) );
AND2_X1 _10629_ ( .A1(_03019_ ), .A2(_03008_ ), .ZN(_00105_ ) );
XOR2_X1 _10630_ ( .A(_03016_ ), .B(_02497_ ), .Z(_03020_ ) );
AND2_X1 _10631_ ( .A1(_03020_ ), .A2(_03008_ ), .ZN(_00106_ ) );
INV_X1 _10632_ ( .A(_03015_ ), .ZN(_03021_ ) );
AND2_X1 _10633_ ( .A1(_03021_ ), .A2(_02589_ ), .ZN(_03022_ ) );
XNOR2_X1 _10634_ ( .A(_03022_ ), .B(_02569_ ), .ZN(_03023_ ) );
NOR2_X1 _10635_ ( .A1(_03023_ ), .A2(_02993_ ), .ZN(_00107_ ) );
AND3_X1 _10636_ ( .A1(_02475_ ), .A2(_02544_ ), .A3(_02584_ ), .ZN(_03024_ ) );
NOR3_X1 _10637_ ( .A1(_03024_ ), .A2(_03015_ ), .A3(_02992_ ), .ZN(_00108_ ) );
NOR2_X1 _10638_ ( .A1(_02888_ ), .A2(_02934_ ), .ZN(_03025_ ) );
NOR2_X1 _10639_ ( .A1(_03025_ ), .A2(_02938_ ), .ZN(_03026_ ) );
XNOR2_X1 _10640_ ( .A(_03026_ ), .B(_02936_ ), .ZN(_03027_ ) );
AND2_X1 _10641_ ( .A1(_03027_ ), .A2(_03008_ ), .ZN(_00109_ ) );
XOR2_X1 _10642_ ( .A(_02888_ ), .B(_02934_ ), .Z(_03028_ ) );
AND2_X1 _10643_ ( .A1(_03028_ ), .A2(_03008_ ), .ZN(_00110_ ) );
OR2_X1 _10644_ ( .A1(_02837_ ), .A2(_02881_ ), .ZN(_03029_ ) );
NAND2_X1 _10645_ ( .A1(_03029_ ), .A2(_02886_ ), .ZN(_03030_ ) );
XNOR2_X1 _10646_ ( .A(_03030_ ), .B(_02859_ ), .ZN(_03031_ ) );
AND2_X1 _10647_ ( .A1(_03031_ ), .A2(_03008_ ), .ZN(_00111_ ) );
XOR2_X1 _10648_ ( .A(_02837_ ), .B(_02881_ ), .Z(_03032_ ) );
AND2_X1 _10649_ ( .A1(_03032_ ), .A2(_03008_ ), .ZN(_00112_ ) );
AND2_X1 _10650_ ( .A1(_02809_ ), .A2(_02810_ ), .ZN(_03033_ ) );
XNOR2_X1 _10651_ ( .A(_02834_ ), .B(\ID_EX_imm [25] ), .ZN(_03034_ ) );
XNOR2_X1 _10652_ ( .A(_03033_ ), .B(_03034_ ), .ZN(_03035_ ) );
NOR2_X1 _10653_ ( .A1(_03035_ ), .A2(_02993_ ), .ZN(_00113_ ) );
OR3_X1 _10654_ ( .A1(_02797_ ), .A2(_02808_ ), .A3(_02164_ ), .ZN(_03036_ ) );
AND3_X1 _10655_ ( .A1(_03036_ ), .A2(_02809_ ), .A3(_03007_ ), .ZN(_00114_ ) );
OAI21_X1 _10656_ ( .A(_02794_ ), .B1(_02996_ ), .B2(_02800_ ), .ZN(_03037_ ) );
NOR2_X1 _10657_ ( .A1(_03037_ ), .A2(_02749_ ), .ZN(_03038_ ) );
NOR2_X1 _10658_ ( .A1(_03038_ ), .A2(_02804_ ), .ZN(_03039_ ) );
XNOR2_X1 _10659_ ( .A(_03039_ ), .B(_02802_ ), .ZN(_03040_ ) );
AND2_X1 _10660_ ( .A1(_03040_ ), .A2(_03008_ ), .ZN(_00115_ ) );
XOR2_X1 _10661_ ( .A(_03037_ ), .B(_02749_ ), .Z(_03041_ ) );
AND2_X1 _10662_ ( .A1(_03041_ ), .A2(_03007_ ), .ZN(_00116_ ) );
INV_X1 _10663_ ( .A(\IF_ID_inst [6] ), .ZN(_03042_ ) );
NOR2_X1 _10664_ ( .A1(_03042_ ), .A2(\IF_ID_inst [12] ), .ZN(_03043_ ) );
AND2_X1 _10665_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03044_ ) );
AND3_X1 _10666_ ( .A1(_03043_ ), .A2(\IF_ID_inst [13] ), .A3(_03044_ ), .ZN(_03045_ ) );
AND2_X1 _10667_ ( .A1(\IF_ID_inst [0] ), .A2(\IF_ID_inst [1] ), .ZN(_03046_ ) );
NOR2_X1 _10668_ ( .A1(\IF_ID_inst [3] ), .A2(\IF_ID_inst [2] ), .ZN(_03047_ ) );
AND2_X2 _10669_ ( .A1(_03046_ ), .A2(_03047_ ), .ZN(_03048_ ) );
CLKBUF_X2 _10670_ ( .A(_03048_ ), .Z(_03049_ ) );
AND2_X1 _10671_ ( .A1(_03045_ ), .A2(_03049_ ), .ZN(_03050_ ) );
AND2_X1 _10672_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03051_ ) );
AND3_X1 _10673_ ( .A1(_03046_ ), .A2(_03051_ ), .A3(_03047_ ), .ZN(_03052_ ) );
CLKBUF_X2 _10674_ ( .A(_03044_ ), .Z(_03053_ ) );
AND2_X2 _10675_ ( .A1(_03052_ ), .A2(_03053_ ), .ZN(_03054_ ) );
NOR2_X1 _10676_ ( .A1(_03050_ ), .A2(_03054_ ), .ZN(_03055_ ) );
BUF_X4 _10677_ ( .A(_03055_ ), .Z(_03056_ ) );
INV_X1 _10678_ ( .A(\IF_ID_inst [31] ), .ZN(_03057_ ) );
BUF_X2 _10679_ ( .A(_03057_ ), .Z(_03058_ ) );
NOR2_X1 _10680_ ( .A1(_02078_ ), .A2(excp_written ), .ZN(_03059_ ) );
INV_X1 _10681_ ( .A(_03059_ ), .ZN(_03060_ ) );
BUF_X4 _10682_ ( .A(_03060_ ), .Z(_03061_ ) );
BUF_X4 _10683_ ( .A(_03061_ ), .Z(_03062_ ) );
NOR3_X1 _10684_ ( .A1(_03056_ ), .A2(_03058_ ), .A3(_03062_ ), .ZN(_00117_ ) );
INV_X1 _10685_ ( .A(\IF_ID_inst [30] ), .ZN(_03063_ ) );
NOR3_X1 _10686_ ( .A1(_03056_ ), .A2(_03063_ ), .A3(_03062_ ), .ZN(_00118_ ) );
INV_X1 _10687_ ( .A(\IF_ID_inst [21] ), .ZN(_03064_ ) );
NOR3_X1 _10688_ ( .A1(_03056_ ), .A2(_03064_ ), .A3(_03062_ ), .ZN(_00119_ ) );
BUF_X4 _10689_ ( .A(_03061_ ), .Z(_03065_ ) );
INV_X1 _10690_ ( .A(_03055_ ), .ZN(_03066_ ) );
INV_X1 _10691_ ( .A(\IF_ID_inst [20] ), .ZN(_03067_ ) );
AOI21_X1 _10692_ ( .A(_03065_ ), .B1(_03066_ ), .B2(_03067_ ), .ZN(_00120_ ) );
INV_X1 _10693_ ( .A(\IF_ID_inst [29] ), .ZN(_03068_ ) );
AOI21_X1 _10694_ ( .A(_03065_ ), .B1(_03066_ ), .B2(_03068_ ), .ZN(_00121_ ) );
INV_X1 _10695_ ( .A(\IF_ID_inst [28] ), .ZN(_03069_ ) );
AOI21_X1 _10696_ ( .A(_03065_ ), .B1(_03066_ ), .B2(_03069_ ), .ZN(_00122_ ) );
INV_X1 _10697_ ( .A(\IF_ID_inst [27] ), .ZN(_03070_ ) );
NOR3_X1 _10698_ ( .A1(_03056_ ), .A2(_03070_ ), .A3(_03062_ ), .ZN(_00123_ ) );
INV_X1 _10699_ ( .A(\IF_ID_inst [26] ), .ZN(_03071_ ) );
AOI21_X1 _10700_ ( .A(_03065_ ), .B1(_03066_ ), .B2(_03071_ ), .ZN(_00124_ ) );
INV_X1 _10701_ ( .A(\IF_ID_inst [25] ), .ZN(_03072_ ) );
NOR3_X1 _10702_ ( .A1(_03056_ ), .A2(_03072_ ), .A3(_03062_ ), .ZN(_00125_ ) );
INV_X1 _10703_ ( .A(\IF_ID_inst [24] ), .ZN(_03073_ ) );
BUF_X4 _10704_ ( .A(_03060_ ), .Z(_03074_ ) );
NOR3_X1 _10705_ ( .A1(_03056_ ), .A2(_03073_ ), .A3(_03074_ ), .ZN(_00126_ ) );
INV_X1 _10706_ ( .A(\IF_ID_inst [23] ), .ZN(_03075_ ) );
NOR3_X1 _10707_ ( .A1(_03056_ ), .A2(_03075_ ), .A3(_03074_ ), .ZN(_00127_ ) );
INV_X1 _10708_ ( .A(\IF_ID_inst [22] ), .ZN(_03076_ ) );
NOR3_X1 _10709_ ( .A1(_03056_ ), .A2(_03076_ ), .A3(_03074_ ), .ZN(_00128_ ) );
BUF_X2 _10710_ ( .A(_03059_ ), .Z(_03077_ ) );
AND2_X1 _10711_ ( .A1(_03077_ ), .A2(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .ZN(_00129_ ) );
AND2_X1 _10712_ ( .A1(_03077_ ), .A2(\myidu.state [2] ), .ZN(_00130_ ) );
INV_X1 _10713_ ( .A(\IF_ID_inst [12] ), .ZN(_03078_ ) );
INV_X1 _10714_ ( .A(\IF_ID_inst [7] ), .ZN(_03079_ ) );
INV_X1 _10715_ ( .A(\IF_ID_inst [15] ), .ZN(_03080_ ) );
AND4_X1 _10716_ ( .A1(_03078_ ), .A2(_03079_ ), .A3(_03080_ ), .A4(\IF_ID_inst [6] ), .ZN(_03081_ ) );
NOR2_X1 _10717_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_03082_ ) );
AND3_X1 _10718_ ( .A1(_03081_ ), .A2(_03053_ ), .A3(_03082_ ), .ZN(_03083_ ) );
BUF_X2 _10719_ ( .A(_03049_ ), .Z(_03084_ ) );
INV_X1 _10720_ ( .A(\IF_ID_inst [11] ), .ZN(_03085_ ) );
INV_X1 _10721_ ( .A(\IF_ID_inst [10] ), .ZN(_03086_ ) );
INV_X1 _10722_ ( .A(\IF_ID_inst [9] ), .ZN(_03087_ ) );
NAND3_X1 _10723_ ( .A1(_03085_ ), .A2(_03086_ ), .A3(_03087_ ), .ZN(_03088_ ) );
NOR2_X1 _10724_ ( .A1(_03088_ ), .A2(\IF_ID_inst [8] ), .ZN(_03089_ ) );
NAND3_X1 _10725_ ( .A1(_03083_ ), .A2(_03084_ ), .A3(_03089_ ), .ZN(_03090_ ) );
NAND2_X1 _10726_ ( .A1(_03057_ ), .A2(\IF_ID_inst [28] ), .ZN(_03091_ ) );
NOR3_X1 _10727_ ( .A1(_03091_ ), .A2(\IF_ID_inst [30] ), .A3(_03068_ ), .ZN(_03092_ ) );
NOR2_X1 _10728_ ( .A1(\IF_ID_inst [23] ), .A2(\IF_ID_inst [22] ), .ZN(_03093_ ) );
AND3_X1 _10729_ ( .A1(_03093_ ), .A2(\IF_ID_inst [21] ), .A3(_03067_ ), .ZN(_03094_ ) );
NOR2_X1 _10730_ ( .A1(\IF_ID_inst [18] ), .A2(\IF_ID_inst [17] ), .ZN(_03095_ ) );
NOR2_X1 _10731_ ( .A1(\IF_ID_inst [19] ), .A2(\IF_ID_inst [16] ), .ZN(_03096_ ) );
AND2_X1 _10732_ ( .A1(_03095_ ), .A2(_03096_ ), .ZN(_03097_ ) );
NOR2_X1 _10733_ ( .A1(\IF_ID_inst [26] ), .A2(\IF_ID_inst [25] ), .ZN(_03098_ ) );
NOR2_X1 _10734_ ( .A1(\IF_ID_inst [27] ), .A2(\IF_ID_inst [24] ), .ZN(_03099_ ) );
AND2_X1 _10735_ ( .A1(_03098_ ), .A2(_03099_ ), .ZN(_03100_ ) );
NAND4_X1 _10736_ ( .A1(_03092_ ), .A2(_03094_ ), .A3(_03097_ ), .A4(_03100_ ), .ZN(_03101_ ) );
NOR2_X1 _10737_ ( .A1(_03090_ ), .A2(_03101_ ), .ZN(_03102_ ) );
INV_X1 _10738_ ( .A(\IF_ID_inst [5] ), .ZN(_03103_ ) );
NOR2_X2 _10739_ ( .A1(_03103_ ), .A2(\IF_ID_inst [4] ), .ZN(_03104_ ) );
AND2_X1 _10740_ ( .A1(_03043_ ), .A2(_03104_ ), .ZN(_03105_ ) );
AND2_X1 _10741_ ( .A1(_03105_ ), .A2(_03049_ ), .ZN(_03106_ ) );
BUF_X2 _10742_ ( .A(_03082_ ), .Z(_03107_ ) );
AND2_X1 _10743_ ( .A1(_03106_ ), .A2(_03107_ ), .ZN(_03108_ ) );
NOR2_X1 _10744_ ( .A1(\IF_ID_inst [4] ), .A2(\IF_ID_inst [5] ), .ZN(_03109_ ) );
AND4_X1 _10745_ ( .A1(\IF_ID_inst [12] ), .A2(_03107_ ), .A3(_03109_ ), .A4(_03042_ ), .ZN(_03110_ ) );
AND3_X2 _10746_ ( .A1(_03046_ ), .A2(\IF_ID_inst [3] ), .A3(\IF_ID_inst [2] ), .ZN(_03111_ ) );
CLKBUF_X2 _10747_ ( .A(_03111_ ), .Z(_03112_ ) );
AND2_X1 _10748_ ( .A1(_03110_ ), .A2(_03112_ ), .ZN(_03113_ ) );
NOR3_X1 _10749_ ( .A1(_03102_ ), .A2(_03108_ ), .A3(_03113_ ), .ZN(_03114_ ) );
NOR2_X1 _10750_ ( .A1(\IF_ID_inst [12] ), .A2(\IF_ID_inst [6] ), .ZN(_03115_ ) );
AND3_X1 _10751_ ( .A1(_03049_ ), .A2(_03104_ ), .A3(_03115_ ), .ZN(_03116_ ) );
INV_X1 _10752_ ( .A(\IF_ID_inst [13] ), .ZN(_03117_ ) );
NOR2_X1 _10753_ ( .A1(_03117_ ), .A2(\IF_ID_inst [14] ), .ZN(_03118_ ) );
AND2_X1 _10754_ ( .A1(_03116_ ), .A2(_03118_ ), .ZN(_03119_ ) );
INV_X1 _10755_ ( .A(_03119_ ), .ZN(_03120_ ) );
NOR2_X1 _10756_ ( .A1(_03078_ ), .A2(\IF_ID_inst [6] ), .ZN(_03121_ ) );
AND3_X1 _10757_ ( .A1(_03049_ ), .A2(_03104_ ), .A3(_03121_ ), .ZN(_03122_ ) );
OAI21_X1 _10758_ ( .A(_03082_ ), .B1(_03116_ ), .B2(_03122_ ), .ZN(_03123_ ) );
AND2_X1 _10759_ ( .A1(_03120_ ), .A2(_03123_ ), .ZN(_03124_ ) );
INV_X1 _10760_ ( .A(_03100_ ), .ZN(_03125_ ) );
NAND4_X1 _10761_ ( .A1(_03063_ ), .A2(_03068_ ), .A3(_03069_ ), .A4(_03057_ ), .ZN(_03126_ ) );
NOR3_X1 _10762_ ( .A1(_03090_ ), .A2(_03125_ ), .A3(_03126_ ), .ZN(_03127_ ) );
AND3_X1 _10763_ ( .A1(_03095_ ), .A2(_03096_ ), .A3(_03093_ ), .ZN(_03128_ ) );
AND3_X1 _10764_ ( .A1(_03128_ ), .A2(_03064_ ), .A3(\IF_ID_inst [20] ), .ZN(_03129_ ) );
NAND2_X1 _10765_ ( .A1(_03127_ ), .A2(_03129_ ), .ZN(_03130_ ) );
AND3_X1 _10766_ ( .A1(_03114_ ), .A2(_03124_ ), .A3(_03130_ ), .ZN(_03131_ ) );
AND2_X1 _10767_ ( .A1(_03052_ ), .A2(_03104_ ), .ZN(_03132_ ) );
AND3_X1 _10768_ ( .A1(_03132_ ), .A2(\IF_ID_inst [13] ), .A3(\IF_ID_inst [14] ), .ZN(_03133_ ) );
AND2_X1 _10769_ ( .A1(_03106_ ), .A2(\IF_ID_inst [14] ), .ZN(_03134_ ) );
AND3_X1 _10770_ ( .A1(_03052_ ), .A2(_03117_ ), .A3(_03104_ ), .ZN(_03135_ ) );
NOR3_X1 _10771_ ( .A1(_03133_ ), .A2(_03134_ ), .A3(_03135_ ), .ZN(_03136_ ) );
AND4_X1 _10772_ ( .A1(\IF_ID_inst [11] ), .A2(_03131_ ), .A3(_03059_ ), .A4(_03136_ ), .ZN(_00131_ ) );
AND4_X1 _10773_ ( .A1(\IF_ID_inst [10] ), .A2(_03131_ ), .A3(_03059_ ), .A4(_03136_ ), .ZN(_00132_ ) );
AND4_X1 _10774_ ( .A1(\IF_ID_inst [9] ), .A2(_03131_ ), .A3(_03059_ ), .A4(_03136_ ), .ZN(_00133_ ) );
AND4_X1 _10775_ ( .A1(\IF_ID_inst [8] ), .A2(_03131_ ), .A3(_03059_ ), .A4(_03136_ ), .ZN(_00134_ ) );
AND4_X1 _10776_ ( .A1(\IF_ID_inst [7] ), .A2(_03131_ ), .A3(_03059_ ), .A4(_03136_ ), .ZN(_00135_ ) );
AND4_X1 _10777_ ( .A1(\IF_ID_inst [6] ), .A2(_03049_ ), .A3(_03079_ ), .A4(_03044_ ), .ZN(_03137_ ) );
NOR4_X1 _10778_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .A3(\IF_ID_inst [12] ), .A4(\IF_ID_inst [15] ), .ZN(_03138_ ) );
AND3_X1 _10779_ ( .A1(_03137_ ), .A2(_03089_ ), .A3(_03138_ ), .ZN(_03139_ ) );
NAND4_X1 _10780_ ( .A1(_03097_ ), .A2(_03064_ ), .A3(\IF_ID_inst [20] ), .A4(_03093_ ), .ZN(_03140_ ) );
NOR3_X1 _10781_ ( .A1(_03140_ ), .A2(_03125_ ), .A3(_03126_ ), .ZN(_03141_ ) );
NAND2_X1 _10782_ ( .A1(_03139_ ), .A2(_03141_ ), .ZN(_03142_ ) );
AND3_X1 _10783_ ( .A1(_03109_ ), .A2(\IF_ID_inst [12] ), .A3(_03042_ ), .ZN(_03143_ ) );
AND2_X1 _10784_ ( .A1(_03112_ ), .A2(_03143_ ), .ZN(_03144_ ) );
NAND2_X1 _10785_ ( .A1(_03144_ ), .A2(_03107_ ), .ZN(_03145_ ) );
NAND2_X1 _10786_ ( .A1(_03142_ ), .A2(_03145_ ), .ZN(_03146_ ) );
AND3_X1 _10787_ ( .A1(_03083_ ), .A2(_03049_ ), .A3(_03089_ ), .ZN(_03147_ ) );
AND4_X1 _10788_ ( .A1(_03097_ ), .A2(_03092_ ), .A3(_03094_ ), .A4(_03100_ ), .ZN(_03148_ ) );
NAND2_X1 _10789_ ( .A1(_03147_ ), .A2(_03148_ ), .ZN(_03149_ ) );
INV_X1 _10790_ ( .A(\IF_ID_inst [2] ), .ZN(_03150_ ) );
NOR2_X1 _10791_ ( .A1(_03150_ ), .A2(\IF_ID_inst [3] ), .ZN(_03151_ ) );
AND2_X1 _10792_ ( .A1(_03151_ ), .A2(_03046_ ), .ZN(_03152_ ) );
INV_X1 _10793_ ( .A(\IF_ID_inst [4] ), .ZN(_03153_ ) );
NOR2_X1 _10794_ ( .A1(_03153_ ), .A2(\IF_ID_inst [6] ), .ZN(_03154_ ) );
AND2_X1 _10795_ ( .A1(_03152_ ), .A2(_03154_ ), .ZN(_03155_ ) );
INV_X1 _10796_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_03156_ ) );
AND2_X2 _10797_ ( .A1(_03104_ ), .A2(_03156_ ), .ZN(_03157_ ) );
AND2_X1 _10798_ ( .A1(_03157_ ), .A2(_03111_ ), .ZN(_03158_ ) );
BUF_X2 _10799_ ( .A(_03158_ ), .Z(_03159_ ) );
NOR2_X1 _10800_ ( .A1(_03155_ ), .A2(_03159_ ), .ZN(_03160_ ) );
NAND2_X1 _10801_ ( .A1(_03149_ ), .A2(_03160_ ), .ZN(_03161_ ) );
INV_X1 _10802_ ( .A(\IF_ID_inst [19] ), .ZN(_03162_ ) );
NOR4_X1 _10803_ ( .A1(_03146_ ), .A2(_03161_ ), .A3(_03162_ ), .A4(_03061_ ), .ZN(_00136_ ) );
INV_X1 _10804_ ( .A(\IF_ID_inst [18] ), .ZN(_03163_ ) );
NOR4_X1 _10805_ ( .A1(_03146_ ), .A2(_03161_ ), .A3(_03163_ ), .A4(_03061_ ), .ZN(_00137_ ) );
INV_X1 _10806_ ( .A(\IF_ID_inst [17] ), .ZN(_03164_ ) );
NOR4_X1 _10807_ ( .A1(_03146_ ), .A2(_03161_ ), .A3(_03164_ ), .A4(_03061_ ), .ZN(_00138_ ) );
AND2_X1 _10808_ ( .A1(_03049_ ), .A2(_03115_ ), .ZN(_03165_ ) );
BUF_X2 _10809_ ( .A(_03165_ ), .Z(_03166_ ) );
NOR2_X1 _10810_ ( .A1(_03153_ ), .A2(\IF_ID_inst [5] ), .ZN(_03167_ ) );
AND2_X2 _10811_ ( .A1(_03166_ ), .A2(_03167_ ), .ZN(_03168_ ) );
AND4_X1 _10812_ ( .A1(\IF_ID_inst [4] ), .A2(_03103_ ), .A3(_03042_ ), .A4(\IF_ID_inst [12] ), .ZN(_03169_ ) );
AND2_X1 _10813_ ( .A1(_03049_ ), .A2(_03169_ ), .ZN(_03170_ ) );
AND2_X1 _10814_ ( .A1(_03170_ ), .A2(\IF_ID_inst [13] ), .ZN(_03171_ ) );
AND3_X1 _10815_ ( .A1(_03043_ ), .A2(_03104_ ), .A3(_03082_ ), .ZN(_03172_ ) );
AND2_X1 _10816_ ( .A1(_03172_ ), .A2(_03152_ ), .ZN(_03173_ ) );
NOR4_X1 _10817_ ( .A1(_03108_ ), .A2(_03168_ ), .A3(_03171_ ), .A4(_03173_ ), .ZN(_03174_ ) );
BUF_X2 _10818_ ( .A(_03170_ ), .Z(_03175_ ) );
NOR3_X1 _10819_ ( .A1(\IF_ID_inst [30] ), .A2(\IF_ID_inst [29] ), .A3(\IF_ID_inst [28] ), .ZN(_03176_ ) );
AND3_X1 _10820_ ( .A1(_03176_ ), .A2(_03070_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03177_ ) );
INV_X1 _10821_ ( .A(\IF_ID_inst [14] ), .ZN(_03178_ ) );
NOR2_X1 _10822_ ( .A1(_03178_ ), .A2(\IF_ID_inst [13] ), .ZN(_03179_ ) );
AND2_X2 _10823_ ( .A1(_03179_ ), .A2(_03098_ ), .ZN(_03180_ ) );
AND2_X2 _10824_ ( .A1(_03177_ ), .A2(_03180_ ), .ZN(_03181_ ) );
NOR2_X1 _10825_ ( .A1(_03063_ ), .A2(\IF_ID_inst [29] ), .ZN(_03182_ ) );
NOR2_X1 _10826_ ( .A1(\IF_ID_inst [28] ), .A2(\IF_ID_inst [27] ), .ZN(_03183_ ) );
AND3_X1 _10827_ ( .A1(_03182_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03183_ ), .ZN(_03184_ ) );
AND2_X1 _10828_ ( .A1(_03184_ ), .A2(_03180_ ), .ZN(_03185_ ) );
OAI21_X1 _10829_ ( .A(_03175_ ), .B1(_03181_ ), .B2(_03185_ ), .ZN(_03186_ ) );
AND2_X1 _10830_ ( .A1(_03165_ ), .A2(_03109_ ), .ZN(_03187_ ) );
AND2_X1 _10831_ ( .A1(_03187_ ), .A2(_03118_ ), .ZN(_03188_ ) );
INV_X1 _10832_ ( .A(_03188_ ), .ZN(_03189_ ) );
AND4_X1 _10833_ ( .A1(_03124_ ), .A2(_03174_ ), .A3(_03186_ ), .A4(_03189_ ), .ZN(_03190_ ) );
NOR2_X1 _10834_ ( .A1(_03146_ ), .A2(_03161_ ), .ZN(_03191_ ) );
AND2_X2 _10835_ ( .A1(_03176_ ), .A2(_03070_ ), .ZN(_03192_ ) );
AND4_X1 _10836_ ( .A1(\IF_ID_inst [13] ), .A2(_03098_ ), .A3(_03178_ ), .A4(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03193_ ) );
AND2_X1 _10837_ ( .A1(_03192_ ), .A2(_03193_ ), .ZN(_03194_ ) );
AND3_X1 _10838_ ( .A1(_03194_ ), .A2(_03053_ ), .A3(_03166_ ), .ZN(_03195_ ) );
AND2_X1 _10839_ ( .A1(_03082_ ), .A2(_03098_ ), .ZN(_03196_ ) );
AND4_X1 _10840_ ( .A1(_03053_ ), .A2(_03166_ ), .A3(_03184_ ), .A4(_03196_ ), .ZN(_03197_ ) );
NOR2_X1 _10841_ ( .A1(_03195_ ), .A2(_03197_ ), .ZN(_03198_ ) );
INV_X1 _10842_ ( .A(_03198_ ), .ZN(_03199_ ) );
AND2_X1 _10843_ ( .A1(_03143_ ), .A2(_03049_ ), .ZN(_03200_ ) );
AND2_X1 _10844_ ( .A1(_03200_ ), .A2(_03117_ ), .ZN(_03201_ ) );
INV_X1 _10845_ ( .A(_03201_ ), .ZN(_03202_ ) );
NAND3_X1 _10846_ ( .A1(_03166_ ), .A2(_03117_ ), .A3(_03109_ ), .ZN(_03203_ ) );
NAND2_X1 _10847_ ( .A1(_03202_ ), .A2(_03203_ ), .ZN(_03204_ ) );
AND3_X1 _10848_ ( .A1(_03175_ ), .A2(_03177_ ), .A3(_03196_ ), .ZN(_03205_ ) );
NOR4_X1 _10849_ ( .A1(_03199_ ), .A2(_03204_ ), .A3(_03066_ ), .A4(_03205_ ), .ZN(_03206_ ) );
AND4_X1 _10850_ ( .A1(_03136_ ), .A2(_03190_ ), .A3(_03191_ ), .A4(_03206_ ), .ZN(_03207_ ) );
AND2_X1 _10851_ ( .A1(_03166_ ), .A2(_03053_ ), .ZN(_03208_ ) );
AND2_X1 _10852_ ( .A1(_03208_ ), .A2(_03181_ ), .ZN(_03209_ ) );
AND2_X2 _10853_ ( .A1(\IF_ID_inst [13] ), .A2(\IF_ID_inst [14] ), .ZN(_03210_ ) );
AND3_X1 _10854_ ( .A1(_03210_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .A3(_03098_ ), .ZN(_03211_ ) );
AND3_X1 _10855_ ( .A1(_03211_ ), .A2(_03070_ ), .A3(_03176_ ), .ZN(_03212_ ) );
NAND3_X1 _10856_ ( .A1(_03212_ ), .A2(_03053_ ), .A3(_03166_ ), .ZN(_03213_ ) );
AND4_X1 _10857_ ( .A1(\IF_ID_inst [4] ), .A2(_03042_ ), .A3(\IF_ID_inst [5] ), .A4(\IF_ID_inst [12] ), .ZN(_03214_ ) );
AND2_X1 _10858_ ( .A1(_03084_ ), .A2(_03214_ ), .ZN(_03215_ ) );
NAND3_X1 _10859_ ( .A1(_03215_ ), .A2(_03192_ ), .A3(_03211_ ), .ZN(_03216_ ) );
NAND2_X1 _10860_ ( .A1(_03213_ ), .A2(_03216_ ), .ZN(_03217_ ) );
AND4_X1 _10861_ ( .A1(_03053_ ), .A2(_03166_ ), .A3(_03177_ ), .A4(_03196_ ), .ZN(_03218_ ) );
NOR3_X1 _10862_ ( .A1(_03209_ ), .A2(_03217_ ), .A3(_03218_ ), .ZN(_03219_ ) );
AND2_X1 _10863_ ( .A1(_03185_ ), .A2(_03215_ ), .ZN(_03220_ ) );
INV_X1 _10864_ ( .A(_03220_ ), .ZN(_03221_ ) );
AND3_X1 _10865_ ( .A1(_03082_ ), .A2(_03098_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03222_ ) );
AND2_X1 _10866_ ( .A1(_03192_ ), .A2(_03222_ ), .ZN(_03223_ ) );
NOR3_X1 _10867_ ( .A1(_03181_ ), .A2(_03194_ ), .A3(_03223_ ), .ZN(_03224_ ) );
INV_X1 _10868_ ( .A(_03215_ ), .ZN(_03225_ ) );
OR2_X1 _10869_ ( .A1(_03224_ ), .A2(_03225_ ), .ZN(_03226_ ) );
AND3_X1 _10870_ ( .A1(_03219_ ), .A2(_03221_ ), .A3(_03226_ ), .ZN(_03227_ ) );
AND2_X2 _10871_ ( .A1(_03207_ ), .A2(_03227_ ), .ZN(_03228_ ) );
XOR2_X1 _10872_ ( .A(\IF_ID_pc [20] ), .B(\myexu.pc_jump [20] ), .Z(_03229_ ) );
XOR2_X1 _10873_ ( .A(\IF_ID_pc [22] ), .B(\myexu.pc_jump [22] ), .Z(_03230_ ) );
XOR2_X1 _10874_ ( .A(\IF_ID_pc [23] ), .B(\myexu.pc_jump [23] ), .Z(_03231_ ) );
XOR2_X1 _10875_ ( .A(\IF_ID_pc [21] ), .B(\myexu.pc_jump [21] ), .Z(_03232_ ) );
OR4_X1 _10876_ ( .A1(_03229_ ), .A2(_03230_ ), .A3(_03231_ ), .A4(_03232_ ), .ZN(_03233_ ) );
XOR2_X1 _10877_ ( .A(\IF_ID_pc [16] ), .B(\myexu.pc_jump [16] ), .Z(_03234_ ) );
XNOR2_X1 _10878_ ( .A(\IF_ID_pc [19] ), .B(\myexu.pc_jump [19] ), .ZN(_03235_ ) );
XNOR2_X1 _10879_ ( .A(\IF_ID_pc [18] ), .B(\myexu.pc_jump [18] ), .ZN(_03236_ ) );
NAND2_X1 _10880_ ( .A1(_03235_ ), .A2(_03236_ ), .ZN(_03237_ ) );
XOR2_X1 _10881_ ( .A(\IF_ID_pc [17] ), .B(\myexu.pc_jump [17] ), .Z(_03238_ ) );
NOR4_X1 _10882_ ( .A1(_03233_ ), .A2(_03234_ ), .A3(_03237_ ), .A4(_03238_ ), .ZN(_03239_ ) );
XNOR2_X1 _10883_ ( .A(\IF_ID_pc [9] ), .B(\myexu.pc_jump [9] ), .ZN(_03240_ ) );
XNOR2_X1 _10884_ ( .A(\IF_ID_pc [8] ), .B(\myexu.pc_jump [8] ), .ZN(_03241_ ) );
XNOR2_X1 _10885_ ( .A(\IF_ID_pc [11] ), .B(\myexu.pc_jump [11] ), .ZN(_03242_ ) );
XNOR2_X1 _10886_ ( .A(\IF_ID_pc [10] ), .B(\myexu.pc_jump [10] ), .ZN(_03243_ ) );
NAND4_X1 _10887_ ( .A1(_03240_ ), .A2(_03241_ ), .A3(_03242_ ), .A4(_03243_ ), .ZN(_03244_ ) );
XNOR2_X1 _10888_ ( .A(\IF_ID_pc [14] ), .B(\myexu.pc_jump [14] ), .ZN(_03245_ ) );
XNOR2_X1 _10889_ ( .A(\IF_ID_pc [15] ), .B(\myexu.pc_jump [15] ), .ZN(_03246_ ) );
NAND2_X1 _10890_ ( .A1(_03245_ ), .A2(_03246_ ), .ZN(_03247_ ) );
XOR2_X1 _10891_ ( .A(\IF_ID_pc [13] ), .B(\myexu.pc_jump [13] ), .Z(_03248_ ) );
XOR2_X1 _10892_ ( .A(\IF_ID_pc [12] ), .B(\myexu.pc_jump [12] ), .Z(_03249_ ) );
NOR4_X1 _10893_ ( .A1(_03244_ ), .A2(_03247_ ), .A3(_03248_ ), .A4(_03249_ ), .ZN(_03250_ ) );
XNOR2_X1 _10894_ ( .A(\myexu.pc_jump [0] ), .B(\IF_ID_pc [0] ), .ZN(_03251_ ) );
XNOR2_X1 _10895_ ( .A(fanout_net_12 ), .B(\myexu.pc_jump [3] ), .ZN(_03252_ ) );
XNOR2_X1 _10896_ ( .A(\myexu.pc_jump [2] ), .B(\IF_ID_pc [2] ), .ZN(_03253_ ) );
XNOR2_X1 _10897_ ( .A(\myexu.pc_jump [1] ), .B(\IF_ID_pc [1] ), .ZN(_03254_ ) );
AND4_X1 _10898_ ( .A1(_03251_ ), .A2(_03252_ ), .A3(_03253_ ), .A4(_03254_ ), .ZN(_03255_ ) );
XNOR2_X1 _10899_ ( .A(\IF_ID_pc [5] ), .B(\myexu.pc_jump [5] ), .ZN(_03256_ ) );
XNOR2_X1 _10900_ ( .A(\IF_ID_pc [7] ), .B(\myexu.pc_jump [7] ), .ZN(_03257_ ) );
XNOR2_X1 _10901_ ( .A(\IF_ID_pc [6] ), .B(\myexu.pc_jump [6] ), .ZN(_03258_ ) );
XNOR2_X1 _10902_ ( .A(fanout_net_16 ), .B(\myexu.pc_jump [4] ), .ZN(_03259_ ) );
AND4_X1 _10903_ ( .A1(_03256_ ), .A2(_03257_ ), .A3(_03258_ ), .A4(_03259_ ), .ZN(_03260_ ) );
AND3_X1 _10904_ ( .A1(_03250_ ), .A2(_03255_ ), .A3(_03260_ ), .ZN(_03261_ ) );
XNOR2_X1 _10905_ ( .A(\IF_ID_pc [24] ), .B(\myexu.pc_jump [24] ), .ZN(_03262_ ) );
XNOR2_X1 _10906_ ( .A(\IF_ID_pc [31] ), .B(\myexu.pc_jump [31] ), .ZN(_03263_ ) );
XNOR2_X1 _10907_ ( .A(\IF_ID_pc [30] ), .B(\myexu.pc_jump [30] ), .ZN(_03264_ ) );
XNOR2_X1 _10908_ ( .A(\IF_ID_pc [28] ), .B(\myexu.pc_jump [28] ), .ZN(_03265_ ) );
XNOR2_X1 _10909_ ( .A(\IF_ID_pc [29] ), .B(\myexu.pc_jump [29] ), .ZN(_03266_ ) );
AND4_X1 _10910_ ( .A1(_03263_ ), .A2(_03264_ ), .A3(_03265_ ), .A4(_03266_ ), .ZN(_03267_ ) );
XNOR2_X1 _10911_ ( .A(\IF_ID_pc [25] ), .B(\myexu.pc_jump [25] ), .ZN(_03268_ ) );
XOR2_X1 _10912_ ( .A(\IF_ID_pc [27] ), .B(\myexu.pc_jump [27] ), .Z(_03269_ ) );
XOR2_X1 _10913_ ( .A(\IF_ID_pc [26] ), .B(\myexu.pc_jump [26] ), .Z(_03270_ ) );
NOR2_X1 _10914_ ( .A1(_03269_ ), .A2(_03270_ ), .ZN(_03271_ ) );
AND4_X1 _10915_ ( .A1(_03262_ ), .A2(_03267_ ), .A3(_03268_ ), .A4(_03271_ ), .ZN(_03272_ ) );
NAND3_X1 _10916_ ( .A1(_03239_ ), .A2(_03261_ ), .A3(_03272_ ), .ZN(_03273_ ) );
AND2_X1 _10917_ ( .A1(_03273_ ), .A2(check_quest ), .ZN(_03274_ ) );
INV_X1 _10918_ ( .A(\myifu.state [1] ), .ZN(_03275_ ) );
NOR2_X1 _10919_ ( .A1(_03275_ ), .A2(fanout_net_49 ), .ZN(_03276_ ) );
INV_X1 _10920_ ( .A(_03276_ ), .ZN(_03277_ ) );
NOR2_X1 _10921_ ( .A1(_03274_ ), .A2(_03277_ ), .ZN(_03278_ ) );
AND2_X2 _10922_ ( .A1(_03278_ ), .A2(IDU_ready_IFU ), .ZN(_03279_ ) );
INV_X1 _10923_ ( .A(_03279_ ), .ZN(_03280_ ) );
BUF_X4 _10924_ ( .A(_03280_ ), .Z(_03281_ ) );
AOI211_X1 _10925_ ( .A(_03228_ ), .B(_03281_ ), .C1(\IF_ID_inst [18] ), .C2(_03191_ ), .ZN(_03282_ ) );
INV_X1 _10926_ ( .A(_03228_ ), .ZN(_03283_ ) );
NAND2_X1 _10927_ ( .A1(_03283_ ), .A2(_03279_ ), .ZN(_03284_ ) );
AOI211_X1 _10928_ ( .A(_03061_ ), .B(_03282_ ), .C1(_02128_ ), .C2(_03284_ ), .ZN(_00139_ ) );
INV_X1 _10929_ ( .A(\IF_ID_inst [16] ), .ZN(_03285_ ) );
NOR4_X1 _10930_ ( .A1(_03146_ ), .A2(_03161_ ), .A3(_03285_ ), .A4(_03061_ ), .ZN(_00140_ ) );
AOI211_X1 _10931_ ( .A(_03228_ ), .B(_03280_ ), .C1(\IF_ID_inst [17] ), .C2(_03191_ ), .ZN(_03286_ ) );
AOI211_X1 _10932_ ( .A(_03061_ ), .B(_03286_ ), .C1(_02135_ ), .C2(_03284_ ), .ZN(_00141_ ) );
NOR4_X1 _10933_ ( .A1(_03146_ ), .A2(_03161_ ), .A3(_03080_ ), .A4(_03061_ ), .ZN(_00142_ ) );
BUF_X4 _10934_ ( .A(_03228_ ), .Z(_03287_ ) );
AOI211_X1 _10935_ ( .A(_03287_ ), .B(_03281_ ), .C1(\IF_ID_inst [16] ), .C2(_03191_ ), .ZN(_03288_ ) );
NOR2_X1 _10936_ ( .A1(_03281_ ), .A2(_03287_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
OAI21_X1 _10937_ ( .A(_03077_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [1] ), .ZN(_03289_ ) );
NOR2_X1 _10938_ ( .A1(_03288_ ), .A2(_03289_ ), .ZN(_00143_ ) );
AND2_X1 _10939_ ( .A1(_03170_ ), .A2(_03118_ ), .ZN(_03290_ ) );
AOI21_X1 _10940_ ( .A(_03290_ ), .B1(_03179_ ), .B2(_03168_ ), .ZN(_03291_ ) );
NAND4_X1 _10941_ ( .A1(_03192_ ), .A2(_03180_ ), .A3(_03084_ ), .A4(_03169_ ), .ZN(_03292_ ) );
INV_X1 _10942_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03293_ ) );
BUF_X2 _10943_ ( .A(_03293_ ), .Z(_03294_ ) );
NOR2_X1 _10944_ ( .A1(_03292_ ), .A2(_03294_ ), .ZN(_03295_ ) );
NAND4_X1 _10945_ ( .A1(_03192_ ), .A2(_03084_ ), .A3(_03196_ ), .A4(_03169_ ), .ZN(_03296_ ) );
NOR2_X1 _10946_ ( .A1(_03296_ ), .A2(_03294_ ), .ZN(_03297_ ) );
NOR2_X1 _10947_ ( .A1(_03295_ ), .A2(_03297_ ), .ZN(_03298_ ) );
AND2_X1 _10948_ ( .A1(_03291_ ), .A2(_03298_ ), .ZN(_03299_ ) );
INV_X1 _10949_ ( .A(_03159_ ), .ZN(_03300_ ) );
NAND2_X1 _10950_ ( .A1(_03168_ ), .A2(_03107_ ), .ZN(_03301_ ) );
OAI21_X1 _10951_ ( .A(_03210_ ), .B1(_03168_ ), .B2(_03175_ ), .ZN(_03302_ ) );
NAND4_X1 _10952_ ( .A1(_03299_ ), .A2(_03300_ ), .A3(_03301_ ), .A4(_03302_ ), .ZN(_03303_ ) );
NAND2_X1 _10953_ ( .A1(_03168_ ), .A2(_03118_ ), .ZN(_03304_ ) );
NAND4_X1 _10954_ ( .A1(_03175_ ), .A2(_03180_ ), .A3(_03182_ ), .A4(_03183_ ), .ZN(_03305_ ) );
OAI21_X1 _10955_ ( .A(_03304_ ), .B1(_03294_ ), .B2(_03305_ ), .ZN(_03306_ ) );
OR4_X2 _10956_ ( .A1(_03155_ ), .A2(_03303_ ), .A3(_03204_ ), .A4(_03306_ ), .ZN(_03307_ ) );
AND4_X1 _10957_ ( .A1(_03097_ ), .A2(_03092_ ), .A3(_03094_ ), .A4(_03100_ ), .ZN(_03308_ ) );
AND3_X1 _10958_ ( .A1(_03084_ ), .A2(_03115_ ), .A3(_03109_ ), .ZN(_03309_ ) );
AOI22_X1 _10959_ ( .A1(_03139_ ), .A2(_03308_ ), .B1(_03118_ ), .B2(_03309_ ), .ZN(_03310_ ) );
AND4_X1 _10960_ ( .A1(_03046_ ), .A2(_03043_ ), .A3(_03104_ ), .A4(_03151_ ), .ZN(_03311_ ) );
NAND2_X1 _10961_ ( .A1(_03311_ ), .A2(_03107_ ), .ZN(_03312_ ) );
AND3_X1 _10962_ ( .A1(_03310_ ), .A2(_03145_ ), .A3(_03312_ ), .ZN(_03313_ ) );
OAI21_X1 _10963_ ( .A(_03054_ ), .B1(_03107_ ), .B2(_03179_ ), .ZN(_03314_ ) );
AND3_X1 _10964_ ( .A1(_03084_ ), .A2(_03053_ ), .A3(_03043_ ), .ZN(_03315_ ) );
OAI21_X1 _10965_ ( .A(_03315_ ), .B1(_03118_ ), .B2(_03210_ ), .ZN(_03316_ ) );
AOI22_X1 _10966_ ( .A1(_03139_ ), .A2(_03141_ ), .B1(\IF_ID_inst [13] ), .B2(_03054_ ), .ZN(_03317_ ) );
NAND4_X1 _10967_ ( .A1(_03313_ ), .A2(_03314_ ), .A3(_03316_ ), .A4(_03317_ ), .ZN(_03318_ ) );
NOR4_X1 _10968_ ( .A1(_03307_ ), .A2(_03073_ ), .A3(_03074_ ), .A4(_03318_ ), .ZN(_00144_ ) );
AOI211_X1 _10969_ ( .A(_03287_ ), .B(_03281_ ), .C1(\IF_ID_inst [15] ), .C2(_03191_ ), .ZN(_03319_ ) );
OAI21_X1 _10970_ ( .A(_03077_ ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .B2(\ID_EX_rs1 [0] ), .ZN(_03320_ ) );
NOR2_X1 _10971_ ( .A1(_03319_ ), .A2(_03320_ ), .ZN(_00145_ ) );
NOR4_X1 _10972_ ( .A1(_03307_ ), .A2(_03075_ ), .A3(_03074_ ), .A4(_03318_ ), .ZN(_00146_ ) );
NOR4_X1 _10973_ ( .A1(_03307_ ), .A2(_03076_ ), .A3(_03074_ ), .A4(_03318_ ), .ZN(_00147_ ) );
NOR2_X1 _10974_ ( .A1(_03307_ ), .A2(_03318_ ), .ZN(_03321_ ) );
AOI211_X1 _10975_ ( .A(_03228_ ), .B(_03280_ ), .C1(\IF_ID_inst [23] ), .C2(_03321_ ), .ZN(_03322_ ) );
INV_X1 _10976_ ( .A(\ID_EX_rs2 [3] ), .ZN(_03323_ ) );
AOI211_X1 _10977_ ( .A(_03061_ ), .B(_03322_ ), .C1(_03323_ ), .C2(_03284_ ), .ZN(_00148_ ) );
NOR4_X1 _10978_ ( .A1(_03307_ ), .A2(_03064_ ), .A3(_03074_ ), .A4(_03318_ ), .ZN(_00149_ ) );
NAND4_X1 _10979_ ( .A1(_03283_ ), .A2(\IF_ID_inst [22] ), .A3(_03279_ ), .A4(_03321_ ), .ZN(_03324_ ) );
OAI21_X1 _10980_ ( .A(\ID_EX_rs2 [2] ), .B1(_03281_ ), .B2(_03287_ ), .ZN(_03325_ ) );
AOI21_X1 _10981_ ( .A(_03065_ ), .B1(_03324_ ), .B2(_03325_ ), .ZN(_00150_ ) );
NOR4_X1 _10982_ ( .A1(_03307_ ), .A2(_03067_ ), .A3(_03074_ ), .A4(_03318_ ), .ZN(_00151_ ) );
NAND4_X1 _10983_ ( .A1(_03283_ ), .A2(\IF_ID_inst [21] ), .A3(_03279_ ), .A4(_03321_ ), .ZN(_03326_ ) );
OAI21_X1 _10984_ ( .A(\ID_EX_rs2 [1] ), .B1(_03281_ ), .B2(_03287_ ), .ZN(_03327_ ) );
AOI21_X1 _10985_ ( .A(_03065_ ), .B1(_03326_ ), .B2(_03327_ ), .ZN(_00152_ ) );
INV_X1 _10986_ ( .A(IDU_valid_EXU ), .ZN(_03328_ ) );
AND3_X1 _10987_ ( .A1(_03113_ ), .A2(_03328_ ), .A3(_03077_ ), .ZN(_00153_ ) );
NAND4_X1 _10988_ ( .A1(_03283_ ), .A2(\IF_ID_inst [20] ), .A3(_03279_ ), .A4(_03321_ ), .ZN(_03329_ ) );
OAI21_X1 _10989_ ( .A(\ID_EX_rs2 [0] ), .B1(_03281_ ), .B2(_03287_ ), .ZN(_03330_ ) );
AOI21_X1 _10990_ ( .A(_03065_ ), .B1(_03329_ ), .B2(_03330_ ), .ZN(_00154_ ) );
OAI21_X1 _10991_ ( .A(_03187_ ), .B1(_03117_ ), .B2(_03178_ ), .ZN(_03331_ ) );
NAND2_X1 _10992_ ( .A1(_03175_ ), .A2(_03210_ ), .ZN(_03332_ ) );
AND3_X1 _10993_ ( .A1(_03175_ ), .A2(\IF_ID_inst [13] ), .A3(_03178_ ), .ZN(_03333_ ) );
INV_X1 _10994_ ( .A(_03333_ ), .ZN(_03334_ ) );
INV_X1 _10995_ ( .A(_03118_ ), .ZN(_03335_ ) );
NAND3_X1 _10996_ ( .A1(_03166_ ), .A2(_03335_ ), .A3(_03167_ ), .ZN(_03336_ ) );
NAND4_X1 _10997_ ( .A1(_03331_ ), .A2(_03332_ ), .A3(_03334_ ), .A4(_03336_ ), .ZN(_03337_ ) );
INV_X1 _10998_ ( .A(_03173_ ), .ZN(_03338_ ) );
NAND3_X1 _10999_ ( .A1(_03304_ ), .A2(_03202_ ), .A3(_03338_ ), .ZN(_03339_ ) );
NOR2_X1 _11000_ ( .A1(_03337_ ), .A2(_03339_ ), .ZN(_03340_ ) );
AND2_X1 _11001_ ( .A1(_03340_ ), .A2(_03055_ ), .ZN(_03341_ ) );
INV_X1 _11002_ ( .A(_03341_ ), .ZN(_03342_ ) );
AND2_X2 _11003_ ( .A1(\ID_EX_typ [6] ), .A2(\ID_EX_typ [5] ), .ZN(_03343_ ) );
INV_X2 _11004_ ( .A(\ID_EX_typ [7] ), .ZN(_03344_ ) );
AND2_X1 _11005_ ( .A1(_03343_ ), .A2(_03344_ ), .ZN(_03345_ ) );
XNOR2_X1 _11006_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [19] ), .ZN(_03346_ ) );
XNOR2_X1 _11007_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [18] ), .ZN(_03347_ ) );
AND3_X1 _11008_ ( .A1(_03345_ ), .A2(_03346_ ), .A3(_03347_ ), .ZN(_03348_ ) );
XNOR2_X1 _11009_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [17] ), .ZN(_03349_ ) );
XNOR2_X1 _11010_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [15] ), .ZN(_03350_ ) );
XNOR2_X1 _11011_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [16] ), .ZN(_03351_ ) );
AND3_X1 _11012_ ( .A1(_03349_ ), .A2(_03350_ ), .A3(_03351_ ), .ZN(_03352_ ) );
NAND2_X1 _11013_ ( .A1(_03348_ ), .A2(_03352_ ), .ZN(_03353_ ) );
XNOR2_X1 _11014_ ( .A(\ID_EX_rd [2] ), .B(\IF_ID_inst [22] ), .ZN(_03354_ ) );
XNOR2_X1 _11015_ ( .A(\ID_EX_rd [3] ), .B(\IF_ID_inst [23] ), .ZN(_03355_ ) );
XNOR2_X1 _11016_ ( .A(\ID_EX_rd [0] ), .B(\IF_ID_inst [20] ), .ZN(_03356_ ) );
AND4_X1 _11017_ ( .A1(_03345_ ), .A2(_03354_ ), .A3(_03355_ ), .A4(_03356_ ), .ZN(_03357_ ) );
XNOR2_X1 _11018_ ( .A(\ID_EX_rd [4] ), .B(\IF_ID_inst [24] ), .ZN(_03358_ ) );
XNOR2_X1 _11019_ ( .A(\ID_EX_rd [1] ), .B(\IF_ID_inst [21] ), .ZN(_03359_ ) );
AND3_X1 _11020_ ( .A1(_03357_ ), .A2(_03358_ ), .A3(_03359_ ), .ZN(_03360_ ) );
INV_X1 _11021_ ( .A(_03360_ ), .ZN(_03361_ ) );
AOI211_X1 _11022_ ( .A(_03161_ ), .B(_03146_ ), .C1(_03353_ ), .C2(_03361_ ), .ZN(_03362_ ) );
OAI211_X1 _11023_ ( .A(IDU_ready_IFU ), .B(_03077_ ), .C1(_03342_ ), .C2(_03362_ ), .ZN(_03363_ ) );
AOI21_X1 _11024_ ( .A(_03341_ ), .B1(_03352_ ), .B2(_03348_ ), .ZN(_03364_ ) );
NOR2_X1 _11025_ ( .A1(_03363_ ), .A2(_03364_ ), .ZN(_00155_ ) );
AND2_X1 _11026_ ( .A1(_03139_ ), .A2(_03308_ ), .ZN(_03365_ ) );
INV_X1 _11027_ ( .A(_03365_ ), .ZN(_03366_ ) );
NOR2_X1 _11028_ ( .A1(_03173_ ), .A2(_03159_ ), .ZN(_03367_ ) );
OAI21_X1 _11029_ ( .A(_03335_ ), .B1(_03106_ ), .B2(_03132_ ), .ZN(_03368_ ) );
AND4_X1 _11030_ ( .A1(_03366_ ), .A2(_03145_ ), .A3(_03367_ ), .A4(_03368_ ), .ZN(_03369_ ) );
AND4_X1 _11031_ ( .A1(_03067_ ), .A2(_03083_ ), .A3(_03084_ ), .A4(_03089_ ), .ZN(_03370_ ) );
NOR2_X1 _11032_ ( .A1(_03125_ ), .A2(_03126_ ), .ZN(_03371_ ) );
AND3_X1 _11033_ ( .A1(_03371_ ), .A2(_03064_ ), .A3(_03128_ ), .ZN(_03372_ ) );
NAND2_X1 _11034_ ( .A1(_03370_ ), .A2(_03372_ ), .ZN(_03373_ ) );
AND2_X1 _11035_ ( .A1(_03373_ ), .A2(_03055_ ), .ZN(_03374_ ) );
AOI21_X1 _11036_ ( .A(_03065_ ), .B1(_03369_ ), .B2(_03374_ ), .ZN(_00156_ ) );
NAND2_X1 _11037_ ( .A1(_03200_ ), .A2(_03107_ ), .ZN(_03375_ ) );
NAND3_X1 _11038_ ( .A1(_03200_ ), .A2(_03117_ ), .A3(\IF_ID_inst [14] ), .ZN(_03376_ ) );
AND4_X1 _11039_ ( .A1(_03124_ ), .A2(_03375_ ), .A3(_03331_ ), .A4(_03376_ ), .ZN(_03377_ ) );
AOI21_X1 _11040_ ( .A(_03065_ ), .B1(_03377_ ), .B2(_03374_ ), .ZN(_00157_ ) );
NAND3_X1 _11041_ ( .A1(_03192_ ), .A2(_03210_ ), .A3(_03098_ ), .ZN(_03378_ ) );
INV_X1 _11042_ ( .A(_03208_ ), .ZN(_03379_ ) );
AOI211_X1 _11043_ ( .A(_03294_ ), .B(_03378_ ), .C1(_03379_ ), .C2(_03225_ ), .ZN(_03380_ ) );
OAI211_X1 _11044_ ( .A(_03053_ ), .B(_03166_ ), .C1(_03181_ ), .C2(_03223_ ), .ZN(_03381_ ) );
OAI21_X1 _11045_ ( .A(_03381_ ), .B1(_03224_ ), .B2(_03225_ ), .ZN(_03382_ ) );
NOR2_X1 _11046_ ( .A1(_03380_ ), .A2(_03382_ ), .ZN(_03383_ ) );
INV_X1 _11047_ ( .A(_03383_ ), .ZN(_03384_ ) );
INV_X1 _11048_ ( .A(_03171_ ), .ZN(_03385_ ) );
NAND2_X1 _11049_ ( .A1(_03385_ ), .A2(_03336_ ), .ZN(_03386_ ) );
AOI22_X1 _11050_ ( .A1(_03370_ ), .A2(_03372_ ), .B1(_03215_ ), .B2(_03185_ ), .ZN(_03387_ ) );
AND2_X1 _11051_ ( .A1(_03184_ ), .A2(_03196_ ), .ZN(_03388_ ) );
OR2_X1 _11052_ ( .A1(_03388_ ), .A2(_03194_ ), .ZN(_03389_ ) );
NAND2_X1 _11053_ ( .A1(_03389_ ), .A2(_03208_ ), .ZN(_03390_ ) );
NAND4_X1 _11054_ ( .A1(_03387_ ), .A2(_03189_ ), .A3(_03390_ ), .A4(_03367_ ), .ZN(_03391_ ) );
NOR4_X1 _11055_ ( .A1(_03384_ ), .A2(_03204_ ), .A3(_03386_ ), .A4(_03391_ ), .ZN(_03392_ ) );
INV_X1 _11056_ ( .A(_03205_ ), .ZN(_03393_ ) );
AND2_X1 _11057_ ( .A1(_03393_ ), .A2(_03186_ ), .ZN(_03394_ ) );
INV_X1 _11058_ ( .A(_03155_ ), .ZN(_03395_ ) );
AND2_X1 _11059_ ( .A1(_03304_ ), .A2(_03395_ ), .ZN(_03396_ ) );
AND2_X1 _11060_ ( .A1(_03394_ ), .A2(_03396_ ), .ZN(_03397_ ) );
AOI21_X1 _11061_ ( .A(_03065_ ), .B1(_03392_ ), .B2(_03397_ ), .ZN(_00158_ ) );
AOI221_X4 _11062_ ( .A(_03113_ ), .B1(\IF_ID_inst [13] ), .B2(_03175_ ), .C1(_03168_ ), .C2(_03335_ ), .ZN(_03398_ ) );
AOI21_X1 _11063_ ( .A(_03062_ ), .B1(_03397_ ), .B2(_03398_ ), .ZN(_00159_ ) );
NOR4_X1 _11064_ ( .A1(_03102_ ), .A2(_03195_ ), .A3(_03197_ ), .A4(_03119_ ), .ZN(_03399_ ) );
AOI21_X1 _11065_ ( .A(_03062_ ), .B1(_03399_ ), .B2(_03396_ ), .ZN(_00160_ ) );
OR2_X1 _11066_ ( .A1(_03188_ ), .A2(_03290_ ), .ZN(_03400_ ) );
OAI21_X1 _11067_ ( .A(_03221_ ), .B1(_03224_ ), .B2(_03225_ ), .ZN(_03401_ ) );
NOR4_X1 _11068_ ( .A1(_03400_ ), .A2(_03401_ ), .A3(_03119_ ), .A4(_03155_ ), .ZN(_03402_ ) );
NAND3_X1 _11069_ ( .A1(_03175_ ), .A2(_03192_ ), .A3(_03222_ ), .ZN(_03403_ ) );
NAND3_X1 _11070_ ( .A1(_03175_ ), .A2(_03180_ ), .A3(_03184_ ), .ZN(_03404_ ) );
NAND4_X1 _11071_ ( .A1(_03177_ ), .A2(_03084_ ), .A3(_03180_ ), .A4(_03169_ ), .ZN(_03405_ ) );
NAND3_X1 _11072_ ( .A1(_03403_ ), .A2(_03404_ ), .A3(_03405_ ), .ZN(_03406_ ) );
AOI221_X4 _11073_ ( .A(_03406_ ), .B1(\IF_ID_inst [13] ), .B2(_03054_ ), .C1(\IF_ID_inst [14] ), .C2(_03132_ ), .ZN(_03407_ ) );
AOI21_X1 _11074_ ( .A(_03062_ ), .B1(_03402_ ), .B2(_03407_ ), .ZN(_00161_ ) );
AND2_X1 _11075_ ( .A1(_03122_ ), .A2(_03107_ ), .ZN(_03408_ ) );
AND3_X1 _11076_ ( .A1(_03042_ ), .A2(\IF_ID_inst [4] ), .A3(\IF_ID_inst [5] ), .ZN(_03409_ ) );
AOI221_X4 _11077_ ( .A(_03408_ ), .B1(_03107_ ), .B2(_03200_ ), .C1(_03152_ ), .C2(_03409_ ), .ZN(_03410_ ) );
INV_X1 _11078_ ( .A(_03209_ ), .ZN(_03411_ ) );
AND4_X1 _11079_ ( .A1(_03120_ ), .A2(_03410_ ), .A3(_03411_ ), .A4(_03376_ ), .ZN(_03412_ ) );
NAND2_X1 _11080_ ( .A1(_03168_ ), .A2(\IF_ID_inst [14] ), .ZN(_03413_ ) );
OAI22_X1 _11081_ ( .A1(_03181_ ), .A2(_03185_ ), .B1(_03215_ ), .B2(_03175_ ), .ZN(_03414_ ) );
AOI22_X1 _11082_ ( .A1(_03106_ ), .A2(\IF_ID_inst [14] ), .B1(_03084_ ), .B2(_03045_ ), .ZN(_03415_ ) );
AND4_X1 _11083_ ( .A1(_03213_ ), .A2(_03413_ ), .A3(_03414_ ), .A4(_03415_ ), .ZN(_03416_ ) );
AOI21_X1 _11084_ ( .A(_03062_ ), .B1(_03412_ ), .B2(_03416_ ), .ZN(_00162_ ) );
OAI211_X1 _11085_ ( .A(_03117_ ), .B(\IF_ID_inst [14] ), .C1(_03168_ ), .C2(_03054_ ), .ZN(_03417_ ) );
AOI21_X1 _11086_ ( .A(_03205_ ), .B1(_03181_ ), .B2(_03208_ ), .ZN(_03418_ ) );
AND3_X1 _11087_ ( .A1(_03130_ ), .A2(_03123_ ), .A3(_03418_ ), .ZN(_03419_ ) );
NAND4_X1 _11088_ ( .A1(_03177_ ), .A2(_03084_ ), .A3(_03214_ ), .A4(_03196_ ), .ZN(_03420_ ) );
AOI221_X4 _11089_ ( .A(_03119_ ), .B1(_03107_ ), .B2(_03132_ ), .C1(\IF_ID_inst [14] ), .C2(_03201_ ), .ZN(_03421_ ) );
AND4_X1 _11090_ ( .A1(_03417_ ), .A2(_03419_ ), .A3(_03420_ ), .A4(_03421_ ), .ZN(_03422_ ) );
INV_X1 _11091_ ( .A(_03133_ ), .ZN(_03423_ ) );
NAND2_X1 _11092_ ( .A1(_03404_ ), .A2(_03332_ ), .ZN(_03424_ ) );
AOI221_X4 _11093_ ( .A(_03424_ ), .B1(\IF_ID_inst [14] ), .B2(_03050_ ), .C1(_03179_ ), .C2(_03187_ ), .ZN(_03425_ ) );
AND3_X1 _11094_ ( .A1(_03215_ ), .A2(_03192_ ), .A3(_03211_ ), .ZN(_03426_ ) );
NOR4_X1 _11095_ ( .A1(_03195_ ), .A2(_03220_ ), .A3(_03426_ ), .A4(_03173_ ), .ZN(_03427_ ) );
OAI21_X1 _11096_ ( .A(_03210_ ), .B1(_03106_ ), .B2(_03054_ ), .ZN(_03428_ ) );
AND4_X1 _11097_ ( .A1(_03423_ ), .A2(_03425_ ), .A3(_03427_ ), .A4(_03428_ ), .ZN(_03429_ ) );
AOI21_X1 _11098_ ( .A(_03062_ ), .B1(_03422_ ), .B2(_03429_ ), .ZN(_00163_ ) );
INV_X1 _11099_ ( .A(fanout_net_49 ), .ZN(_03430_ ) );
BUF_X4 _11100_ ( .A(_03430_ ), .Z(_03431_ ) );
NAND4_X1 _11101_ ( .A1(_03273_ ), .A2(check_quest ), .A3(\myexu.pc_jump [0] ), .A4(_03431_ ), .ZN(_03432_ ) );
NAND2_X1 _11102_ ( .A1(\mtvec [0] ), .A2(fanout_net_49 ), .ZN(_03433_ ) );
AOI21_X1 _11103_ ( .A(fanout_net_2 ), .B1(_03432_ ), .B2(_03433_ ), .ZN(_00167_ ) );
INV_X1 _11104_ ( .A(_03274_ ), .ZN(_03434_ ) );
BUF_X4 _11105_ ( .A(_03434_ ), .Z(_03435_ ) );
AND4_X2 _11106_ ( .A1(\IF_ID_inst [31] ), .A2(_03153_ ), .A3(_03156_ ), .A4(\IF_ID_inst [5] ), .ZN(_03436_ ) );
AND2_X1 _11107_ ( .A1(_03048_ ), .A2(_03436_ ), .ZN(_03437_ ) );
BUF_X4 _11108_ ( .A(_03437_ ), .Z(_03438_ ) );
AND2_X1 _11109_ ( .A1(_03438_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03439_ ) );
CLKBUF_X2 _11110_ ( .A(_03157_ ), .Z(_03440_ ) );
OAI211_X1 _11111_ ( .A(_03440_ ), .B(\IF_ID_inst [31] ), .C1(_03112_ ), .C2(_03048_ ), .ZN(_03441_ ) );
NOR2_X1 _11112_ ( .A1(_03439_ ), .A2(_03441_ ), .ZN(_03442_ ) );
BUF_X4 _11113_ ( .A(_03442_ ), .Z(_03443_ ) );
BUF_X4 _11114_ ( .A(_03443_ ), .Z(_03444_ ) );
XNOR2_X1 _11115_ ( .A(_03444_ ), .B(_01856_ ), .ZN(_03445_ ) );
INV_X1 _11116_ ( .A(_03445_ ), .ZN(_03446_ ) );
AND3_X1 _11117_ ( .A1(_03440_ ), .A2(_03112_ ), .A3(\IF_ID_inst [18] ), .ZN(_03447_ ) );
MUX2_X1 _11118_ ( .A(_03447_ ), .B(_03294_ ), .S(_03438_ ), .Z(_03448_ ) );
XNOR2_X1 _11119_ ( .A(_03448_ ), .B(_01986_ ), .ZN(_03449_ ) );
AND2_X1 _11120_ ( .A1(_03159_ ), .A2(\IF_ID_inst [20] ), .ZN(_03450_ ) );
INV_X1 _11121_ ( .A(_03450_ ), .ZN(_03451_ ) );
INV_X1 _11122_ ( .A(_03437_ ), .ZN(_03452_ ) );
OAI21_X1 _11123_ ( .A(_03451_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .B2(_03452_ ), .ZN(_03453_ ) );
AND2_X1 _11124_ ( .A1(_03453_ ), .A2(\IF_ID_pc [11] ), .ZN(_03454_ ) );
AND2_X1 _11125_ ( .A1(_03159_ ), .A2(\IF_ID_inst [29] ), .ZN(_03455_ ) );
INV_X1 _11126_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03456_ ) );
AOI21_X1 _11127_ ( .A(_03455_ ), .B1(_03456_ ), .B2(_03437_ ), .ZN(_03457_ ) );
XNOR2_X1 _11128_ ( .A(_03457_ ), .B(\IF_ID_pc [9] ), .ZN(_03458_ ) );
INV_X1 _11129_ ( .A(_03458_ ), .ZN(_03459_ ) );
NAND3_X1 _11130_ ( .A1(_03157_ ), .A2(_03111_ ), .A3(\IF_ID_inst [24] ), .ZN(_03460_ ) );
INV_X1 _11131_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03461_ ) );
NAND3_X1 _11132_ ( .A1(_03048_ ), .A2(_03436_ ), .A3(_03461_ ), .ZN(_03462_ ) );
NAND2_X1 _11133_ ( .A1(_03460_ ), .A2(_03462_ ), .ZN(_03463_ ) );
NAND2_X1 _11134_ ( .A1(_03463_ ), .A2(fanout_net_16 ), .ZN(_03464_ ) );
NAND3_X1 _11135_ ( .A1(_03157_ ), .A2(_03111_ ), .A3(\IF_ID_inst [23] ), .ZN(_03465_ ) );
INV_X1 _11136_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03466_ ) );
NAND3_X1 _11137_ ( .A1(_03048_ ), .A2(_03436_ ), .A3(_03466_ ), .ZN(_03467_ ) );
NAND2_X1 _11138_ ( .A1(_03465_ ), .A2(_03467_ ), .ZN(_03468_ ) );
INV_X1 _11139_ ( .A(_03468_ ), .ZN(_03469_ ) );
OR2_X1 _11140_ ( .A1(_03469_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03470_ ) );
NAND3_X1 _11141_ ( .A1(_03157_ ), .A2(_03111_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_03471_ ) );
NAND3_X1 _11142_ ( .A1(_03048_ ), .A2(_03436_ ), .A3(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03472_ ) );
AND3_X1 _11143_ ( .A1(_03471_ ), .A2(\IF_ID_pc [2] ), .A3(_03472_ ), .ZN(_03473_ ) );
AOI21_X1 _11144_ ( .A(\IF_ID_pc [2] ), .B1(_03471_ ), .B2(_03472_ ), .ZN(_03474_ ) );
NOR2_X1 _11145_ ( .A1(_03473_ ), .A2(_03474_ ), .ZN(_03475_ ) );
NAND3_X1 _11146_ ( .A1(_03157_ ), .A2(_03111_ ), .A3(\IF_ID_inst [21] ), .ZN(_03476_ ) );
INV_X1 _11147_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ), .ZN(_03477_ ) );
NAND3_X1 _11148_ ( .A1(_03048_ ), .A2(_03436_ ), .A3(_03477_ ), .ZN(_03478_ ) );
NAND2_X1 _11149_ ( .A1(_03476_ ), .A2(_03478_ ), .ZN(_03479_ ) );
AND2_X1 _11150_ ( .A1(_03479_ ), .A2(\IF_ID_pc [1] ), .ZN(_03480_ ) );
AND2_X1 _11151_ ( .A1(_03475_ ), .A2(_03480_ ), .ZN(_03481_ ) );
NOR2_X1 _11152_ ( .A1(_03481_ ), .A2(_03473_ ), .ZN(_03482_ ) );
XNOR2_X1 _11153_ ( .A(_03468_ ), .B(fanout_net_12 ), .ZN(_03483_ ) );
OAI211_X1 _11154_ ( .A(_03464_ ), .B(_03470_ ), .C1(_03482_ ), .C2(_03483_ ), .ZN(_03484_ ) );
INV_X1 _11155_ ( .A(fanout_net_16 ), .ZN(_03485_ ) );
NAND3_X1 _11156_ ( .A1(_03460_ ), .A2(_03485_ ), .A3(_03462_ ), .ZN(_03486_ ) );
NAND2_X1 _11157_ ( .A1(_03484_ ), .A2(_03486_ ), .ZN(_03487_ ) );
AND2_X1 _11158_ ( .A1(_03158_ ), .A2(\IF_ID_inst [25] ), .ZN(_03488_ ) );
INV_X1 _11159_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .ZN(_03489_ ) );
AND3_X1 _11160_ ( .A1(_03048_ ), .A2(_03436_ ), .A3(_03489_ ), .ZN(_03490_ ) );
NOR2_X1 _11161_ ( .A1(_03488_ ), .A2(_03490_ ), .ZN(_03491_ ) );
XOR2_X1 _11162_ ( .A(_03491_ ), .B(\IF_ID_pc [5] ), .Z(_03492_ ) );
NOR2_X1 _11163_ ( .A1(_03487_ ), .A2(_03492_ ), .ZN(_03493_ ) );
NOR2_X1 _11164_ ( .A1(_03491_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_03494_ ) );
NOR2_X2 _11165_ ( .A1(_03493_ ), .A2(_03494_ ), .ZN(_03495_ ) );
INV_X1 _11166_ ( .A(\IF_ID_pc [6] ), .ZN(_03496_ ) );
AND2_X1 _11167_ ( .A1(_03159_ ), .A2(\IF_ID_inst [26] ), .ZN(_03497_ ) );
INV_X1 _11168_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03498_ ) );
AOI21_X1 _11169_ ( .A(_03497_ ), .B1(_03498_ ), .B2(_03437_ ), .ZN(_03499_ ) );
OAI21_X1 _11170_ ( .A(_03495_ ), .B1(_03496_ ), .B2(_03499_ ), .ZN(_03500_ ) );
INV_X1 _11171_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_03501_ ) );
AND3_X1 _11172_ ( .A1(_03048_ ), .A2(_03436_ ), .A3(_03501_ ), .ZN(_03502_ ) );
AOI21_X1 _11173_ ( .A(_03502_ ), .B1(\IF_ID_inst [27] ), .B2(_03159_ ), .ZN(_03503_ ) );
XNOR2_X1 _11174_ ( .A(_03503_ ), .B(\IF_ID_pc [7] ), .ZN(_03504_ ) );
NAND2_X1 _11175_ ( .A1(_03499_ ), .A2(_03496_ ), .ZN(_03505_ ) );
AND3_X2 _11176_ ( .A1(_03500_ ), .A2(_03504_ ), .A3(_03505_ ), .ZN(_03506_ ) );
NOR2_X1 _11177_ ( .A1(_03503_ ), .A2(_01869_ ), .ZN(_03507_ ) );
AND2_X1 _11178_ ( .A1(_03159_ ), .A2(\IF_ID_inst [28] ), .ZN(_03508_ ) );
INV_X1 _11179_ ( .A(_03508_ ), .ZN(_03509_ ) );
OAI21_X1 _11180_ ( .A(_03509_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .B2(_03452_ ), .ZN(_03510_ ) );
OAI22_X1 _11181_ ( .A1(_03506_ ), .A2(_03507_ ), .B1(\IF_ID_pc [8] ), .B2(_03510_ ), .ZN(_03511_ ) );
NAND2_X1 _11182_ ( .A1(_03510_ ), .A2(\IF_ID_pc [8] ), .ZN(_03512_ ) );
AOI21_X1 _11183_ ( .A(_03459_ ), .B1(_03511_ ), .B2(_03512_ ), .ZN(_03513_ ) );
NOR2_X1 _11184_ ( .A1(_03457_ ), .A2(_01794_ ), .ZN(_03514_ ) );
NOR2_X1 _11185_ ( .A1(_03513_ ), .A2(_03514_ ), .ZN(_03515_ ) );
INV_X1 _11186_ ( .A(\IF_ID_pc [10] ), .ZN(_03516_ ) );
AND2_X1 _11187_ ( .A1(_03159_ ), .A2(\IF_ID_inst [30] ), .ZN(_03517_ ) );
INV_X1 _11188_ ( .A(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_03518_ ) );
AOI21_X1 _11189_ ( .A(_03517_ ), .B1(_03518_ ), .B2(_03438_ ), .ZN(_03519_ ) );
OAI21_X1 _11190_ ( .A(_03515_ ), .B1(_03516_ ), .B2(_03519_ ), .ZN(_03520_ ) );
INV_X1 _11191_ ( .A(\IF_ID_pc [11] ), .ZN(_03521_ ) );
XNOR2_X1 _11192_ ( .A(_03453_ ), .B(_03521_ ), .ZN(_03522_ ) );
AND2_X1 _11193_ ( .A1(_03519_ ), .A2(_03516_ ), .ZN(_03523_ ) );
INV_X1 _11194_ ( .A(_03523_ ), .ZN(_03524_ ) );
AND3_X1 _11195_ ( .A1(_03520_ ), .A2(_03522_ ), .A3(_03524_ ), .ZN(_03525_ ) );
AND3_X1 _11196_ ( .A1(_03440_ ), .A2(_03112_ ), .A3(\IF_ID_inst [12] ), .ZN(_03526_ ) );
MUX2_X1 _11197_ ( .A(_03526_ ), .B(_03294_ ), .S(_03438_ ), .Z(_03527_ ) );
AOI211_X2 _11198_ ( .A(_03454_ ), .B(_03525_ ), .C1(\IF_ID_pc [12] ), .C2(_03527_ ), .ZN(_03528_ ) );
NOR2_X1 _11199_ ( .A1(_03527_ ), .A2(\IF_ID_pc [12] ), .ZN(_03529_ ) );
NOR2_X1 _11200_ ( .A1(_03528_ ), .A2(_03529_ ), .ZN(_03530_ ) );
NAND3_X1 _11201_ ( .A1(_03440_ ), .A2(_03111_ ), .A3(\IF_ID_inst [16] ), .ZN(_03531_ ) );
MUX2_X1 _11202_ ( .A(_03531_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .S(_03438_ ), .Z(_03532_ ) );
XNOR2_X1 _11203_ ( .A(_03532_ ), .B(_02004_ ), .ZN(_03533_ ) );
AND3_X1 _11204_ ( .A1(_03440_ ), .A2(_03111_ ), .A3(\IF_ID_inst [15] ), .ZN(_03534_ ) );
MUX2_X1 _11205_ ( .A(_03534_ ), .B(_03293_ ), .S(_03438_ ), .Z(_03535_ ) );
XNOR2_X1 _11206_ ( .A(_03535_ ), .B(\IF_ID_pc [15] ), .ZN(_03536_ ) );
NOR2_X1 _11207_ ( .A1(_03533_ ), .A2(_03536_ ), .ZN(_03537_ ) );
NAND3_X1 _11208_ ( .A1(_03440_ ), .A2(_03112_ ), .A3(\IF_ID_inst [14] ), .ZN(_03538_ ) );
MUX2_X1 _11209_ ( .A(_03538_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .S(_03438_ ), .Z(_03539_ ) );
XNOR2_X1 _11210_ ( .A(_03539_ ), .B(\IF_ID_pc [14] ), .ZN(_03540_ ) );
AND3_X1 _11211_ ( .A1(_03440_ ), .A2(_03112_ ), .A3(\IF_ID_inst [13] ), .ZN(_03541_ ) );
MUX2_X1 _11212_ ( .A(_03541_ ), .B(_03293_ ), .S(_03438_ ), .Z(_03542_ ) );
INV_X1 _11213_ ( .A(\IF_ID_pc [13] ), .ZN(_03543_ ) );
XNOR2_X1 _11214_ ( .A(_03542_ ), .B(_03543_ ), .ZN(_03544_ ) );
NAND4_X1 _11215_ ( .A1(_03530_ ), .A2(_03537_ ), .A3(_03540_ ), .A4(_03544_ ), .ZN(_03545_ ) );
AND2_X1 _11216_ ( .A1(_03535_ ), .A2(\IF_ID_pc [15] ), .ZN(_03546_ ) );
INV_X1 _11217_ ( .A(_03546_ ), .ZN(_03547_ ) );
OR2_X1 _11218_ ( .A1(_03533_ ), .A2(_03547_ ), .ZN(_03548_ ) );
OAI21_X1 _11219_ ( .A(_03548_ ), .B1(_02004_ ), .B2(_03532_ ), .ZN(_03549_ ) );
AND2_X1 _11220_ ( .A1(_03542_ ), .A2(\IF_ID_pc [13] ), .ZN(_03550_ ) );
NAND2_X1 _11221_ ( .A1(_03540_ ), .A2(_03550_ ), .ZN(_03551_ ) );
INV_X1 _11222_ ( .A(\IF_ID_pc [14] ), .ZN(_03552_ ) );
OAI21_X1 _11223_ ( .A(_03551_ ), .B1(_03552_ ), .B2(_03539_ ), .ZN(_03553_ ) );
AOI21_X1 _11224_ ( .A(_03549_ ), .B1(_03553_ ), .B2(_03537_ ), .ZN(_03554_ ) );
NAND2_X1 _11225_ ( .A1(_03545_ ), .A2(_03554_ ), .ZN(_03555_ ) );
NAND3_X1 _11226_ ( .A1(_03440_ ), .A2(_03112_ ), .A3(\IF_ID_inst [17] ), .ZN(_03556_ ) );
MUX2_X1 _11227_ ( .A(_03556_ ), .B(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .S(_03438_ ), .Z(_03557_ ) );
XNOR2_X1 _11228_ ( .A(_03557_ ), .B(\IF_ID_pc [17] ), .ZN(_03558_ ) );
AND3_X1 _11229_ ( .A1(_03440_ ), .A2(_03112_ ), .A3(\IF_ID_inst [19] ), .ZN(_03559_ ) );
MUX2_X1 _11230_ ( .A(_03559_ ), .B(_03294_ ), .S(_03438_ ), .Z(_03560_ ) );
XNOR2_X1 _11231_ ( .A(_03560_ ), .B(_02001_ ), .ZN(_03561_ ) );
XNOR2_X1 _11232_ ( .A(_03442_ ), .B(_01863_ ), .ZN(_03562_ ) );
AND2_X1 _11233_ ( .A1(_03561_ ), .A2(_03562_ ), .ZN(_03563_ ) );
AND4_X1 _11234_ ( .A1(_03449_ ), .A2(_03555_ ), .A3(_03558_ ), .A4(_03563_ ), .ZN(_03564_ ) );
AND2_X1 _11235_ ( .A1(_03560_ ), .A2(\IF_ID_pc [19] ), .ZN(_03565_ ) );
AND2_X1 _11236_ ( .A1(_03562_ ), .A2(_03565_ ), .ZN(_03566_ ) );
AOI21_X1 _11237_ ( .A(_03566_ ), .B1(\IF_ID_pc [20] ), .B2(_03442_ ), .ZN(_03567_ ) );
NOR2_X1 _11238_ ( .A1(_03557_ ), .A2(_01759_ ), .ZN(_03568_ ) );
AND2_X1 _11239_ ( .A1(_03449_ ), .A2(_03568_ ), .ZN(_03569_ ) );
AOI21_X1 _11240_ ( .A(_03569_ ), .B1(\IF_ID_pc [18] ), .B2(_03448_ ), .ZN(_03570_ ) );
INV_X1 _11241_ ( .A(_03563_ ), .ZN(_03571_ ) );
OAI21_X1 _11242_ ( .A(_03567_ ), .B1(_03570_ ), .B2(_03571_ ), .ZN(_03572_ ) );
OR2_X4 _11243_ ( .A1(_03564_ ), .A2(_03572_ ), .ZN(_03573_ ) );
XNOR2_X1 _11244_ ( .A(_03442_ ), .B(_01955_ ), .ZN(_03574_ ) );
XNOR2_X1 _11245_ ( .A(_03442_ ), .B(_01898_ ), .ZN(_03575_ ) );
AND2_X1 _11246_ ( .A1(_03574_ ), .A2(_03575_ ), .ZN(_03576_ ) );
XNOR2_X1 _11247_ ( .A(_03442_ ), .B(\IF_ID_pc [21] ), .ZN(_03577_ ) );
XNOR2_X1 _11248_ ( .A(_03443_ ), .B(\IF_ID_pc [22] ), .ZN(_03578_ ) );
NOR2_X1 _11249_ ( .A1(_03577_ ), .A2(_03578_ ), .ZN(_03579_ ) );
AND3_X1 _11250_ ( .A1(_03573_ ), .A2(_03576_ ), .A3(_03579_ ), .ZN(_03580_ ) );
AND2_X1 _11251_ ( .A1(_03443_ ), .A2(\IF_ID_pc [22] ), .ZN(_03581_ ) );
AND2_X1 _11252_ ( .A1(_03443_ ), .A2(\IF_ID_pc [21] ), .ZN(_03582_ ) );
OAI21_X1 _11253_ ( .A(_03576_ ), .B1(_03581_ ), .B2(_03582_ ), .ZN(_03583_ ) );
NAND2_X1 _11254_ ( .A1(_03443_ ), .A2(\IF_ID_pc [24] ), .ZN(_03584_ ) );
NAND2_X1 _11255_ ( .A1(_03443_ ), .A2(\IF_ID_pc [23] ), .ZN(_03585_ ) );
NAND3_X1 _11256_ ( .A1(_03583_ ), .A2(_03584_ ), .A3(_03585_ ), .ZN(_03586_ ) );
NOR2_X1 _11257_ ( .A1(_03580_ ), .A2(_03586_ ), .ZN(_03587_ ) );
INV_X1 _11258_ ( .A(_03587_ ), .ZN(_03588_ ) );
XNOR2_X1 _11259_ ( .A(_03443_ ), .B(_01975_ ), .ZN(_03589_ ) );
XNOR2_X1 _11260_ ( .A(_03443_ ), .B(_01889_ ), .ZN(_03590_ ) );
XNOR2_X1 _11261_ ( .A(_03443_ ), .B(_01830_ ), .ZN(_03591_ ) );
XNOR2_X1 _11262_ ( .A(_03443_ ), .B(_01949_ ), .ZN(_03592_ ) );
AND2_X1 _11263_ ( .A1(_03591_ ), .A2(_03592_ ), .ZN(_03593_ ) );
NAND4_X2 _11264_ ( .A1(_03588_ ), .A2(_03589_ ), .A3(_03590_ ), .A4(_03593_ ), .ZN(_03594_ ) );
OAI21_X1 _11265_ ( .A(_03444_ ), .B1(\IF_ID_pc [26] ), .B2(\IF_ID_pc [25] ), .ZN(_03595_ ) );
INV_X1 _11266_ ( .A(_03595_ ), .ZN(_03596_ ) );
NAND3_X1 _11267_ ( .A1(_03589_ ), .A2(_03590_ ), .A3(_03596_ ), .ZN(_03597_ ) );
NAND2_X1 _11268_ ( .A1(_03444_ ), .A2(\IF_ID_pc [28] ), .ZN(_03598_ ) );
NAND2_X1 _11269_ ( .A1(_03444_ ), .A2(\IF_ID_pc [27] ), .ZN(_03599_ ) );
AND3_X1 _11270_ ( .A1(_03597_ ), .A2(_03598_ ), .A3(_03599_ ), .ZN(_03600_ ) );
AOI21_X1 _11271_ ( .A(_03446_ ), .B1(_03594_ ), .B2(_03600_ ), .ZN(_03601_ ) );
NOR3_X1 _11272_ ( .A1(_03439_ ), .A2(_01856_ ), .A3(_03441_ ), .ZN(_03602_ ) );
OR2_X2 _11273_ ( .A1(_03601_ ), .A2(_03602_ ), .ZN(_03603_ ) );
XNOR2_X1 _11274_ ( .A(_03444_ ), .B(_01982_ ), .ZN(_03604_ ) );
OAI21_X1 _11275_ ( .A(_03435_ ), .B1(_03603_ ), .B2(_03604_ ), .ZN(_03605_ ) );
AOI21_X1 _11276_ ( .A(_03605_ ), .B1(_03603_ ), .B2(_03604_ ), .ZN(_03606_ ) );
BUF_X2 _11277_ ( .A(_03274_ ), .Z(_03607_ ) );
BUF_X4 _11278_ ( .A(_03607_ ), .Z(_03608_ ) );
AOI211_X1 _11279_ ( .A(fanout_net_49 ), .B(_03606_ ), .C1(\myexu.pc_jump [30] ), .C2(_03608_ ), .ZN(_03609_ ) );
BUF_X4 _11280_ ( .A(_03431_ ), .Z(_03610_ ) );
NOR2_X1 _11281_ ( .A1(_03610_ ), .A2(\mtvec [30] ), .ZN(_03611_ ) );
NOR3_X1 _11282_ ( .A1(_03609_ ), .A2(fanout_net_2 ), .A3(_03611_ ), .ZN(_00168_ ) );
XNOR2_X1 _11283_ ( .A(_03573_ ), .B(_03577_ ), .ZN(_03612_ ) );
MUX2_X1 _11284_ ( .A(\myexu.pc_jump [21] ), .B(_03612_ ), .S(_03435_ ), .Z(_03613_ ) );
MUX2_X1 _11285_ ( .A(\mtvec [21] ), .B(_03613_ ), .S(_03431_ ), .Z(_03614_ ) );
AND2_X1 _11286_ ( .A1(_03614_ ), .A2(_01564_ ), .ZN(_00169_ ) );
INV_X1 _11287_ ( .A(_03561_ ), .ZN(_03615_ ) );
INV_X1 _11288_ ( .A(_03558_ ), .ZN(_03616_ ) );
AOI21_X1 _11289_ ( .A(_03616_ ), .B1(_03545_ ), .B2(_03554_ ), .ZN(_03617_ ) );
NAND2_X1 _11290_ ( .A1(_03617_ ), .A2(_03449_ ), .ZN(_03618_ ) );
AOI21_X1 _11291_ ( .A(_03615_ ), .B1(_03618_ ), .B2(_03570_ ), .ZN(_03619_ ) );
OR3_X1 _11292_ ( .A1(_03619_ ), .A2(_03565_ ), .A3(_03562_ ), .ZN(_03620_ ) );
OAI21_X1 _11293_ ( .A(_03562_ ), .B1(_03619_ ), .B2(_03565_ ), .ZN(_03621_ ) );
AND3_X1 _11294_ ( .A1(_03620_ ), .A2(_03435_ ), .A3(_03621_ ), .ZN(_03622_ ) );
AOI211_X1 _11295_ ( .A(fanout_net_49 ), .B(_03622_ ), .C1(\myexu.pc_jump [20] ), .C2(_03608_ ), .ZN(_03623_ ) );
NOR2_X1 _11296_ ( .A1(_03610_ ), .A2(\mtvec [20] ), .ZN(_03624_ ) );
NOR3_X1 _11297_ ( .A1(_03623_ ), .A2(fanout_net_2 ), .A3(_03624_ ), .ZN(_00170_ ) );
AND2_X1 _11298_ ( .A1(_03618_ ), .A2(_03570_ ), .ZN(_03625_ ) );
OAI21_X1 _11299_ ( .A(_03435_ ), .B1(_03625_ ), .B2(_03615_ ), .ZN(_03626_ ) );
AOI21_X1 _11300_ ( .A(_03626_ ), .B1(_03615_ ), .B2(_03625_ ), .ZN(_03627_ ) );
AOI211_X1 _11301_ ( .A(fanout_net_49 ), .B(_03627_ ), .C1(\myexu.pc_jump [19] ), .C2(_03608_ ), .ZN(_03628_ ) );
NOR2_X1 _11302_ ( .A1(_03610_ ), .A2(\mtvec [19] ), .ZN(_03629_ ) );
NOR3_X1 _11303_ ( .A1(_03628_ ), .A2(fanout_net_2 ), .A3(_03629_ ), .ZN(_00171_ ) );
OR3_X1 _11304_ ( .A1(_03617_ ), .A2(_03449_ ), .A3(_03568_ ), .ZN(_03630_ ) );
OAI21_X1 _11305_ ( .A(_03449_ ), .B1(_03617_ ), .B2(_03568_ ), .ZN(_03631_ ) );
AND3_X1 _11306_ ( .A1(_03630_ ), .A2(_03435_ ), .A3(_03631_ ), .ZN(_03632_ ) );
AOI211_X1 _11307_ ( .A(fanout_net_49 ), .B(_03632_ ), .C1(\myexu.pc_jump [18] ), .C2(_03608_ ), .ZN(_03633_ ) );
NOR2_X1 _11308_ ( .A1(_03610_ ), .A2(\mtvec [18] ), .ZN(_03634_ ) );
NOR3_X1 _11309_ ( .A1(_03633_ ), .A2(fanout_net_2 ), .A3(_03634_ ), .ZN(_00172_ ) );
BUF_X4 _11310_ ( .A(_03435_ ), .Z(_03635_ ) );
BUF_X4 _11311_ ( .A(_03635_ ), .Z(_03636_ ) );
AND3_X1 _11312_ ( .A1(_03545_ ), .A2(_03554_ ), .A3(_03616_ ), .ZN(_03637_ ) );
OAI21_X1 _11313_ ( .A(_03636_ ), .B1(_03637_ ), .B2(_03617_ ), .ZN(_03638_ ) );
BUF_X4 _11314_ ( .A(_03431_ ), .Z(_03639_ ) );
BUF_X4 _11315_ ( .A(_03635_ ), .Z(_03640_ ) );
OAI211_X1 _11316_ ( .A(_03638_ ), .B(_03639_ ), .C1(\myexu.pc_jump [17] ), .C2(_03640_ ), .ZN(_03641_ ) );
NAND2_X1 _11317_ ( .A1(\mtvec [17] ), .A2(fanout_net_49 ), .ZN(_03642_ ) );
AOI21_X1 _11318_ ( .A(fanout_net_2 ), .B1(_03641_ ), .B2(_03642_ ), .ZN(_00173_ ) );
INV_X1 _11319_ ( .A(_03540_ ), .ZN(_03643_ ) );
INV_X1 _11320_ ( .A(_03544_ ), .ZN(_03644_ ) );
NOR4_X1 _11321_ ( .A1(_03528_ ), .A2(_03643_ ), .A3(_03644_ ), .A4(_03529_ ), .ZN(_03645_ ) );
NOR2_X1 _11322_ ( .A1(_03645_ ), .A2(_03553_ ), .ZN(_03646_ ) );
NOR2_X1 _11323_ ( .A1(_03646_ ), .A2(_03536_ ), .ZN(_03647_ ) );
NOR2_X1 _11324_ ( .A1(_03647_ ), .A2(_03546_ ), .ZN(_03648_ ) );
XOR2_X1 _11325_ ( .A(_03648_ ), .B(_03533_ ), .Z(_03649_ ) );
MUX2_X1 _11326_ ( .A(\myexu.pc_jump [16] ), .B(_03649_ ), .S(_03434_ ), .Z(_03650_ ) );
MUX2_X1 _11327_ ( .A(\mtvec [16] ), .B(_03650_ ), .S(_03430_ ), .Z(_03651_ ) );
AND2_X1 _11328_ ( .A1(_03651_ ), .A2(_01564_ ), .ZN(_00174_ ) );
AND2_X1 _11329_ ( .A1(_03646_ ), .A2(_03536_ ), .ZN(_03652_ ) );
OAI21_X1 _11330_ ( .A(_03635_ ), .B1(_03652_ ), .B2(_03647_ ), .ZN(_03653_ ) );
OAI211_X1 _11331_ ( .A(_03653_ ), .B(_03639_ ), .C1(\myexu.pc_jump [15] ), .C2(_03640_ ), .ZN(_03654_ ) );
NAND2_X1 _11332_ ( .A1(\mtvec [15] ), .A2(fanout_net_49 ), .ZN(_03655_ ) );
AOI21_X1 _11333_ ( .A(fanout_net_2 ), .B1(_03654_ ), .B2(_03655_ ), .ZN(_00175_ ) );
NOR2_X1 _11334_ ( .A1(_03431_ ), .A2(\mtvec [14] ), .ZN(_03656_ ) );
NOR3_X1 _11335_ ( .A1(_03528_ ), .A2(_03644_ ), .A3(_03529_ ), .ZN(_03657_ ) );
OR3_X1 _11336_ ( .A1(_03657_ ), .A2(_03550_ ), .A3(_03540_ ), .ZN(_03658_ ) );
OAI21_X1 _11337_ ( .A(_03540_ ), .B1(_03657_ ), .B2(_03550_ ), .ZN(_03659_ ) );
NAND3_X1 _11338_ ( .A1(_03658_ ), .A2(_03640_ ), .A3(_03659_ ), .ZN(_03660_ ) );
AOI21_X1 _11339_ ( .A(fanout_net_49 ), .B1(_03608_ ), .B2(\myexu.pc_jump [14] ), .ZN(_03661_ ) );
AOI211_X1 _11340_ ( .A(fanout_net_2 ), .B(_03656_ ), .C1(_03660_ ), .C2(_03661_ ), .ZN(_00176_ ) );
NOR2_X1 _11341_ ( .A1(_03530_ ), .A2(_03544_ ), .ZN(_03662_ ) );
OAI21_X1 _11342_ ( .A(_03635_ ), .B1(_03662_ ), .B2(_03657_ ), .ZN(_03663_ ) );
OAI211_X1 _11343_ ( .A(_03663_ ), .B(_03639_ ), .C1(\myexu.pc_jump [13] ), .C2(_03640_ ), .ZN(_03664_ ) );
NAND2_X1 _11344_ ( .A1(\mtvec [13] ), .A2(fanout_net_49 ), .ZN(_03665_ ) );
AOI21_X1 _11345_ ( .A(fanout_net_2 ), .B1(_03664_ ), .B2(_03665_ ), .ZN(_00177_ ) );
NOR2_X1 _11346_ ( .A1(_03525_ ), .A2(_03454_ ), .ZN(_03666_ ) );
INV_X1 _11347_ ( .A(_03666_ ), .ZN(_03667_ ) );
XNOR2_X1 _11348_ ( .A(_03527_ ), .B(_01849_ ), .ZN(_03668_ ) );
OAI21_X1 _11349_ ( .A(_03435_ ), .B1(_03667_ ), .B2(_03668_ ), .ZN(_03669_ ) );
AOI21_X1 _11350_ ( .A(_03669_ ), .B1(_03667_ ), .B2(_03668_ ), .ZN(_03670_ ) );
AOI211_X1 _11351_ ( .A(fanout_net_49 ), .B(_03670_ ), .C1(\myexu.pc_jump [12] ), .C2(_03608_ ), .ZN(_03671_ ) );
NOR2_X1 _11352_ ( .A1(_03610_ ), .A2(\mtvec [12] ), .ZN(_03672_ ) );
NOR3_X1 _11353_ ( .A1(_03671_ ), .A2(fanout_net_2 ), .A3(_03672_ ), .ZN(_00178_ ) );
AND3_X1 _11354_ ( .A1(_03594_ ), .A2(_03600_ ), .A3(_03445_ ), .ZN(_03673_ ) );
AOI21_X1 _11355_ ( .A(_03445_ ), .B1(_03594_ ), .B2(_03600_ ), .ZN(_03674_ ) );
OR3_X1 _11356_ ( .A1(_03673_ ), .A2(_03674_ ), .A3(_03607_ ), .ZN(_03675_ ) );
OAI211_X1 _11357_ ( .A(_03675_ ), .B(_03639_ ), .C1(\myexu.pc_jump [29] ), .C2(_03640_ ), .ZN(_03676_ ) );
NAND2_X1 _11358_ ( .A1(\mtvec [29] ), .A2(fanout_net_49 ), .ZN(_03677_ ) );
AOI21_X1 _11359_ ( .A(fanout_net_2 ), .B1(_03676_ ), .B2(_03677_ ), .ZN(_00179_ ) );
AOI21_X1 _11360_ ( .A(_03522_ ), .B1(_03520_ ), .B2(_03524_ ), .ZN(_03678_ ) );
OAI21_X1 _11361_ ( .A(_03635_ ), .B1(_03525_ ), .B2(_03678_ ), .ZN(_03679_ ) );
OAI211_X1 _11362_ ( .A(_03679_ ), .B(_03639_ ), .C1(\myexu.pc_jump [11] ), .C2(_03640_ ), .ZN(_03680_ ) );
NAND2_X1 _11363_ ( .A1(\mtvec [11] ), .A2(fanout_net_49 ), .ZN(_03681_ ) );
AOI21_X1 _11364_ ( .A(fanout_net_2 ), .B1(_03680_ ), .B2(_03681_ ), .ZN(_00180_ ) );
INV_X1 _11365_ ( .A(_03515_ ), .ZN(_03682_ ) );
XNOR2_X1 _11366_ ( .A(_03519_ ), .B(\IF_ID_pc [10] ), .ZN(_03683_ ) );
OAI21_X1 _11367_ ( .A(_03435_ ), .B1(_03682_ ), .B2(_03683_ ), .ZN(_03684_ ) );
AOI21_X1 _11368_ ( .A(_03684_ ), .B1(_03682_ ), .B2(_03683_ ), .ZN(_03685_ ) );
AOI211_X1 _11369_ ( .A(fanout_net_49 ), .B(_03685_ ), .C1(\myexu.pc_jump [10] ), .C2(_03608_ ), .ZN(_03686_ ) );
NOR2_X1 _11370_ ( .A1(_03610_ ), .A2(\mtvec [10] ), .ZN(_03687_ ) );
NOR3_X1 _11371_ ( .A1(_03686_ ), .A2(fanout_net_2 ), .A3(_03687_ ), .ZN(_00181_ ) );
AND3_X1 _11372_ ( .A1(_03511_ ), .A2(_03512_ ), .A3(_03459_ ), .ZN(_03688_ ) );
OAI21_X1 _11373_ ( .A(_03635_ ), .B1(_03688_ ), .B2(_03513_ ), .ZN(_03689_ ) );
OAI211_X1 _11374_ ( .A(_03689_ ), .B(_03639_ ), .C1(\myexu.pc_jump [9] ), .C2(_03640_ ), .ZN(_03690_ ) );
NAND2_X1 _11375_ ( .A1(\mtvec [9] ), .A2(fanout_net_49 ), .ZN(_03691_ ) );
AOI21_X1 _11376_ ( .A(fanout_net_2 ), .B1(_03690_ ), .B2(_03691_ ), .ZN(_00182_ ) );
NOR2_X1 _11377_ ( .A1(_03506_ ), .A2(_03507_ ), .ZN(_03692_ ) );
XNOR2_X1 _11378_ ( .A(_03510_ ), .B(\IF_ID_pc [8] ), .ZN(_03693_ ) );
OR2_X1 _11379_ ( .A1(_03692_ ), .A2(_03693_ ), .ZN(_03694_ ) );
AOI21_X1 _11380_ ( .A(_03607_ ), .B1(_03692_ ), .B2(_03693_ ), .ZN(_03695_ ) );
AOI221_X4 _11381_ ( .A(fanout_net_49 ), .B1(\myexu.pc_jump [8] ), .B2(_03607_ ), .C1(_03694_ ), .C2(_03695_ ), .ZN(_03696_ ) );
NOR2_X1 _11382_ ( .A1(_03610_ ), .A2(\mtvec [8] ), .ZN(_03697_ ) );
NOR3_X1 _11383_ ( .A1(_03696_ ), .A2(fanout_net_2 ), .A3(_03697_ ), .ZN(_00183_ ) );
AOI21_X1 _11384_ ( .A(_03504_ ), .B1(_03500_ ), .B2(_03505_ ), .ZN(_03698_ ) );
OAI21_X1 _11385_ ( .A(_03635_ ), .B1(_03506_ ), .B2(_03698_ ), .ZN(_03699_ ) );
OAI211_X1 _11386_ ( .A(_03699_ ), .B(_03639_ ), .C1(\myexu.pc_jump [7] ), .C2(_03636_ ), .ZN(_03700_ ) );
NAND2_X1 _11387_ ( .A1(\mtvec [7] ), .A2(fanout_net_49 ), .ZN(_03701_ ) );
AOI21_X1 _11388_ ( .A(fanout_net_2 ), .B1(_03700_ ), .B2(_03701_ ), .ZN(_00184_ ) );
NOR2_X1 _11389_ ( .A1(_03431_ ), .A2(\mtvec [6] ), .ZN(_03702_ ) );
XNOR2_X1 _11390_ ( .A(_03499_ ), .B(_03496_ ), .ZN(_03703_ ) );
AOI21_X1 _11391_ ( .A(_03607_ ), .B1(_03495_ ), .B2(_03703_ ), .ZN(_03704_ ) );
OAI21_X1 _11392_ ( .A(_03704_ ), .B1(_03495_ ), .B2(_03703_ ), .ZN(_03705_ ) );
AOI21_X1 _11393_ ( .A(fanout_net_49 ), .B1(_03608_ ), .B2(\myexu.pc_jump [6] ), .ZN(_03706_ ) );
AOI211_X1 _11394_ ( .A(fanout_net_2 ), .B(_03702_ ), .C1(_03705_ ), .C2(_03706_ ), .ZN(_00185_ ) );
AND2_X1 _11395_ ( .A1(_03487_ ), .A2(_03492_ ), .ZN(_03707_ ) );
OAI21_X1 _11396_ ( .A(_03635_ ), .B1(_03707_ ), .B2(_03493_ ), .ZN(_03708_ ) );
OAI211_X1 _11397_ ( .A(_03708_ ), .B(_03639_ ), .C1(\myexu.pc_jump [5] ), .C2(_03636_ ), .ZN(_03709_ ) );
NAND2_X1 _11398_ ( .A1(\mtvec [5] ), .A2(fanout_net_49 ), .ZN(_03710_ ) );
AOI21_X1 _11399_ ( .A(fanout_net_2 ), .B1(_03709_ ), .B2(_03710_ ), .ZN(_00186_ ) );
OR2_X1 _11400_ ( .A1(_03482_ ), .A2(_03483_ ), .ZN(_03711_ ) );
AND2_X1 _11401_ ( .A1(_03464_ ), .A2(_03486_ ), .ZN(_03712_ ) );
AND3_X1 _11402_ ( .A1(_03711_ ), .A2(_03470_ ), .A3(_03712_ ), .ZN(_03713_ ) );
AOI21_X1 _11403_ ( .A(_03712_ ), .B1(_03711_ ), .B2(_03470_ ), .ZN(_03714_ ) );
OR3_X1 _11404_ ( .A1(_03713_ ), .A2(_03714_ ), .A3(_03607_ ), .ZN(_03715_ ) );
OAI211_X1 _11405_ ( .A(_03715_ ), .B(_03430_ ), .C1(\myexu.pc_jump [4] ), .C2(_03435_ ), .ZN(_03716_ ) );
NAND2_X1 _11406_ ( .A1(\mtvec [4] ), .A2(fanout_net_49 ), .ZN(_03717_ ) );
AOI21_X1 _11407_ ( .A(fanout_net_2 ), .B1(_03716_ ), .B2(_03717_ ), .ZN(_00187_ ) );
AND2_X1 _11408_ ( .A1(_03434_ ), .A2(_03711_ ), .ZN(_03718_ ) );
NAND2_X1 _11409_ ( .A1(_03482_ ), .A2(_03483_ ), .ZN(_03719_ ) );
AOI22_X1 _11410_ ( .A1(_03718_ ), .A2(_03719_ ), .B1(\myexu.pc_jump [3] ), .B2(_03607_ ), .ZN(_03720_ ) );
NOR2_X1 _11411_ ( .A1(_03720_ ), .A2(fanout_net_49 ), .ZN(_03721_ ) );
AOI21_X1 _11412_ ( .A(_03721_ ), .B1(\mtvec [3] ), .B2(fanout_net_49 ), .ZN(_03722_ ) );
NOR2_X1 _11413_ ( .A1(_03722_ ), .A2(fanout_net_2 ), .ZN(_00188_ ) );
AND2_X1 _11414_ ( .A1(IDU_ready_IFU ), .A2(\myifu.state [1] ), .ZN(\myifu.pc_$_SDFFE_PP1P__Q_E ) );
AND3_X1 _11415_ ( .A1(_03716_ ), .A2(_03717_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_03723_ ) );
BUF_X2 _11416_ ( .A(_03485_ ), .Z(_03724_ ) );
BUF_X4 _11417_ ( .A(_03724_ ), .Z(_03725_ ) );
BUF_X2 _11418_ ( .A(_03725_ ), .Z(_03726_ ) );
INV_X1 _11419_ ( .A(\myifu.pc_$_SDFFE_PP1P__Q_E ), .ZN(_03727_ ) );
AOI211_X1 _11420_ ( .A(fanout_net_2 ), .B(_03723_ ), .C1(_03726_ ), .C2(_03727_ ), .ZN(_00189_ ) );
XNOR2_X1 _11421_ ( .A(_03475_ ), .B(_03480_ ), .ZN(_03728_ ) );
AND3_X1 _11422_ ( .A1(_03239_ ), .A2(_03261_ ), .A3(_03272_ ), .ZN(_03729_ ) );
INV_X1 _11423_ ( .A(check_quest ), .ZN(_03730_ ) );
OAI21_X1 _11424_ ( .A(_03728_ ), .B1(_03729_ ), .B2(_03730_ ), .ZN(_03731_ ) );
OAI211_X1 _11425_ ( .A(_03610_ ), .B(_03731_ ), .C1(_03640_ ), .C2(\myexu.pc_jump [2] ), .ZN(_03732_ ) );
NAND2_X1 _11426_ ( .A1(\mtvec [2] ), .A2(fanout_net_49 ), .ZN(_03733_ ) );
AOI21_X1 _11427_ ( .A(fanout_net_2 ), .B1(_03732_ ), .B2(_03733_ ), .ZN(_00190_ ) );
AOI211_X1 _11428_ ( .A(_03727_ ), .B(_03721_ ), .C1(\mtvec [3] ), .C2(fanout_net_49 ), .ZN(_03734_ ) );
INV_X1 _11429_ ( .A(fanout_net_12 ), .ZN(_03735_ ) );
BUF_X4 _11430_ ( .A(_03735_ ), .Z(_03736_ ) );
BUF_X2 _11431_ ( .A(_03736_ ), .Z(_03737_ ) );
AOI211_X1 _11432_ ( .A(fanout_net_2 ), .B(_03734_ ), .C1(_03737_ ), .C2(_03727_ ), .ZN(_00191_ ) );
AND2_X1 _11433_ ( .A1(_03588_ ), .A2(_03593_ ), .ZN(_03738_ ) );
OAI21_X1 _11434_ ( .A(_03590_ ), .B1(_03738_ ), .B2(_03596_ ), .ZN(_03739_ ) );
AND3_X1 _11435_ ( .A1(_03739_ ), .A2(_03589_ ), .A3(_03599_ ), .ZN(_03740_ ) );
AOI21_X1 _11436_ ( .A(_03589_ ), .B1(_03739_ ), .B2(_03599_ ), .ZN(_03741_ ) );
OR3_X1 _11437_ ( .A1(_03740_ ), .A2(_03741_ ), .A3(_03607_ ), .ZN(_03742_ ) );
OAI211_X1 _11438_ ( .A(_03742_ ), .B(_03639_ ), .C1(\myexu.pc_jump [28] ), .C2(_03636_ ), .ZN(_03743_ ) );
NAND2_X1 _11439_ ( .A1(\mtvec [28] ), .A2(fanout_net_49 ), .ZN(_03744_ ) );
AOI21_X1 _11440_ ( .A(fanout_net_2 ), .B1(_03743_ ), .B2(_03744_ ), .ZN(_00192_ ) );
XNOR2_X1 _11441_ ( .A(_03479_ ), .B(\IF_ID_pc [1] ), .ZN(_03745_ ) );
AOI21_X1 _11442_ ( .A(_03745_ ), .B1(_03273_ ), .B2(check_quest ), .ZN(_03746_ ) );
AOI211_X1 _11443_ ( .A(fanout_net_49 ), .B(_03746_ ), .C1(\myexu.pc_jump [1] ), .C2(_03608_ ), .ZN(_03747_ ) );
NOR2_X1 _11444_ ( .A1(_03610_ ), .A2(\mtvec [1] ), .ZN(_03748_ ) );
NOR3_X1 _11445_ ( .A1(_03747_ ), .A2(fanout_net_2 ), .A3(_03748_ ), .ZN(_00193_ ) );
NOR2_X1 _11446_ ( .A1(_03738_ ), .A2(_03596_ ), .ZN(_03749_ ) );
XOR2_X1 _11447_ ( .A(_03749_ ), .B(_03590_ ), .Z(_03750_ ) );
NAND2_X1 _11448_ ( .A1(_03750_ ), .A2(_03636_ ), .ZN(_03751_ ) );
OAI211_X1 _11449_ ( .A(_03751_ ), .B(_03639_ ), .C1(\myexu.pc_jump [27] ), .C2(_03636_ ), .ZN(_03752_ ) );
NAND2_X1 _11450_ ( .A1(\mtvec [27] ), .A2(fanout_net_49 ), .ZN(_03753_ ) );
AOI21_X1 _11451_ ( .A(fanout_net_2 ), .B1(_03752_ ), .B2(_03753_ ), .ZN(_00194_ ) );
AND2_X1 _11452_ ( .A1(_03588_ ), .A2(_03592_ ), .ZN(_03754_ ) );
AND2_X1 _11453_ ( .A1(_03444_ ), .A2(\IF_ID_pc [25] ), .ZN(_03755_ ) );
OR3_X1 _11454_ ( .A1(_03754_ ), .A2(_03755_ ), .A3(_03591_ ), .ZN(_03756_ ) );
OAI21_X1 _11455_ ( .A(_03591_ ), .B1(_03754_ ), .B2(_03755_ ), .ZN(_03757_ ) );
AND3_X1 _11456_ ( .A1(_03756_ ), .A2(_03435_ ), .A3(_03757_ ), .ZN(_03758_ ) );
AOI211_X1 _11457_ ( .A(fanout_net_49 ), .B(_03758_ ), .C1(\myexu.pc_jump [26] ), .C2(_03607_ ), .ZN(_03759_ ) );
NOR2_X1 _11458_ ( .A1(_03610_ ), .A2(\mtvec [26] ), .ZN(_03760_ ) );
NOR3_X1 _11459_ ( .A1(_03759_ ), .A2(fanout_net_2 ), .A3(_03760_ ), .ZN(_00195_ ) );
NOR3_X1 _11460_ ( .A1(_03580_ ), .A2(_03586_ ), .A3(_03592_ ), .ZN(_03761_ ) );
OAI21_X1 _11461_ ( .A(_03635_ ), .B1(_03754_ ), .B2(_03761_ ), .ZN(_03762_ ) );
OAI211_X1 _11462_ ( .A(_03762_ ), .B(_03431_ ), .C1(\myexu.pc_jump [25] ), .C2(_03636_ ), .ZN(_03763_ ) );
NAND2_X1 _11463_ ( .A1(\mtvec [25] ), .A2(fanout_net_49 ), .ZN(_03764_ ) );
AOI21_X1 _11464_ ( .A(fanout_net_2 ), .B1(_03763_ ), .B2(_03764_ ), .ZN(_00196_ ) );
OAI21_X1 _11465_ ( .A(_03579_ ), .B1(_03564_ ), .B2(_03572_ ), .ZN(_03765_ ) );
OAI21_X1 _11466_ ( .A(_03444_ ), .B1(\IF_ID_pc [22] ), .B2(\IF_ID_pc [21] ), .ZN(_03766_ ) );
NAND2_X1 _11467_ ( .A1(_03765_ ), .A2(_03766_ ), .ZN(_03767_ ) );
NAND2_X1 _11468_ ( .A1(_03767_ ), .A2(_03575_ ), .ZN(_03768_ ) );
AND3_X1 _11469_ ( .A1(_03768_ ), .A2(_03574_ ), .A3(_03585_ ), .ZN(_03769_ ) );
AOI21_X1 _11470_ ( .A(_03574_ ), .B1(_03768_ ), .B2(_03585_ ), .ZN(_03770_ ) );
OR3_X1 _11471_ ( .A1(_03769_ ), .A2(_03770_ ), .A3(_03607_ ), .ZN(_03771_ ) );
OAI211_X1 _11472_ ( .A(_03771_ ), .B(_03431_ ), .C1(\myexu.pc_jump [24] ), .C2(_03636_ ), .ZN(_03772_ ) );
NAND2_X1 _11473_ ( .A1(\mtvec [24] ), .A2(\myifu.to_reset ), .ZN(_03773_ ) );
AOI21_X1 _11474_ ( .A(fanout_net_3 ), .B1(_03772_ ), .B2(_03773_ ), .ZN(_00197_ ) );
XNOR2_X1 _11475_ ( .A(_03767_ ), .B(_03575_ ), .ZN(_03774_ ) );
NAND2_X1 _11476_ ( .A1(_03774_ ), .A2(_03636_ ), .ZN(_03775_ ) );
OAI211_X1 _11477_ ( .A(_03775_ ), .B(_03431_ ), .C1(\myexu.pc_jump [23] ), .C2(_03636_ ), .ZN(_03776_ ) );
NAND2_X1 _11478_ ( .A1(\mtvec [23] ), .A2(\myifu.to_reset ), .ZN(_03777_ ) );
AOI21_X1 _11479_ ( .A(fanout_net_3 ), .B1(_03776_ ), .B2(_03777_ ), .ZN(_00198_ ) );
INV_X1 _11480_ ( .A(_03573_ ), .ZN(_03778_ ) );
NOR2_X1 _11481_ ( .A1(_03778_ ), .A2(_03577_ ), .ZN(_03779_ ) );
NOR2_X1 _11482_ ( .A1(_03779_ ), .A2(_03582_ ), .ZN(_03780_ ) );
XOR2_X1 _11483_ ( .A(_03780_ ), .B(_03578_ ), .Z(_03781_ ) );
MUX2_X1 _11484_ ( .A(\myexu.pc_jump [22] ), .B(_03781_ ), .S(_03434_ ), .Z(_03782_ ) );
MUX2_X1 _11485_ ( .A(\mtvec [22] ), .B(_03782_ ), .S(_03430_ ), .Z(_03783_ ) );
AND2_X1 _11486_ ( .A1(_03783_ ), .A2(_01564_ ), .ZN(_00199_ ) );
NAND2_X1 _11487_ ( .A1(\mtvec [31] ), .A2(\myifu.to_reset ), .ZN(_03784_ ) );
OAI22_X1 _11488_ ( .A1(_03601_ ), .A2(_03602_ ), .B1(\IF_ID_pc [30] ), .B2(_03444_ ), .ZN(_03785_ ) );
NAND2_X1 _11489_ ( .A1(_03444_ ), .A2(\IF_ID_pc [30] ), .ZN(_03786_ ) );
NAND2_X1 _11490_ ( .A1(_03785_ ), .A2(_03786_ ), .ZN(_03787_ ) );
XNOR2_X1 _11491_ ( .A(_03444_ ), .B(\IF_ID_pc [31] ), .ZN(_03788_ ) );
OAI21_X1 _11492_ ( .A(_03635_ ), .B1(_03787_ ), .B2(_03788_ ), .ZN(_03789_ ) );
AOI21_X1 _11493_ ( .A(_03789_ ), .B1(_03787_ ), .B2(_03788_ ), .ZN(_03790_ ) );
OAI21_X1 _11494_ ( .A(_03431_ ), .B1(_03640_ ), .B2(\myexu.pc_jump [31] ), .ZN(_03791_ ) );
OAI211_X1 _11495_ ( .A(_01735_ ), .B(_03784_ ), .C1(_03790_ ), .C2(_03791_ ), .ZN(_00200_ ) );
INV_X1 _11496_ ( .A(\myifu.tmp_offset [2] ), .ZN(_03792_ ) );
OR2_X1 _11497_ ( .A1(_02061_ ), .A2(\myclint.state_r_$_NOT__A_Y ), .ZN(_03793_ ) );
NAND2_X1 _11498_ ( .A1(_02062_ ), .A2(io_master_rvalid ), .ZN(_03794_ ) );
NAND2_X2 _11499_ ( .A1(_03793_ ), .A2(_03794_ ), .ZN(_03795_ ) );
BUF_X4 _11500_ ( .A(_01956_ ), .Z(_03796_ ) );
NOR2_X1 _11501_ ( .A1(\io_master_rresp [1] ), .A2(\io_master_rresp [0] ), .ZN(_03797_ ) );
NOR2_X1 _11502_ ( .A1(\io_master_rid [3] ), .A2(\io_master_rid [2] ), .ZN(_03798_ ) );
INV_X1 _11503_ ( .A(\io_master_rid [1] ), .ZN(_03799_ ) );
NAND4_X1 _11504_ ( .A1(_03797_ ), .A2(_03798_ ), .A3(_03799_ ), .A4(\io_master_rid [0] ), .ZN(_03800_ ) );
AOI21_X1 _11505_ ( .A(_03796_ ), .B1(_02062_ ), .B2(_03800_ ), .ZN(_03801_ ) );
AND2_X2 _11506_ ( .A1(_03795_ ), .A2(_03801_ ), .ZN(_03802_ ) );
INV_X1 _11507_ ( .A(_03802_ ), .ZN(_03803_ ) );
NOR2_X1 _11508_ ( .A1(_02060_ ), .A2(io_master_rlast ), .ZN(_03804_ ) );
OAI211_X1 _11509_ ( .A(_01682_ ), .B(_03792_ ), .C1(_03803_ ), .C2(_03804_ ), .ZN(_03805_ ) );
INV_X1 _11510_ ( .A(_03805_ ), .ZN(_00201_ ) );
NOR3_X1 _11511_ ( .A1(fanout_net_3 ), .A2(\myifu.state [1] ), .A3(\myifu.state [2] ), .ZN(_00202_ ) );
AND3_X1 _11512_ ( .A1(_02076_ ), .A2(_03275_ ), .A3(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_03806_ ) );
INV_X1 _11513_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .ZN(_03807_ ) );
MUX2_X1 _11514_ ( .A(_02076_ ), .B(_03807_ ), .S(\myifu.to_reset ), .Z(_03808_ ) );
AOI211_X1 _11515_ ( .A(fanout_net_3 ), .B(_03806_ ), .C1(_03808_ ), .C2(\myifu.state [1] ), .ZN(_00203_ ) );
AND3_X1 _11516_ ( .A1(fanout_net_5 ), .A2(_01682_ ), .A3(\EX_LS_pc [2] ), .ZN(_00204_ ) );
AND2_X1 _11517_ ( .A1(fanout_net_5 ), .A2(_01456_ ), .ZN(_03809_ ) );
BUF_X2 _11518_ ( .A(_03809_ ), .Z(_03810_ ) );
AND2_X1 _11519_ ( .A1(_03810_ ), .A2(\mylsu.state [3] ), .ZN(_00205_ ) );
BUF_X2 _11520_ ( .A(_02035_ ), .Z(_03811_ ) );
AOI21_X1 _11521_ ( .A(\LS_WB_waddr_csreg [11] ), .B1(_03811_ ), .B2(\EX_LS_flag [2] ), .ZN(_03812_ ) );
NOR2_X1 _11522_ ( .A1(_02046_ ), .A2(_02037_ ), .ZN(_03813_ ) );
NAND2_X1 _11523_ ( .A1(_02034_ ), .A2(\EX_LS_flag [2] ), .ZN(_03814_ ) );
NAND2_X1 _11524_ ( .A1(_02150_ ), .A2(_03814_ ), .ZN(_03815_ ) );
AND2_X1 _11525_ ( .A1(_02152_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_03816_ ) );
NOR2_X1 _11526_ ( .A1(_03815_ ), .A2(_03816_ ), .ZN(_03817_ ) );
INV_X1 _11527_ ( .A(_03817_ ), .ZN(_03818_ ) );
OR2_X2 _11528_ ( .A1(_03813_ ), .A2(_03818_ ), .ZN(_03819_ ) );
BUF_X4 _11529_ ( .A(_03819_ ), .Z(_03820_ ) );
INV_X1 _11530_ ( .A(\EX_LS_dest_csreg_mem [11] ), .ZN(_03821_ ) );
AND2_X1 _11531_ ( .A1(_02035_ ), .A2(\EX_LS_flag [2] ), .ZN(_03822_ ) );
BUF_X2 _11532_ ( .A(_03822_ ), .Z(_03823_ ) );
BUF_X4 _11533_ ( .A(_03823_ ), .Z(_03824_ ) );
AOI211_X1 _11534_ ( .A(_03812_ ), .B(_03820_ ), .C1(_03821_ ), .C2(_03824_ ), .ZN(_00206_ ) );
NOR2_X1 _11535_ ( .A1(_03813_ ), .A2(_03816_ ), .ZN(_03825_ ) );
AND2_X1 _11536_ ( .A1(_03825_ ), .A2(_02018_ ), .ZN(_03826_ ) );
INV_X1 _11537_ ( .A(_03826_ ), .ZN(_03827_ ) );
NAND3_X1 _11538_ ( .A1(_03811_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(\EX_LS_flag [2] ), .ZN(_03828_ ) );
BUF_X4 _11539_ ( .A(_01945_ ), .Z(_03829_ ) );
NAND2_X1 _11540_ ( .A1(_03829_ ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_03830_ ) );
AOI21_X1 _11541_ ( .A(_03827_ ), .B1(_03828_ ), .B2(_03830_ ), .ZN(_00207_ ) );
NAND3_X1 _11542_ ( .A1(_03811_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(\EX_LS_flag [2] ), .ZN(_03831_ ) );
NAND2_X1 _11543_ ( .A1(_03829_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_03832_ ) );
AOI21_X1 _11544_ ( .A(_03827_ ), .B1(_03831_ ), .B2(_03832_ ), .ZN(_00208_ ) );
NAND3_X1 _11545_ ( .A1(_03811_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(\EX_LS_flag [2] ), .ZN(_03833_ ) );
NAND2_X1 _11546_ ( .A1(_03829_ ), .A2(\LS_WB_waddr_csreg [5] ), .ZN(_03834_ ) );
AOI21_X1 _11547_ ( .A(_03827_ ), .B1(_03833_ ), .B2(_03834_ ), .ZN(_00209_ ) );
NAND3_X1 _11548_ ( .A1(_03811_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(\EX_LS_flag [2] ), .ZN(_03835_ ) );
NAND2_X1 _11549_ ( .A1(_03829_ ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_03836_ ) );
AOI21_X1 _11550_ ( .A(_03827_ ), .B1(_03835_ ), .B2(_03836_ ), .ZN(_00210_ ) );
NAND3_X1 _11551_ ( .A1(_03811_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(\EX_LS_flag [2] ), .ZN(_03837_ ) );
NAND2_X1 _11552_ ( .A1(_03829_ ), .A2(\LS_WB_waddr_csreg [3] ), .ZN(_03838_ ) );
AOI21_X1 _11553_ ( .A(_03827_ ), .B1(_03837_ ), .B2(_03838_ ), .ZN(_00211_ ) );
NAND3_X1 _11554_ ( .A1(_03811_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(\EX_LS_flag [2] ), .ZN(_03839_ ) );
NAND2_X1 _11555_ ( .A1(_03829_ ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_03840_ ) );
AOI21_X1 _11556_ ( .A(_03827_ ), .B1(_03839_ ), .B2(_03840_ ), .ZN(_00212_ ) );
NAND3_X1 _11557_ ( .A1(_03811_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(\EX_LS_flag [2] ), .ZN(_03841_ ) );
NAND2_X1 _11558_ ( .A1(_03829_ ), .A2(\LS_WB_waddr_csreg [1] ), .ZN(_03842_ ) );
AOI21_X1 _11559_ ( .A(_03827_ ), .B1(_03841_ ), .B2(_03842_ ), .ZN(_00213_ ) );
INV_X1 _11560_ ( .A(\EX_LS_dest_csreg_mem [9] ), .ZN(_03843_ ) );
INV_X1 _11561_ ( .A(\EX_LS_flag [0] ), .ZN(_03844_ ) );
AND4_X1 _11562_ ( .A1(_03843_ ), .A2(_03844_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03845_ ) );
NOR2_X1 _11563_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [9] ), .ZN(_03846_ ) );
OAI211_X1 _11564_ ( .A(_03825_ ), .B(_02018_ ), .C1(_03845_ ), .C2(_03846_ ), .ZN(_00214_ ) );
INV_X1 _11565_ ( .A(\EX_LS_dest_csreg_mem [8] ), .ZN(_03847_ ) );
AND4_X1 _11566_ ( .A1(_03847_ ), .A2(_03844_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03848_ ) );
NOR2_X1 _11567_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_03849_ ) );
OAI211_X1 _11568_ ( .A(_03825_ ), .B(_02018_ ), .C1(_03848_ ), .C2(_03849_ ), .ZN(_00215_ ) );
INV_X1 _11569_ ( .A(\EX_LS_dest_csreg_mem [6] ), .ZN(_03850_ ) );
AND4_X1 _11570_ ( .A1(_03850_ ), .A2(_03844_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03851_ ) );
NOR2_X1 _11571_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_03852_ ) );
OAI211_X1 _11572_ ( .A(_03825_ ), .B(_02018_ ), .C1(_03851_ ), .C2(_03852_ ), .ZN(_00216_ ) );
INV_X1 _11573_ ( .A(fanout_net_7 ), .ZN(_03853_ ) );
AND4_X1 _11574_ ( .A1(_03853_ ), .A2(_03844_ ), .A3(\EX_LS_flag [2] ), .A4(\EX_LS_flag [1] ), .ZN(_03854_ ) );
NOR2_X1 _11575_ ( .A1(\EX_LS_flag [2] ), .A2(\LS_WB_waddr_csreg [0] ), .ZN(_03855_ ) );
OAI211_X1 _11576_ ( .A(_03825_ ), .B(_02018_ ), .C1(_03854_ ), .C2(_03855_ ), .ZN(_00217_ ) );
INV_X1 _11577_ ( .A(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(_03856_ ) );
AND2_X1 _11578_ ( .A1(_03809_ ), .A2(_03856_ ), .ZN(_03857_ ) );
NOR2_X1 _11579_ ( .A1(\mylsu.state [3] ), .A2(\mylsu.state [1] ), .ZN(_03858_ ) );
NAND2_X1 _11580_ ( .A1(_03857_ ), .A2(_03858_ ), .ZN(_03859_ ) );
OAI211_X1 _11581_ ( .A(_02034_ ), .B(_02083_ ), .C1(_02080_ ), .C2(_02081_ ), .ZN(_03860_ ) );
AND2_X1 _11582_ ( .A1(_03860_ ), .A2(\EX_LS_flag [2] ), .ZN(_03861_ ) );
NOR3_X1 _11583_ ( .A1(_02019_ ), .A2(_02032_ ), .A3(_03861_ ), .ZN(_03862_ ) );
AOI21_X1 _11584_ ( .A(_03859_ ), .B1(_03825_ ), .B2(_03862_ ), .ZN(_00218_ ) );
INV_X1 _11585_ ( .A(_03811_ ), .ZN(_03863_ ) );
AOI21_X1 _11586_ ( .A(_02074_ ), .B1(_03861_ ), .B2(_03863_ ), .ZN(_03864_ ) );
AOI21_X1 _11587_ ( .A(_03859_ ), .B1(_03864_ ), .B2(_03825_ ), .ZN(_00219_ ) );
INV_X1 _11588_ ( .A(_02082_ ), .ZN(_03865_ ) );
AND2_X1 _11589_ ( .A1(_01944_ ), .A2(\EX_LS_flag [2] ), .ZN(_03866_ ) );
NAND3_X1 _11590_ ( .A1(_03865_ ), .A2(_02083_ ), .A3(_03866_ ), .ZN(_03867_ ) );
NOR2_X1 _11591_ ( .A1(_03867_ ), .A2(_03859_ ), .ZN(_00220_ ) );
INV_X1 _11592_ ( .A(_03813_ ), .ZN(_03868_ ) );
BUF_X4 _11593_ ( .A(_03868_ ), .Z(_03869_ ) );
AOI21_X1 _11594_ ( .A(_03859_ ), .B1(_03869_ ), .B2(_02033_ ), .ZN(_00221_ ) );
AOI21_X1 _11595_ ( .A(_03859_ ), .B1(_03825_ ), .B2(_03867_ ), .ZN(_00222_ ) );
AND3_X1 _11596_ ( .A1(_02056_ ), .A2(\myclint.rvalid ), .A3(_02059_ ), .ZN(_03870_ ) );
INV_X1 _11597_ ( .A(_03870_ ), .ZN(_03871_ ) );
OAI21_X1 _11598_ ( .A(_03871_ ), .B1(_02060_ ), .B2(io_master_arready ), .ZN(_03872_ ) );
INV_X1 _11599_ ( .A(_01979_ ), .ZN(_03873_ ) );
BUF_X4 _11600_ ( .A(_03873_ ), .Z(_03874_ ) );
NOR2_X1 _11601_ ( .A1(_03872_ ), .A2(_03874_ ), .ZN(_03875_ ) );
NOR3_X1 _11602_ ( .A1(_02084_ ), .A2(_02035_ ), .A3(_01945_ ), .ZN(_03876_ ) );
OAI21_X1 _11603_ ( .A(_03876_ ), .B1(_02082_ ), .B2(\EX_LS_flag [1] ), .ZN(_03877_ ) );
OAI21_X1 _11604_ ( .A(_02016_ ), .B1(_03875_ ), .B2(_03877_ ), .ZN(_03878_ ) );
INV_X1 _11605_ ( .A(_02032_ ), .ZN(_03879_ ) );
NAND3_X1 _11606_ ( .A1(_03878_ ), .A2(_02017_ ), .A3(_03879_ ), .ZN(_03880_ ) );
INV_X1 _11607_ ( .A(_02038_ ), .ZN(_03881_ ) );
NAND3_X1 _11608_ ( .A1(_03880_ ), .A2(_03881_ ), .A3(_03877_ ), .ZN(_03882_ ) );
INV_X1 _11609_ ( .A(_02045_ ), .ZN(_03883_ ) );
INV_X1 _11610_ ( .A(_03816_ ), .ZN(_03884_ ) );
AND4_X1 _11611_ ( .A1(EXU_valid_LSU ), .A2(_03882_ ), .A3(_03883_ ), .A4(_03884_ ), .ZN(_03885_ ) );
AND3_X1 _11612_ ( .A1(_03885_ ), .A2(_03810_ ), .A3(_03858_ ), .ZN(_00223_ ) );
INV_X1 _11613_ ( .A(_00205_ ), .ZN(_03886_ ) );
AND4_X1 _11614_ ( .A1(_01456_ ), .A2(fanout_net_5 ), .A3(EXU_valid_LSU ), .A4(_03858_ ), .ZN(_03887_ ) );
NOR2_X1 _11615_ ( .A1(_03844_ ), .A2(\EX_LS_flag [1] ), .ZN(_03888_ ) );
OAI21_X1 _11616_ ( .A(_03887_ ), .B1(_03888_ ), .B2(_03824_ ), .ZN(_03889_ ) );
OAI21_X1 _11617_ ( .A(_03886_ ), .B1(_02038_ ), .B2(_03889_ ), .ZN(_00224_ ) );
INV_X1 _11618_ ( .A(\mysc.state [2] ), .ZN(_03890_ ) );
NOR2_X1 _11619_ ( .A1(_03890_ ), .A2(fanout_net_3 ), .ZN(_00225_ ) );
AND3_X1 _11620_ ( .A1(_01457_ ), .A2(\LS_WB_wen_csreg [6] ), .A3(\LS_WB_wen_csreg [7] ), .ZN(_00094_ ) );
AND2_X1 _11621_ ( .A1(_02049_ ), .A2(\myifu.myicache.valid_data_in ), .ZN(_03891_ ) );
CLKBUF_X2 _11622_ ( .A(_03891_ ), .Z(\myifu.wen_$_ANDNOT__A_Y ) );
NOR2_X2 _11623_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .ZN(_03892_ ) );
BUF_X2 _11624_ ( .A(_03892_ ), .Z(_03893_ ) );
AND3_X1 _11625_ ( .A1(_02049_ ), .A2(_03893_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(_00164_ ) );
AND3_X1 _11626_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_03726_ ), .A3(fanout_net_12 ), .ZN(_00165_ ) );
AND3_X1 _11627_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(fanout_net_16 ), .A3(_03737_ ), .ZN(_00166_ ) );
CLKBUF_X2 _11628_ ( .A(_02012_ ), .Z(_03894_ ) );
CLKBUF_X2 _11629_ ( .A(_03894_ ), .Z(\io_master_arburst [0] ) );
CLKBUF_X2 _11630_ ( .A(_01971_ ), .Z(_03895_ ) );
NOR3_X1 _11631_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .A3(fanout_net_20 ), .ZN(_03896_ ) );
BUF_X4 _11632_ ( .A(_03874_ ), .Z(_03897_ ) );
BUF_X4 _11633_ ( .A(_03897_ ), .Z(_03898_ ) );
BUF_X4 _11634_ ( .A(_03898_ ), .Z(_03899_ ) );
INV_X1 _11635_ ( .A(\mylsu.araddr_tmp [1] ), .ZN(_03900_ ) );
INV_X1 _11636_ ( .A(_01973_ ), .ZN(_03901_ ) );
AOI211_X1 _11637_ ( .A(_03896_ ), .B(_03899_ ), .C1(_03900_ ), .C2(_03901_ ), .ZN(\io_master_araddr [1] ) );
NOR3_X1 _11638_ ( .A1(_03895_ ), .A2(fanout_net_7 ), .A3(fanout_net_20 ), .ZN(_03902_ ) );
INV_X1 _11639_ ( .A(\mylsu.araddr_tmp [0] ), .ZN(_03903_ ) );
AOI211_X1 _11640_ ( .A(_03902_ ), .B(_03899_ ), .C1(_03903_ ), .C2(_03901_ ), .ZN(\io_master_araddr [0] ) );
OAI221_X1 _11641_ ( .A(\IF_ID_pc [15] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01930_ ), .C2(_01931_ ), .ZN(_03904_ ) );
OR3_X1 _11642_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [15] ), .A3(fanout_net_20 ), .ZN(_03905_ ) );
BUF_X4 _11643_ ( .A(_01973_ ), .Z(_03906_ ) );
OAI211_X1 _11644_ ( .A(_01961_ ), .B(_03905_ ), .C1(\mylsu.araddr_tmp [15] ), .C2(_03906_ ), .ZN(_03907_ ) );
OAI21_X1 _11645_ ( .A(_03904_ ), .B1(\io_master_arburst [0] ), .B2(_03907_ ), .ZN(\io_master_araddr [15] ) );
OR3_X1 _11646_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [14] ), .A3(fanout_net_20 ), .ZN(_03908_ ) );
OAI21_X1 _11647_ ( .A(_03908_ ), .B1(_03906_ ), .B2(\mylsu.araddr_tmp [14] ), .ZN(_03909_ ) );
BUF_X4 _11648_ ( .A(_03796_ ), .Z(_03910_ ) );
BUF_X4 _11649_ ( .A(_03910_ ), .Z(_03911_ ) );
OAI22_X1 _11650_ ( .A1(_03899_ ), .A2(_03909_ ), .B1(_03552_ ), .B2(_03911_ ), .ZN(\io_master_araddr [14] ) );
OAI221_X1 _11651_ ( .A(\IF_ID_pc [5] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01930_ ), .C2(_01931_ ), .ZN(_03912_ ) );
OR3_X1 _11652_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [5] ), .A3(fanout_net_20 ), .ZN(_03913_ ) );
OAI211_X1 _11653_ ( .A(_01961_ ), .B(_03913_ ), .C1(\mylsu.araddr_tmp [5] ), .C2(_03906_ ), .ZN(_03914_ ) );
OAI21_X1 _11654_ ( .A(_03912_ ), .B1(\io_master_arburst [0] ), .B2(_03914_ ), .ZN(\io_master_araddr [5] ) );
OR3_X1 _11655_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [4] ), .A3(fanout_net_20 ), .ZN(_03915_ ) );
OAI21_X1 _11656_ ( .A(_03915_ ), .B1(_03906_ ), .B2(\mylsu.araddr_tmp [4] ), .ZN(_03916_ ) );
BUF_X2 _11657_ ( .A(_03796_ ), .Z(_03917_ ) );
OAI22_X1 _11658_ ( .A1(_03899_ ), .A2(_03916_ ), .B1(_03726_ ), .B2(_03917_ ), .ZN(\io_master_araddr [4] ) );
OAI221_X1 _11659_ ( .A(fanout_net_12 ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01930_ ), .C2(_01931_ ), .ZN(_03918_ ) );
OR3_X1 _11660_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [3] ), .A3(fanout_net_20 ), .ZN(_03919_ ) );
OAI211_X1 _11661_ ( .A(_01961_ ), .B(_03919_ ), .C1(\mylsu.araddr_tmp [3] ), .C2(_03906_ ), .ZN(_03920_ ) );
OAI21_X1 _11662_ ( .A(_03918_ ), .B1(\io_master_arburst [0] ), .B2(_03920_ ), .ZN(\io_master_araddr [3] ) );
OAI221_X1 _11663_ ( .A(\IF_ID_pc [13] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01930_ ), .C2(_01931_ ), .ZN(_03921_ ) );
OR3_X1 _11664_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [13] ), .A3(fanout_net_20 ), .ZN(_03922_ ) );
OAI211_X1 _11665_ ( .A(_01961_ ), .B(_03922_ ), .C1(\mylsu.araddr_tmp [13] ), .C2(_03906_ ), .ZN(_03923_ ) );
OAI21_X1 _11666_ ( .A(_03921_ ), .B1(\io_master_arburst [0] ), .B2(_03923_ ), .ZN(\io_master_araddr [13] ) );
OAI221_X1 _11667_ ( .A(\IF_ID_pc [12] ), .B1(\myminixbar.state [2] ), .B2(\myminixbar.state [0] ), .C1(_01930_ ), .C2(_01931_ ), .ZN(_03924_ ) );
OR3_X1 _11668_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [12] ), .A3(fanout_net_20 ), .ZN(_03925_ ) );
OAI211_X1 _11669_ ( .A(_01961_ ), .B(_03925_ ), .C1(\mylsu.araddr_tmp [12] ), .C2(_03906_ ), .ZN(_03926_ ) );
OAI21_X1 _11670_ ( .A(_03924_ ), .B1(\io_master_arburst [0] ), .B2(_03926_ ), .ZN(\io_master_araddr [12] ) );
NAND4_X1 _11671_ ( .A1(_01942_ ), .A2(_03821_ ), .A3(_01944_ ), .A4(_01945_ ), .ZN(_03927_ ) );
OAI21_X1 _11672_ ( .A(_03927_ ), .B1(_03906_ ), .B2(\mylsu.araddr_tmp [11] ), .ZN(_03928_ ) );
OAI22_X1 _11673_ ( .A1(_03899_ ), .A2(_03928_ ), .B1(_03521_ ), .B2(_03917_ ), .ZN(\io_master_araddr [11] ) );
OR3_X1 _11674_ ( .A1(_03895_ ), .A2(\EX_LS_dest_csreg_mem [10] ), .A3(fanout_net_20 ), .ZN(_03929_ ) );
OAI21_X1 _11675_ ( .A(_03929_ ), .B1(_03906_ ), .B2(\mylsu.araddr_tmp [10] ), .ZN(_03930_ ) );
OAI22_X1 _11676_ ( .A1(_03899_ ), .A2(_03930_ ), .B1(_03516_ ), .B2(_03917_ ), .ZN(\io_master_araddr [10] ) );
NAND4_X1 _11677_ ( .A1(_01942_ ), .A2(_03843_ ), .A3(_01944_ ), .A4(_01945_ ), .ZN(_03931_ ) );
OAI21_X1 _11678_ ( .A(_03931_ ), .B1(_03906_ ), .B2(\mylsu.araddr_tmp [9] ), .ZN(_03932_ ) );
OAI22_X1 _11679_ ( .A1(_03899_ ), .A2(_03932_ ), .B1(_01794_ ), .B2(_03917_ ), .ZN(\io_master_araddr [9] ) );
NOR3_X1 _11680_ ( .A1(_01971_ ), .A2(_03847_ ), .A3(fanout_net_20 ), .ZN(_03933_ ) );
AOI21_X1 _11681_ ( .A(_03933_ ), .B1(_03901_ ), .B2(\mylsu.araddr_tmp [8] ), .ZN(_03934_ ) );
NOR2_X1 _11682_ ( .A1(_03934_ ), .A2(_01939_ ), .ZN(_03935_ ) );
MUX2_X1 _11683_ ( .A(_03935_ ), .B(\IF_ID_pc [8] ), .S(_03894_ ), .Z(\io_master_araddr [8] ) );
NOR2_X1 _11684_ ( .A1(_01973_ ), .A2(\mylsu.araddr_tmp [7] ), .ZN(_03936_ ) );
NOR3_X1 _11685_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [7] ), .A3(fanout_net_20 ), .ZN(_03937_ ) );
NOR3_X1 _11686_ ( .A1(_01939_ ), .A2(_03936_ ), .A3(_03937_ ), .ZN(_03938_ ) );
MUX2_X1 _11687_ ( .A(_03938_ ), .B(\IF_ID_pc [7] ), .S(_03894_ ), .Z(\io_master_araddr [7] ) );
NOR3_X1 _11688_ ( .A1(_03895_ ), .A2(_03850_ ), .A3(fanout_net_20 ), .ZN(_03939_ ) );
AOI21_X1 _11689_ ( .A(_03939_ ), .B1(_03901_ ), .B2(\mylsu.araddr_tmp [6] ), .ZN(_03940_ ) );
OAI22_X1 _11690_ ( .A1(_03899_ ), .A2(_03940_ ), .B1(_03496_ ), .B2(_03917_ ), .ZN(\io_master_araddr [6] ) );
OR3_X1 _11691_ ( .A1(_01971_ ), .A2(\EX_LS_dest_csreg_mem [2] ), .A3(fanout_net_20 ), .ZN(_03941_ ) );
OAI211_X1 _11692_ ( .A(_01961_ ), .B(_03941_ ), .C1(\mylsu.araddr_tmp [2] ), .C2(_01973_ ), .ZN(_03942_ ) );
NOR2_X1 _11693_ ( .A1(_01964_ ), .A2(_03942_ ), .ZN(_03943_ ) );
BUF_X4 _11694_ ( .A(_03943_ ), .Z(_03944_ ) );
BUF_X4 _11695_ ( .A(_03944_ ), .Z(_03945_ ) );
BUF_X2 _11696_ ( .A(_03945_ ), .Z(\io_master_araddr [2] ) );
CLKBUF_X2 _11697_ ( .A(_01979_ ), .Z(\io_master_arid [1] ) );
AND3_X1 _11698_ ( .A1(_03917_ ), .A2(\EX_LS_typ [3] ), .A3(_01961_ ), .ZN(\io_master_arsize [2] ) );
AND3_X1 _11699_ ( .A1(_03917_ ), .A2(\EX_LS_typ [1] ), .A3(_01961_ ), .ZN(\io_master_arsize [0] ) );
OAI22_X1 _11700_ ( .A1(_01932_ ), .A2(_01933_ ), .B1(_02022_ ), .B2(_01939_ ), .ZN(\io_master_arsize [1] ) );
AOI211_X1 _11701_ ( .A(_02063_ ), .B(_02064_ ), .C1(_02056_ ), .C2(_02059_ ), .ZN(io_master_arvalid ) );
AND2_X1 _11702_ ( .A1(\mylsu.state [0] ), .A2(EXU_valid_LSU ), .ZN(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ) );
AND2_X1 _11703_ ( .A1(_02036_ ), .A2(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_03946_ ) );
BUF_X4 _11704_ ( .A(_03946_ ), .Z(_03947_ ) );
BUF_X4 _11705_ ( .A(_03947_ ), .Z(_03948_ ) );
MUX2_X1 _11706_ ( .A(\mylsu.awaddr_tmp [31] ), .B(\EX_LS_dest_csreg_mem [31] ), .S(_03948_ ), .Z(\io_master_awaddr [31] ) );
MUX2_X1 _11707_ ( .A(\mylsu.awaddr_tmp [30] ), .B(\EX_LS_dest_csreg_mem [30] ), .S(_03948_ ), .Z(\io_master_awaddr [30] ) );
MUX2_X1 _11708_ ( .A(\mylsu.awaddr_tmp [21] ), .B(\EX_LS_dest_csreg_mem [21] ), .S(_03948_ ), .Z(\io_master_awaddr [21] ) );
MUX2_X1 _11709_ ( .A(\mylsu.awaddr_tmp [20] ), .B(\EX_LS_dest_csreg_mem [20] ), .S(_03948_ ), .Z(\io_master_awaddr [20] ) );
MUX2_X1 _11710_ ( .A(\mylsu.awaddr_tmp [19] ), .B(\EX_LS_dest_csreg_mem [19] ), .S(_03948_ ), .Z(\io_master_awaddr [19] ) );
MUX2_X1 _11711_ ( .A(\mylsu.awaddr_tmp [18] ), .B(\EX_LS_dest_csreg_mem [18] ), .S(_03948_ ), .Z(\io_master_awaddr [18] ) );
MUX2_X1 _11712_ ( .A(\mylsu.awaddr_tmp [17] ), .B(\EX_LS_dest_csreg_mem [17] ), .S(_03948_ ), .Z(\io_master_awaddr [17] ) );
MUX2_X1 _11713_ ( .A(\mylsu.awaddr_tmp [16] ), .B(\EX_LS_dest_csreg_mem [16] ), .S(_03948_ ), .Z(\io_master_awaddr [16] ) );
BUF_X4 _11714_ ( .A(_03947_ ), .Z(_03949_ ) );
MUX2_X1 _11715_ ( .A(\mylsu.awaddr_tmp [15] ), .B(\EX_LS_dest_csreg_mem [15] ), .S(_03949_ ), .Z(\io_master_awaddr [15] ) );
MUX2_X1 _11716_ ( .A(\mylsu.awaddr_tmp [14] ), .B(\EX_LS_dest_csreg_mem [14] ), .S(_03949_ ), .Z(\io_master_awaddr [14] ) );
MUX2_X1 _11717_ ( .A(\mylsu.awaddr_tmp [13] ), .B(\EX_LS_dest_csreg_mem [13] ), .S(_03949_ ), .Z(\io_master_awaddr [13] ) );
MUX2_X1 _11718_ ( .A(\mylsu.awaddr_tmp [12] ), .B(\EX_LS_dest_csreg_mem [12] ), .S(_03949_ ), .Z(\io_master_awaddr [12] ) );
MUX2_X1 _11719_ ( .A(\mylsu.awaddr_tmp [29] ), .B(\EX_LS_dest_csreg_mem [29] ), .S(_03949_ ), .Z(\io_master_awaddr [29] ) );
MUX2_X1 _11720_ ( .A(\mylsu.awaddr_tmp [11] ), .B(\EX_LS_dest_csreg_mem [11] ), .S(_03949_ ), .Z(\io_master_awaddr [11] ) );
MUX2_X1 _11721_ ( .A(\mylsu.awaddr_tmp [10] ), .B(\EX_LS_dest_csreg_mem [10] ), .S(_03949_ ), .Z(\io_master_awaddr [10] ) );
MUX2_X1 _11722_ ( .A(\mylsu.awaddr_tmp [9] ), .B(\EX_LS_dest_csreg_mem [9] ), .S(_03949_ ), .Z(\io_master_awaddr [9] ) );
MUX2_X1 _11723_ ( .A(\mylsu.awaddr_tmp [8] ), .B(\EX_LS_dest_csreg_mem [8] ), .S(_03949_ ), .Z(\io_master_awaddr [8] ) );
MUX2_X1 _11724_ ( .A(\mylsu.awaddr_tmp [7] ), .B(\EX_LS_dest_csreg_mem [7] ), .S(_03949_ ), .Z(\io_master_awaddr [7] ) );
BUF_X4 _11725_ ( .A(_03947_ ), .Z(_03950_ ) );
MUX2_X1 _11726_ ( .A(\mylsu.awaddr_tmp [6] ), .B(\EX_LS_dest_csreg_mem [6] ), .S(_03950_ ), .Z(\io_master_awaddr [6] ) );
MUX2_X1 _11727_ ( .A(\mylsu.awaddr_tmp [5] ), .B(\EX_LS_dest_csreg_mem [5] ), .S(_03950_ ), .Z(\io_master_awaddr [5] ) );
MUX2_X1 _11728_ ( .A(\mylsu.awaddr_tmp [4] ), .B(\EX_LS_dest_csreg_mem [4] ), .S(_03950_ ), .Z(\io_master_awaddr [4] ) );
MUX2_X1 _11729_ ( .A(\mylsu.awaddr_tmp [3] ), .B(\EX_LS_dest_csreg_mem [3] ), .S(_03950_ ), .Z(\io_master_awaddr [3] ) );
MUX2_X1 _11730_ ( .A(\mylsu.awaddr_tmp [2] ), .B(\EX_LS_dest_csreg_mem [2] ), .S(_03950_ ), .Z(\io_master_awaddr [2] ) );
MUX2_X1 _11731_ ( .A(\mylsu.awaddr_tmp [28] ), .B(\EX_LS_dest_csreg_mem [28] ), .S(_03950_ ), .Z(\io_master_awaddr [28] ) );
MUX2_X1 _11732_ ( .A(\mylsu.awaddr_tmp [1] ), .B(\EX_LS_dest_csreg_mem [1] ), .S(_03950_ ), .Z(\io_master_awaddr [1] ) );
MUX2_X1 _11733_ ( .A(\mylsu.awaddr_tmp [0] ), .B(fanout_net_7 ), .S(_03950_ ), .Z(\io_master_awaddr [0] ) );
MUX2_X1 _11734_ ( .A(\mylsu.awaddr_tmp [27] ), .B(\EX_LS_dest_csreg_mem [27] ), .S(_03950_ ), .Z(\io_master_awaddr [27] ) );
MUX2_X1 _11735_ ( .A(\mylsu.awaddr_tmp [26] ), .B(\EX_LS_dest_csreg_mem [26] ), .S(_03950_ ), .Z(\io_master_awaddr [26] ) );
MUX2_X1 _11736_ ( .A(\mylsu.awaddr_tmp [25] ), .B(\EX_LS_dest_csreg_mem [25] ), .S(_03947_ ), .Z(\io_master_awaddr [25] ) );
MUX2_X1 _11737_ ( .A(\mylsu.awaddr_tmp [24] ), .B(\EX_LS_dest_csreg_mem [24] ), .S(_03947_ ), .Z(\io_master_awaddr [24] ) );
MUX2_X1 _11738_ ( .A(\mylsu.awaddr_tmp [23] ), .B(\EX_LS_dest_csreg_mem [23] ), .S(_03947_ ), .Z(\io_master_awaddr [23] ) );
MUX2_X1 _11739_ ( .A(\mylsu.awaddr_tmp [22] ), .B(\EX_LS_dest_csreg_mem [22] ), .S(_03947_ ), .Z(\io_master_awaddr [22] ) );
NAND3_X1 _11740_ ( .A1(_02030_ ), .A2(_03844_ ), .A3(\EX_LS_flag [1] ), .ZN(_03951_ ) );
NOR2_X1 _11741_ ( .A1(_03951_ ), .A2(\EX_LS_flag [2] ), .ZN(_03952_ ) );
AND4_X1 _11742_ ( .A1(\EX_LS_typ [1] ), .A2(_03952_ ), .A3(\EX_LS_typ [0] ), .A4(_02025_ ), .ZN(\io_master_awsize [0] ) );
NAND3_X1 _11743_ ( .A1(_03952_ ), .A2(\EX_LS_typ [0] ), .A3(_02025_ ), .ZN(\io_master_awsize [1] ) );
NAND3_X1 _11744_ ( .A1(_02033_ ), .A2(_02046_ ), .A3(_03948_ ), .ZN(_03953_ ) );
INV_X1 _11745_ ( .A(\mylsu.state [4] ), .ZN(_03954_ ) );
NAND2_X1 _11746_ ( .A1(_03953_ ), .A2(_03954_ ), .ZN(io_master_awvalid ) );
INV_X1 _11747_ ( .A(\mylsu.state [2] ), .ZN(_03955_ ) );
INV_X1 _11748_ ( .A(\mylsu.state [1] ), .ZN(_03956_ ) );
NAND4_X1 _11749_ ( .A1(_03953_ ), .A2(_03955_ ), .A3(_03954_ ), .A4(_03956_ ), .ZN(io_master_bready ) );
NOR3_X1 _11750_ ( .A1(_01938_ ), .A2(\mylsu.state [1] ), .A3(\mylsu.state [0] ), .ZN(_03957_ ) );
INV_X1 _11751_ ( .A(\mylsu.state [3] ), .ZN(_03958_ ) );
BUF_X2 _11752_ ( .A(_03958_ ), .Z(_03959_ ) );
NAND3_X1 _11753_ ( .A1(_02056_ ), .A2(\io_master_arid [1] ), .A3(_02059_ ), .ZN(_03960_ ) );
NOR2_X1 _11754_ ( .A1(_03799_ ), .A2(\io_master_rid [0] ), .ZN(_03961_ ) );
NAND4_X1 _11755_ ( .A1(_03961_ ), .A2(io_master_rlast ), .A3(_03797_ ), .A4(_03798_ ), .ZN(_03962_ ) );
OAI21_X1 _11756_ ( .A(_03960_ ), .B1(_03898_ ), .B2(_03962_ ), .ZN(_03963_ ) );
AOI21_X1 _11757_ ( .A(_03959_ ), .B1(_03795_ ), .B2(_03963_ ), .ZN(_03964_ ) );
NOR2_X1 _11758_ ( .A1(\io_master_bresp [1] ), .A2(\io_master_bresp [0] ), .ZN(_03965_ ) );
AND2_X1 _11759_ ( .A1(_03965_ ), .A2(io_master_bvalid ), .ZN(_03966_ ) );
NAND2_X1 _11760_ ( .A1(\io_master_bid [1] ), .A2(\io_master_bid [0] ), .ZN(_03967_ ) );
NOR3_X1 _11761_ ( .A1(_03967_ ), .A2(\io_master_bid [3] ), .A3(\io_master_bid [2] ), .ZN(_03968_ ) );
NAND2_X1 _11762_ ( .A1(_03966_ ), .A2(_03968_ ), .ZN(_03969_ ) );
AOI211_X1 _11763_ ( .A(_03957_ ), .B(_03964_ ), .C1(\mylsu.state [1] ), .C2(_03969_ ), .ZN(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ) );
AOI211_X1 _11764_ ( .A(_02048_ ), .B(_02051_ ), .C1(_02056_ ), .C2(_02059_ ), .ZN(io_master_rready ) );
MUX2_X1 _11765_ ( .A(\EX_LS_result_csreg_mem [15] ), .B(\EX_LS_result_csreg_mem [7] ), .S(fanout_net_7 ), .Z(_03970_ ) );
INV_X1 _11766_ ( .A(\EX_LS_dest_csreg_mem [1] ), .ZN(_03971_ ) );
CLKBUF_X2 _11767_ ( .A(_03971_ ), .Z(_03972_ ) );
AND2_X1 _11768_ ( .A1(_03970_ ), .A2(_03972_ ), .ZN(\io_master_wdata [15] ) );
MUX2_X1 _11769_ ( .A(\EX_LS_result_csreg_mem [14] ), .B(\EX_LS_result_csreg_mem [6] ), .S(fanout_net_7 ), .Z(_03973_ ) );
AND2_X1 _11770_ ( .A1(_03973_ ), .A2(_03972_ ), .ZN(\io_master_wdata [14] ) );
INV_X1 _11771_ ( .A(\EX_LS_result_csreg_mem [5] ), .ZN(_03974_ ) );
NOR3_X1 _11772_ ( .A1(_03974_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [5] ) );
INV_X1 _11773_ ( .A(\EX_LS_result_csreg_mem [4] ), .ZN(_03975_ ) );
NOR3_X1 _11774_ ( .A1(_03975_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [4] ) );
INV_X1 _11775_ ( .A(\EX_LS_result_csreg_mem [3] ), .ZN(_03976_ ) );
NOR3_X1 _11776_ ( .A1(_03976_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [3] ) );
INV_X1 _11777_ ( .A(\EX_LS_result_csreg_mem [2] ), .ZN(_03977_ ) );
NOR3_X1 _11778_ ( .A1(_03977_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [2] ) );
INV_X1 _11779_ ( .A(\EX_LS_result_csreg_mem [1] ), .ZN(_03978_ ) );
NOR3_X1 _11780_ ( .A1(_03978_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [1] ) );
INV_X1 _11781_ ( .A(\EX_LS_result_csreg_mem [0] ), .ZN(_03979_ ) );
NOR3_X1 _11782_ ( .A1(_03979_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [0] ) );
MUX2_X1 _11783_ ( .A(\EX_LS_result_csreg_mem [13] ), .B(\EX_LS_result_csreg_mem [5] ), .S(fanout_net_7 ), .Z(_03980_ ) );
AND2_X1 _11784_ ( .A1(_03980_ ), .A2(_03972_ ), .ZN(\io_master_wdata [13] ) );
MUX2_X1 _11785_ ( .A(\EX_LS_result_csreg_mem [12] ), .B(\EX_LS_result_csreg_mem [4] ), .S(fanout_net_7 ), .Z(_03981_ ) );
AND2_X1 _11786_ ( .A1(_03981_ ), .A2(_03972_ ), .ZN(\io_master_wdata [12] ) );
MUX2_X1 _11787_ ( .A(\EX_LS_result_csreg_mem [11] ), .B(\EX_LS_result_csreg_mem [3] ), .S(fanout_net_7 ), .Z(_03982_ ) );
AND2_X1 _11788_ ( .A1(_03982_ ), .A2(_03972_ ), .ZN(\io_master_wdata [11] ) );
MUX2_X1 _11789_ ( .A(\EX_LS_result_csreg_mem [10] ), .B(\EX_LS_result_csreg_mem [2] ), .S(fanout_net_7 ), .Z(_03983_ ) );
AND2_X1 _11790_ ( .A1(_03983_ ), .A2(_03972_ ), .ZN(\io_master_wdata [10] ) );
MUX2_X1 _11791_ ( .A(\EX_LS_result_csreg_mem [9] ), .B(\EX_LS_result_csreg_mem [1] ), .S(fanout_net_7 ), .Z(_03984_ ) );
AND2_X1 _11792_ ( .A1(_03984_ ), .A2(_03972_ ), .ZN(\io_master_wdata [9] ) );
MUX2_X1 _11793_ ( .A(\EX_LS_result_csreg_mem [8] ), .B(\EX_LS_result_csreg_mem [0] ), .S(fanout_net_7 ), .Z(_03985_ ) );
AND2_X1 _11794_ ( .A1(_03985_ ), .A2(_03972_ ), .ZN(\io_master_wdata [8] ) );
INV_X1 _11795_ ( .A(\EX_LS_result_csreg_mem [7] ), .ZN(_03986_ ) );
NOR3_X1 _11796_ ( .A1(_03986_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [7] ) );
INV_X1 _11797_ ( .A(\EX_LS_result_csreg_mem [6] ), .ZN(_03987_ ) );
NOR3_X1 _11798_ ( .A1(_03987_ ), .A2(fanout_net_7 ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wdata [6] ) );
MUX2_X1 _11799_ ( .A(\EX_LS_result_csreg_mem [31] ), .B(\EX_LS_result_csreg_mem [23] ), .S(fanout_net_7 ), .Z(_03988_ ) );
MUX2_X1 _11800_ ( .A(_03988_ ), .B(_03970_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [31] ) );
MUX2_X1 _11801_ ( .A(\EX_LS_result_csreg_mem [30] ), .B(\EX_LS_result_csreg_mem [22] ), .S(fanout_net_7 ), .Z(_03989_ ) );
MUX2_X1 _11802_ ( .A(_03989_ ), .B(_03973_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [30] ) );
NOR2_X1 _11803_ ( .A1(_03971_ ), .A2(fanout_net_7 ), .ZN(_03990_ ) );
INV_X1 _11804_ ( .A(_03990_ ), .ZN(_03991_ ) );
OAI21_X1 _11805_ ( .A(_03971_ ), .B1(_03853_ ), .B2(\EX_LS_result_csreg_mem [13] ), .ZN(_03992_ ) );
NOR2_X1 _11806_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [21] ), .ZN(_03993_ ) );
OAI22_X1 _11807_ ( .A1(_03991_ ), .A2(_03974_ ), .B1(_03992_ ), .B2(_03993_ ), .ZN(\io_master_wdata [21] ) );
OAI21_X1 _11808_ ( .A(_03971_ ), .B1(_03853_ ), .B2(\EX_LS_result_csreg_mem [12] ), .ZN(_03994_ ) );
NOR2_X1 _11809_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [20] ), .ZN(_03995_ ) );
OAI22_X1 _11810_ ( .A1(_03991_ ), .A2(_03975_ ), .B1(_03994_ ), .B2(_03995_ ), .ZN(\io_master_wdata [20] ) );
OAI21_X1 _11811_ ( .A(_03971_ ), .B1(_03853_ ), .B2(\EX_LS_result_csreg_mem [11] ), .ZN(_03996_ ) );
NOR2_X1 _11812_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [19] ), .ZN(_03997_ ) );
OAI22_X1 _11813_ ( .A1(_03991_ ), .A2(_03976_ ), .B1(_03996_ ), .B2(_03997_ ), .ZN(\io_master_wdata [19] ) );
INV_X1 _11814_ ( .A(\EX_LS_result_csreg_mem [18] ), .ZN(_03998_ ) );
INV_X1 _11815_ ( .A(\EX_LS_result_csreg_mem [10] ), .ZN(_03999_ ) );
MUX2_X1 _11816_ ( .A(_03998_ ), .B(_03999_ ), .S(fanout_net_7 ), .Z(_04000_ ) );
OAI22_X1 _11817_ ( .A1(_04000_ ), .A2(\EX_LS_dest_csreg_mem [1] ), .B1(_03991_ ), .B2(_03977_ ), .ZN(\io_master_wdata [18] ) );
OAI21_X1 _11818_ ( .A(_03971_ ), .B1(_03853_ ), .B2(\EX_LS_result_csreg_mem [9] ), .ZN(_04001_ ) );
NOR2_X1 _11819_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [17] ), .ZN(_04002_ ) );
OAI22_X1 _11820_ ( .A1(_03991_ ), .A2(_03978_ ), .B1(_04001_ ), .B2(_04002_ ), .ZN(\io_master_wdata [17] ) );
OAI21_X1 _11821_ ( .A(_03971_ ), .B1(_03853_ ), .B2(\EX_LS_result_csreg_mem [8] ), .ZN(_04003_ ) );
NOR2_X1 _11822_ ( .A1(fanout_net_7 ), .A2(\EX_LS_result_csreg_mem [16] ), .ZN(_04004_ ) );
OAI22_X1 _11823_ ( .A1(_03991_ ), .A2(_03979_ ), .B1(_04003_ ), .B2(_04004_ ), .ZN(\io_master_wdata [16] ) );
MUX2_X1 _11824_ ( .A(\EX_LS_result_csreg_mem [29] ), .B(\EX_LS_result_csreg_mem [21] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04005_ ) );
MUX2_X1 _11825_ ( .A(_04005_ ), .B(_03980_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [29] ) );
MUX2_X1 _11826_ ( .A(\EX_LS_result_csreg_mem [28] ), .B(\EX_LS_result_csreg_mem [20] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04006_ ) );
MUX2_X1 _11827_ ( .A(_04006_ ), .B(_03981_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [28] ) );
MUX2_X1 _11828_ ( .A(\EX_LS_result_csreg_mem [27] ), .B(\EX_LS_result_csreg_mem [19] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04007_ ) );
MUX2_X1 _11829_ ( .A(_04007_ ), .B(_03982_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [27] ) );
MUX2_X1 _11830_ ( .A(\EX_LS_result_csreg_mem [26] ), .B(\EX_LS_result_csreg_mem [18] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04008_ ) );
MUX2_X1 _11831_ ( .A(_04008_ ), .B(_03983_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [26] ) );
MUX2_X1 _11832_ ( .A(\EX_LS_result_csreg_mem [25] ), .B(\EX_LS_result_csreg_mem [17] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04009_ ) );
MUX2_X1 _11833_ ( .A(_04009_ ), .B(_03984_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [25] ) );
MUX2_X1 _11834_ ( .A(\EX_LS_result_csreg_mem [24] ), .B(\EX_LS_result_csreg_mem [16] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04010_ ) );
MUX2_X1 _11835_ ( .A(_04010_ ), .B(_03985_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wdata [24] ) );
OAI21_X1 _11836_ ( .A(_03971_ ), .B1(_03853_ ), .B2(\EX_LS_result_csreg_mem [15] ), .ZN(_04011_ ) );
NOR2_X1 _11837_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [23] ), .ZN(_04012_ ) );
OAI22_X1 _11838_ ( .A1(_03991_ ), .A2(_03986_ ), .B1(_04011_ ), .B2(_04012_ ), .ZN(\io_master_wdata [23] ) );
OAI21_X1 _11839_ ( .A(_03971_ ), .B1(_03853_ ), .B2(\EX_LS_result_csreg_mem [14] ), .ZN(_04013_ ) );
NOR2_X1 _11840_ ( .A1(\EX_LS_dest_csreg_mem [0] ), .A2(\EX_LS_result_csreg_mem [22] ), .ZN(_04014_ ) );
OAI22_X1 _11841_ ( .A1(_03991_ ), .A2(_03987_ ), .B1(_04013_ ), .B2(_04014_ ), .ZN(\io_master_wdata [22] ) );
NAND2_X1 _11842_ ( .A1(_02036_ ), .A2(EXU_valid_LSU ), .ZN(_04015_ ) );
INV_X1 _11843_ ( .A(io_master_awready ), .ZN(_04016_ ) );
INV_X1 _11844_ ( .A(io_master_wready ), .ZN(_04017_ ) );
AOI211_X1 _11845_ ( .A(io_master_wready_$_NOR__B_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ), .B(_04015_ ), .C1(_04016_ ), .C2(_04017_ ), .ZN(_04018_ ) );
AND4_X1 _11846_ ( .A1(_03881_ ), .A2(_04018_ ), .A3(_03883_ ), .A4(_03810_ ), .ZN(io_master_wready_$_NOR__B_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _11847_ ( .A(\EX_LS_typ [1] ), .B(\EX_LS_typ [0] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04019_ ) );
AND2_X1 _11848_ ( .A1(_04019_ ), .A2(_03972_ ), .ZN(\io_master_wstrb [1] ) );
NOR3_X1 _11849_ ( .A1(_02020_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_dest_csreg_mem [1] ), .ZN(\io_master_wstrb [0] ) );
MUX2_X1 _11850_ ( .A(\EX_LS_typ [3] ), .B(\EX_LS_typ [2] ), .S(\EX_LS_dest_csreg_mem [0] ), .Z(_04020_ ) );
MUX2_X1 _11851_ ( .A(_04020_ ), .B(_04019_ ), .S(\EX_LS_dest_csreg_mem [1] ), .Z(\io_master_wstrb [3] ) );
NAND3_X1 _11852_ ( .A1(_03972_ ), .A2(\EX_LS_dest_csreg_mem [0] ), .A3(\EX_LS_typ [1] ), .ZN(_04021_ ) );
OAI221_X1 _11853_ ( .A(_04021_ ), .B1(_02042_ ), .B2(_02022_ ), .C1(_03991_ ), .C2(_02020_ ), .ZN(\io_master_wstrb [2] ) );
NAND2_X1 _11854_ ( .A1(_03953_ ), .A2(_03955_ ), .ZN(io_master_wvalid ) );
MUX2_X1 _11855_ ( .A(\LS_WB_wdata_csreg [2] ), .B(\LS_WB_wen_csreg [2] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _11856_ ( .A(\LS_WB_wdata_csreg [1] ), .B(\LS_WB_wen_csreg [1] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _11857_ ( .A(\LS_WB_wdata_csreg [0] ), .B(\LS_WB_wen_csreg [0] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _11858_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\LS_WB_wen_csreg [3] ), .S(\LS_WB_wen_csreg [6] ), .Z(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ) );
AND3_X1 _11859_ ( .A1(_01457_ ), .A2(\LS_WB_wen_csreg [7] ), .A3(\LS_WB_waddr_csreg [2] ), .ZN(_04022_ ) );
NOR2_X1 _11860_ ( .A1(\LS_WB_waddr_csreg [5] ), .A2(\LS_WB_waddr_csreg [4] ), .ZN(_04023_ ) );
INV_X1 _11861_ ( .A(\LS_WB_waddr_csreg [7] ), .ZN(_04024_ ) );
INV_X1 _11862_ ( .A(\LS_WB_waddr_csreg [6] ), .ZN(_04025_ ) );
AND3_X1 _11863_ ( .A1(_04023_ ), .A2(_04024_ ), .A3(_04025_ ), .ZN(_04026_ ) );
OR2_X1 _11864_ ( .A1(\LS_WB_waddr_csreg [11] ), .A2(\LS_WB_waddr_csreg [10] ), .ZN(_04027_ ) );
NAND2_X1 _11865_ ( .A1(\LS_WB_waddr_csreg [9] ), .A2(\LS_WB_waddr_csreg [8] ), .ZN(_04028_ ) );
NOR2_X1 _11866_ ( .A1(_04027_ ), .A2(_04028_ ), .ZN(_04029_ ) );
INV_X1 _11867_ ( .A(\LS_WB_waddr_csreg [0] ), .ZN(_04030_ ) );
NOR3_X1 _11868_ ( .A1(_04030_ ), .A2(\LS_WB_waddr_csreg [1] ), .A3(\LS_WB_waddr_csreg [3] ), .ZN(_04031_ ) );
AND4_X1 _11869_ ( .A1(_04022_ ), .A2(_04026_ ), .A3(_04029_ ), .A4(_04031_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ) );
AND2_X1 _11870_ ( .A1(_01456_ ), .A2(\LS_WB_wen_csreg [7] ), .ZN(_04032_ ) );
NOR2_X1 _11871_ ( .A1(\LS_WB_waddr_csreg [3] ), .A2(\LS_WB_waddr_csreg [2] ), .ZN(_04033_ ) );
AND3_X1 _11872_ ( .A1(_04029_ ), .A2(_04032_ ), .A3(_04033_ ), .ZN(_04034_ ) );
INV_X1 _11873_ ( .A(\LS_WB_waddr_csreg [1] ), .ZN(_04035_ ) );
NAND2_X1 _11874_ ( .A1(_04023_ ), .A2(\LS_WB_waddr_csreg [6] ), .ZN(_04036_ ) );
NOR2_X1 _11875_ ( .A1(_04036_ ), .A2(\LS_WB_waddr_csreg [7] ), .ZN(_04037_ ) );
AND4_X1 _11876_ ( .A1(\LS_WB_waddr_csreg [0] ), .A2(_04034_ ), .A3(_04035_ ), .A4(_04037_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ) );
AND4_X1 _11877_ ( .A1(_04030_ ), .A2(_04029_ ), .A3(\LS_WB_waddr_csreg [1] ), .A4(_04033_ ), .ZN(_04038_ ) );
AND3_X1 _11878_ ( .A1(_04038_ ), .A2(_04032_ ), .A3(_04037_ ), .ZN(_04039_ ) );
OR2_X1 _11879_ ( .A1(_04039_ ), .A2(_00094_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_OR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
AND4_X1 _11880_ ( .A1(_04030_ ), .A2(_04034_ ), .A3(_04035_ ), .A4(_04026_ ), .ZN(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _11881_ ( .A(_02047_ ), .ZN(_04040_ ) );
AOI21_X1 _11882_ ( .A(exception_quest_IDU ), .B1(_03865_ ), .B2(_02083_ ), .ZN(_04041_ ) );
NOR2_X1 _11883_ ( .A1(_04040_ ), .A2(_04041_ ), .ZN(_04042_ ) );
BUF_X4 _11884_ ( .A(_04042_ ), .Z(_04043_ ) );
MUX2_X1 _11885_ ( .A(\EX_LS_pc [21] ), .B(\ID_EX_pc [21] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ) );
MUX2_X1 _11886_ ( .A(\EX_LS_pc [20] ), .B(\ID_EX_pc [20] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _11887_ ( .A(\EX_LS_pc [19] ), .B(\ID_EX_pc [19] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _11888_ ( .A(\EX_LS_pc [18] ), .B(\ID_EX_pc [18] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ) );
MUX2_X1 _11889_ ( .A(\EX_LS_pc [17] ), .B(\ID_EX_pc [17] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ) );
MUX2_X1 _11890_ ( .A(\EX_LS_pc [16] ), .B(\ID_EX_pc [16] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _11891_ ( .A(\EX_LS_pc [15] ), .B(\ID_EX_pc [15] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ) );
MUX2_X1 _11892_ ( .A(\EX_LS_pc [14] ), .B(\ID_EX_pc [14] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _11893_ ( .A(\EX_LS_pc [13] ), .B(\ID_EX_pc [13] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _11894_ ( .A(\EX_LS_pc [12] ), .B(\ID_EX_pc [12] ), .S(_04043_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ) );
BUF_X4 _11895_ ( .A(_04042_ ), .Z(_04044_ ) );
MUX2_X1 _11896_ ( .A(\EX_LS_pc [30] ), .B(\ID_EX_pc [30] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _11897_ ( .A(\EX_LS_pc [11] ), .B(\ID_EX_pc [11] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _11898_ ( .A(\EX_LS_pc [10] ), .B(\ID_EX_pc [10] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ) );
MUX2_X1 _11899_ ( .A(\EX_LS_pc [9] ), .B(\ID_EX_pc [9] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ) );
MUX2_X1 _11900_ ( .A(\EX_LS_pc [8] ), .B(\ID_EX_pc [8] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ) );
MUX2_X1 _11901_ ( .A(\EX_LS_pc [7] ), .B(\ID_EX_pc [7] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ) );
MUX2_X1 _11902_ ( .A(\EX_LS_pc [6] ), .B(\ID_EX_pc [6] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _11903_ ( .A(\EX_LS_pc [5] ), .B(\ID_EX_pc [5] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ) );
MUX2_X1 _11904_ ( .A(\EX_LS_pc [4] ), .B(\ID_EX_pc [4] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _11905_ ( .A(\EX_LS_pc [3] ), .B(\ID_EX_pc [3] ), .S(_04044_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ) );
BUF_X4 _11906_ ( .A(_04042_ ), .Z(_04045_ ) );
MUX2_X1 _11907_ ( .A(\EX_LS_pc [2] ), .B(\ID_EX_pc [2] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _11908_ ( .A(\EX_LS_pc [29] ), .B(\ID_EX_pc [29] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ) );
MUX2_X1 _11909_ ( .A(\EX_LS_pc [1] ), .B(\ID_EX_pc [1] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ) );
MUX2_X1 _11910_ ( .A(\EX_LS_pc [0] ), .B(\ID_EX_pc [0] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _11911_ ( .A(\EX_LS_pc [28] ), .B(\ID_EX_pc [28] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ) );
MUX2_X1 _11912_ ( .A(\EX_LS_pc [27] ), .B(\ID_EX_pc [27] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _11913_ ( .A(\EX_LS_pc [26] ), .B(\ID_EX_pc [26] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ) );
MUX2_X1 _11914_ ( .A(\EX_LS_pc [25] ), .B(\ID_EX_pc [25] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _11915_ ( .A(\EX_LS_pc [24] ), .B(\ID_EX_pc [24] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _11916_ ( .A(\EX_LS_pc [23] ), .B(\ID_EX_pc [23] ), .S(_04045_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _11917_ ( .A(\EX_LS_pc [22] ), .B(\ID_EX_pc [22] ), .S(_04042_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _11918_ ( .A(\EX_LS_pc [31] ), .B(\ID_EX_pc [31] ), .S(_04042_ ), .Z(\myec.mepc_tmp_$_DFFE_PP__Q_D ) );
INV_X1 _11919_ ( .A(_02076_ ), .ZN(_04046_ ) );
NOR4_X1 _11920_ ( .A1(_04040_ ), .A2(exception_quest_IDU ), .A3(_04046_ ), .A4(_04041_ ), .ZN(_04047_ ) );
XNOR2_X1 _11921_ ( .A(\mepc [30] ), .B(\myec.mepc_tmp [30] ), .ZN(_04048_ ) );
XNOR2_X1 _11922_ ( .A(\mepc [31] ), .B(\myec.mepc_tmp [31] ), .ZN(_04049_ ) );
XNOR2_X1 _11923_ ( .A(\mepc [28] ), .B(\myec.mepc_tmp [28] ), .ZN(_04050_ ) );
XNOR2_X1 _11924_ ( .A(\mepc [29] ), .B(\myec.mepc_tmp [29] ), .ZN(_04051_ ) );
AND4_X1 _11925_ ( .A1(_04048_ ), .A2(_04049_ ), .A3(_04050_ ), .A4(_04051_ ), .ZN(_04052_ ) );
XNOR2_X1 _11926_ ( .A(\mepc [24] ), .B(\myec.mepc_tmp [24] ), .ZN(_04053_ ) );
XNOR2_X1 _11927_ ( .A(\mepc [26] ), .B(\myec.mepc_tmp [26] ), .ZN(_04054_ ) );
XNOR2_X1 _11928_ ( .A(\mepc [27] ), .B(\myec.mepc_tmp [27] ), .ZN(_04055_ ) );
XNOR2_X1 _11929_ ( .A(\mepc [25] ), .B(\myec.mepc_tmp [25] ), .ZN(_04056_ ) );
AND4_X1 _11930_ ( .A1(_04053_ ), .A2(_04054_ ), .A3(_04055_ ), .A4(_04056_ ), .ZN(_04057_ ) );
XNOR2_X1 _11931_ ( .A(\mepc [20] ), .B(\myec.mepc_tmp [20] ), .ZN(_04058_ ) );
XNOR2_X1 _11932_ ( .A(\mepc [22] ), .B(\myec.mepc_tmp [22] ), .ZN(_04059_ ) );
XNOR2_X1 _11933_ ( .A(\mepc [23] ), .B(\myec.mepc_tmp [23] ), .ZN(_04060_ ) );
XNOR2_X1 _11934_ ( .A(\mepc [21] ), .B(\myec.mepc_tmp [21] ), .ZN(_04061_ ) );
AND4_X1 _11935_ ( .A1(_04058_ ), .A2(_04059_ ), .A3(_04060_ ), .A4(_04061_ ), .ZN(_04062_ ) );
XNOR2_X1 _11936_ ( .A(\mepc [18] ), .B(\myec.mepc_tmp [18] ), .ZN(_04063_ ) );
XNOR2_X1 _11937_ ( .A(\mepc [16] ), .B(\myec.mepc_tmp [16] ), .ZN(_04064_ ) );
XNOR2_X1 _11938_ ( .A(\mepc [19] ), .B(\myec.mepc_tmp [19] ), .ZN(_04065_ ) );
XNOR2_X1 _11939_ ( .A(\mepc [17] ), .B(\myec.mepc_tmp [17] ), .ZN(_04066_ ) );
AND4_X1 _11940_ ( .A1(_04063_ ), .A2(_04064_ ), .A3(_04065_ ), .A4(_04066_ ), .ZN(_04067_ ) );
AND4_X1 _11941_ ( .A1(_04052_ ), .A2(_04057_ ), .A3(_04062_ ), .A4(_04067_ ), .ZN(_04068_ ) );
XNOR2_X1 _11942_ ( .A(\mepc [12] ), .B(\myec.mepc_tmp [12] ), .ZN(_04069_ ) );
XNOR2_X1 _11943_ ( .A(\mepc [14] ), .B(\myec.mepc_tmp [14] ), .ZN(_04070_ ) );
XNOR2_X1 _11944_ ( .A(\mepc [15] ), .B(\myec.mepc_tmp [15] ), .ZN(_04071_ ) );
XNOR2_X1 _11945_ ( .A(\mepc [13] ), .B(\myec.mepc_tmp [13] ), .ZN(_04072_ ) );
AND4_X1 _11946_ ( .A1(_04069_ ), .A2(_04070_ ), .A3(_04071_ ), .A4(_04072_ ), .ZN(_04073_ ) );
XNOR2_X1 _11947_ ( .A(\mepc [8] ), .B(\myec.mepc_tmp [8] ), .ZN(_04074_ ) );
XNOR2_X1 _11948_ ( .A(\mepc [10] ), .B(\myec.mepc_tmp [10] ), .ZN(_04075_ ) );
XNOR2_X1 _11949_ ( .A(\mepc [11] ), .B(\myec.mepc_tmp [11] ), .ZN(_04076_ ) );
XNOR2_X1 _11950_ ( .A(\mepc [9] ), .B(\myec.mepc_tmp [9] ), .ZN(_04077_ ) );
AND4_X1 _11951_ ( .A1(_04074_ ), .A2(_04075_ ), .A3(_04076_ ), .A4(_04077_ ), .ZN(_04078_ ) );
XNOR2_X1 _11952_ ( .A(\mepc [6] ), .B(\myec.mepc_tmp [6] ), .ZN(_04079_ ) );
XNOR2_X1 _11953_ ( .A(\mepc [4] ), .B(\myec.mepc_tmp [4] ), .ZN(_04080_ ) );
XNOR2_X1 _11954_ ( .A(\mepc [7] ), .B(\myec.mepc_tmp [7] ), .ZN(_04081_ ) );
XNOR2_X1 _11955_ ( .A(\mepc [5] ), .B(\myec.mepc_tmp [5] ), .ZN(_04082_ ) );
AND4_X1 _11956_ ( .A1(_04079_ ), .A2(_04080_ ), .A3(_04081_ ), .A4(_04082_ ), .ZN(_04083_ ) );
XNOR2_X1 _11957_ ( .A(\mepc [2] ), .B(\myec.mepc_tmp [2] ), .ZN(_04084_ ) );
XNOR2_X1 _11958_ ( .A(\mepc [3] ), .B(\myec.mepc_tmp [3] ), .ZN(_04085_ ) );
XNOR2_X1 _11959_ ( .A(\mepc [1] ), .B(\myec.mepc_tmp [1] ), .ZN(_04086_ ) );
XNOR2_X1 _11960_ ( .A(\mepc [0] ), .B(\myec.mepc_tmp [0] ), .ZN(_04087_ ) );
AND4_X1 _11961_ ( .A1(_04084_ ), .A2(_04085_ ), .A3(_04086_ ), .A4(_04087_ ), .ZN(_04088_ ) );
AND4_X1 _11962_ ( .A1(_04073_ ), .A2(_04078_ ), .A3(_04083_ ), .A4(_04088_ ), .ZN(_04089_ ) );
NAND4_X1 _11963_ ( .A1(_04068_ ), .A2(_04089_ ), .A3(excp_written ), .A4(_04046_ ), .ZN(_04090_ ) );
AOI21_X1 _11964_ ( .A(_04047_ ), .B1(_04046_ ), .B2(_04090_ ), .ZN(\myec.state_$_SDFFE_PP0P__Q_E ) );
NAND2_X1 _11965_ ( .A1(_01941_ ), .A2(IDU_valid_EXU ), .ZN(_04091_ ) );
NOR2_X1 _11966_ ( .A1(_03730_ ), .A2(check_assert ), .ZN(_04092_ ) );
INV_X1 _11967_ ( .A(_04092_ ), .ZN(_04093_ ) );
NOR2_X1 _11968_ ( .A1(_03344_ ), .A2(\ID_EX_typ [6] ), .ZN(_04094_ ) );
INV_X1 _11969_ ( .A(_04094_ ), .ZN(_04095_ ) );
AOI211_X1 _11970_ ( .A(fanout_net_3 ), .B(_04091_ ), .C1(_04093_ ), .C2(_04095_ ), .ZN(_04096_ ) );
INV_X2 _11971_ ( .A(\ID_EX_typ [5] ), .ZN(_04097_ ) );
NAND3_X1 _11972_ ( .A1(_04094_ ), .A2(fanout_net_11 ), .A3(_04097_ ), .ZN(_04098_ ) );
NAND2_X1 _11973_ ( .A1(_04096_ ), .A2(_04098_ ), .ZN(_04099_ ) );
AND3_X1 _11974_ ( .A1(_04094_ ), .A2(\myexu.check_quest_$_DFF_PP0__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .A3(\ID_EX_typ [5] ), .ZN(_04100_ ) );
OAI21_X1 _11975_ ( .A(_01457_ ), .B1(_03328_ ), .B2(EXU_valid_LSU ), .ZN(\myifu.check_assert_$_ORNOT__A_Y_$_MUX__A_S_$_OR__A_Y_$_ANDNOT__A_B_$_NOR__B_Y ) );
OAI22_X1 _11976_ ( .A1(_04099_ ), .A2(_04100_ ), .B1(_04093_ ), .B2(\myifu.check_assert_$_ORNOT__A_Y_$_MUX__A_S_$_OR__A_Y_$_ANDNOT__A_B_$_NOR__B_Y ), .ZN(\myexu.check_quest_$_DFF_PP0__Q_D ) );
XOR2_X1 _11977_ ( .A(_02286_ ), .B(_02309_ ), .Z(_04101_ ) );
NAND2_X1 _11978_ ( .A1(_04101_ ), .A2(_03007_ ), .ZN(_04102_ ) );
INV_X1 _11979_ ( .A(\ID_EX_csr [1] ), .ZN(_04103_ ) );
AND2_X1 _11980_ ( .A1(_02991_ ), .A2(_04097_ ), .ZN(_04104_ ) );
BUF_X4 _11981_ ( .A(_04104_ ), .Z(_04105_ ) );
INV_X1 _11982_ ( .A(_04105_ ), .ZN(_04106_ ) );
BUF_X4 _11983_ ( .A(_04106_ ), .Z(_04107_ ) );
BUF_X4 _11984_ ( .A(_04107_ ), .Z(_04108_ ) );
OAI21_X1 _11985_ ( .A(_04102_ ), .B1(_04103_ ), .B2(_04108_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ) );
AND2_X1 _11986_ ( .A1(_02306_ ), .A2(_02308_ ), .ZN(_04109_ ) );
BUF_X4 _11987_ ( .A(_04109_ ), .Z(_04110_ ) );
XNOR2_X1 _11988_ ( .A(_04110_ ), .B(\ID_EX_imm [0] ), .ZN(_04111_ ) );
INV_X1 _11989_ ( .A(\ID_EX_csr [0] ), .ZN(_04112_ ) );
BUF_X4 _11990_ ( .A(_04105_ ), .Z(_04113_ ) );
BUF_X4 _11991_ ( .A(_04113_ ), .Z(_04114_ ) );
AOI22_X1 _11992_ ( .A1(_04111_ ), .A2(_03008_ ), .B1(_04112_ ), .B2(_04114_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ) );
AOI21_X1 _11993_ ( .A(_02583_ ), .B1(_02378_ ), .B2(_02474_ ), .ZN(_04115_ ) );
XOR2_X1 _11994_ ( .A(_04115_ ), .B(_02423_ ), .Z(_04116_ ) );
NAND2_X1 _11995_ ( .A1(_04116_ ), .A2(_03007_ ), .ZN(_04117_ ) );
INV_X1 _11996_ ( .A(\ID_EX_csr [10] ), .ZN(_04118_ ) );
OAI21_X1 _11997_ ( .A(_04117_ ), .B1(_04118_ ), .B2(_04108_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ) );
OAI21_X1 _11998_ ( .A(_02450_ ), .B1(_02373_ ), .B2(_02377_ ), .ZN(_04119_ ) );
AND2_X1 _11999_ ( .A1(_04119_ ), .A2(_02579_ ), .ZN(_04120_ ) );
XNOR2_X1 _12000_ ( .A(_04120_ ), .B(_02473_ ), .ZN(_04121_ ) );
INV_X1 _12001_ ( .A(\ID_EX_csr [9] ), .ZN(_04122_ ) );
AOI22_X1 _12002_ ( .A1(_04121_ ), .A2(_03008_ ), .B1(_04122_ ), .B2(_04114_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ) );
XNOR2_X1 _12003_ ( .A(_02378_ ), .B(_02451_ ), .ZN(_04123_ ) );
NOR2_X1 _12004_ ( .A1(_04123_ ), .A2(_02992_ ), .ZN(_04124_ ) );
INV_X1 _12005_ ( .A(\ID_EX_csr [8] ), .ZN(_04125_ ) );
BUF_X4 _12006_ ( .A(_04105_ ), .Z(_04126_ ) );
BUF_X4 _12007_ ( .A(_04126_ ), .Z(_04127_ ) );
AOI21_X1 _12008_ ( .A(_04124_ ), .B1(_04125_ ), .B2(_04127_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ) );
OR2_X1 _12009_ ( .A1(_02324_ ), .A2(_02372_ ), .ZN(_04128_ ) );
NAND2_X1 _12010_ ( .A1(_04128_ ), .A2(_02374_ ), .ZN(_04129_ ) );
XNOR2_X1 _12011_ ( .A(_04129_ ), .B(_02346_ ), .ZN(_04130_ ) );
AND2_X2 _12012_ ( .A1(_03343_ ), .A2(\ID_EX_typ [7] ), .ZN(_04131_ ) );
INV_X1 _12013_ ( .A(_04131_ ), .ZN(_04132_ ) );
BUF_X4 _12014_ ( .A(_04132_ ), .Z(_04133_ ) );
AND2_X1 _12015_ ( .A1(_04130_ ), .A2(_04133_ ), .ZN(_04134_ ) );
BUF_X4 _12016_ ( .A(_04106_ ), .Z(_04135_ ) );
MUX2_X1 _12017_ ( .A(\ID_EX_csr [7] ), .B(_04134_ ), .S(_04135_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ) );
XOR2_X1 _12018_ ( .A(_02324_ ), .B(_02372_ ), .Z(_04136_ ) );
NOR2_X1 _12019_ ( .A1(_04136_ ), .A2(_02992_ ), .ZN(_04137_ ) );
INV_X1 _12020_ ( .A(\ID_EX_csr [6] ), .ZN(_04138_ ) );
AOI21_X1 _12021_ ( .A(_04137_ ), .B1(_04138_ ), .B2(_04127_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ) );
INV_X1 _12022_ ( .A(_02322_ ), .ZN(_04139_ ) );
NAND2_X1 _12023_ ( .A1(_04139_ ), .A2(_02211_ ), .ZN(_04140_ ) );
XNOR2_X1 _12024_ ( .A(_04140_ ), .B(_02323_ ), .ZN(_04141_ ) );
INV_X1 _12025_ ( .A(\ID_EX_csr [5] ), .ZN(_04142_ ) );
OAI22_X1 _12026_ ( .A1(_04141_ ), .A2(_02993_ ), .B1(_04142_ ), .B2(_04108_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ) );
XNOR2_X1 _12027_ ( .A(_02317_ ), .B(_02321_ ), .ZN(_04143_ ) );
NAND2_X1 _12028_ ( .A1(_04143_ ), .A2(_03007_ ), .ZN(_04144_ ) );
INV_X1 _12029_ ( .A(\ID_EX_csr [4] ), .ZN(_04145_ ) );
OAI21_X1 _12030_ ( .A(_04144_ ), .B1(_04145_ ), .B2(_04108_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ) );
AOI21_X1 _12031_ ( .A(_02261_ ), .B1(_02310_ ), .B2(_02284_ ), .ZN(_04146_ ) );
OR2_X1 _12032_ ( .A1(_04146_ ), .A2(_02312_ ), .ZN(_04147_ ) );
XNOR2_X1 _12033_ ( .A(_04147_ ), .B(_02237_ ), .ZN(_04148_ ) );
NAND2_X1 _12034_ ( .A1(_04148_ ), .A2(_03007_ ), .ZN(_04149_ ) );
INV_X1 _12035_ ( .A(\ID_EX_csr [3] ), .ZN(_04150_ ) );
OAI21_X1 _12036_ ( .A(_04149_ ), .B1(_04150_ ), .B2(_04108_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ) );
AND3_X1 _12037_ ( .A1(_02310_ ), .A2(_02284_ ), .A3(_02261_ ), .ZN(_04151_ ) );
NOR3_X1 _12038_ ( .A1(_04151_ ), .A2(_04146_ ), .A3(_04131_ ), .ZN(_04152_ ) );
MUX2_X1 _12039_ ( .A(\ID_EX_csr [2] ), .B(_04152_ ), .S(_04135_ ), .Z(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ) );
NOR2_X1 _12040_ ( .A1(_04115_ ), .A2(_02423_ ), .ZN(_04153_ ) );
AND2_X1 _12041_ ( .A1(_02422_ ), .A2(\ID_EX_imm [10] ), .ZN(_04154_ ) );
OR2_X1 _12042_ ( .A1(_04153_ ), .A2(_04154_ ), .ZN(_04155_ ) );
XNOR2_X1 _12043_ ( .A(_04155_ ), .B(_02400_ ), .ZN(_04156_ ) );
NAND2_X1 _12044_ ( .A1(_04156_ ), .A2(_03007_ ), .ZN(_04157_ ) );
INV_X1 _12045_ ( .A(\ID_EX_csr [11] ), .ZN(_04158_ ) );
OAI21_X1 _12046_ ( .A(_04157_ ), .B1(_04158_ ), .B2(_04108_ ), .ZN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ) );
AND2_X1 _12047_ ( .A1(_01735_ ), .A2(\ID_EX_rd [3] ), .ZN(\myexu.dest_reg_$_DFFE_PP0P__Q_1_D ) );
AND2_X1 _12048_ ( .A1(_01735_ ), .A2(\ID_EX_rd [2] ), .ZN(\myexu.dest_reg_$_DFFE_PP0P__Q_2_D ) );
AND2_X1 _12049_ ( .A1(_01735_ ), .A2(\ID_EX_rd [1] ), .ZN(\myexu.dest_reg_$_DFFE_PP0P__Q_3_D ) );
AND2_X1 _12050_ ( .A1(_01735_ ), .A2(\ID_EX_rd [0] ), .ZN(\myexu.dest_reg_$_DFFE_PP0P__Q_4_D ) );
AND2_X1 _12051_ ( .A1(_01735_ ), .A2(\ID_EX_rd [4] ), .ZN(\myexu.dest_reg_$_DFFE_PP0P__Q_D ) );
INV_X2 _12052_ ( .A(fanout_net_10 ), .ZN(_04159_ ) );
BUF_X4 _12053_ ( .A(_04159_ ), .Z(_04160_ ) );
AOI22_X1 _12054_ ( .A1(\EX_LS_dest_csreg_mem [9] ), .A2(_04122_ ), .B1(_04125_ ), .B2(\EX_LS_dest_csreg_mem [8] ), .ZN(_04161_ ) );
AOI22_X1 _12055_ ( .A1(_03843_ ), .A2(\ID_EX_csr [9] ), .B1(_03847_ ), .B2(\ID_EX_csr [8] ), .ZN(_04162_ ) );
XNOR2_X1 _12056_ ( .A(\EX_LS_dest_csreg_mem [11] ), .B(\ID_EX_csr [11] ), .ZN(_04163_ ) );
AND4_X1 _12057_ ( .A1(_03823_ ), .A2(_04161_ ), .A3(_04162_ ), .A4(_04163_ ), .ZN(_04164_ ) );
XNOR2_X1 _12058_ ( .A(\EX_LS_dest_csreg_mem [4] ), .B(\ID_EX_csr [4] ), .ZN(_04165_ ) );
XNOR2_X1 _12059_ ( .A(\EX_LS_dest_csreg_mem [1] ), .B(\ID_EX_csr [1] ), .ZN(_04166_ ) );
XNOR2_X1 _12060_ ( .A(\EX_LS_dest_csreg_mem [5] ), .B(\ID_EX_csr [5] ), .ZN(_04167_ ) );
XNOR2_X1 _12061_ ( .A(\EX_LS_dest_csreg_mem [0] ), .B(\ID_EX_csr [0] ), .ZN(_04168_ ) );
AND4_X1 _12062_ ( .A1(_04165_ ), .A2(_04166_ ), .A3(_04167_ ), .A4(_04168_ ), .ZN(_04169_ ) );
NAND2_X1 _12063_ ( .A1(_04164_ ), .A2(_04169_ ), .ZN(_04170_ ) );
BUF_X2 _12064_ ( .A(_04170_ ), .Z(_04171_ ) );
BUF_X2 _12065_ ( .A(_04171_ ), .Z(_04172_ ) );
XNOR2_X1 _12066_ ( .A(\EX_LS_dest_csreg_mem [10] ), .B(\ID_EX_csr [10] ), .ZN(_04173_ ) );
XNOR2_X1 _12067_ ( .A(\EX_LS_dest_csreg_mem [7] ), .B(\ID_EX_csr [7] ), .ZN(_04174_ ) );
XNOR2_X1 _12068_ ( .A(\EX_LS_dest_csreg_mem [6] ), .B(\ID_EX_csr [6] ), .ZN(_04175_ ) );
AND3_X1 _12069_ ( .A1(_04173_ ), .A2(_04174_ ), .A3(_04175_ ), .ZN(_04176_ ) );
XNOR2_X1 _12070_ ( .A(\EX_LS_dest_csreg_mem [3] ), .B(\ID_EX_csr [3] ), .ZN(_04177_ ) );
XNOR2_X1 _12071_ ( .A(\EX_LS_dest_csreg_mem [2] ), .B(\ID_EX_csr [2] ), .ZN(_04178_ ) );
NAND3_X1 _12072_ ( .A1(_04176_ ), .A2(_04177_ ), .A3(_04178_ ), .ZN(_04179_ ) );
BUF_X2 _12073_ ( .A(_04179_ ), .Z(_04180_ ) );
BUF_X2 _12074_ ( .A(_04180_ ), .Z(_04181_ ) );
NOR3_X1 _12075_ ( .A1(_04172_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_04181_ ), .ZN(_04182_ ) );
AND2_X1 _12076_ ( .A1(\ID_EX_csr [9] ), .A2(\ID_EX_csr [8] ), .ZN(_04183_ ) );
NAND3_X1 _12077_ ( .A1(_04183_ ), .A2(\ID_EX_csr [10] ), .A3(\ID_EX_csr [11] ), .ZN(_04184_ ) );
NOR2_X1 _12078_ ( .A1(\ID_EX_csr [7] ), .A2(\ID_EX_csr [6] ), .ZN(_04185_ ) );
NAND3_X1 _12079_ ( .A1(_04185_ ), .A2(_04142_ ), .A3(\ID_EX_csr [4] ), .ZN(_04186_ ) );
NOR2_X1 _12080_ ( .A1(_04184_ ), .A2(_04186_ ), .ZN(_04187_ ) );
NOR2_X1 _12081_ ( .A1(_04112_ ), .A2(\ID_EX_csr [1] ), .ZN(_04188_ ) );
NOR2_X1 _12082_ ( .A1(\ID_EX_csr [3] ), .A2(\ID_EX_csr [2] ), .ZN(_04189_ ) );
AND2_X1 _12083_ ( .A1(_04188_ ), .A2(_04189_ ), .ZN(_04190_ ) );
BUF_X2 _12084_ ( .A(_04190_ ), .Z(_04191_ ) );
AND2_X1 _12085_ ( .A1(_04187_ ), .A2(_04191_ ), .ZN(_04192_ ) );
INV_X1 _12086_ ( .A(_04192_ ), .ZN(_04193_ ) );
NOR2_X1 _12087_ ( .A1(_04103_ ), .A2(\ID_EX_csr [0] ), .ZN(_04194_ ) );
AND2_X1 _12088_ ( .A1(_04194_ ), .A2(_04189_ ), .ZN(_04195_ ) );
BUF_X4 _12089_ ( .A(_04195_ ), .Z(_04196_ ) );
AND2_X1 _12090_ ( .A1(_04187_ ), .A2(_04196_ ), .ZN(_04197_ ) );
INV_X1 _12091_ ( .A(_04197_ ), .ZN(_04198_ ) );
NOR2_X1 _12092_ ( .A1(_04138_ ), .A2(\ID_EX_csr [7] ), .ZN(_04199_ ) );
BUF_X4 _12093_ ( .A(_04199_ ), .Z(_04200_ ) );
NOR2_X1 _12094_ ( .A1(\ID_EX_csr [5] ), .A2(\ID_EX_csr [4] ), .ZN(_04201_ ) );
AND4_X2 _12095_ ( .A1(_04189_ ), .A2(_04194_ ), .A3(_04200_ ), .A4(_04201_ ), .ZN(_04202_ ) );
BUF_X2 _12096_ ( .A(_04202_ ), .Z(_04203_ ) );
NAND3_X1 _12097_ ( .A1(_04158_ ), .A2(\ID_EX_csr [9] ), .A3(\ID_EX_csr [8] ), .ZN(_04204_ ) );
NOR2_X1 _12098_ ( .A1(_04204_ ), .A2(\ID_EX_csr [10] ), .ZN(_04205_ ) );
BUF_X2 _12099_ ( .A(_04205_ ), .Z(_04206_ ) );
BUF_X2 _12100_ ( .A(_04206_ ), .Z(_04207_ ) );
NAND3_X1 _12101_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][20] ), .A3(_04207_ ), .ZN(_04208_ ) );
NAND3_X1 _12102_ ( .A1(_04193_ ), .A2(_04198_ ), .A3(_04208_ ), .ZN(_04209_ ) );
NOR2_X1 _12103_ ( .A1(_04170_ ), .A2(_04179_ ), .ZN(_04210_ ) );
NOR2_X1 _12104_ ( .A1(_04209_ ), .A2(_04210_ ), .ZN(_04211_ ) );
AND3_X2 _12105_ ( .A1(_04205_ ), .A2(_04185_ ), .A3(_04201_ ), .ZN(_04212_ ) );
BUF_X4 _12106_ ( .A(_04212_ ), .Z(_04213_ ) );
BUF_X2 _12107_ ( .A(_04213_ ), .Z(_04214_ ) );
AND3_X1 _12108_ ( .A1(_04188_ ), .A2(_04150_ ), .A3(\ID_EX_csr [2] ), .ZN(_04215_ ) );
BUF_X4 _12109_ ( .A(_04215_ ), .Z(_04216_ ) );
BUF_X4 _12110_ ( .A(_04216_ ), .Z(_04217_ ) );
BUF_X4 _12111_ ( .A(_04217_ ), .Z(_04218_ ) );
NAND3_X1 _12112_ ( .A1(_04214_ ), .A2(\mtvec [20] ), .A3(_04218_ ), .ZN(_04219_ ) );
AND3_X1 _12113_ ( .A1(_04189_ ), .A2(_04103_ ), .A3(_04112_ ), .ZN(_04220_ ) );
BUF_X4 _12114_ ( .A(_04220_ ), .Z(_04221_ ) );
BUF_X4 _12115_ ( .A(_04221_ ), .Z(_04222_ ) );
BUF_X2 _12116_ ( .A(_04222_ ), .Z(_04223_ ) );
NAND3_X1 _12117_ ( .A1(_04214_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_04223_ ), .ZN(_04224_ ) );
AND4_X1 _12118_ ( .A1(_04188_ ), .A2(_04199_ ), .A3(_04189_ ), .A4(_04201_ ), .ZN(_04225_ ) );
BUF_X2 _12119_ ( .A(_04225_ ), .Z(_04226_ ) );
NAND3_X1 _12120_ ( .A1(_04226_ ), .A2(\mepc [20] ), .A3(_04207_ ), .ZN(_04227_ ) );
AND3_X1 _12121_ ( .A1(_04219_ ), .A2(_04224_ ), .A3(_04227_ ), .ZN(_04228_ ) );
AOI211_X1 _12122_ ( .A(_04160_ ), .B(_04182_ ), .C1(_04211_ ), .C2(_04228_ ), .ZN(_04229_ ) );
AND3_X1 _12123_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_pc [3] ), .A3(\ID_EX_pc [2] ), .ZN(_04230_ ) );
AND2_X1 _12124_ ( .A1(_04230_ ), .A2(\ID_EX_pc [5] ), .ZN(_04231_ ) );
AND3_X1 _12125_ ( .A1(_04231_ ), .A2(\ID_EX_pc [7] ), .A3(\ID_EX_pc [6] ), .ZN(_04232_ ) );
AND2_X1 _12126_ ( .A1(_04232_ ), .A2(\ID_EX_pc [8] ), .ZN(_04233_ ) );
AND2_X2 _12127_ ( .A1(_04233_ ), .A2(\ID_EX_pc [9] ), .ZN(_04234_ ) );
AND2_X1 _12128_ ( .A1(\ID_EX_pc [19] ), .A2(\ID_EX_pc [18] ), .ZN(_04235_ ) );
AND2_X1 _12129_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_pc [10] ), .ZN(_04236_ ) );
AND3_X1 _12130_ ( .A1(_04236_ ), .A2(\ID_EX_pc [13] ), .A3(\ID_EX_pc [12] ), .ZN(_04237_ ) );
AND2_X1 _12131_ ( .A1(\ID_EX_pc [15] ), .A2(\ID_EX_pc [14] ), .ZN(_04238_ ) );
AND4_X1 _12132_ ( .A1(\ID_EX_pc [17] ), .A2(_04237_ ), .A3(\ID_EX_pc [16] ), .A4(_04238_ ), .ZN(_04239_ ) );
AND3_X1 _12133_ ( .A1(_04234_ ), .A2(_04235_ ), .A3(_04239_ ), .ZN(_04240_ ) );
XNOR2_X1 _12134_ ( .A(_04240_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_04241_ ) );
XOR2_X1 _12135_ ( .A(\ID_EX_pc [8] ), .B(\ID_EX_imm [8] ), .Z(_04242_ ) );
AND2_X1 _12136_ ( .A1(\ID_EX_pc [9] ), .A2(\ID_EX_imm [9] ), .ZN(_04243_ ) );
NOR2_X1 _12137_ ( .A1(\ID_EX_pc [9] ), .A2(\ID_EX_imm [9] ), .ZN(_04244_ ) );
NOR2_X1 _12138_ ( .A1(_04243_ ), .A2(_04244_ ), .ZN(_04245_ ) );
AND2_X1 _12139_ ( .A1(_04242_ ), .A2(_04245_ ), .ZN(_04246_ ) );
XOR2_X1 _12140_ ( .A(\ID_EX_pc [10] ), .B(\ID_EX_imm [10] ), .Z(_04247_ ) );
AND2_X1 _12141_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_imm [11] ), .ZN(_04248_ ) );
NOR2_X1 _12142_ ( .A1(\ID_EX_pc [11] ), .A2(\ID_EX_imm [11] ), .ZN(_04249_ ) );
NOR2_X1 _12143_ ( .A1(_04248_ ), .A2(_04249_ ), .ZN(_04250_ ) );
AND3_X1 _12144_ ( .A1(_04246_ ), .A2(_04247_ ), .A3(_04250_ ), .ZN(_04251_ ) );
XOR2_X1 _12145_ ( .A(\ID_EX_pc [15] ), .B(\ID_EX_imm [15] ), .Z(_04252_ ) );
XOR2_X1 _12146_ ( .A(\ID_EX_pc [14] ), .B(\ID_EX_imm [14] ), .Z(_04253_ ) );
AND2_X1 _12147_ ( .A1(_04252_ ), .A2(_04253_ ), .ZN(_04254_ ) );
XOR2_X1 _12148_ ( .A(\ID_EX_pc [12] ), .B(\ID_EX_imm [12] ), .Z(_04255_ ) );
XOR2_X1 _12149_ ( .A(\ID_EX_pc [13] ), .B(\ID_EX_imm [13] ), .Z(_04256_ ) );
AND2_X1 _12150_ ( .A1(_04255_ ), .A2(_04256_ ), .ZN(_04257_ ) );
AND2_X1 _12151_ ( .A1(_04254_ ), .A2(_04257_ ), .ZN(_04258_ ) );
NOR2_X1 _12152_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04259_ ) );
AND2_X1 _12153_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_04260_ ) );
INV_X1 _12154_ ( .A(_04260_ ), .ZN(_04261_ ) );
XOR2_X1 _12155_ ( .A(\ID_EX_pc [1] ), .B(\ID_EX_imm [1] ), .Z(_04262_ ) );
AND2_X1 _12156_ ( .A1(\ID_EX_pc [0] ), .A2(\ID_EX_imm [0] ), .ZN(_04263_ ) );
NAND2_X1 _12157_ ( .A1(_04262_ ), .A2(_04263_ ), .ZN(_04264_ ) );
INV_X1 _12158_ ( .A(\ID_EX_pc [1] ), .ZN(_04265_ ) );
OAI21_X1 _12159_ ( .A(_04264_ ), .B1(_04265_ ), .B2(_02285_ ), .ZN(_04266_ ) );
XOR2_X1 _12160_ ( .A(\ID_EX_pc [2] ), .B(\ID_EX_imm [2] ), .Z(_04267_ ) );
NAND2_X1 _12161_ ( .A1(_04266_ ), .A2(_04267_ ), .ZN(_04268_ ) );
NAND2_X1 _12162_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_04269_ ) );
NAND2_X1 _12163_ ( .A1(\ID_EX_pc [2] ), .A2(\ID_EX_imm [2] ), .ZN(_04270_ ) );
NAND3_X1 _12164_ ( .A1(_04268_ ), .A2(_04269_ ), .A3(_04270_ ), .ZN(_04271_ ) );
OR2_X1 _12165_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_imm [3] ), .ZN(_04272_ ) );
XOR2_X1 _12166_ ( .A(\ID_EX_pc [4] ), .B(\ID_EX_imm [4] ), .Z(_04273_ ) );
AND3_X1 _12167_ ( .A1(_04271_ ), .A2(_04272_ ), .A3(_04273_ ), .ZN(_04274_ ) );
AND2_X1 _12168_ ( .A1(\ID_EX_pc [4] ), .A2(\ID_EX_imm [4] ), .ZN(_04275_ ) );
NOR2_X1 _12169_ ( .A1(_04274_ ), .A2(_04275_ ), .ZN(_04276_ ) );
NOR2_X1 _12170_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_imm [5] ), .ZN(_04277_ ) );
OAI21_X1 _12171_ ( .A(_04261_ ), .B1(_04276_ ), .B2(_04277_ ), .ZN(_04278_ ) );
XOR2_X1 _12172_ ( .A(\ID_EX_pc [6] ), .B(\ID_EX_imm [6] ), .Z(_04279_ ) );
NAND2_X1 _12173_ ( .A1(_04278_ ), .A2(_04279_ ), .ZN(_04280_ ) );
NAND2_X1 _12174_ ( .A1(\ID_EX_pc [6] ), .A2(\ID_EX_imm [6] ), .ZN(_04281_ ) );
AOI21_X1 _12175_ ( .A(_04259_ ), .B1(_04280_ ), .B2(_04281_ ), .ZN(_04282_ ) );
AND2_X1 _12176_ ( .A1(\ID_EX_pc [7] ), .A2(\ID_EX_imm [7] ), .ZN(_04283_ ) );
OAI211_X1 _12177_ ( .A(_04251_ ), .B(_04258_ ), .C1(_04282_ ), .C2(_04283_ ), .ZN(_04284_ ) );
AND2_X1 _12178_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_04285_ ) );
NAND2_X1 _12179_ ( .A1(_04252_ ), .A2(_04285_ ), .ZN(_04286_ ) );
INV_X1 _12180_ ( .A(\ID_EX_pc [15] ), .ZN(_04287_ ) );
OAI21_X1 _12181_ ( .A(_04286_ ), .B1(_04287_ ), .B2(_02586_ ), .ZN(_04288_ ) );
AND2_X1 _12182_ ( .A1(\ID_EX_pc [12] ), .A2(\ID_EX_imm [12] ), .ZN(_04289_ ) );
AND2_X1 _12183_ ( .A1(_04256_ ), .A2(_04289_ ), .ZN(_04290_ ) );
AOI21_X1 _12184_ ( .A(_04290_ ), .B1(\ID_EX_pc [13] ), .B2(\ID_EX_imm [13] ), .ZN(_04291_ ) );
INV_X1 _12185_ ( .A(_04291_ ), .ZN(_04292_ ) );
INV_X1 _12186_ ( .A(_04247_ ), .ZN(_04293_ ) );
INV_X1 _12187_ ( .A(_04244_ ), .ZN(_04294_ ) );
AND2_X1 _12188_ ( .A1(\ID_EX_pc [8] ), .A2(\ID_EX_imm [8] ), .ZN(_04295_ ) );
AOI21_X1 _12189_ ( .A(_04243_ ), .B1(_04294_ ), .B2(_04295_ ), .ZN(_04296_ ) );
NOR4_X1 _12190_ ( .A1(_04293_ ), .A2(_04296_ ), .A3(_04248_ ), .A4(_04249_ ), .ZN(_04297_ ) );
AND2_X1 _12191_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_imm [10] ), .ZN(_04298_ ) );
AND2_X1 _12192_ ( .A1(_04250_ ), .A2(_04298_ ), .ZN(_04299_ ) );
OR3_X1 _12193_ ( .A1(_04297_ ), .A2(_04248_ ), .A3(_04299_ ), .ZN(_04300_ ) );
AOI221_X4 _12194_ ( .A(_04288_ ), .B1(_04254_ ), .B2(_04292_ ), .C1(_04300_ ), .C2(_04258_ ), .ZN(_04301_ ) );
NAND2_X1 _12195_ ( .A1(_04284_ ), .A2(_04301_ ), .ZN(_04302_ ) );
XOR2_X1 _12196_ ( .A(\ID_EX_pc [19] ), .B(\ID_EX_imm [19] ), .Z(_04303_ ) );
XOR2_X1 _12197_ ( .A(\ID_EX_pc [18] ), .B(\ID_EX_imm [18] ), .Z(_04304_ ) );
XOR2_X1 _12198_ ( .A(\ID_EX_pc [16] ), .B(\ID_EX_imm [16] ), .Z(_04305_ ) );
AND2_X1 _12199_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_imm [17] ), .ZN(_04306_ ) );
NOR2_X1 _12200_ ( .A1(\ID_EX_pc [17] ), .A2(\ID_EX_imm [17] ), .ZN(_04307_ ) );
NOR2_X1 _12201_ ( .A1(_04306_ ), .A2(_04307_ ), .ZN(_04308_ ) );
AND2_X1 _12202_ ( .A1(_04305_ ), .A2(_04308_ ), .ZN(_04309_ ) );
NAND4_X1 _12203_ ( .A1(_04302_ ), .A2(_04303_ ), .A3(_04304_ ), .A4(_04309_ ), .ZN(_04310_ ) );
AND2_X1 _12204_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_04311_ ) );
AND2_X1 _12205_ ( .A1(_04303_ ), .A2(_04311_ ), .ZN(_04312_ ) );
AOI21_X1 _12206_ ( .A(_04312_ ), .B1(\ID_EX_pc [19] ), .B2(\ID_EX_imm [19] ), .ZN(_04313_ ) );
AND2_X1 _12207_ ( .A1(\ID_EX_pc [16] ), .A2(\ID_EX_imm [16] ), .ZN(_04314_ ) );
AND2_X1 _12208_ ( .A1(_04308_ ), .A2(_04314_ ), .ZN(_04315_ ) );
OAI211_X1 _12209_ ( .A(_04303_ ), .B(_04304_ ), .C1(_04315_ ), .C2(_04306_ ), .ZN(_04316_ ) );
AND2_X1 _12210_ ( .A1(_04313_ ), .A2(_04316_ ), .ZN(_04317_ ) );
NAND2_X1 _12211_ ( .A1(_04310_ ), .A2(_04317_ ), .ZN(_04318_ ) );
XOR2_X1 _12212_ ( .A(\ID_EX_pc [20] ), .B(\ID_EX_imm [20] ), .Z(_04319_ ) );
INV_X1 _12213_ ( .A(_04319_ ), .ZN(_04320_ ) );
XNOR2_X1 _12214_ ( .A(_04318_ ), .B(_04320_ ), .ZN(_04321_ ) );
NOR2_X1 _12215_ ( .A1(fanout_net_8 ), .A2(\ID_EX_typ [1] ), .ZN(_04322_ ) );
AND2_X1 _12216_ ( .A1(_04322_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_04323_ ) );
INV_X1 _12217_ ( .A(_04323_ ), .ZN(_04324_ ) );
XOR2_X1 _12218_ ( .A(\EX_LS_dest_reg [0] ), .B(\ID_EX_rs2 [0] ), .Z(_04325_ ) );
AND2_X1 _12219_ ( .A1(_02130_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_04326_ ) );
OR4_X4 _12220_ ( .A1(_02154_ ), .A2(_02133_ ), .A3(_04325_ ), .A4(_04326_ ), .ZN(_04327_ ) );
BUF_X8 _12221_ ( .A(_04327_ ), .Z(_04328_ ) );
BUF_X4 _12222_ ( .A(_04328_ ), .Z(_04329_ ) );
BUF_X2 _12223_ ( .A(_04329_ ), .Z(_04330_ ) );
XNOR2_X1 _12224_ ( .A(\EX_LS_dest_reg [4] ), .B(\ID_EX_rs2 [4] ), .ZN(_04331_ ) );
NAND2_X1 _12225_ ( .A1(_03323_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_04332_ ) );
AND3_X4 _12226_ ( .A1(_04331_ ), .A2(\myidu.fc_disenable_$_NOT__A_Y ), .A3(_04332_ ), .ZN(_04333_ ) );
OR2_X1 _12227_ ( .A1(_03323_ ), .A2(\EX_LS_dest_reg [3] ), .ZN(_04334_ ) );
OR2_X1 _12228_ ( .A1(_02130_ ), .A2(\ID_EX_rs2 [1] ), .ZN(_04335_ ) );
XNOR2_X1 _12229_ ( .A(\EX_LS_dest_reg [2] ), .B(\ID_EX_rs2 [2] ), .ZN(_04336_ ) );
NAND4_X4 _12230_ ( .A1(_04333_ ), .A2(_04334_ ), .A3(_04335_ ), .A4(_04336_ ), .ZN(_04337_ ) );
CLKBUF_X2 _12231_ ( .A(_04337_ ), .Z(_04338_ ) );
CLKBUF_X2 _12232_ ( .A(_04338_ ), .Z(_04339_ ) );
BUF_X2 _12233_ ( .A(_04339_ ), .Z(_04340_ ) );
OR3_X1 _12234_ ( .A1(_04330_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04340_ ), .ZN(_04341_ ) );
INV_X1 _12235_ ( .A(fanout_net_47 ), .ZN(_04342_ ) );
BUF_X4 _12236_ ( .A(_04342_ ), .Z(_04343_ ) );
BUF_X4 _12237_ ( .A(_04343_ ), .Z(_04344_ ) );
INV_X2 _12238_ ( .A(fanout_net_35 ), .ZN(_04345_ ) );
BUF_X4 _12239_ ( .A(_04345_ ), .Z(_04346_ ) );
BUF_X4 _12240_ ( .A(_04346_ ), .Z(_04347_ ) );
BUF_X4 _12241_ ( .A(_04347_ ), .Z(_04348_ ) );
BUF_X4 _12242_ ( .A(_04348_ ), .Z(_04349_ ) );
OR2_X1 _12243_ ( .A1(_04349_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04350_ ) );
OAI211_X1 _12244_ ( .A(_04350_ ), .B(fanout_net_43 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04351_ ) );
INV_X1 _12245_ ( .A(fanout_net_46 ), .ZN(_04352_ ) );
BUF_X4 _12246_ ( .A(_04352_ ), .Z(_04353_ ) );
BUF_X4 _12247_ ( .A(_04353_ ), .Z(_04354_ ) );
BUF_X4 _12248_ ( .A(_04354_ ), .Z(_04355_ ) );
BUF_X4 _12249_ ( .A(_04355_ ), .Z(_04356_ ) );
OR2_X1 _12250_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04357_ ) );
INV_X1 _12251_ ( .A(fanout_net_43 ), .ZN(_04358_ ) );
BUF_X4 _12252_ ( .A(_04358_ ), .Z(_04359_ ) );
BUF_X4 _12253_ ( .A(_04359_ ), .Z(_04360_ ) );
BUF_X4 _12254_ ( .A(_04360_ ), .Z(_04361_ ) );
BUF_X4 _12255_ ( .A(_04361_ ), .Z(_04362_ ) );
BUF_X4 _12256_ ( .A(_04362_ ), .Z(_04363_ ) );
BUF_X4 _12257_ ( .A(_04349_ ), .Z(_04364_ ) );
OAI211_X1 _12258_ ( .A(_04357_ ), .B(_04363_ ), .C1(_04364_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04365_ ) );
NAND3_X1 _12259_ ( .A1(_04351_ ), .A2(_04356_ ), .A3(_04365_ ), .ZN(_04366_ ) );
MUX2_X1 _12260_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04367_ ) );
MUX2_X1 _12261_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04368_ ) );
MUX2_X1 _12262_ ( .A(_04367_ ), .B(_04368_ ), .S(_04363_ ), .Z(_04369_ ) );
BUF_X4 _12263_ ( .A(_04356_ ), .Z(_04370_ ) );
OAI211_X1 _12264_ ( .A(_04344_ ), .B(_04366_ ), .C1(_04369_ ), .C2(_04370_ ), .ZN(_04371_ ) );
OR2_X1 _12265_ ( .A1(_04349_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04372_ ) );
OAI211_X1 _12266_ ( .A(_04372_ ), .B(_04363_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04373_ ) );
OR2_X1 _12267_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04374_ ) );
OAI211_X1 _12268_ ( .A(_04374_ ), .B(fanout_net_43 ), .C1(_04349_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04375_ ) );
NAND3_X1 _12269_ ( .A1(_04373_ ), .A2(fanout_net_46 ), .A3(_04375_ ), .ZN(_04376_ ) );
MUX2_X1 _12270_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04377_ ) );
MUX2_X1 _12271_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04378_ ) );
MUX2_X1 _12272_ ( .A(_04377_ ), .B(_04378_ ), .S(fanout_net_43 ), .Z(_04379_ ) );
OAI211_X1 _12273_ ( .A(fanout_net_47 ), .B(_04376_ ), .C1(_04379_ ), .C2(fanout_net_46 ), .ZN(_04380_ ) );
BUF_X2 _12274_ ( .A(_04330_ ), .Z(_04381_ ) );
BUF_X2 _12275_ ( .A(_04340_ ), .Z(_04382_ ) );
OAI211_X1 _12276_ ( .A(_04371_ ), .B(_04380_ ), .C1(_04381_ ), .C2(_04382_ ), .ZN(_04383_ ) );
NAND2_X1 _12277_ ( .A1(_04341_ ), .A2(_04383_ ), .ZN(_04384_ ) );
XNOR2_X1 _12278_ ( .A(_02909_ ), .B(_04384_ ), .ZN(_04385_ ) );
OR3_X1 _12279_ ( .A1(_04381_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04382_ ), .ZN(_04386_ ) );
OR2_X1 _12280_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04387_ ) );
BUF_X4 _12281_ ( .A(_04363_ ), .Z(_04388_ ) );
BUF_X4 _12282_ ( .A(_04364_ ), .Z(_04389_ ) );
OAI211_X1 _12283_ ( .A(_04387_ ), .B(_04388_ ), .C1(_04389_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04390_ ) );
OR2_X1 _12284_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04391_ ) );
OAI211_X1 _12285_ ( .A(_04391_ ), .B(fanout_net_43 ), .C1(_04389_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04392_ ) );
NAND3_X1 _12286_ ( .A1(_04390_ ), .A2(_04392_ ), .A3(_04370_ ), .ZN(_04393_ ) );
MUX2_X1 _12287_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04394_ ) );
MUX2_X1 _12288_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04395_ ) );
MUX2_X1 _12289_ ( .A(_04394_ ), .B(_04395_ ), .S(_04388_ ), .Z(_04396_ ) );
OAI211_X1 _12290_ ( .A(_04344_ ), .B(_04393_ ), .C1(_04396_ ), .C2(_04370_ ), .ZN(_04397_ ) );
OR2_X1 _12291_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04398_ ) );
OAI211_X1 _12292_ ( .A(_04398_ ), .B(fanout_net_43 ), .C1(_04389_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04399_ ) );
NAND2_X1 _12293_ ( .A1(_02922_ ), .A2(fanout_net_35 ), .ZN(_04400_ ) );
OAI211_X1 _12294_ ( .A(_04400_ ), .B(_04388_ ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04401_ ) );
NAND3_X1 _12295_ ( .A1(_04399_ ), .A2(_04401_ ), .A3(fanout_net_46 ), .ZN(_04402_ ) );
MUX2_X1 _12296_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04403_ ) );
MUX2_X1 _12297_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04404_ ) );
MUX2_X1 _12298_ ( .A(_04403_ ), .B(_04404_ ), .S(fanout_net_43 ), .Z(_04405_ ) );
OAI211_X1 _12299_ ( .A(fanout_net_47 ), .B(_04402_ ), .C1(_04405_ ), .C2(fanout_net_46 ), .ZN(_04406_ ) );
OAI211_X1 _12300_ ( .A(_04397_ ), .B(_04406_ ), .C1(_04381_ ), .C2(_04382_ ), .ZN(_04407_ ) );
NAND2_X1 _12301_ ( .A1(_04386_ ), .A2(_04407_ ), .ZN(_04408_ ) );
XNOR2_X1 _12302_ ( .A(_02933_ ), .B(_04408_ ), .ZN(_04409_ ) );
AND2_X1 _12303_ ( .A1(_04385_ ), .A2(_04409_ ), .ZN(_04410_ ) );
NOR2_X1 _12304_ ( .A1(_04327_ ), .A2(_04337_ ), .ZN(_04411_ ) );
OR2_X1 _12305_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04412_ ) );
OAI211_X1 _12306_ ( .A(_04412_ ), .B(_04388_ ), .C1(_04389_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04413_ ) );
NAND2_X1 _12307_ ( .A1(_02969_ ), .A2(fanout_net_35 ), .ZN(_04414_ ) );
OAI211_X1 _12308_ ( .A(_04414_ ), .B(fanout_net_43 ), .C1(fanout_net_35 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04415_ ) );
NAND3_X1 _12309_ ( .A1(_04413_ ), .A2(_04415_ ), .A3(_04370_ ), .ZN(_04416_ ) );
MUX2_X1 _12310_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04417_ ) );
MUX2_X1 _12311_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04418_ ) );
MUX2_X1 _12312_ ( .A(_04417_ ), .B(_04418_ ), .S(_04388_ ), .Z(_04419_ ) );
OAI211_X1 _12313_ ( .A(_04344_ ), .B(_04416_ ), .C1(_04419_ ), .C2(_04370_ ), .ZN(_04420_ ) );
OR2_X1 _12314_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04421_ ) );
OAI211_X1 _12315_ ( .A(_04421_ ), .B(fanout_net_43 ), .C1(_04389_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04422_ ) );
OR2_X1 _12316_ ( .A1(fanout_net_35 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04423_ ) );
OAI211_X1 _12317_ ( .A(_04423_ ), .B(_04388_ ), .C1(_04389_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04424_ ) );
NAND3_X1 _12318_ ( .A1(_04422_ ), .A2(_04424_ ), .A3(fanout_net_46 ), .ZN(_04425_ ) );
MUX2_X1 _12319_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04426_ ) );
MUX2_X1 _12320_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04427_ ) );
MUX2_X1 _12321_ ( .A(_04426_ ), .B(_04427_ ), .S(fanout_net_43 ), .Z(_04428_ ) );
OAI211_X1 _12322_ ( .A(fanout_net_47 ), .B(_04425_ ), .C1(_04428_ ), .C2(fanout_net_46 ), .ZN(_04429_ ) );
AOI21_X1 _12323_ ( .A(_04411_ ), .B1(_04420_ ), .B2(_04429_ ), .ZN(_04430_ ) );
AND2_X1 _12324_ ( .A1(_04411_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04431_ ) );
NOR2_X1 _12325_ ( .A1(_04430_ ), .A2(_04431_ ), .ZN(_04432_ ) );
XNOR2_X1 _12326_ ( .A(_04432_ ), .B(_02987_ ), .ZN(_04433_ ) );
OR3_X1 _12327_ ( .A1(_04381_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_B ), .A3(_04382_ ), .ZN(_04434_ ) );
OR2_X1 _12328_ ( .A1(_04364_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04435_ ) );
OAI211_X1 _12329_ ( .A(_04435_ ), .B(fanout_net_43 ), .C1(fanout_net_35 ), .C2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04436_ ) );
OR2_X1 _12330_ ( .A1(fanout_net_35 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04437_ ) );
OAI211_X1 _12331_ ( .A(_04437_ ), .B(_04388_ ), .C1(_04389_ ), .C2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04438_ ) );
NAND3_X1 _12332_ ( .A1(_04436_ ), .A2(fanout_net_46 ), .A3(_04438_ ), .ZN(_04439_ ) );
MUX2_X1 _12333_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_35 ), .Z(_04440_ ) );
MUX2_X1 _12334_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04441_ ) );
MUX2_X1 _12335_ ( .A(_04440_ ), .B(_04441_ ), .S(_04388_ ), .Z(_04442_ ) );
OAI211_X1 _12336_ ( .A(_04344_ ), .B(_04439_ ), .C1(_04442_ ), .C2(fanout_net_46 ), .ZN(_04443_ ) );
NOR2_X1 _12337_ ( .A1(_04389_ ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04444_ ) );
OAI21_X1 _12338_ ( .A(fanout_net_43 ), .B1(fanout_net_36 ), .B2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04445_ ) );
NOR2_X1 _12339_ ( .A1(fanout_net_36 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04446_ ) );
OAI21_X1 _12340_ ( .A(_04388_ ), .B1(_04389_ ), .B2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04447_ ) );
OAI221_X1 _12341_ ( .A(_04370_ ), .B1(_04444_ ), .B2(_04445_ ), .C1(_04446_ ), .C2(_04447_ ), .ZN(_04448_ ) );
MUX2_X1 _12342_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04449_ ) );
MUX2_X1 _12343_ ( .A(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04450_ ) );
MUX2_X1 _12344_ ( .A(_04449_ ), .B(_04450_ ), .S(fanout_net_43 ), .Z(_04451_ ) );
OAI211_X1 _12345_ ( .A(fanout_net_47 ), .B(_04448_ ), .C1(_04451_ ), .C2(_04370_ ), .ZN(_04452_ ) );
OAI211_X1 _12346_ ( .A(_04443_ ), .B(_04452_ ), .C1(_04381_ ), .C2(_04382_ ), .ZN(_04453_ ) );
NAND2_X1 _12347_ ( .A1(_04434_ ), .A2(_04453_ ), .ZN(_04454_ ) );
XOR2_X1 _12348_ ( .A(_02961_ ), .B(_04454_ ), .Z(_04455_ ) );
AND3_X1 _12349_ ( .A1(_04410_ ), .A2(_04433_ ), .A3(_04455_ ), .ZN(_04456_ ) );
INV_X1 _12350_ ( .A(\EX_LS_result_reg [27] ), .ZN(_04457_ ) );
OR3_X1 _12351_ ( .A1(_04381_ ), .A2(_04457_ ), .A3(_04382_ ), .ZN(_04458_ ) );
OR2_X1 _12352_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04459_ ) );
OAI211_X1 _12353_ ( .A(_04459_ ), .B(_04363_ ), .C1(_04364_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04460_ ) );
OR2_X1 _12354_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04461_ ) );
OAI211_X1 _12355_ ( .A(_04461_ ), .B(fanout_net_43 ), .C1(_04364_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04462_ ) );
NAND3_X1 _12356_ ( .A1(_04460_ ), .A2(_04462_ ), .A3(fanout_net_46 ), .ZN(_04463_ ) );
MUX2_X1 _12357_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04464_ ) );
MUX2_X1 _12358_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04465_ ) );
MUX2_X1 _12359_ ( .A(_04464_ ), .B(_04465_ ), .S(_04363_ ), .Z(_04466_ ) );
OAI211_X1 _12360_ ( .A(_04344_ ), .B(_04463_ ), .C1(_04466_ ), .C2(fanout_net_46 ), .ZN(_04467_ ) );
NOR2_X1 _12361_ ( .A1(_04364_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04468_ ) );
OAI21_X1 _12362_ ( .A(fanout_net_43 ), .B1(fanout_net_36 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04469_ ) );
NOR2_X1 _12363_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04470_ ) );
OAI21_X1 _12364_ ( .A(_04363_ ), .B1(_04364_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04471_ ) );
OAI221_X1 _12365_ ( .A(_04356_ ), .B1(_04468_ ), .B2(_04469_ ), .C1(_04470_ ), .C2(_04471_ ), .ZN(_04472_ ) );
MUX2_X1 _12366_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04473_ ) );
MUX2_X1 _12367_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04474_ ) );
MUX2_X1 _12368_ ( .A(_04473_ ), .B(_04474_ ), .S(fanout_net_43 ), .Z(_04475_ ) );
OAI211_X1 _12369_ ( .A(fanout_net_47 ), .B(_04472_ ), .C1(_04475_ ), .C2(_04370_ ), .ZN(_04476_ ) );
OAI211_X1 _12370_ ( .A(_04467_ ), .B(_04476_ ), .C1(_04381_ ), .C2(_04382_ ), .ZN(_04477_ ) );
NAND2_X1 _12371_ ( .A1(_04458_ ), .A2(_04477_ ), .ZN(_04478_ ) );
INV_X1 _12372_ ( .A(_04478_ ), .ZN(_04479_ ) );
XNOR2_X1 _12373_ ( .A(_02858_ ), .B(_04479_ ), .ZN(_04480_ ) );
OR3_X1 _12374_ ( .A1(_04330_ ), .A2(\EX_LS_result_reg [26] ), .A3(_04340_ ), .ZN(_04481_ ) );
BUF_X4 _12375_ ( .A(_04353_ ), .Z(_04482_ ) );
BUF_X4 _12376_ ( .A(_04482_ ), .Z(_04483_ ) );
BUF_X2 _12377_ ( .A(_04346_ ), .Z(_04484_ ) );
BUF_X4 _12378_ ( .A(_04484_ ), .Z(_04485_ ) );
NOR2_X1 _12379_ ( .A1(_04485_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04486_ ) );
OAI21_X1 _12380_ ( .A(fanout_net_43 ), .B1(fanout_net_36 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04487_ ) );
NOR2_X1 _12381_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04488_ ) );
BUF_X4 _12382_ ( .A(_04360_ ), .Z(_04489_ ) );
BUF_X4 _12383_ ( .A(_04489_ ), .Z(_04490_ ) );
OAI21_X1 _12384_ ( .A(_04490_ ), .B1(_04485_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04491_ ) );
OAI221_X1 _12385_ ( .A(_04483_ ), .B1(_04486_ ), .B2(_04487_ ), .C1(_04488_ ), .C2(_04491_ ), .ZN(_04492_ ) );
MUX2_X1 _12386_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04493_ ) );
MUX2_X1 _12387_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04494_ ) );
MUX2_X1 _12388_ ( .A(_04493_ ), .B(_04494_ ), .S(fanout_net_43 ), .Z(_04495_ ) );
OAI211_X1 _12389_ ( .A(fanout_net_47 ), .B(_04492_ ), .C1(_04495_ ), .C2(_04356_ ), .ZN(_04496_ ) );
OR2_X1 _12390_ ( .A1(_04348_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04497_ ) );
OAI211_X1 _12391_ ( .A(_04497_ ), .B(_04490_ ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04498_ ) );
OR2_X1 _12392_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04499_ ) );
OAI211_X1 _12393_ ( .A(_04499_ ), .B(fanout_net_43 ), .C1(_04349_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04500_ ) );
NAND3_X1 _12394_ ( .A1(_04498_ ), .A2(fanout_net_46 ), .A3(_04500_ ), .ZN(_04501_ ) );
MUX2_X1 _12395_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04502_ ) );
MUX2_X1 _12396_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04503_ ) );
MUX2_X1 _12397_ ( .A(_04502_ ), .B(_04503_ ), .S(_04490_ ), .Z(_04504_ ) );
OAI211_X1 _12398_ ( .A(_04344_ ), .B(_04501_ ), .C1(_04504_ ), .C2(fanout_net_46 ), .ZN(_04505_ ) );
NAND2_X1 _12399_ ( .A1(_04496_ ), .A2(_04505_ ), .ZN(_04506_ ) );
OAI21_X1 _12400_ ( .A(_04506_ ), .B1(_04340_ ), .B2(_04330_ ), .ZN(_04507_ ) );
AND2_X1 _12401_ ( .A1(_04481_ ), .A2(_04507_ ), .ZN(_04508_ ) );
NOR2_X1 _12402_ ( .A1(_02885_ ), .A2(_04508_ ), .ZN(_04509_ ) );
AND4_X1 _12403_ ( .A1(_02860_ ), .A2(_04481_ ), .A3(_02879_ ), .A4(_04507_ ), .ZN(_04510_ ) );
NOR3_X1 _12404_ ( .A1(_04480_ ), .A2(_04509_ ), .A3(_04510_ ), .ZN(_04511_ ) );
OR3_X1 _12405_ ( .A1(_04330_ ), .A2(\EX_LS_result_reg [24] ), .A3(_04340_ ), .ZN(_04512_ ) );
OR2_X1 _12406_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04513_ ) );
OAI211_X1 _12407_ ( .A(_04513_ ), .B(_04490_ ), .C1(_04349_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04514_ ) );
NOR2_X1 _12408_ ( .A1(_04349_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04515_ ) );
OAI21_X1 _12409_ ( .A(fanout_net_43 ), .B1(fanout_net_36 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04516_ ) );
OAI211_X1 _12410_ ( .A(_04514_ ), .B(_04356_ ), .C1(_04515_ ), .C2(_04516_ ), .ZN(_04517_ ) );
MUX2_X1 _12411_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04518_ ) );
MUX2_X1 _12412_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04519_ ) );
MUX2_X1 _12413_ ( .A(_04518_ ), .B(_04519_ ), .S(_04490_ ), .Z(_04520_ ) );
OAI211_X1 _12414_ ( .A(_04344_ ), .B(_04517_ ), .C1(_04520_ ), .C2(_04356_ ), .ZN(_04521_ ) );
OR2_X1 _12415_ ( .A1(fanout_net_36 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04522_ ) );
OAI211_X1 _12416_ ( .A(_04522_ ), .B(fanout_net_43 ), .C1(_04349_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04523_ ) );
NAND2_X1 _12417_ ( .A1(_02113_ ), .A2(fanout_net_36 ), .ZN(_04524_ ) );
OAI211_X1 _12418_ ( .A(_04524_ ), .B(_04490_ ), .C1(fanout_net_36 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04525_ ) );
NAND3_X1 _12419_ ( .A1(_04523_ ), .A2(_04525_ ), .A3(_04356_ ), .ZN(_04526_ ) );
MUX2_X1 _12420_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04527_ ) );
MUX2_X1 _12421_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_36 ), .Z(_04528_ ) );
MUX2_X1 _12422_ ( .A(_04527_ ), .B(_04528_ ), .S(_04490_ ), .Z(_04529_ ) );
OAI211_X1 _12423_ ( .A(fanout_net_47 ), .B(_04526_ ), .C1(_04529_ ), .C2(_04356_ ), .ZN(_04530_ ) );
NAND2_X1 _12424_ ( .A1(_04521_ ), .A2(_04530_ ), .ZN(_04531_ ) );
OAI21_X1 _12425_ ( .A(_04531_ ), .B1(_04382_ ), .B2(_04381_ ), .ZN(_04532_ ) );
AND2_X1 _12426_ ( .A1(_04512_ ), .A2(_04532_ ), .ZN(_04533_ ) );
XNOR2_X1 _12427_ ( .A(_02162_ ), .B(_04533_ ), .ZN(_04534_ ) );
INV_X1 _12428_ ( .A(\EX_LS_result_reg [25] ), .ZN(_04535_ ) );
OR3_X1 _12429_ ( .A1(_04381_ ), .A2(_04535_ ), .A3(_04382_ ), .ZN(_04536_ ) );
OR2_X1 _12430_ ( .A1(fanout_net_37 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04537_ ) );
OAI211_X1 _12431_ ( .A(_04537_ ), .B(_04388_ ), .C1(_04389_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04538_ ) );
OR2_X1 _12432_ ( .A1(fanout_net_37 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04539_ ) );
OAI211_X1 _12433_ ( .A(_04539_ ), .B(fanout_net_43 ), .C1(_04364_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04540_ ) );
NAND3_X1 _12434_ ( .A1(_04538_ ), .A2(_04540_ ), .A3(fanout_net_46 ), .ZN(_04541_ ) );
MUX2_X1 _12435_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04542_ ) );
MUX2_X1 _12436_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04543_ ) );
MUX2_X1 _12437_ ( .A(_04542_ ), .B(_04543_ ), .S(_04363_ ), .Z(_04544_ ) );
OAI211_X1 _12438_ ( .A(_04344_ ), .B(_04541_ ), .C1(_04544_ ), .C2(fanout_net_46 ), .ZN(_04545_ ) );
NOR2_X1 _12439_ ( .A1(_04364_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04546_ ) );
OAI21_X1 _12440_ ( .A(fanout_net_43 ), .B1(fanout_net_37 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04547_ ) );
NOR2_X1 _12441_ ( .A1(fanout_net_37 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04548_ ) );
OAI21_X1 _12442_ ( .A(_04363_ ), .B1(_04364_ ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04549_ ) );
OAI221_X1 _12443_ ( .A(_04370_ ), .B1(_04546_ ), .B2(_04547_ ), .C1(_04548_ ), .C2(_04549_ ), .ZN(_04550_ ) );
MUX2_X1 _12444_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04551_ ) );
MUX2_X1 _12445_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_37 ), .Z(_04552_ ) );
MUX2_X1 _12446_ ( .A(_04551_ ), .B(_04552_ ), .S(fanout_net_43 ), .Z(_04553_ ) );
OAI211_X1 _12447_ ( .A(fanout_net_47 ), .B(_04550_ ), .C1(_04553_ ), .C2(_04370_ ), .ZN(_04554_ ) );
OAI211_X1 _12448_ ( .A(_04545_ ), .B(_04554_ ), .C1(_04381_ ), .C2(_04382_ ), .ZN(_04555_ ) );
NAND2_X1 _12449_ ( .A1(_04536_ ), .A2(_04555_ ), .ZN(_04556_ ) );
XNOR2_X1 _12450_ ( .A(_02834_ ), .B(_04556_ ), .ZN(_04557_ ) );
AND2_X1 _12451_ ( .A1(_04534_ ), .A2(_04557_ ), .ZN(_04558_ ) );
AND3_X1 _12452_ ( .A1(_04456_ ), .A2(_04511_ ), .A3(_04558_ ), .ZN(_04559_ ) );
BUF_X4 _12453_ ( .A(_04328_ ), .Z(_04560_ ) );
OR3_X1 _12454_ ( .A1(_04560_ ), .A2(\EX_LS_result_reg [22] ), .A3(_04339_ ), .ZN(_04561_ ) );
BUF_X4 _12455_ ( .A(_04343_ ), .Z(_04562_ ) );
OR2_X1 _12456_ ( .A1(_04347_ ), .A2(\myreg.Reg[1][22] ), .ZN(_04563_ ) );
BUF_X4 _12457_ ( .A(_04361_ ), .Z(_04564_ ) );
OAI211_X1 _12458_ ( .A(_04563_ ), .B(_04564_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[0][22] ), .ZN(_04565_ ) );
OR2_X1 _12459_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][22] ), .ZN(_04566_ ) );
OAI211_X1 _12460_ ( .A(_04566_ ), .B(fanout_net_43 ), .C1(_04348_ ), .C2(\myreg.Reg[3][22] ), .ZN(_04567_ ) );
NAND3_X1 _12461_ ( .A1(_04565_ ), .A2(_04355_ ), .A3(_04567_ ), .ZN(_04568_ ) );
MUX2_X1 _12462_ ( .A(\myreg.Reg[6][22] ), .B(\myreg.Reg[7][22] ), .S(fanout_net_37 ), .Z(_04569_ ) );
MUX2_X1 _12463_ ( .A(\myreg.Reg[4][22] ), .B(\myreg.Reg[5][22] ), .S(fanout_net_37 ), .Z(_04570_ ) );
MUX2_X1 _12464_ ( .A(_04569_ ), .B(_04570_ ), .S(_04489_ ), .Z(_04571_ ) );
OAI211_X1 _12465_ ( .A(_04562_ ), .B(_04568_ ), .C1(_04571_ ), .C2(_04483_ ), .ZN(_04572_ ) );
OR2_X1 _12466_ ( .A1(_04347_ ), .A2(\myreg.Reg[13][22] ), .ZN(_04573_ ) );
OAI211_X1 _12467_ ( .A(_04573_ ), .B(_04564_ ), .C1(fanout_net_37 ), .C2(\myreg.Reg[12][22] ), .ZN(_04574_ ) );
OR2_X1 _12468_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[14][22] ), .ZN(_04575_ ) );
OAI211_X1 _12469_ ( .A(_04575_ ), .B(fanout_net_43 ), .C1(_04348_ ), .C2(\myreg.Reg[15][22] ), .ZN(_04576_ ) );
NAND3_X1 _12470_ ( .A1(_04574_ ), .A2(fanout_net_46 ), .A3(_04576_ ), .ZN(_04577_ ) );
MUX2_X1 _12471_ ( .A(\myreg.Reg[8][22] ), .B(\myreg.Reg[9][22] ), .S(fanout_net_37 ), .Z(_04578_ ) );
MUX2_X1 _12472_ ( .A(\myreg.Reg[10][22] ), .B(\myreg.Reg[11][22] ), .S(fanout_net_37 ), .Z(_04579_ ) );
MUX2_X1 _12473_ ( .A(_04578_ ), .B(_04579_ ), .S(fanout_net_43 ), .Z(_04580_ ) );
OAI211_X1 _12474_ ( .A(fanout_net_47 ), .B(_04577_ ), .C1(_04580_ ), .C2(fanout_net_46 ), .ZN(_04581_ ) );
BUF_X2 _12475_ ( .A(_04328_ ), .Z(_04582_ ) );
BUF_X2 _12476_ ( .A(_04338_ ), .Z(_04583_ ) );
OAI211_X1 _12477_ ( .A(_04572_ ), .B(_04581_ ), .C1(_04582_ ), .C2(_04583_ ), .ZN(_04584_ ) );
NAND2_X1 _12478_ ( .A1(_04561_ ), .A2(_04584_ ), .ZN(_04585_ ) );
XOR2_X1 _12479_ ( .A(_02748_ ), .B(_04585_ ), .Z(_04586_ ) );
OR3_X1 _12480_ ( .A1(_04328_ ), .A2(\EX_LS_result_reg [23] ), .A3(_04338_ ), .ZN(_04587_ ) );
OR2_X1 _12481_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[8][23] ), .ZN(_04588_ ) );
BUF_X2 _12482_ ( .A(_04346_ ), .Z(_04589_ ) );
OAI211_X1 _12483_ ( .A(_04588_ ), .B(_04361_ ), .C1(_04589_ ), .C2(\myreg.Reg[9][23] ), .ZN(_04590_ ) );
OR2_X1 _12484_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[10][23] ), .ZN(_04591_ ) );
OAI211_X1 _12485_ ( .A(_04591_ ), .B(fanout_net_43 ), .C1(_04589_ ), .C2(\myreg.Reg[11][23] ), .ZN(_04592_ ) );
NAND3_X1 _12486_ ( .A1(_04590_ ), .A2(_04592_ ), .A3(_04354_ ), .ZN(_04593_ ) );
MUX2_X1 _12487_ ( .A(\myreg.Reg[14][23] ), .B(\myreg.Reg[15][23] ), .S(fanout_net_37 ), .Z(_04594_ ) );
MUX2_X1 _12488_ ( .A(\myreg.Reg[12][23] ), .B(\myreg.Reg[13][23] ), .S(fanout_net_37 ), .Z(_04595_ ) );
MUX2_X1 _12489_ ( .A(_04594_ ), .B(_04595_ ), .S(_04360_ ), .Z(_04596_ ) );
OAI211_X1 _12490_ ( .A(fanout_net_47 ), .B(_04593_ ), .C1(_04596_ ), .C2(_04482_ ), .ZN(_04597_ ) );
OAI21_X1 _12491_ ( .A(_04360_ ), .B1(_04347_ ), .B2(\myreg.Reg[1][23] ), .ZN(_04598_ ) );
NOR2_X1 _12492_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[0][23] ), .ZN(_04599_ ) );
NOR2_X1 _12493_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][23] ), .ZN(_04600_ ) );
OAI21_X1 _12494_ ( .A(fanout_net_43 ), .B1(_04347_ ), .B2(\myreg.Reg[3][23] ), .ZN(_04601_ ) );
OAI221_X1 _12495_ ( .A(_04353_ ), .B1(_04598_ ), .B2(_04599_ ), .C1(_04600_ ), .C2(_04601_ ), .ZN(_04602_ ) );
MUX2_X1 _12496_ ( .A(\myreg.Reg[6][23] ), .B(\myreg.Reg[7][23] ), .S(fanout_net_37 ), .Z(_04603_ ) );
MUX2_X1 _12497_ ( .A(\myreg.Reg[4][23] ), .B(\myreg.Reg[5][23] ), .S(fanout_net_37 ), .Z(_04604_ ) );
MUX2_X1 _12498_ ( .A(_04603_ ), .B(_04604_ ), .S(_04360_ ), .Z(_04605_ ) );
OAI211_X1 _12499_ ( .A(_04343_ ), .B(_04602_ ), .C1(_04605_ ), .C2(_04482_ ), .ZN(_04606_ ) );
OAI211_X1 _12500_ ( .A(_04597_ ), .B(_04606_ ), .C1(_04329_ ), .C2(_04339_ ), .ZN(_04607_ ) );
NAND2_X1 _12501_ ( .A1(_04587_ ), .A2(_04607_ ), .ZN(_04608_ ) );
XOR2_X1 _12502_ ( .A(_02726_ ), .B(_04608_ ), .Z(_04609_ ) );
AND2_X1 _12503_ ( .A1(_04586_ ), .A2(_04609_ ), .ZN(_04610_ ) );
OR3_X2 _12504_ ( .A1(_04329_ ), .A2(\EX_LS_result_reg [21] ), .A3(_04339_ ), .ZN(_04611_ ) );
OR2_X1 _12505_ ( .A1(\myreg.Reg[0][21] ), .A2(fanout_net_37 ), .ZN(_04612_ ) );
BUF_X4 _12506_ ( .A(_04347_ ), .Z(_04613_ ) );
OAI211_X1 _12507_ ( .A(_04612_ ), .B(_04489_ ), .C1(\myreg.Reg[1][21] ), .C2(_04613_ ), .ZN(_04614_ ) );
OR2_X1 _12508_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[2][21] ), .ZN(_04615_ ) );
OAI211_X1 _12509_ ( .A(_04615_ ), .B(fanout_net_43 ), .C1(_04613_ ), .C2(\myreg.Reg[3][21] ), .ZN(_04616_ ) );
NAND3_X1 _12510_ ( .A1(_04614_ ), .A2(_04616_ ), .A3(_04482_ ), .ZN(_04617_ ) );
MUX2_X1 _12511_ ( .A(\myreg.Reg[6][21] ), .B(\myreg.Reg[7][21] ), .S(fanout_net_37 ), .Z(_04618_ ) );
MUX2_X1 _12512_ ( .A(\myreg.Reg[4][21] ), .B(\myreg.Reg[5][21] ), .S(fanout_net_37 ), .Z(_04619_ ) );
BUF_X4 _12513_ ( .A(_04360_ ), .Z(_04620_ ) );
MUX2_X1 _12514_ ( .A(_04618_ ), .B(_04619_ ), .S(_04620_ ), .Z(_04621_ ) );
BUF_X4 _12515_ ( .A(_04354_ ), .Z(_04622_ ) );
OAI211_X1 _12516_ ( .A(_04562_ ), .B(_04617_ ), .C1(_04621_ ), .C2(_04622_ ), .ZN(_04623_ ) );
OR2_X1 _12517_ ( .A1(_04347_ ), .A2(\myreg.Reg[15][21] ), .ZN(_04624_ ) );
OAI211_X1 _12518_ ( .A(_04624_ ), .B(fanout_net_44 ), .C1(fanout_net_37 ), .C2(\myreg.Reg[14][21] ), .ZN(_04625_ ) );
OR2_X1 _12519_ ( .A1(fanout_net_37 ), .A2(\myreg.Reg[12][21] ), .ZN(_04626_ ) );
OAI211_X1 _12520_ ( .A(_04626_ ), .B(_04620_ ), .C1(_04613_ ), .C2(\myreg.Reg[13][21] ), .ZN(_04627_ ) );
NAND3_X1 _12521_ ( .A1(_04625_ ), .A2(fanout_net_46 ), .A3(_04627_ ), .ZN(_04628_ ) );
MUX2_X1 _12522_ ( .A(\myreg.Reg[8][21] ), .B(\myreg.Reg[9][21] ), .S(fanout_net_38 ), .Z(_04629_ ) );
MUX2_X1 _12523_ ( .A(\myreg.Reg[10][21] ), .B(\myreg.Reg[11][21] ), .S(fanout_net_38 ), .Z(_04630_ ) );
MUX2_X1 _12524_ ( .A(_04629_ ), .B(_04630_ ), .S(fanout_net_44 ), .Z(_04631_ ) );
OAI211_X1 _12525_ ( .A(fanout_net_47 ), .B(_04628_ ), .C1(_04631_ ), .C2(fanout_net_46 ), .ZN(_04632_ ) );
OAI211_X1 _12526_ ( .A(_04623_ ), .B(_04632_ ), .C1(_04582_ ), .C2(_04583_ ), .ZN(_04633_ ) );
NAND2_X1 _12527_ ( .A1(_04611_ ), .A2(_04633_ ), .ZN(_04634_ ) );
AND2_X1 _12528_ ( .A1(_02793_ ), .A2(_04634_ ), .ZN(_04635_ ) );
NOR2_X1 _12529_ ( .A1(_02793_ ), .A2(_04634_ ), .ZN(_04636_ ) );
NOR2_X1 _12530_ ( .A1(_04635_ ), .A2(_04636_ ), .ZN(_04637_ ) );
BUF_X2 _12531_ ( .A(_04338_ ), .Z(_04638_ ) );
OR3_X1 _12532_ ( .A1(_04560_ ), .A2(\EX_LS_result_reg [20] ), .A3(_04638_ ), .ZN(_04639_ ) );
OR2_X1 _12533_ ( .A1(_04589_ ), .A2(\myreg.Reg[1][20] ), .ZN(_04640_ ) );
OAI211_X1 _12534_ ( .A(_04640_ ), .B(_04362_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[0][20] ), .ZN(_04641_ ) );
OR2_X1 _12535_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[2][20] ), .ZN(_04642_ ) );
OAI211_X1 _12536_ ( .A(_04642_ ), .B(fanout_net_44 ), .C1(_04348_ ), .C2(\myreg.Reg[3][20] ), .ZN(_04643_ ) );
NAND3_X1 _12537_ ( .A1(_04641_ ), .A2(_04355_ ), .A3(_04643_ ), .ZN(_04644_ ) );
MUX2_X1 _12538_ ( .A(\myreg.Reg[6][20] ), .B(\myreg.Reg[7][20] ), .S(fanout_net_38 ), .Z(_04645_ ) );
MUX2_X1 _12539_ ( .A(\myreg.Reg[4][20] ), .B(\myreg.Reg[5][20] ), .S(fanout_net_38 ), .Z(_04646_ ) );
MUX2_X1 _12540_ ( .A(_04645_ ), .B(_04646_ ), .S(_04564_ ), .Z(_04647_ ) );
OAI211_X1 _12541_ ( .A(_04562_ ), .B(_04644_ ), .C1(_04647_ ), .C2(_04483_ ), .ZN(_04648_ ) );
OR2_X1 _12542_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[14][20] ), .ZN(_04649_ ) );
OAI211_X1 _12543_ ( .A(_04649_ ), .B(fanout_net_44 ), .C1(_04348_ ), .C2(\myreg.Reg[15][20] ), .ZN(_04650_ ) );
OR2_X1 _12544_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[12][20] ), .ZN(_04651_ ) );
OAI211_X1 _12545_ ( .A(_04651_ ), .B(_04564_ ), .C1(_04348_ ), .C2(\myreg.Reg[13][20] ), .ZN(_04652_ ) );
NAND3_X1 _12546_ ( .A1(_04650_ ), .A2(_04652_ ), .A3(fanout_net_46 ), .ZN(_04653_ ) );
MUX2_X1 _12547_ ( .A(\myreg.Reg[8][20] ), .B(\myreg.Reg[9][20] ), .S(fanout_net_38 ), .Z(_04654_ ) );
MUX2_X1 _12548_ ( .A(\myreg.Reg[10][20] ), .B(\myreg.Reg[11][20] ), .S(fanout_net_38 ), .Z(_04655_ ) );
MUX2_X1 _12549_ ( .A(_04654_ ), .B(_04655_ ), .S(fanout_net_44 ), .Z(_04656_ ) );
OAI211_X1 _12550_ ( .A(fanout_net_47 ), .B(_04653_ ), .C1(_04656_ ), .C2(fanout_net_46 ), .ZN(_04657_ ) );
OAI211_X1 _12551_ ( .A(_04648_ ), .B(_04657_ ), .C1(_04582_ ), .C2(_04583_ ), .ZN(_04658_ ) );
NAND2_X1 _12552_ ( .A1(_04639_ ), .A2(_04658_ ), .ZN(_04659_ ) );
XOR2_X1 _12553_ ( .A(_02770_ ), .B(_04659_ ), .Z(_04660_ ) );
AND3_X1 _12554_ ( .A1(_04610_ ), .A2(_04637_ ), .A3(_04660_ ), .ZN(_04661_ ) );
OR3_X1 _12555_ ( .A1(_04329_ ), .A2(\EX_LS_result_reg [18] ), .A3(_04339_ ), .ZN(_04662_ ) );
OR2_X1 _12556_ ( .A1(_04347_ ), .A2(\myreg.Reg[1][18] ), .ZN(_04663_ ) );
OAI211_X1 _12557_ ( .A(_04663_ ), .B(_04489_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[0][18] ), .ZN(_04664_ ) );
OR2_X1 _12558_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[2][18] ), .ZN(_04665_ ) );
OAI211_X1 _12559_ ( .A(_04665_ ), .B(fanout_net_44 ), .C1(_04613_ ), .C2(\myreg.Reg[3][18] ), .ZN(_04666_ ) );
NAND3_X1 _12560_ ( .A1(_04664_ ), .A2(_04482_ ), .A3(_04666_ ), .ZN(_04667_ ) );
MUX2_X1 _12561_ ( .A(\myreg.Reg[6][18] ), .B(\myreg.Reg[7][18] ), .S(fanout_net_38 ), .Z(_04668_ ) );
MUX2_X1 _12562_ ( .A(\myreg.Reg[4][18] ), .B(\myreg.Reg[5][18] ), .S(fanout_net_38 ), .Z(_04669_ ) );
MUX2_X1 _12563_ ( .A(_04668_ ), .B(_04669_ ), .S(_04620_ ), .Z(_04670_ ) );
OAI211_X1 _12564_ ( .A(_04562_ ), .B(_04667_ ), .C1(_04670_ ), .C2(_04622_ ), .ZN(_04671_ ) );
OR2_X1 _12565_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[14][18] ), .ZN(_04672_ ) );
OAI211_X1 _12566_ ( .A(_04672_ ), .B(fanout_net_44 ), .C1(_04613_ ), .C2(\myreg.Reg[15][18] ), .ZN(_04673_ ) );
OR2_X1 _12567_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[12][18] ), .ZN(_04674_ ) );
OAI211_X1 _12568_ ( .A(_04674_ ), .B(_04489_ ), .C1(_04613_ ), .C2(\myreg.Reg[13][18] ), .ZN(_04675_ ) );
NAND3_X1 _12569_ ( .A1(_04673_ ), .A2(_04675_ ), .A3(fanout_net_46 ), .ZN(_04676_ ) );
MUX2_X1 _12570_ ( .A(\myreg.Reg[8][18] ), .B(\myreg.Reg[9][18] ), .S(fanout_net_38 ), .Z(_04677_ ) );
MUX2_X1 _12571_ ( .A(\myreg.Reg[10][18] ), .B(\myreg.Reg[11][18] ), .S(fanout_net_38 ), .Z(_04678_ ) );
MUX2_X1 _12572_ ( .A(_04677_ ), .B(_04678_ ), .S(fanout_net_44 ), .Z(_04679_ ) );
OAI211_X1 _12573_ ( .A(fanout_net_47 ), .B(_04676_ ), .C1(_04679_ ), .C2(fanout_net_46 ), .ZN(_04680_ ) );
OAI211_X1 _12574_ ( .A(_04671_ ), .B(_04680_ ), .C1(_04582_ ), .C2(_04583_ ), .ZN(_04681_ ) );
NAND2_X1 _12575_ ( .A1(_04662_ ), .A2(_04681_ ), .ZN(_04682_ ) );
XOR2_X1 _12576_ ( .A(_02642_ ), .B(_04682_ ), .Z(_04683_ ) );
OR3_X1 _12577_ ( .A1(_04328_ ), .A2(\EX_LS_result_reg [19] ), .A3(_04338_ ), .ZN(_04684_ ) );
OR2_X1 _12578_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[0][19] ), .ZN(_04685_ ) );
CLKBUF_X2 _12579_ ( .A(_04346_ ), .Z(_04686_ ) );
BUF_X2 _12580_ ( .A(_04686_ ), .Z(_04687_ ) );
OAI211_X1 _12581_ ( .A(_04685_ ), .B(_04620_ ), .C1(_04687_ ), .C2(\myreg.Reg[1][19] ), .ZN(_04688_ ) );
OR2_X1 _12582_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[2][19] ), .ZN(_04689_ ) );
OAI211_X1 _12583_ ( .A(_04689_ ), .B(fanout_net_44 ), .C1(_04687_ ), .C2(\myreg.Reg[3][19] ), .ZN(_04690_ ) );
NAND3_X1 _12584_ ( .A1(_04688_ ), .A2(_04690_ ), .A3(_04354_ ), .ZN(_04691_ ) );
MUX2_X1 _12585_ ( .A(\myreg.Reg[6][19] ), .B(\myreg.Reg[7][19] ), .S(fanout_net_38 ), .Z(_04692_ ) );
MUX2_X1 _12586_ ( .A(\myreg.Reg[4][19] ), .B(\myreg.Reg[5][19] ), .S(fanout_net_38 ), .Z(_04693_ ) );
MUX2_X1 _12587_ ( .A(_04692_ ), .B(_04693_ ), .S(_04361_ ), .Z(_04694_ ) );
OAI211_X1 _12588_ ( .A(_04343_ ), .B(_04691_ ), .C1(_04694_ ), .C2(_04355_ ), .ZN(_04695_ ) );
OR2_X1 _12589_ ( .A1(_04686_ ), .A2(\myreg.Reg[13][19] ), .ZN(_04696_ ) );
BUF_X4 _12590_ ( .A(_04360_ ), .Z(_04697_ ) );
OAI211_X1 _12591_ ( .A(_04696_ ), .B(_04697_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[12][19] ), .ZN(_04698_ ) );
OR2_X1 _12592_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[14][19] ), .ZN(_04699_ ) );
OAI211_X1 _12593_ ( .A(_04699_ ), .B(fanout_net_44 ), .C1(_04484_ ), .C2(\myreg.Reg[15][19] ), .ZN(_04700_ ) );
NAND3_X1 _12594_ ( .A1(_04698_ ), .A2(fanout_net_46 ), .A3(_04700_ ), .ZN(_04701_ ) );
MUX2_X1 _12595_ ( .A(\myreg.Reg[8][19] ), .B(\myreg.Reg[9][19] ), .S(fanout_net_38 ), .Z(_04702_ ) );
MUX2_X1 _12596_ ( .A(\myreg.Reg[10][19] ), .B(\myreg.Reg[11][19] ), .S(fanout_net_38 ), .Z(_04703_ ) );
MUX2_X1 _12597_ ( .A(_04702_ ), .B(_04703_ ), .S(fanout_net_44 ), .Z(_04704_ ) );
OAI211_X1 _12598_ ( .A(fanout_net_47 ), .B(_04701_ ), .C1(_04704_ ), .C2(fanout_net_46 ), .ZN(_04705_ ) );
OAI211_X1 _12599_ ( .A(_04695_ ), .B(_04705_ ), .C1(_04560_ ), .C2(_04638_ ), .ZN(_04706_ ) );
NAND2_X1 _12600_ ( .A1(_04684_ ), .A2(_04706_ ), .ZN(_04707_ ) );
INV_X1 _12601_ ( .A(_04707_ ), .ZN(_04708_ ) );
XNOR2_X1 _12602_ ( .A(_02618_ ), .B(_04708_ ), .ZN(_04709_ ) );
AND2_X1 _12603_ ( .A1(_04683_ ), .A2(_04709_ ), .ZN(_04710_ ) );
OR3_X1 _12604_ ( .A1(_04329_ ), .A2(\EX_LS_result_reg [17] ), .A3(_04339_ ), .ZN(_04711_ ) );
OR2_X1 _12605_ ( .A1(_04686_ ), .A2(\myreg.Reg[1][17] ), .ZN(_04712_ ) );
OAI211_X1 _12606_ ( .A(_04712_ ), .B(_04489_ ), .C1(fanout_net_38 ), .C2(\myreg.Reg[0][17] ), .ZN(_04713_ ) );
OR2_X1 _12607_ ( .A1(fanout_net_38 ), .A2(\myreg.Reg[2][17] ), .ZN(_04714_ ) );
OAI211_X1 _12608_ ( .A(_04714_ ), .B(fanout_net_44 ), .C1(_04687_ ), .C2(\myreg.Reg[3][17] ), .ZN(_04715_ ) );
NAND3_X1 _12609_ ( .A1(_04713_ ), .A2(_04482_ ), .A3(_04715_ ), .ZN(_04716_ ) );
MUX2_X1 _12610_ ( .A(\myreg.Reg[6][17] ), .B(\myreg.Reg[7][17] ), .S(fanout_net_38 ), .Z(_04717_ ) );
MUX2_X1 _12611_ ( .A(\myreg.Reg[4][17] ), .B(\myreg.Reg[5][17] ), .S(fanout_net_38 ), .Z(_04718_ ) );
MUX2_X1 _12612_ ( .A(_04717_ ), .B(_04718_ ), .S(_04697_ ), .Z(_04719_ ) );
OAI211_X1 _12613_ ( .A(_04343_ ), .B(_04716_ ), .C1(_04719_ ), .C2(_04622_ ), .ZN(_04720_ ) );
OR2_X1 _12614_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[14][17] ), .ZN(_04721_ ) );
OAI211_X1 _12615_ ( .A(_04721_ ), .B(fanout_net_44 ), .C1(_04613_ ), .C2(\myreg.Reg[15][17] ), .ZN(_04722_ ) );
OR2_X1 _12616_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[12][17] ), .ZN(_04723_ ) );
OAI211_X1 _12617_ ( .A(_04723_ ), .B(_04620_ ), .C1(_04687_ ), .C2(\myreg.Reg[13][17] ), .ZN(_04724_ ) );
NAND3_X1 _12618_ ( .A1(_04722_ ), .A2(_04724_ ), .A3(fanout_net_46 ), .ZN(_04725_ ) );
MUX2_X1 _12619_ ( .A(\myreg.Reg[8][17] ), .B(\myreg.Reg[9][17] ), .S(fanout_net_39 ), .Z(_04726_ ) );
MUX2_X1 _12620_ ( .A(\myreg.Reg[10][17] ), .B(\myreg.Reg[11][17] ), .S(fanout_net_39 ), .Z(_04727_ ) );
MUX2_X1 _12621_ ( .A(_04726_ ), .B(_04727_ ), .S(fanout_net_44 ), .Z(_04728_ ) );
OAI211_X1 _12622_ ( .A(fanout_net_47 ), .B(_04725_ ), .C1(_04728_ ), .C2(fanout_net_46 ), .ZN(_04729_ ) );
OAI211_X1 _12623_ ( .A(_04720_ ), .B(_04729_ ), .C1(_04560_ ), .C2(_04638_ ), .ZN(_04730_ ) );
NAND2_X1 _12624_ ( .A1(_04711_ ), .A2(_04730_ ), .ZN(_04731_ ) );
XOR2_X1 _12625_ ( .A(_02688_ ), .B(_04731_ ), .Z(_04732_ ) );
OR3_X1 _12626_ ( .A1(_04330_ ), .A2(\EX_LS_result_reg [16] ), .A3(_04340_ ), .ZN(_04733_ ) );
OR2_X1 _12627_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[4][16] ), .ZN(_04734_ ) );
OAI211_X1 _12628_ ( .A(_04734_ ), .B(_04490_ ), .C1(_04349_ ), .C2(\myreg.Reg[5][16] ), .ZN(_04735_ ) );
OR2_X1 _12629_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[6][16] ), .ZN(_04736_ ) );
OAI211_X1 _12630_ ( .A(_04736_ ), .B(fanout_net_44 ), .C1(_04349_ ), .C2(\myreg.Reg[7][16] ), .ZN(_04737_ ) );
NAND3_X1 _12631_ ( .A1(_04735_ ), .A2(_04737_ ), .A3(fanout_net_46 ), .ZN(_04738_ ) );
MUX2_X1 _12632_ ( .A(\myreg.Reg[2][16] ), .B(\myreg.Reg[3][16] ), .S(fanout_net_39 ), .Z(_04739_ ) );
MUX2_X1 _12633_ ( .A(\myreg.Reg[0][16] ), .B(\myreg.Reg[1][16] ), .S(fanout_net_39 ), .Z(_04740_ ) );
MUX2_X1 _12634_ ( .A(_04739_ ), .B(_04740_ ), .S(_04490_ ), .Z(_04741_ ) );
OAI211_X1 _12635_ ( .A(_04344_ ), .B(_04738_ ), .C1(_04741_ ), .C2(fanout_net_46 ), .ZN(_04742_ ) );
NOR2_X1 _12636_ ( .A1(_04485_ ), .A2(\myreg.Reg[11][16] ), .ZN(_04743_ ) );
OAI21_X1 _12637_ ( .A(fanout_net_44 ), .B1(fanout_net_39 ), .B2(\myreg.Reg[10][16] ), .ZN(_04744_ ) );
NOR2_X1 _12638_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[8][16] ), .ZN(_04745_ ) );
OAI21_X1 _12639_ ( .A(_04490_ ), .B1(_04485_ ), .B2(\myreg.Reg[9][16] ), .ZN(_04746_ ) );
OAI221_X1 _12640_ ( .A(_04483_ ), .B1(_04743_ ), .B2(_04744_ ), .C1(_04745_ ), .C2(_04746_ ), .ZN(_04747_ ) );
MUX2_X1 _12641_ ( .A(\myreg.Reg[12][16] ), .B(\myreg.Reg[13][16] ), .S(fanout_net_39 ), .Z(_04748_ ) );
MUX2_X1 _12642_ ( .A(\myreg.Reg[14][16] ), .B(\myreg.Reg[15][16] ), .S(fanout_net_39 ), .Z(_04749_ ) );
MUX2_X1 _12643_ ( .A(_04748_ ), .B(_04749_ ), .S(fanout_net_44 ), .Z(_04750_ ) );
OAI211_X1 _12644_ ( .A(fanout_net_47 ), .B(_04747_ ), .C1(_04750_ ), .C2(_04356_ ), .ZN(_04751_ ) );
OAI211_X1 _12645_ ( .A(_04742_ ), .B(_04751_ ), .C1(_04330_ ), .C2(_04340_ ), .ZN(_04752_ ) );
NAND2_X1 _12646_ ( .A1(_04733_ ), .A2(_04752_ ), .ZN(_04753_ ) );
XOR2_X1 _12647_ ( .A(_02666_ ), .B(_04753_ ), .Z(_04754_ ) );
AND2_X1 _12648_ ( .A1(_04732_ ), .A2(_04754_ ), .ZN(_04755_ ) );
AND2_X1 _12649_ ( .A1(_04710_ ), .A2(_04755_ ), .ZN(_04756_ ) );
AND2_X1 _12650_ ( .A1(_04661_ ), .A2(_04756_ ), .ZN(_04757_ ) );
OR3_X4 _12651_ ( .A1(_04329_ ), .A2(\EX_LS_result_reg [6] ), .A3(_04339_ ), .ZN(_04758_ ) );
OR2_X1 _12652_ ( .A1(_04347_ ), .A2(\myreg.Reg[5][6] ), .ZN(_04759_ ) );
OAI211_X1 _12653_ ( .A(_04759_ ), .B(_04489_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[4][6] ), .ZN(_04760_ ) );
OR2_X1 _12654_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[6][6] ), .ZN(_04761_ ) );
OAI211_X1 _12655_ ( .A(_04761_ ), .B(fanout_net_44 ), .C1(_04613_ ), .C2(\myreg.Reg[7][6] ), .ZN(_04762_ ) );
NAND3_X1 _12656_ ( .A1(_04760_ ), .A2(fanout_net_46 ), .A3(_04762_ ), .ZN(_04763_ ) );
MUX2_X1 _12657_ ( .A(\myreg.Reg[2][6] ), .B(\myreg.Reg[3][6] ), .S(fanout_net_39 ), .Z(_04764_ ) );
MUX2_X1 _12658_ ( .A(\myreg.Reg[0][6] ), .B(\myreg.Reg[1][6] ), .S(fanout_net_39 ), .Z(_04765_ ) );
MUX2_X1 _12659_ ( .A(_04764_ ), .B(_04765_ ), .S(_04620_ ), .Z(_04766_ ) );
OAI211_X1 _12660_ ( .A(_04562_ ), .B(_04763_ ), .C1(_04766_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04767_ ) );
NOR2_X1 _12661_ ( .A1(_04687_ ), .A2(\myreg.Reg[11][6] ), .ZN(_04768_ ) );
OAI21_X1 _12662_ ( .A(fanout_net_44 ), .B1(fanout_net_39 ), .B2(\myreg.Reg[10][6] ), .ZN(_04769_ ) );
NOR2_X1 _12663_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[8][6] ), .ZN(_04770_ ) );
OAI21_X1 _12664_ ( .A(_04620_ ), .B1(_04687_ ), .B2(\myreg.Reg[9][6] ), .ZN(_04771_ ) );
OAI221_X1 _12665_ ( .A(_04482_ ), .B1(_04768_ ), .B2(_04769_ ), .C1(_04770_ ), .C2(_04771_ ), .ZN(_04772_ ) );
MUX2_X1 _12666_ ( .A(\myreg.Reg[12][6] ), .B(\myreg.Reg[13][6] ), .S(fanout_net_39 ), .Z(_04773_ ) );
MUX2_X1 _12667_ ( .A(\myreg.Reg[14][6] ), .B(\myreg.Reg[15][6] ), .S(fanout_net_39 ), .Z(_04774_ ) );
MUX2_X1 _12668_ ( .A(_04773_ ), .B(_04774_ ), .S(fanout_net_44 ), .Z(_04775_ ) );
OAI211_X1 _12669_ ( .A(fanout_net_47 ), .B(_04772_ ), .C1(_04775_ ), .C2(_04622_ ), .ZN(_04776_ ) );
OAI211_X1 _12670_ ( .A(_04767_ ), .B(_04776_ ), .C1(_04582_ ), .C2(_04583_ ), .ZN(_04777_ ) );
NAND2_X1 _12671_ ( .A1(_04758_ ), .A2(_04777_ ), .ZN(_04778_ ) );
XNOR2_X1 _12672_ ( .A(_02371_ ), .B(_04778_ ), .ZN(_04779_ ) );
OR3_X4 _12673_ ( .A1(_04329_ ), .A2(\EX_LS_result_reg [7] ), .A3(_04339_ ), .ZN(_04780_ ) );
OR2_X1 _12674_ ( .A1(_04686_ ), .A2(\myreg.Reg[1][7] ), .ZN(_04781_ ) );
OAI211_X1 _12675_ ( .A(_04781_ ), .B(_04489_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[0][7] ), .ZN(_04782_ ) );
OR2_X1 _12676_ ( .A1(_04686_ ), .A2(\myreg.Reg[3][7] ), .ZN(_04783_ ) );
OAI211_X1 _12677_ ( .A(_04783_ ), .B(fanout_net_44 ), .C1(fanout_net_39 ), .C2(\myreg.Reg[2][7] ), .ZN(_04784_ ) );
NAND3_X1 _12678_ ( .A1(_04782_ ), .A2(_04784_ ), .A3(_04482_ ), .ZN(_04785_ ) );
MUX2_X1 _12679_ ( .A(\myreg.Reg[6][7] ), .B(\myreg.Reg[7][7] ), .S(fanout_net_39 ), .Z(_04786_ ) );
MUX2_X1 _12680_ ( .A(\myreg.Reg[4][7] ), .B(\myreg.Reg[5][7] ), .S(fanout_net_39 ), .Z(_04787_ ) );
MUX2_X1 _12681_ ( .A(_04786_ ), .B(_04787_ ), .S(_04620_ ), .Z(_04788_ ) );
OAI211_X1 _12682_ ( .A(_04562_ ), .B(_04785_ ), .C1(_04788_ ), .C2(_04622_ ), .ZN(_04789_ ) );
OR2_X1 _12683_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[14][7] ), .ZN(_04790_ ) );
OAI211_X1 _12684_ ( .A(_04790_ ), .B(fanout_net_44 ), .C1(_04613_ ), .C2(\myreg.Reg[15][7] ), .ZN(_04791_ ) );
OR2_X1 _12685_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[12][7] ), .ZN(_04792_ ) );
OAI211_X1 _12686_ ( .A(_04792_ ), .B(_04620_ ), .C1(_04687_ ), .C2(\myreg.Reg[13][7] ), .ZN(_04793_ ) );
NAND3_X1 _12687_ ( .A1(_04791_ ), .A2(_04793_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04794_ ) );
MUX2_X1 _12688_ ( .A(\myreg.Reg[8][7] ), .B(\myreg.Reg[9][7] ), .S(fanout_net_39 ), .Z(_04795_ ) );
MUX2_X1 _12689_ ( .A(\myreg.Reg[10][7] ), .B(\myreg.Reg[11][7] ), .S(fanout_net_39 ), .Z(_04796_ ) );
MUX2_X1 _12690_ ( .A(_04795_ ), .B(_04796_ ), .S(fanout_net_44 ), .Z(_04797_ ) );
OAI211_X1 _12691_ ( .A(fanout_net_47 ), .B(_04794_ ), .C1(_04797_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04798_ ) );
OAI211_X1 _12692_ ( .A(_04789_ ), .B(_04798_ ), .C1(_04560_ ), .C2(_04638_ ), .ZN(_04799_ ) );
NAND2_X1 _12693_ ( .A1(_04780_ ), .A2(_04799_ ), .ZN(_04800_ ) );
XNOR2_X1 _12694_ ( .A(_02345_ ), .B(_04800_ ), .ZN(_04801_ ) );
NOR2_X1 _12695_ ( .A1(_04779_ ), .A2(_04801_ ), .ZN(_04802_ ) );
OR2_X1 _12696_ ( .A1(_04484_ ), .A2(\myreg.Reg[9][4] ), .ZN(_04803_ ) );
OAI211_X1 _12697_ ( .A(_04803_ ), .B(_04362_ ), .C1(fanout_net_39 ), .C2(\myreg.Reg[8][4] ), .ZN(_04804_ ) );
OR2_X1 _12698_ ( .A1(fanout_net_39 ), .A2(\myreg.Reg[10][4] ), .ZN(_04805_ ) );
OAI211_X1 _12699_ ( .A(_04805_ ), .B(fanout_net_44 ), .C1(_04485_ ), .C2(\myreg.Reg[11][4] ), .ZN(_04806_ ) );
NAND3_X1 _12700_ ( .A1(_04804_ ), .A2(_04622_ ), .A3(_04806_ ), .ZN(_04807_ ) );
MUX2_X1 _12701_ ( .A(\myreg.Reg[14][4] ), .B(\myreg.Reg[15][4] ), .S(fanout_net_40 ), .Z(_04808_ ) );
MUX2_X1 _12702_ ( .A(\myreg.Reg[12][4] ), .B(\myreg.Reg[13][4] ), .S(fanout_net_40 ), .Z(_04809_ ) );
MUX2_X1 _12703_ ( .A(_04808_ ), .B(_04809_ ), .S(_04362_ ), .Z(_04810_ ) );
OAI211_X1 _12704_ ( .A(fanout_net_47 ), .B(_04807_ ), .C1(_04810_ ), .C2(_04483_ ), .ZN(_04811_ ) );
MUX2_X1 _12705_ ( .A(\myreg.Reg[0][4] ), .B(\myreg.Reg[1][4] ), .S(fanout_net_40 ), .Z(_04812_ ) );
AND2_X1 _12706_ ( .A1(_04812_ ), .A2(_04564_ ), .ZN(_04813_ ) );
MUX2_X1 _12707_ ( .A(\myreg.Reg[2][4] ), .B(\myreg.Reg[3][4] ), .S(fanout_net_40 ), .Z(_04814_ ) );
AOI211_X1 _12708_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_04813_ ), .C1(fanout_net_44 ), .C2(_04814_ ), .ZN(_04815_ ) );
MUX2_X1 _12709_ ( .A(\myreg.Reg[6][4] ), .B(\myreg.Reg[7][4] ), .S(fanout_net_40 ), .Z(_04816_ ) );
MUX2_X1 _12710_ ( .A(\myreg.Reg[4][4] ), .B(\myreg.Reg[5][4] ), .S(fanout_net_40 ), .Z(_04817_ ) );
MUX2_X1 _12711_ ( .A(_04816_ ), .B(_04817_ ), .S(_04489_ ), .Z(_04818_ ) );
OAI21_X1 _12712_ ( .A(_04562_ ), .B1(_04818_ ), .B2(_04483_ ), .ZN(_04819_ ) );
OAI221_X2 _12713_ ( .A(_04811_ ), .B1(_04815_ ), .B2(_04819_ ), .C1(_04330_ ), .C2(_04340_ ), .ZN(_04820_ ) );
OR3_X4 _12714_ ( .A1(_04582_ ), .A2(\EX_LS_result_reg [4] ), .A3(_04583_ ), .ZN(_04821_ ) );
NAND2_X1 _12715_ ( .A1(_04820_ ), .A2(_04821_ ), .ZN(_04822_ ) );
XOR2_X1 _12716_ ( .A(_02319_ ), .B(_04822_ ), .Z(_04823_ ) );
OR3_X1 _12717_ ( .A1(_04328_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .A3(_04338_ ), .ZN(_04824_ ) );
NAND2_X1 _12718_ ( .A1(_02166_ ), .A2(fanout_net_40 ), .ZN(_04825_ ) );
OAI211_X1 _12719_ ( .A(_04825_ ), .B(_04361_ ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04826_ ) );
NAND2_X1 _12720_ ( .A1(_02169_ ), .A2(fanout_net_40 ), .ZN(_04827_ ) );
OAI211_X1 _12721_ ( .A(_04827_ ), .B(fanout_net_44 ), .C1(fanout_net_40 ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04828_ ) );
NAND3_X1 _12722_ ( .A1(_04826_ ), .A2(_04828_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04829_ ) );
MUX2_X1 _12723_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04830_ ) );
MUX2_X1 _12724_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04831_ ) );
MUX2_X1 _12725_ ( .A(_04830_ ), .B(_04831_ ), .S(_04360_ ), .Z(_04832_ ) );
OAI211_X1 _12726_ ( .A(_04343_ ), .B(_04829_ ), .C1(_04832_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04833_ ) );
NOR2_X1 _12727_ ( .A1(_04347_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04834_ ) );
OAI21_X1 _12728_ ( .A(fanout_net_44 ), .B1(fanout_net_40 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04835_ ) );
MUX2_X1 _12729_ ( .A(_02179_ ), .B(_02180_ ), .S(fanout_net_40 ), .Z(_04836_ ) );
OAI221_X1 _12730_ ( .A(_04354_ ), .B1(_04834_ ), .B2(_04835_ ), .C1(_04836_ ), .C2(fanout_net_44 ), .ZN(_04837_ ) );
MUX2_X1 _12731_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04838_ ) );
MUX2_X1 _12732_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04839_ ) );
MUX2_X1 _12733_ ( .A(_04838_ ), .B(_04839_ ), .S(fanout_net_44 ), .Z(_04840_ ) );
OAI211_X1 _12734_ ( .A(fanout_net_47 ), .B(_04837_ ), .C1(_04840_ ), .C2(_04482_ ), .ZN(_04841_ ) );
OAI211_X1 _12735_ ( .A(_04833_ ), .B(_04841_ ), .C1(_04329_ ), .C2(_04339_ ), .ZN(_04842_ ) );
NAND2_X2 _12736_ ( .A1(_04824_ ), .A2(_04842_ ), .ZN(_04843_ ) );
XNOR2_X1 _12737_ ( .A(_02188_ ), .B(_04843_ ), .ZN(_04844_ ) );
AND3_X1 _12738_ ( .A1(_04802_ ), .A2(_04823_ ), .A3(_04844_ ), .ZN(_04845_ ) );
OR3_X1 _12739_ ( .A1(_04327_ ), .A2(\EX_LS_result_reg [2] ), .A3(_04337_ ), .ZN(_04846_ ) );
OR2_X1 _12740_ ( .A1(_04345_ ), .A2(\myreg.Reg[1][2] ), .ZN(_04847_ ) );
OAI211_X1 _12741_ ( .A(_04847_ ), .B(_04359_ ), .C1(fanout_net_40 ), .C2(\myreg.Reg[0][2] ), .ZN(_04848_ ) );
OR2_X1 _12742_ ( .A1(fanout_net_40 ), .A2(\myreg.Reg[2][2] ), .ZN(_04849_ ) );
OAI211_X1 _12743_ ( .A(_04849_ ), .B(fanout_net_44 ), .C1(_04346_ ), .C2(\myreg.Reg[3][2] ), .ZN(_04850_ ) );
NAND3_X1 _12744_ ( .A1(_04848_ ), .A2(_04353_ ), .A3(_04850_ ), .ZN(_04851_ ) );
MUX2_X1 _12745_ ( .A(\myreg.Reg[6][2] ), .B(\myreg.Reg[7][2] ), .S(fanout_net_40 ), .Z(_04852_ ) );
MUX2_X1 _12746_ ( .A(\myreg.Reg[4][2] ), .B(\myreg.Reg[5][2] ), .S(fanout_net_40 ), .Z(_04853_ ) );
MUX2_X1 _12747_ ( .A(_04852_ ), .B(_04853_ ), .S(_04359_ ), .Z(_04854_ ) );
OAI211_X1 _12748_ ( .A(_04342_ ), .B(_04851_ ), .C1(_04854_ ), .C2(_04353_ ), .ZN(_04855_ ) );
OR2_X1 _12749_ ( .A1(_04345_ ), .A2(\myreg.Reg[13][2] ), .ZN(_04856_ ) );
OAI211_X1 _12750_ ( .A(_04856_ ), .B(_04359_ ), .C1(fanout_net_40 ), .C2(\myreg.Reg[12][2] ), .ZN(_04857_ ) );
OR2_X1 _12751_ ( .A1(fanout_net_40 ), .A2(\myreg.Reg[14][2] ), .ZN(_04858_ ) );
OAI211_X1 _12752_ ( .A(_04858_ ), .B(fanout_net_45 ), .C1(_04346_ ), .C2(\myreg.Reg[15][2] ), .ZN(_04859_ ) );
NAND3_X1 _12753_ ( .A1(_04857_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04859_ ), .ZN(_04860_ ) );
MUX2_X1 _12754_ ( .A(\myreg.Reg[8][2] ), .B(\myreg.Reg[9][2] ), .S(fanout_net_40 ), .Z(_04861_ ) );
MUX2_X1 _12755_ ( .A(\myreg.Reg[10][2] ), .B(\myreg.Reg[11][2] ), .S(fanout_net_40 ), .Z(_04862_ ) );
MUX2_X1 _12756_ ( .A(_04861_ ), .B(_04862_ ), .S(fanout_net_45 ), .Z(_04863_ ) );
OAI211_X1 _12757_ ( .A(fanout_net_47 ), .B(_04860_ ), .C1(_04863_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04864_ ) );
OAI211_X1 _12758_ ( .A(_04855_ ), .B(_04864_ ), .C1(_04328_ ), .C2(_04338_ ), .ZN(_04865_ ) );
NAND2_X1 _12759_ ( .A1(_04846_ ), .A2(_04865_ ), .ZN(_04866_ ) );
XOR2_X1 _12760_ ( .A(_02258_ ), .B(_04866_ ), .Z(_04867_ ) );
OR2_X1 _12761_ ( .A1(fanout_net_40 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04868_ ) );
OAI211_X1 _12762_ ( .A(_04868_ ), .B(_04360_ ), .C1(_04686_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04869_ ) );
OR2_X1 _12763_ ( .A1(fanout_net_40 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04870_ ) );
OAI211_X1 _12764_ ( .A(_04870_ ), .B(fanout_net_45 ), .C1(_04346_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04871_ ) );
NAND3_X1 _12765_ ( .A1(_04869_ ), .A2(_04871_ ), .A3(_04353_ ), .ZN(_04872_ ) );
MUX2_X1 _12766_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04873_ ) );
MUX2_X1 _12767_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_40 ), .Z(_04874_ ) );
MUX2_X1 _12768_ ( .A(_04873_ ), .B(_04874_ ), .S(_04359_ ), .Z(_04875_ ) );
OAI211_X1 _12769_ ( .A(_04342_ ), .B(_04872_ ), .C1(_04875_ ), .C2(_04353_ ), .ZN(_04876_ ) );
OR2_X1 _12770_ ( .A1(fanout_net_40 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_04877_ ) );
OAI211_X1 _12771_ ( .A(_04877_ ), .B(fanout_net_45 ), .C1(_04346_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ), .ZN(_04878_ ) );
OR2_X1 _12772_ ( .A1(fanout_net_40 ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .ZN(_04879_ ) );
OAI211_X1 _12773_ ( .A(_04879_ ), .B(_04360_ ), .C1(_04346_ ), .C2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_04880_ ) );
NAND3_X1 _12774_ ( .A1(_04878_ ), .A2(_04880_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04881_ ) );
MUX2_X1 _12775_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .S(fanout_net_41 ), .Z(_04882_ ) );
MUX2_X1 _12776_ ( .A(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ), .B(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ), .S(fanout_net_41 ), .Z(_04883_ ) );
MUX2_X1 _12777_ ( .A(_04882_ ), .B(_04883_ ), .S(fanout_net_45 ), .Z(_04884_ ) );
OAI211_X1 _12778_ ( .A(fanout_net_47 ), .B(_04881_ ), .C1(_04884_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04885_ ) );
AOI21_X1 _12779_ ( .A(_04411_ ), .B1(_04876_ ), .B2(_04885_ ), .ZN(_04886_ ) );
AND2_X1 _12780_ ( .A1(_04411_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_04887_ ) );
NOR2_X2 _12781_ ( .A1(_04886_ ), .A2(_04887_ ), .ZN(_04888_ ) );
XNOR2_X1 _12782_ ( .A(_04888_ ), .B(_02235_ ), .ZN(_04889_ ) );
AND2_X1 _12783_ ( .A1(_04867_ ), .A2(_04889_ ), .ZN(_04890_ ) );
AND4_X1 _12784_ ( .A1(_04559_ ), .A2(_04757_ ), .A3(_04845_ ), .A4(_04890_ ), .ZN(_04891_ ) );
OR3_X1 _12785_ ( .A1(_04328_ ), .A2(\EX_LS_result_reg [10] ), .A3(_04338_ ), .ZN(_04892_ ) );
OR2_X1 _12786_ ( .A1(_04686_ ), .A2(\myreg.Reg[7][10] ), .ZN(_04893_ ) );
OAI211_X1 _12787_ ( .A(_04893_ ), .B(fanout_net_45 ), .C1(fanout_net_41 ), .C2(\myreg.Reg[6][10] ), .ZN(_04894_ ) );
OR2_X1 _12788_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[4][10] ), .ZN(_04895_ ) );
OAI211_X1 _12789_ ( .A(_04895_ ), .B(_04697_ ), .C1(_04687_ ), .C2(\myreg.Reg[5][10] ), .ZN(_04896_ ) );
NAND3_X1 _12790_ ( .A1(_04894_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04896_ ), .ZN(_04897_ ) );
MUX2_X1 _12791_ ( .A(\myreg.Reg[2][10] ), .B(\myreg.Reg[3][10] ), .S(fanout_net_41 ), .Z(_04898_ ) );
MUX2_X1 _12792_ ( .A(\myreg.Reg[0][10] ), .B(\myreg.Reg[1][10] ), .S(fanout_net_41 ), .Z(_04899_ ) );
MUX2_X1 _12793_ ( .A(_04898_ ), .B(_04899_ ), .S(_04697_ ), .Z(_04900_ ) );
OAI211_X1 _12794_ ( .A(_04343_ ), .B(_04897_ ), .C1(_04900_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04901_ ) );
NOR2_X1 _12795_ ( .A1(_04484_ ), .A2(\myreg.Reg[11][10] ), .ZN(_04902_ ) );
OAI21_X1 _12796_ ( .A(fanout_net_45 ), .B1(fanout_net_41 ), .B2(\myreg.Reg[10][10] ), .ZN(_04903_ ) );
NOR2_X1 _12797_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[8][10] ), .ZN(_04904_ ) );
OAI21_X1 _12798_ ( .A(_04697_ ), .B1(_04484_ ), .B2(\myreg.Reg[9][10] ), .ZN(_04905_ ) );
OAI221_X1 _12799_ ( .A(_04354_ ), .B1(_04902_ ), .B2(_04903_ ), .C1(_04904_ ), .C2(_04905_ ), .ZN(_04906_ ) );
MUX2_X1 _12800_ ( .A(\myreg.Reg[12][10] ), .B(\myreg.Reg[13][10] ), .S(fanout_net_41 ), .Z(_04907_ ) );
MUX2_X1 _12801_ ( .A(\myreg.Reg[14][10] ), .B(\myreg.Reg[15][10] ), .S(fanout_net_41 ), .Z(_04908_ ) );
MUX2_X1 _12802_ ( .A(_04907_ ), .B(_04908_ ), .S(fanout_net_45 ), .Z(_04909_ ) );
OAI211_X1 _12803_ ( .A(fanout_net_47 ), .B(_04906_ ), .C1(_04909_ ), .C2(_04355_ ), .ZN(_04910_ ) );
OAI211_X1 _12804_ ( .A(_04901_ ), .B(_04910_ ), .C1(_04560_ ), .C2(_04638_ ), .ZN(_04911_ ) );
NAND2_X1 _12805_ ( .A1(_04892_ ), .A2(_04911_ ), .ZN(_04912_ ) );
XOR2_X1 _12806_ ( .A(_02422_ ), .B(_04912_ ), .Z(_04913_ ) );
OR3_X1 _12807_ ( .A1(_04328_ ), .A2(\EX_LS_result_reg [11] ), .A3(_04338_ ), .ZN(_04914_ ) );
OR2_X1 _12808_ ( .A1(_04686_ ), .A2(\myreg.Reg[5][11] ), .ZN(_04915_ ) );
OAI211_X1 _12809_ ( .A(_04915_ ), .B(_04697_ ), .C1(fanout_net_41 ), .C2(\myreg.Reg[4][11] ), .ZN(_04916_ ) );
OR2_X1 _12810_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[6][11] ), .ZN(_04917_ ) );
OAI211_X1 _12811_ ( .A(_04917_ ), .B(fanout_net_45 ), .C1(_04484_ ), .C2(\myreg.Reg[7][11] ), .ZN(_04918_ ) );
NAND3_X1 _12812_ ( .A1(_04916_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04918_ ), .ZN(_04919_ ) );
MUX2_X1 _12813_ ( .A(\myreg.Reg[2][11] ), .B(\myreg.Reg[3][11] ), .S(fanout_net_41 ), .Z(_04920_ ) );
MUX2_X1 _12814_ ( .A(\myreg.Reg[0][11] ), .B(\myreg.Reg[1][11] ), .S(fanout_net_41 ), .Z(_04921_ ) );
MUX2_X1 _12815_ ( .A(_04920_ ), .B(_04921_ ), .S(_04361_ ), .Z(_04922_ ) );
OAI211_X1 _12816_ ( .A(_04343_ ), .B(_04919_ ), .C1(_04922_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04923_ ) );
NOR2_X1 _12817_ ( .A1(_04589_ ), .A2(\myreg.Reg[11][11] ), .ZN(_04924_ ) );
OAI21_X1 _12818_ ( .A(fanout_net_45 ), .B1(fanout_net_41 ), .B2(\myreg.Reg[10][11] ), .ZN(_04925_ ) );
NOR2_X1 _12819_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[8][11] ), .ZN(_04926_ ) );
OAI21_X1 _12820_ ( .A(_04361_ ), .B1(_04589_ ), .B2(\myreg.Reg[9][11] ), .ZN(_04927_ ) );
OAI221_X1 _12821_ ( .A(_04354_ ), .B1(_04924_ ), .B2(_04925_ ), .C1(_04926_ ), .C2(_04927_ ), .ZN(_04928_ ) );
MUX2_X1 _12822_ ( .A(\myreg.Reg[12][11] ), .B(\myreg.Reg[13][11] ), .S(fanout_net_41 ), .Z(_04929_ ) );
MUX2_X1 _12823_ ( .A(\myreg.Reg[14][11] ), .B(\myreg.Reg[15][11] ), .S(fanout_net_41 ), .Z(_04930_ ) );
MUX2_X1 _12824_ ( .A(_04929_ ), .B(_04930_ ), .S(fanout_net_45 ), .Z(_04931_ ) );
OAI211_X1 _12825_ ( .A(fanout_net_47 ), .B(_04928_ ), .C1(_04931_ ), .C2(_04355_ ), .ZN(_04932_ ) );
OAI211_X1 _12826_ ( .A(_04923_ ), .B(_04932_ ), .C1(_04329_ ), .C2(_04638_ ), .ZN(_04933_ ) );
NAND2_X1 _12827_ ( .A1(_04914_ ), .A2(_04933_ ), .ZN(_04934_ ) );
INV_X1 _12828_ ( .A(_04934_ ), .ZN(_04935_ ) );
XNOR2_X1 _12829_ ( .A(_02399_ ), .B(_04935_ ), .ZN(_04936_ ) );
AND2_X1 _12830_ ( .A1(_04913_ ), .A2(_04936_ ), .ZN(_04937_ ) );
OR2_X1 _12831_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[8][9] ), .ZN(_04938_ ) );
OAI211_X1 _12832_ ( .A(_04938_ ), .B(_04362_ ), .C1(_04485_ ), .C2(\myreg.Reg[9][9] ), .ZN(_04939_ ) );
OR2_X1 _12833_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[10][9] ), .ZN(_04940_ ) );
OAI211_X1 _12834_ ( .A(_04940_ ), .B(fanout_net_45 ), .C1(_04485_ ), .C2(\myreg.Reg[11][9] ), .ZN(_04941_ ) );
NAND3_X1 _12835_ ( .A1(_04939_ ), .A2(_04941_ ), .A3(_04622_ ), .ZN(_04942_ ) );
MUX2_X1 _12836_ ( .A(\myreg.Reg[14][9] ), .B(\myreg.Reg[15][9] ), .S(fanout_net_41 ), .Z(_04943_ ) );
MUX2_X1 _12837_ ( .A(\myreg.Reg[12][9] ), .B(\myreg.Reg[13][9] ), .S(fanout_net_41 ), .Z(_04944_ ) );
MUX2_X1 _12838_ ( .A(_04943_ ), .B(_04944_ ), .S(_04564_ ), .Z(_04945_ ) );
OAI211_X1 _12839_ ( .A(fanout_net_47 ), .B(_04942_ ), .C1(_04945_ ), .C2(_04483_ ), .ZN(_04946_ ) );
MUX2_X1 _12840_ ( .A(\myreg.Reg[2][9] ), .B(\myreg.Reg[3][9] ), .S(fanout_net_41 ), .Z(_04947_ ) );
AND2_X1 _12841_ ( .A1(_04947_ ), .A2(fanout_net_45 ), .ZN(_04948_ ) );
MUX2_X1 _12842_ ( .A(\myreg.Reg[0][9] ), .B(\myreg.Reg[1][9] ), .S(fanout_net_41 ), .Z(_04949_ ) );
AOI211_X1 _12843_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .B(_04948_ ), .C1(_04363_ ), .C2(_04949_ ), .ZN(_04950_ ) );
MUX2_X1 _12844_ ( .A(\myreg.Reg[6][9] ), .B(\myreg.Reg[7][9] ), .S(fanout_net_41 ), .Z(_04951_ ) );
MUX2_X1 _12845_ ( .A(\myreg.Reg[4][9] ), .B(\myreg.Reg[5][9] ), .S(fanout_net_41 ), .Z(_04952_ ) );
MUX2_X1 _12846_ ( .A(_04951_ ), .B(_04952_ ), .S(_04489_ ), .Z(_04953_ ) );
OAI21_X1 _12847_ ( .A(_04562_ ), .B1(_04953_ ), .B2(_04622_ ), .ZN(_04954_ ) );
OAI221_X1 _12848_ ( .A(_04946_ ), .B1(_04950_ ), .B2(_04954_ ), .C1(_04582_ ), .C2(_04583_ ), .ZN(_04955_ ) );
OR3_X1 _12849_ ( .A1(_04560_ ), .A2(\EX_LS_result_reg [9] ), .A3(_04638_ ), .ZN(_04956_ ) );
NAND2_X1 _12850_ ( .A1(_04955_ ), .A2(_04956_ ), .ZN(_04957_ ) );
AND2_X1 _12851_ ( .A1(_02472_ ), .A2(_04957_ ), .ZN(_04958_ ) );
NOR2_X1 _12852_ ( .A1(_02472_ ), .A2(_04957_ ), .ZN(_04959_ ) );
NOR2_X1 _12853_ ( .A1(_04958_ ), .A2(_04959_ ), .ZN(_04960_ ) );
OR3_X1 _12854_ ( .A1(_04582_ ), .A2(\EX_LS_result_reg [8] ), .A3(_04583_ ), .ZN(_04961_ ) );
OR2_X1 _12855_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[0][8] ), .ZN(_04962_ ) );
OAI211_X1 _12856_ ( .A(_04962_ ), .B(_04362_ ), .C1(_04485_ ), .C2(\myreg.Reg[1][8] ), .ZN(_04963_ ) );
OR2_X1 _12857_ ( .A1(fanout_net_41 ), .A2(\myreg.Reg[2][8] ), .ZN(_04964_ ) );
OAI211_X1 _12858_ ( .A(_04964_ ), .B(fanout_net_45 ), .C1(_04485_ ), .C2(\myreg.Reg[3][8] ), .ZN(_04965_ ) );
NAND3_X1 _12859_ ( .A1(_04963_ ), .A2(_04965_ ), .A3(_04483_ ), .ZN(_04966_ ) );
MUX2_X1 _12860_ ( .A(\myreg.Reg[6][8] ), .B(\myreg.Reg[7][8] ), .S(fanout_net_41 ), .Z(_04967_ ) );
MUX2_X1 _12861_ ( .A(\myreg.Reg[4][8] ), .B(\myreg.Reg[5][8] ), .S(fanout_net_41 ), .Z(_04968_ ) );
MUX2_X1 _12862_ ( .A(_04967_ ), .B(_04968_ ), .S(_04362_ ), .Z(_04969_ ) );
OAI211_X1 _12863_ ( .A(_04344_ ), .B(_04966_ ), .C1(_04969_ ), .C2(_04356_ ), .ZN(_04970_ ) );
OR2_X1 _12864_ ( .A1(_04687_ ), .A2(\myreg.Reg[15][8] ), .ZN(_04971_ ) );
OAI211_X1 _12865_ ( .A(_04971_ ), .B(fanout_net_45 ), .C1(fanout_net_42 ), .C2(\myreg.Reg[14][8] ), .ZN(_04972_ ) );
OR2_X1 _12866_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[12][8] ), .ZN(_04973_ ) );
OAI211_X1 _12867_ ( .A(_04973_ ), .B(_04362_ ), .C1(_04485_ ), .C2(\myreg.Reg[13][8] ), .ZN(_04974_ ) );
NAND3_X1 _12868_ ( .A1(_04972_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_04974_ ), .ZN(_04975_ ) );
MUX2_X1 _12869_ ( .A(\myreg.Reg[8][8] ), .B(\myreg.Reg[9][8] ), .S(fanout_net_42 ), .Z(_04976_ ) );
MUX2_X1 _12870_ ( .A(\myreg.Reg[10][8] ), .B(\myreg.Reg[11][8] ), .S(fanout_net_42 ), .Z(_04977_ ) );
MUX2_X1 _12871_ ( .A(_04976_ ), .B(_04977_ ), .S(fanout_net_45 ), .Z(_04978_ ) );
OAI211_X1 _12872_ ( .A(fanout_net_47 ), .B(_04975_ ), .C1(_04978_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04979_ ) );
OAI211_X1 _12873_ ( .A(_04970_ ), .B(_04979_ ), .C1(_04330_ ), .C2(_04340_ ), .ZN(_04980_ ) );
NAND2_X1 _12874_ ( .A1(_04961_ ), .A2(_04980_ ), .ZN(_04981_ ) );
XOR2_X1 _12875_ ( .A(_02448_ ), .B(_04981_ ), .Z(_04982_ ) );
AND3_X1 _12876_ ( .A1(_04937_ ), .A2(_04960_ ), .A3(_04982_ ), .ZN(_04983_ ) );
OR3_X4 _12877_ ( .A1(_04582_ ), .A2(\EX_LS_result_reg [14] ), .A3(_04583_ ), .ZN(_04984_ ) );
OR2_X1 _12878_ ( .A1(_04484_ ), .A2(\myreg.Reg[1][14] ), .ZN(_04985_ ) );
OAI211_X1 _12879_ ( .A(_04985_ ), .B(_04362_ ), .C1(fanout_net_42 ), .C2(\myreg.Reg[0][14] ), .ZN(_04986_ ) );
OR2_X1 _12880_ ( .A1(_04589_ ), .A2(\myreg.Reg[3][14] ), .ZN(_04987_ ) );
OAI211_X1 _12881_ ( .A(_04987_ ), .B(fanout_net_45 ), .C1(fanout_net_42 ), .C2(\myreg.Reg[2][14] ), .ZN(_04988_ ) );
NAND3_X1 _12882_ ( .A1(_04986_ ), .A2(_04988_ ), .A3(_04622_ ), .ZN(_04989_ ) );
MUX2_X1 _12883_ ( .A(\myreg.Reg[6][14] ), .B(\myreg.Reg[7][14] ), .S(fanout_net_42 ), .Z(_04990_ ) );
MUX2_X1 _12884_ ( .A(\myreg.Reg[4][14] ), .B(\myreg.Reg[5][14] ), .S(fanout_net_42 ), .Z(_04991_ ) );
MUX2_X1 _12885_ ( .A(_04990_ ), .B(_04991_ ), .S(_04564_ ), .Z(_04992_ ) );
OAI211_X1 _12886_ ( .A(_04562_ ), .B(_04989_ ), .C1(_04992_ ), .C2(_04483_ ), .ZN(_04993_ ) );
OR2_X1 _12887_ ( .A1(_04484_ ), .A2(\myreg.Reg[15][14] ), .ZN(_04994_ ) );
OAI211_X1 _12888_ ( .A(_04994_ ), .B(fanout_net_45 ), .C1(fanout_net_42 ), .C2(\myreg.Reg[14][14] ), .ZN(_04995_ ) );
OR2_X1 _12889_ ( .A1(_04589_ ), .A2(\myreg.Reg[13][14] ), .ZN(_04996_ ) );
OAI211_X1 _12890_ ( .A(_04996_ ), .B(_04362_ ), .C1(fanout_net_42 ), .C2(\myreg.Reg[12][14] ), .ZN(_04997_ ) );
NAND3_X1 _12891_ ( .A1(_04995_ ), .A2(_04997_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_04998_ ) );
MUX2_X1 _12892_ ( .A(\myreg.Reg[8][14] ), .B(\myreg.Reg[9][14] ), .S(fanout_net_42 ), .Z(_04999_ ) );
MUX2_X1 _12893_ ( .A(\myreg.Reg[10][14] ), .B(\myreg.Reg[11][14] ), .S(fanout_net_42 ), .Z(_05000_ ) );
MUX2_X1 _12894_ ( .A(_04999_ ), .B(_05000_ ), .S(fanout_net_45 ), .Z(_05001_ ) );
OAI211_X1 _12895_ ( .A(fanout_net_47 ), .B(_04998_ ), .C1(_05001_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05002_ ) );
OAI211_X1 _12896_ ( .A(_04993_ ), .B(_05002_ ), .C1(_04330_ ), .C2(_04340_ ), .ZN(_05003_ ) );
NAND2_X1 _12897_ ( .A1(_04984_ ), .A2(_05003_ ), .ZN(_05004_ ) );
XOR2_X1 _12898_ ( .A(_02592_ ), .B(_05004_ ), .Z(_05005_ ) );
OR3_X4 _12899_ ( .A1(_04329_ ), .A2(\EX_LS_result_reg [15] ), .A3(_04339_ ), .ZN(_05006_ ) );
OR2_X1 _12900_ ( .A1(_04686_ ), .A2(\myreg.Reg[9][15] ), .ZN(_05007_ ) );
OAI211_X1 _12901_ ( .A(_05007_ ), .B(_04620_ ), .C1(fanout_net_42 ), .C2(\myreg.Reg[8][15] ), .ZN(_05008_ ) );
OR2_X1 _12902_ ( .A1(_04686_ ), .A2(\myreg.Reg[11][15] ), .ZN(_05009_ ) );
OAI211_X1 _12903_ ( .A(_05009_ ), .B(fanout_net_45 ), .C1(fanout_net_42 ), .C2(\myreg.Reg[10][15] ), .ZN(_05010_ ) );
NAND3_X1 _12904_ ( .A1(_05008_ ), .A2(_05010_ ), .A3(_04482_ ), .ZN(_05011_ ) );
MUX2_X1 _12905_ ( .A(\myreg.Reg[14][15] ), .B(\myreg.Reg[15][15] ), .S(fanout_net_42 ), .Z(_05012_ ) );
MUX2_X1 _12906_ ( .A(\myreg.Reg[12][15] ), .B(\myreg.Reg[13][15] ), .S(fanout_net_42 ), .Z(_05013_ ) );
MUX2_X1 _12907_ ( .A(_05012_ ), .B(_05013_ ), .S(_04697_ ), .Z(_05014_ ) );
OAI211_X1 _12908_ ( .A(fanout_net_47 ), .B(_05011_ ), .C1(_05014_ ), .C2(_04622_ ), .ZN(_05015_ ) );
OR2_X1 _12909_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[0][15] ), .ZN(_05016_ ) );
OAI211_X1 _12910_ ( .A(_05016_ ), .B(_04697_ ), .C1(_04484_ ), .C2(\myreg.Reg[1][15] ), .ZN(_05017_ ) );
NOR2_X1 _12911_ ( .A1(_04613_ ), .A2(\myreg.Reg[3][15] ), .ZN(_05018_ ) );
OAI21_X1 _12912_ ( .A(fanout_net_45 ), .B1(fanout_net_42 ), .B2(\myreg.Reg[2][15] ), .ZN(_05019_ ) );
OAI211_X1 _12913_ ( .A(_05017_ ), .B(_04354_ ), .C1(_05018_ ), .C2(_05019_ ), .ZN(_05020_ ) );
MUX2_X1 _12914_ ( .A(\myreg.Reg[6][15] ), .B(\myreg.Reg[7][15] ), .S(fanout_net_42 ), .Z(_05021_ ) );
MUX2_X1 _12915_ ( .A(\myreg.Reg[4][15] ), .B(\myreg.Reg[5][15] ), .S(fanout_net_42 ), .Z(_05022_ ) );
MUX2_X1 _12916_ ( .A(_05021_ ), .B(_05022_ ), .S(_04697_ ), .Z(_05023_ ) );
OAI211_X1 _12917_ ( .A(_04343_ ), .B(_05020_ ), .C1(_05023_ ), .C2(_04355_ ), .ZN(_05024_ ) );
OAI211_X1 _12918_ ( .A(_05015_ ), .B(_05024_ ), .C1(_04560_ ), .C2(_04638_ ), .ZN(_05025_ ) );
NAND2_X1 _12919_ ( .A1(_05006_ ), .A2(_05025_ ), .ZN(_05026_ ) );
INV_X1 _12920_ ( .A(_05026_ ), .ZN(_05027_ ) );
XNOR2_X1 _12921_ ( .A(_02518_ ), .B(_05027_ ), .ZN(_05028_ ) );
AND2_X1 _12922_ ( .A1(_05005_ ), .A2(_05028_ ), .ZN(_05029_ ) );
OR3_X1 _12923_ ( .A1(_04560_ ), .A2(\EX_LS_result_reg [12] ), .A3(_04638_ ), .ZN(_05030_ ) );
OR2_X1 _12924_ ( .A1(_04589_ ), .A2(\myreg.Reg[1][12] ), .ZN(_05031_ ) );
OAI211_X1 _12925_ ( .A(_05031_ ), .B(_04564_ ), .C1(fanout_net_42 ), .C2(\myreg.Reg[0][12] ), .ZN(_05032_ ) );
OR2_X1 _12926_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[2][12] ), .ZN(_05033_ ) );
OAI211_X1 _12927_ ( .A(_05033_ ), .B(fanout_net_45 ), .C1(_04348_ ), .C2(\myreg.Reg[3][12] ), .ZN(_05034_ ) );
NAND3_X1 _12928_ ( .A1(_05032_ ), .A2(_04355_ ), .A3(_05034_ ), .ZN(_05035_ ) );
MUX2_X1 _12929_ ( .A(\myreg.Reg[6][12] ), .B(\myreg.Reg[7][12] ), .S(fanout_net_42 ), .Z(_05036_ ) );
MUX2_X1 _12930_ ( .A(\myreg.Reg[4][12] ), .B(\myreg.Reg[5][12] ), .S(fanout_net_42 ), .Z(_05037_ ) );
MUX2_X1 _12931_ ( .A(_05036_ ), .B(_05037_ ), .S(_04564_ ), .Z(_05038_ ) );
OAI211_X1 _12932_ ( .A(_04562_ ), .B(_05035_ ), .C1(_05038_ ), .C2(_04483_ ), .ZN(_05039_ ) );
OR2_X1 _12933_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[14][12] ), .ZN(_05040_ ) );
OAI211_X1 _12934_ ( .A(_05040_ ), .B(fanout_net_45 ), .C1(_04348_ ), .C2(\myreg.Reg[15][12] ), .ZN(_05041_ ) );
OR2_X1 _12935_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[12][12] ), .ZN(_05042_ ) );
OAI211_X1 _12936_ ( .A(_05042_ ), .B(_04564_ ), .C1(_04348_ ), .C2(\myreg.Reg[13][12] ), .ZN(_05043_ ) );
NAND3_X1 _12937_ ( .A1(_05041_ ), .A2(_05043_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05044_ ) );
MUX2_X1 _12938_ ( .A(\myreg.Reg[8][12] ), .B(\myreg.Reg[9][12] ), .S(fanout_net_42 ), .Z(_05045_ ) );
MUX2_X1 _12939_ ( .A(\myreg.Reg[10][12] ), .B(\myreg.Reg[11][12] ), .S(fanout_net_42 ), .Z(_05046_ ) );
MUX2_X1 _12940_ ( .A(_05045_ ), .B(_05046_ ), .S(fanout_net_45 ), .Z(_05047_ ) );
OAI211_X1 _12941_ ( .A(fanout_net_47 ), .B(_05044_ ), .C1(_05047_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05048_ ) );
OAI211_X1 _12942_ ( .A(_05039_ ), .B(_05048_ ), .C1(_04582_ ), .C2(_04583_ ), .ZN(_05049_ ) );
NAND2_X1 _12943_ ( .A1(_05030_ ), .A2(_05049_ ), .ZN(_05050_ ) );
XOR2_X1 _12944_ ( .A(_02588_ ), .B(_05050_ ), .Z(_05051_ ) );
OR3_X1 _12945_ ( .A1(_04328_ ), .A2(\EX_LS_result_reg [13] ), .A3(_04338_ ), .ZN(_05052_ ) );
OR2_X1 _12946_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[8][13] ), .ZN(_05053_ ) );
OAI211_X1 _12947_ ( .A(_05053_ ), .B(_04697_ ), .C1(_04687_ ), .C2(\myreg.Reg[9][13] ), .ZN(_05054_ ) );
OR2_X1 _12948_ ( .A1(fanout_net_42 ), .A2(\myreg.Reg[10][13] ), .ZN(_05055_ ) );
OAI211_X1 _12949_ ( .A(_05055_ ), .B(fanout_net_45 ), .C1(_04484_ ), .C2(\myreg.Reg[11][13] ), .ZN(_05056_ ) );
NAND3_X1 _12950_ ( .A1(_05054_ ), .A2(_05056_ ), .A3(_04354_ ), .ZN(_05057_ ) );
MUX2_X1 _12951_ ( .A(\myreg.Reg[14][13] ), .B(\myreg.Reg[15][13] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05058_ ) );
MUX2_X1 _12952_ ( .A(\myreg.Reg[12][13] ), .B(\myreg.Reg[13][13] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05059_ ) );
MUX2_X1 _12953_ ( .A(_05058_ ), .B(_05059_ ), .S(_04361_ ), .Z(_05060_ ) );
OAI211_X1 _12954_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05057_ ), .C1(_05060_ ), .C2(_04355_ ), .ZN(_05061_ ) );
OR2_X1 _12955_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[0][13] ), .ZN(_05062_ ) );
OAI211_X1 _12956_ ( .A(_05062_ ), .B(_04361_ ), .C1(_04589_ ), .C2(\myreg.Reg[1][13] ), .ZN(_05063_ ) );
NOR2_X1 _12957_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[2][13] ), .ZN(_05064_ ) );
OAI21_X1 _12958_ ( .A(fanout_net_45 ), .B1(_04589_ ), .B2(\myreg.Reg[3][13] ), .ZN(_05065_ ) );
OAI211_X1 _12959_ ( .A(_05063_ ), .B(_04354_ ), .C1(_05064_ ), .C2(_05065_ ), .ZN(_05066_ ) );
MUX2_X1 _12960_ ( .A(\myreg.Reg[6][13] ), .B(\myreg.Reg[7][13] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05067_ ) );
MUX2_X1 _12961_ ( .A(\myreg.Reg[4][13] ), .B(\myreg.Reg[5][13] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05068_ ) );
MUX2_X1 _12962_ ( .A(_05067_ ), .B(_05068_ ), .S(_04361_ ), .Z(_05069_ ) );
OAI211_X1 _12963_ ( .A(_04343_ ), .B(_05066_ ), .C1(_05069_ ), .C2(_04355_ ), .ZN(_05070_ ) );
OAI211_X1 _12964_ ( .A(_05061_ ), .B(_05070_ ), .C1(_04560_ ), .C2(_04638_ ), .ZN(_05071_ ) );
NAND2_X1 _12965_ ( .A1(_05052_ ), .A2(_05071_ ), .ZN(_05072_ ) );
AND2_X1 _12966_ ( .A1(_02565_ ), .A2(_05072_ ), .ZN(_05073_ ) );
NOR2_X1 _12967_ ( .A1(_02565_ ), .A2(_05072_ ), .ZN(_05074_ ) );
NOR2_X1 _12968_ ( .A1(_05073_ ), .A2(_05074_ ), .ZN(_05075_ ) );
AND2_X1 _12969_ ( .A1(_05051_ ), .A2(_05075_ ), .ZN(_05076_ ) );
AND2_X1 _12970_ ( .A1(_05029_ ), .A2(_05076_ ), .ZN(_05077_ ) );
AND2_X1 _12971_ ( .A1(_04983_ ), .A2(_05077_ ), .ZN(_05078_ ) );
OR3_X4 _12972_ ( .A1(_04327_ ), .A2(\EX_LS_result_reg [1] ), .A3(_04337_ ), .ZN(_05079_ ) );
OR2_X1 _12973_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[0][1] ), .ZN(_05080_ ) );
OAI211_X1 _12974_ ( .A(_05080_ ), .B(_04359_ ), .C1(_04346_ ), .C2(\myreg.Reg[1][1] ), .ZN(_05081_ ) );
OR2_X1 _12975_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[2][1] ), .ZN(_05082_ ) );
OAI211_X1 _12976_ ( .A(_05082_ ), .B(fanout_net_45 ), .C1(_04345_ ), .C2(\myreg.Reg[3][1] ), .ZN(_05083_ ) );
NAND3_X1 _12977_ ( .A1(_05081_ ), .A2(_05083_ ), .A3(_04353_ ), .ZN(_05084_ ) );
MUX2_X1 _12978_ ( .A(\myreg.Reg[6][1] ), .B(\myreg.Reg[7][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05085_ ) );
MUX2_X1 _12979_ ( .A(\myreg.Reg[4][1] ), .B(\myreg.Reg[5][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05086_ ) );
MUX2_X1 _12980_ ( .A(_05085_ ), .B(_05086_ ), .S(_04359_ ), .Z(_05087_ ) );
OAI211_X1 _12981_ ( .A(_04342_ ), .B(_05084_ ), .C1(_05087_ ), .C2(_04353_ ), .ZN(_05088_ ) );
OR2_X1 _12982_ ( .A1(_04345_ ), .A2(\myreg.Reg[13][1] ), .ZN(_05089_ ) );
OAI211_X1 _12983_ ( .A(_05089_ ), .B(_04359_ ), .C1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .C2(\myreg.Reg[12][1] ), .ZN(_05090_ ) );
OR2_X1 _12984_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[14][1] ), .ZN(_05091_ ) );
OAI211_X1 _12985_ ( .A(_05091_ ), .B(fanout_net_45 ), .C1(_04345_ ), .C2(\myreg.Reg[15][1] ), .ZN(_05092_ ) );
NAND3_X1 _12986_ ( .A1(_05090_ ), .A2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .A3(_05092_ ), .ZN(_05093_ ) );
MUX2_X1 _12987_ ( .A(\myreg.Reg[8][1] ), .B(\myreg.Reg[9][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05094_ ) );
MUX2_X1 _12988_ ( .A(\myreg.Reg[10][1] ), .B(\myreg.Reg[11][1] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05095_ ) );
MUX2_X1 _12989_ ( .A(_05094_ ), .B(_05095_ ), .S(fanout_net_45 ), .Z(_05096_ ) );
OAI211_X1 _12990_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05093_ ), .C1(_05096_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05097_ ) );
OAI211_X1 _12991_ ( .A(_05088_ ), .B(_05097_ ), .C1(_04327_ ), .C2(_04337_ ), .ZN(_05098_ ) );
NAND2_X2 _12992_ ( .A1(_05079_ ), .A2(_05098_ ), .ZN(_05099_ ) );
XOR2_X1 _12993_ ( .A(_02282_ ), .B(_05099_ ), .Z(_05100_ ) );
OR3_X4 _12994_ ( .A1(_04327_ ), .A2(\EX_LS_result_reg [0] ), .A3(_04337_ ), .ZN(_05101_ ) );
OR2_X1 _12995_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[4][0] ), .ZN(_05102_ ) );
OAI211_X1 _12996_ ( .A(_05102_ ), .B(_04359_ ), .C1(_04345_ ), .C2(\myreg.Reg[5][0] ), .ZN(_05103_ ) );
OR2_X1 _12997_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[6][0] ), .ZN(_05104_ ) );
OAI211_X1 _12998_ ( .A(_05104_ ), .B(fanout_net_45 ), .C1(_04345_ ), .C2(\myreg.Reg[7][0] ), .ZN(_05105_ ) );
NAND3_X1 _12999_ ( .A1(_05103_ ), .A2(_05105_ ), .A3(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05106_ ) );
MUX2_X1 _13000_ ( .A(\myreg.Reg[2][0] ), .B(\myreg.Reg[3][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05107_ ) );
MUX2_X1 _13001_ ( .A(\myreg.Reg[0][0] ), .B(\myreg.Reg[1][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05108_ ) );
MUX2_X1 _13002_ ( .A(_05107_ ), .B(_05108_ ), .S(_04359_ ), .Z(_05109_ ) );
OAI211_X1 _13003_ ( .A(_04342_ ), .B(_05106_ ), .C1(_05109_ ), .C2(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .ZN(_05110_ ) );
NOR2_X1 _13004_ ( .A1(_04345_ ), .A2(\myreg.Reg[11][0] ), .ZN(_05111_ ) );
OAI21_X1 _13005_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .B1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .B2(\myreg.Reg[10][0] ), .ZN(_05112_ ) );
NOR2_X1 _13006_ ( .A1(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .A2(\myreg.Reg[8][0] ), .ZN(_05113_ ) );
OAI21_X1 _13007_ ( .A(_04358_ ), .B1(_04345_ ), .B2(\myreg.Reg[9][0] ), .ZN(_05114_ ) );
OAI221_X1 _13008_ ( .A(_04352_ ), .B1(_05111_ ), .B2(_05112_ ), .C1(_05113_ ), .C2(_05114_ ), .ZN(_05115_ ) );
MUX2_X1 _13009_ ( .A(\myreg.Reg[12][0] ), .B(\myreg.Reg[13][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05116_ ) );
MUX2_X1 _13010_ ( .A(\myreg.Reg[14][0] ), .B(\myreg.Reg[15][0] ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(_05117_ ) );
MUX2_X1 _13011_ ( .A(_05116_ ), .B(_05117_ ), .S(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(_05118_ ) );
OAI211_X1 _13012_ ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .B(_05115_ ), .C1(_05118_ ), .C2(_04353_ ), .ZN(_05119_ ) );
OAI211_X1 _13013_ ( .A(_05110_ ), .B(_05119_ ), .C1(_04327_ ), .C2(_04337_ ), .ZN(_05120_ ) );
NAND2_X2 _13014_ ( .A1(_05101_ ), .A2(_05120_ ), .ZN(_05121_ ) );
OR2_X1 _13015_ ( .A1(_04110_ ), .A2(_05121_ ), .ZN(_05122_ ) );
NAND2_X1 _13016_ ( .A1(_05100_ ), .A2(_05122_ ), .ZN(_05123_ ) );
AOI21_X1 _13017_ ( .A(_05123_ ), .B1(_04110_ ), .B2(_05121_ ), .ZN(_05124_ ) );
AND3_X1 _13018_ ( .A1(_04891_ ), .A2(_05078_ ), .A3(_05124_ ), .ZN(_05125_ ) );
INV_X1 _13019_ ( .A(fanout_net_8 ), .ZN(_05126_ ) );
NOR2_X1 _13020_ ( .A1(_05126_ ), .A2(\ID_EX_typ [1] ), .ZN(_05127_ ) );
AND2_X2 _13021_ ( .A1(_05127_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05128_ ) );
INV_X1 _13022_ ( .A(_05128_ ), .ZN(_05129_ ) );
INV_X1 _13023_ ( .A(fanout_net_11 ), .ZN(_05130_ ) );
BUF_X4 _13024_ ( .A(_05130_ ), .Z(_05131_ ) );
BUF_X2 _13025_ ( .A(_05131_ ), .Z(_05132_ ) );
BUF_X2 _13026_ ( .A(_05132_ ), .Z(_05133_ ) );
NAND2_X1 _13027_ ( .A1(_04384_ ), .A2(_05133_ ), .ZN(_05134_ ) );
NAND2_X1 _13028_ ( .A1(_02939_ ), .A2(fanout_net_11 ), .ZN(_05135_ ) );
NAND2_X1 _13029_ ( .A1(_05134_ ), .A2(_05135_ ), .ZN(_05136_ ) );
INV_X1 _13030_ ( .A(_02909_ ), .ZN(_05137_ ) );
XNOR2_X1 _13031_ ( .A(_05136_ ), .B(_05137_ ), .ZN(_05138_ ) );
NAND3_X1 _13032_ ( .A1(_04386_ ), .A2(_05133_ ), .A3(_04407_ ), .ZN(_05139_ ) );
NAND2_X1 _13033_ ( .A1(fanout_net_11 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_1_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05140_ ) );
AND2_X2 _13034_ ( .A1(_05139_ ), .A2(_05140_ ), .ZN(_05141_ ) );
OR3_X1 _13035_ ( .A1(_05138_ ), .A2(_02937_ ), .A3(_05141_ ), .ZN(_05142_ ) );
OAI21_X1 _13036_ ( .A(_05142_ ), .B1(_05137_ ), .B2(_05136_ ), .ZN(_05143_ ) );
NAND3_X1 _13037_ ( .A1(_04434_ ), .A2(_05133_ ), .A3(_04453_ ), .ZN(_05144_ ) );
NAND2_X1 _13038_ ( .A1(fanout_net_11 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B ), .ZN(_05145_ ) );
AND2_X2 _13039_ ( .A1(_05144_ ), .A2(_05145_ ), .ZN(_05146_ ) );
XNOR2_X1 _13040_ ( .A(_05146_ ), .B(_02962_ ), .ZN(_05147_ ) );
NAND2_X1 _13041_ ( .A1(_04432_ ), .A2(_05133_ ), .ZN(_05148_ ) );
OR2_X1 _13042_ ( .A1(_05133_ ), .A2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_05149_ ) );
AOI21_X1 _13043_ ( .A(_02987_ ), .B1(_05148_ ), .B2(_05149_ ), .ZN(_05150_ ) );
AND3_X1 _13044_ ( .A1(_05148_ ), .A2(_02987_ ), .A3(_05149_ ), .ZN(_05151_ ) );
NOR3_X1 _13045_ ( .A1(_05147_ ), .A2(_05150_ ), .A3(_05151_ ), .ZN(_05152_ ) );
AND2_X1 _13046_ ( .A1(_05143_ ), .A2(_05152_ ), .ZN(_05153_ ) );
INV_X1 _13047_ ( .A(_05153_ ), .ZN(_05154_ ) );
NOR2_X1 _13048_ ( .A1(_05151_ ), .A2(_05150_ ), .ZN(_05155_ ) );
NOR2_X1 _13049_ ( .A1(_05146_ ), .A2(_02962_ ), .ZN(_05156_ ) );
NAND2_X1 _13050_ ( .A1(_05155_ ), .A2(_05156_ ), .ZN(_05157_ ) );
NAND2_X1 _13051_ ( .A1(_05148_ ), .A2(_05149_ ), .ZN(_05158_ ) );
INV_X1 _13052_ ( .A(_05158_ ), .ZN(_05159_ ) );
OAI211_X1 _13053_ ( .A(_05154_ ), .B(_05157_ ), .C1(_02988_ ), .C2(_05159_ ), .ZN(_05160_ ) );
BUF_X4 _13054_ ( .A(_05131_ ), .Z(_05161_ ) );
NAND2_X1 _13055_ ( .A1(_04608_ ), .A2(_05161_ ), .ZN(_05162_ ) );
OR2_X1 _13056_ ( .A1(_05131_ ), .A2(\ID_EX_imm [23] ), .ZN(_05163_ ) );
NAND2_X2 _13057_ ( .A1(_05162_ ), .A2(_05163_ ), .ZN(_05164_ ) );
NOR2_X1 _13058_ ( .A1(_05164_ ), .A2(_02806_ ), .ZN(_05165_ ) );
AOI21_X1 _13059_ ( .A(_02726_ ), .B1(_05162_ ), .B2(_05163_ ), .ZN(_05166_ ) );
NOR2_X2 _13060_ ( .A1(_05165_ ), .A2(_05166_ ), .ZN(_05167_ ) );
INV_X1 _13061_ ( .A(_02748_ ), .ZN(_05168_ ) );
NAND3_X1 _13062_ ( .A1(_04561_ ), .A2(_05161_ ), .A3(_04584_ ), .ZN(_05169_ ) );
NAND2_X1 _13063_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [22] ), .ZN(_05170_ ) );
AND2_X4 _13064_ ( .A1(_05169_ ), .A2(_05170_ ), .ZN(_05171_ ) );
INV_X1 _13065_ ( .A(_05171_ ), .ZN(_05172_ ) );
NOR3_X1 _13066_ ( .A1(_05167_ ), .A2(_05168_ ), .A3(_05172_ ), .ZN(_05173_ ) );
XNOR2_X1 _13067_ ( .A(_05171_ ), .B(_02748_ ), .ZN(_05174_ ) );
NOR2_X2 _13068_ ( .A1(_05167_ ), .A2(_05174_ ), .ZN(_05175_ ) );
NAND3_X1 _13069_ ( .A1(_04639_ ), .A2(_05132_ ), .A3(_04658_ ), .ZN(_05176_ ) );
NAND2_X1 _13070_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [20] ), .ZN(_05177_ ) );
AND2_X2 _13071_ ( .A1(_05176_ ), .A2(_05177_ ), .ZN(_05178_ ) );
XNOR2_X1 _13072_ ( .A(_05178_ ), .B(_02770_ ), .ZN(_05179_ ) );
INV_X1 _13073_ ( .A(_05179_ ), .ZN(_05180_ ) );
NAND3_X1 _13074_ ( .A1(_04611_ ), .A2(_05161_ ), .A3(_04633_ ), .ZN(_05181_ ) );
NAND2_X1 _13075_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [21] ), .ZN(_05182_ ) );
AND2_X4 _13076_ ( .A1(_05181_ ), .A2(_05182_ ), .ZN(_05183_ ) );
XNOR2_X1 _13077_ ( .A(_05183_ ), .B(_02793_ ), .ZN(_05184_ ) );
INV_X1 _13078_ ( .A(_05184_ ), .ZN(_05185_ ) );
AND3_X2 _13079_ ( .A1(_05175_ ), .A2(_05180_ ), .A3(_05185_ ), .ZN(_05186_ ) );
NAND3_X1 _13080_ ( .A1(_04662_ ), .A2(_05161_ ), .A3(_04681_ ), .ZN(_05187_ ) );
NAND2_X1 _13081_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [18] ), .ZN(_05188_ ) );
AND2_X1 _13082_ ( .A1(_05187_ ), .A2(_05188_ ), .ZN(_05189_ ) );
XNOR2_X1 _13083_ ( .A(_05189_ ), .B(_02642_ ), .ZN(_05190_ ) );
NAND3_X1 _13084_ ( .A1(_04684_ ), .A2(_05161_ ), .A3(_04706_ ), .ZN(_05191_ ) );
NAND2_X1 _13085_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [19] ), .ZN(_05192_ ) );
AND2_X1 _13086_ ( .A1(_05191_ ), .A2(_05192_ ), .ZN(_05193_ ) );
XNOR2_X2 _13087_ ( .A(_05193_ ), .B(_02618_ ), .ZN(_05194_ ) );
NOR2_X2 _13088_ ( .A1(_05190_ ), .A2(_05194_ ), .ZN(_05195_ ) );
NAND3_X1 _13089_ ( .A1(_04711_ ), .A2(_05161_ ), .A3(_04730_ ), .ZN(_05196_ ) );
NAND2_X1 _13090_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [17] ), .ZN(_05197_ ) );
AND2_X1 _13091_ ( .A1(_05196_ ), .A2(_05197_ ), .ZN(_05198_ ) );
XNOR2_X1 _13092_ ( .A(_05198_ ), .B(_02688_ ), .ZN(_05199_ ) );
INV_X1 _13093_ ( .A(_02665_ ), .ZN(_05200_ ) );
NAND3_X1 _13094_ ( .A1(_04733_ ), .A2(_04752_ ), .A3(_05132_ ), .ZN(_05201_ ) );
NAND2_X1 _13095_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [16] ), .ZN(_05202_ ) );
AND2_X2 _13096_ ( .A1(_05201_ ), .A2(_05202_ ), .ZN(_05203_ ) );
INV_X1 _13097_ ( .A(_05203_ ), .ZN(_05204_ ) );
NOR3_X1 _13098_ ( .A1(_05199_ ), .A2(_05200_ ), .A3(_05204_ ), .ZN(_05205_ ) );
AND3_X1 _13099_ ( .A1(_02688_ ), .A2(_05197_ ), .A3(_05196_ ), .ZN(_05206_ ) );
OAI21_X1 _13100_ ( .A(_05195_ ), .B1(_05205_ ), .B2(_05206_ ), .ZN(_05207_ ) );
NAND3_X1 _13101_ ( .A1(_02618_ ), .A2(_05192_ ), .A3(_05191_ ), .ZN(_05208_ ) );
NAND2_X1 _13102_ ( .A1(_05207_ ), .A2(_05208_ ), .ZN(_05209_ ) );
INV_X1 _13103_ ( .A(_02642_ ), .ZN(_05210_ ) );
INV_X1 _13104_ ( .A(_05189_ ), .ZN(_05211_ ) );
NOR3_X1 _13105_ ( .A1(_05194_ ), .A2(_05210_ ), .A3(_05211_ ), .ZN(_05212_ ) );
OAI21_X2 _13106_ ( .A(_05186_ ), .B1(_05209_ ), .B2(_05212_ ), .ZN(_05213_ ) );
AND3_X1 _13107_ ( .A1(_05185_ ), .A2(_02770_ ), .A3(_05178_ ), .ZN(_05214_ ) );
AND3_X1 _13108_ ( .A1(_02793_ ), .A2(_05182_ ), .A3(_05181_ ), .ZN(_05215_ ) );
OAI21_X1 _13109_ ( .A(_05175_ ), .B1(_05214_ ), .B2(_05215_ ), .ZN(_05216_ ) );
INV_X1 _13110_ ( .A(_05164_ ), .ZN(_05217_ ) );
OAI211_X1 _13111_ ( .A(_05213_ ), .B(_05216_ ), .C1(_02806_ ), .C2(_05217_ ), .ZN(_05218_ ) );
NAND3_X1 _13112_ ( .A1(_04984_ ), .A2(_05132_ ), .A3(_05003_ ), .ZN(_05219_ ) );
NAND2_X1 _13113_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [14] ), .ZN(_05220_ ) );
AND2_X2 _13114_ ( .A1(_05219_ ), .A2(_05220_ ), .ZN(_05221_ ) );
XNOR2_X2 _13115_ ( .A(_05221_ ), .B(_02592_ ), .ZN(_05222_ ) );
NAND3_X1 _13116_ ( .A1(_05006_ ), .A2(_05161_ ), .A3(_05025_ ), .ZN(_05223_ ) );
NAND2_X1 _13117_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [15] ), .ZN(_05224_ ) );
AND2_X4 _13118_ ( .A1(_05223_ ), .A2(_05224_ ), .ZN(_05225_ ) );
XNOR2_X1 _13119_ ( .A(_05225_ ), .B(_02518_ ), .ZN(_05226_ ) );
NOR2_X2 _13120_ ( .A1(_05222_ ), .A2(_05226_ ), .ZN(_05227_ ) );
INV_X1 _13121_ ( .A(_05227_ ), .ZN(_05228_ ) );
NAND3_X1 _13122_ ( .A1(_05052_ ), .A2(_05131_ ), .A3(_05071_ ), .ZN(_05229_ ) );
NAND2_X1 _13123_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [13] ), .ZN(_05230_ ) );
NAND2_X1 _13124_ ( .A1(_05229_ ), .A2(_05230_ ), .ZN(_05231_ ) );
AND2_X1 _13125_ ( .A1(_05231_ ), .A2(_02565_ ), .ZN(_05232_ ) );
NOR2_X1 _13126_ ( .A1(_05231_ ), .A2(_02565_ ), .ZN(_05233_ ) );
NOR2_X4 _13127_ ( .A1(_05232_ ), .A2(_05233_ ), .ZN(_05234_ ) );
NAND3_X1 _13128_ ( .A1(_05030_ ), .A2(_05132_ ), .A3(_05049_ ), .ZN(_05235_ ) );
NAND2_X1 _13129_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [12] ), .ZN(_05236_ ) );
AND2_X1 _13130_ ( .A1(_05235_ ), .A2(_05236_ ), .ZN(_05237_ ) );
XNOR2_X1 _13131_ ( .A(_05237_ ), .B(_02588_ ), .ZN(_05238_ ) );
NOR3_X2 _13132_ ( .A1(_05228_ ), .A2(_05234_ ), .A3(_05238_ ), .ZN(_05239_ ) );
NAND3_X1 _13133_ ( .A1(_04892_ ), .A2(_04911_ ), .A3(_05131_ ), .ZN(_05240_ ) );
NAND2_X1 _13134_ ( .A1(\ID_EX_imm [10] ), .A2(fanout_net_11 ), .ZN(_05241_ ) );
AND2_X1 _13135_ ( .A1(_05240_ ), .A2(_05241_ ), .ZN(_05242_ ) );
XNOR2_X1 _13136_ ( .A(_05242_ ), .B(_02422_ ), .ZN(_05243_ ) );
NAND3_X1 _13137_ ( .A1(_04914_ ), .A2(_05131_ ), .A3(_04933_ ), .ZN(_05244_ ) );
NAND2_X1 _13138_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [11] ), .ZN(_05245_ ) );
AND2_X2 _13139_ ( .A1(_05244_ ), .A2(_05245_ ), .ZN(_05246_ ) );
XNOR2_X2 _13140_ ( .A(_05246_ ), .B(_02399_ ), .ZN(_05247_ ) );
NOR2_X1 _13141_ ( .A1(_05243_ ), .A2(_05247_ ), .ZN(_05248_ ) );
NAND3_X1 _13142_ ( .A1(_04955_ ), .A2(_04956_ ), .A3(_05132_ ), .ZN(_05249_ ) );
NAND2_X1 _13143_ ( .A1(\ID_EX_imm [9] ), .A2(fanout_net_11 ), .ZN(_05250_ ) );
AND2_X4 _13144_ ( .A1(_05249_ ), .A2(_05250_ ), .ZN(_05251_ ) );
XNOR2_X1 _13145_ ( .A(_05251_ ), .B(_02472_ ), .ZN(_05252_ ) );
INV_X1 _13146_ ( .A(_05252_ ), .ZN(_05253_ ) );
NAND3_X1 _13147_ ( .A1(_04961_ ), .A2(_05132_ ), .A3(_04980_ ), .ZN(_05254_ ) );
NAND2_X1 _13148_ ( .A1(\ID_EX_imm [8] ), .A2(fanout_net_11 ), .ZN(_05255_ ) );
AND2_X1 _13149_ ( .A1(_05254_ ), .A2(_05255_ ), .ZN(_05256_ ) );
XNOR2_X1 _13150_ ( .A(_05256_ ), .B(_02448_ ), .ZN(_05257_ ) );
INV_X1 _13151_ ( .A(_05257_ ), .ZN(_05258_ ) );
AND3_X1 _13152_ ( .A1(_05248_ ), .A2(_05253_ ), .A3(_05258_ ), .ZN(_05259_ ) );
NAND2_X1 _13153_ ( .A1(_04888_ ), .A2(_05131_ ), .ZN(_05260_ ) );
NAND2_X1 _13154_ ( .A1(_02236_ ), .A2(fanout_net_11 ), .ZN(_05261_ ) );
NAND2_X2 _13155_ ( .A1(_05260_ ), .A2(_05261_ ), .ZN(_05262_ ) );
XNOR2_X1 _13156_ ( .A(_05262_ ), .B(_02315_ ), .ZN(_05263_ ) );
NAND3_X1 _13157_ ( .A1(_04846_ ), .A2(_05131_ ), .A3(_04865_ ), .ZN(_05264_ ) );
NAND2_X1 _13158_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [2] ), .ZN(_05265_ ) );
AND2_X1 _13159_ ( .A1(_05264_ ), .A2(_05265_ ), .ZN(_05266_ ) );
BUF_X4 _13160_ ( .A(_05266_ ), .Z(_05267_ ) );
XNOR2_X1 _13161_ ( .A(_05267_ ), .B(_02258_ ), .ZN(_05268_ ) );
NAND2_X1 _13162_ ( .A1(_05099_ ), .A2(_05131_ ), .ZN(_05269_ ) );
NAND2_X1 _13163_ ( .A1(_02285_ ), .A2(fanout_net_11 ), .ZN(_05270_ ) );
NAND2_X2 _13164_ ( .A1(_05269_ ), .A2(_05270_ ), .ZN(_05271_ ) );
XNOR2_X1 _13165_ ( .A(_05271_ ), .B(_02282_ ), .ZN(_05272_ ) );
NAND2_X2 _13166_ ( .A1(_05121_ ), .A2(_05130_ ), .ZN(_05273_ ) );
OR2_X1 _13167_ ( .A1(_05130_ ), .A2(\ID_EX_imm [0] ), .ZN(_05274_ ) );
NAND2_X4 _13168_ ( .A1(_05273_ ), .A2(_05274_ ), .ZN(_05275_ ) );
NOR2_X1 _13169_ ( .A1(_05275_ ), .A2(_04110_ ), .ZN(_05276_ ) );
OR2_X1 _13170_ ( .A1(_05272_ ), .A2(_05276_ ), .ZN(_05277_ ) );
NAND2_X1 _13171_ ( .A1(_05271_ ), .A2(_02282_ ), .ZN(_05278_ ) );
AOI211_X1 _13172_ ( .A(_05263_ ), .B(_05268_ ), .C1(_05277_ ), .C2(_05278_ ), .ZN(_05279_ ) );
AND3_X1 _13173_ ( .A1(_05260_ ), .A2(_02235_ ), .A3(_05261_ ), .ZN(_05280_ ) );
INV_X1 _13174_ ( .A(_02258_ ), .ZN(_05281_ ) );
INV_X1 _13175_ ( .A(_05267_ ), .ZN(_05282_ ) );
NOR3_X1 _13176_ ( .A1(_05263_ ), .A2(_05281_ ), .A3(_05282_ ), .ZN(_05283_ ) );
OR3_X1 _13177_ ( .A1(_05279_ ), .A2(_05280_ ), .A3(_05283_ ), .ZN(_05284_ ) );
NAND3_X1 _13178_ ( .A1(_04820_ ), .A2(_04821_ ), .A3(_05132_ ), .ZN(_05285_ ) );
NAND2_X1 _13179_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [4] ), .ZN(_05286_ ) );
AND2_X2 _13180_ ( .A1(_05285_ ), .A2(_05286_ ), .ZN(_05287_ ) );
XNOR2_X1 _13181_ ( .A(_05287_ ), .B(_02319_ ), .ZN(_05288_ ) );
NAND2_X1 _13182_ ( .A1(_04843_ ), .A2(_05161_ ), .ZN(_05289_ ) );
OR2_X1 _13183_ ( .A1(_05131_ ), .A2(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_05290_ ) );
NAND2_X4 _13184_ ( .A1(_05289_ ), .A2(_05290_ ), .ZN(_05291_ ) );
XNOR2_X1 _13185_ ( .A(_05291_ ), .B(_02213_ ), .ZN(_05292_ ) );
NAND3_X1 _13186_ ( .A1(_04780_ ), .A2(_05161_ ), .A3(_04799_ ), .ZN(_05293_ ) );
NAND2_X1 _13187_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [7] ), .ZN(_05294_ ) );
AND2_X4 _13188_ ( .A1(_05293_ ), .A2(_05294_ ), .ZN(_05295_ ) );
XNOR2_X1 _13189_ ( .A(_05295_ ), .B(_02345_ ), .ZN(_05296_ ) );
NAND3_X1 _13190_ ( .A1(_04758_ ), .A2(_04777_ ), .A3(_05161_ ), .ZN(_05297_ ) );
NAND2_X1 _13191_ ( .A1(\ID_EX_imm [6] ), .A2(fanout_net_11 ), .ZN(_05298_ ) );
AND2_X4 _13192_ ( .A1(_05297_ ), .A2(_05298_ ), .ZN(_05299_ ) );
XNOR2_X1 _13193_ ( .A(_05299_ ), .B(_02371_ ), .ZN(_05300_ ) );
NOR4_X2 _13194_ ( .A1(_05288_ ), .A2(_05292_ ), .A3(_05296_ ), .A4(_05300_ ), .ZN(_05301_ ) );
AND2_X1 _13195_ ( .A1(_05284_ ), .A2(_05301_ ), .ZN(_05302_ ) );
INV_X1 _13196_ ( .A(_05296_ ), .ZN(_05303_ ) );
INV_X1 _13197_ ( .A(_05300_ ), .ZN(_05304_ ) );
INV_X1 _13198_ ( .A(_02319_ ), .ZN(_05305_ ) );
INV_X1 _13199_ ( .A(_05287_ ), .ZN(_05306_ ) );
NOR3_X1 _13200_ ( .A1(_05292_ ), .A2(_05305_ ), .A3(_05306_ ), .ZN(_05307_ ) );
AND3_X1 _13201_ ( .A1(_05289_ ), .A2(_02188_ ), .A3(_05290_ ), .ZN(_05308_ ) );
OAI211_X1 _13202_ ( .A(_05303_ ), .B(_05304_ ), .C1(_05307_ ), .C2(_05308_ ), .ZN(_05309_ ) );
NAND3_X1 _13203_ ( .A1(_05303_ ), .A2(_02371_ ), .A3(_05299_ ), .ZN(_05310_ ) );
INV_X1 _13204_ ( .A(_05295_ ), .ZN(_05311_ ) );
OAI211_X1 _13205_ ( .A(_05309_ ), .B(_05310_ ), .C1(_02376_ ), .C2(_05311_ ), .ZN(_05312_ ) );
OAI211_X1 _13206_ ( .A(_05239_ ), .B(_05259_ ), .C1(_05302_ ), .C2(_05312_ ), .ZN(_05313_ ) );
INV_X1 _13207_ ( .A(_02543_ ), .ZN(_05314_ ) );
INV_X1 _13208_ ( .A(_05237_ ), .ZN(_05315_ ) );
NOR3_X1 _13209_ ( .A1(_05234_ ), .A2(_05314_ ), .A3(_05315_ ), .ZN(_05316_ ) );
AND3_X1 _13210_ ( .A1(_02565_ ), .A2(_05230_ ), .A3(_05229_ ), .ZN(_05317_ ) );
OAI21_X1 _13211_ ( .A(_05227_ ), .B1(_05316_ ), .B2(_05317_ ), .ZN(_05318_ ) );
INV_X1 _13212_ ( .A(_05226_ ), .ZN(_05319_ ) );
NAND3_X1 _13213_ ( .A1(_05319_ ), .A2(_02592_ ), .A3(_05221_ ), .ZN(_05320_ ) );
NAND3_X1 _13214_ ( .A1(_02518_ ), .A2(_05224_ ), .A3(_05223_ ), .ZN(_05321_ ) );
AND3_X1 _13215_ ( .A1(_05318_ ), .A2(_05320_ ), .A3(_05321_ ), .ZN(_05322_ ) );
INV_X1 _13216_ ( .A(_02448_ ), .ZN(_05323_ ) );
INV_X1 _13217_ ( .A(_05256_ ), .ZN(_05324_ ) );
NOR3_X1 _13218_ ( .A1(_05252_ ), .A2(_05323_ ), .A3(_05324_ ), .ZN(_05325_ ) );
AND3_X1 _13219_ ( .A1(_02472_ ), .A2(_05249_ ), .A3(_05250_ ), .ZN(_05326_ ) );
OAI21_X1 _13220_ ( .A(_05248_ ), .B1(_05325_ ), .B2(_05326_ ), .ZN(_05327_ ) );
NAND3_X1 _13221_ ( .A1(_02399_ ), .A2(_05245_ ), .A3(_05244_ ), .ZN(_05328_ ) );
NAND2_X1 _13222_ ( .A1(_05327_ ), .A2(_05328_ ), .ZN(_05329_ ) );
INV_X1 _13223_ ( .A(_05242_ ), .ZN(_05330_ ) );
NOR3_X1 _13224_ ( .A1(_05247_ ), .A2(_02574_ ), .A3(_05330_ ), .ZN(_05331_ ) );
OAI21_X1 _13225_ ( .A(_05239_ ), .B1(_05329_ ), .B2(_05331_ ), .ZN(_05332_ ) );
NAND3_X1 _13226_ ( .A1(_05313_ ), .A2(_05322_ ), .A3(_05332_ ), .ZN(_05333_ ) );
NAND4_X1 _13227_ ( .A1(_05175_ ), .A2(_05195_ ), .A3(_05180_ ), .A4(_05185_ ), .ZN(_05334_ ) );
XNOR2_X1 _13228_ ( .A(_05203_ ), .B(_02666_ ), .ZN(_05335_ ) );
NOR3_X1 _13229_ ( .A1(_05334_ ), .A2(_05199_ ), .A3(_05335_ ), .ZN(_05336_ ) );
AOI211_X1 _13230_ ( .A(_05173_ ), .B(_05218_ ), .C1(_05333_ ), .C2(_05336_ ), .ZN(_05337_ ) );
NAND3_X1 _13231_ ( .A1(_04458_ ), .A2(_05132_ ), .A3(_04477_ ), .ZN(_05338_ ) );
NAND2_X1 _13232_ ( .A1(_02883_ ), .A2(fanout_net_11 ), .ZN(_05339_ ) );
NAND2_X1 _13233_ ( .A1(_05338_ ), .A2(_05339_ ), .ZN(_05340_ ) );
XNOR2_X1 _13234_ ( .A(_05340_ ), .B(_02858_ ), .ZN(_05341_ ) );
OR2_X1 _13235_ ( .A1(_04508_ ), .A2(fanout_net_11 ), .ZN(_05342_ ) );
OR2_X1 _13236_ ( .A1(_05132_ ), .A2(\ID_EX_imm [26] ), .ZN(_05343_ ) );
NAND2_X1 _13237_ ( .A1(_05342_ ), .A2(_05343_ ), .ZN(_05344_ ) );
NOR2_X1 _13238_ ( .A1(_05344_ ), .A2(_02885_ ), .ZN(_05345_ ) );
INV_X1 _13239_ ( .A(_05345_ ), .ZN(_05346_ ) );
AOI21_X1 _13240_ ( .A(_02880_ ), .B1(_05342_ ), .B2(_05343_ ), .ZN(_05347_ ) );
INV_X1 _13241_ ( .A(_05347_ ), .ZN(_05348_ ) );
AOI21_X1 _13242_ ( .A(_05341_ ), .B1(_05346_ ), .B2(_05348_ ), .ZN(_05349_ ) );
AOI21_X1 _13243_ ( .A(fanout_net_11 ), .B1(_04536_ ), .B2(_04555_ ), .ZN(_05350_ ) );
AND2_X1 _13244_ ( .A1(fanout_net_11 ), .A2(\ID_EX_imm [25] ), .ZN(_05351_ ) );
NOR2_X1 _13245_ ( .A1(_05350_ ), .A2(_05351_ ), .ZN(_05352_ ) );
XNOR2_X1 _13246_ ( .A(_05352_ ), .B(_02834_ ), .ZN(_05353_ ) );
INV_X1 _13247_ ( .A(_05353_ ), .ZN(_05354_ ) );
OR2_X1 _13248_ ( .A1(_04533_ ), .A2(\ID_EX_typ [4] ), .ZN(_05355_ ) );
NAND2_X1 _13249_ ( .A1(_02163_ ), .A2(\ID_EX_typ [4] ), .ZN(_05356_ ) );
NAND2_X1 _13250_ ( .A1(_05355_ ), .A2(_05356_ ), .ZN(_05357_ ) );
INV_X1 _13251_ ( .A(_02162_ ), .ZN(_05358_ ) );
NOR2_X1 _13252_ ( .A1(_05357_ ), .A2(_05358_ ), .ZN(_05359_ ) );
AOI21_X1 _13253_ ( .A(_02162_ ), .B1(_05355_ ), .B2(_05356_ ), .ZN(_05360_ ) );
NOR2_X1 _13254_ ( .A1(_05359_ ), .A2(_05360_ ), .ZN(_05361_ ) );
INV_X1 _13255_ ( .A(_05361_ ), .ZN(_05362_ ) );
NAND3_X1 _13256_ ( .A1(_05349_ ), .A2(_05354_ ), .A3(_05362_ ), .ZN(_05363_ ) );
OR2_X1 _13257_ ( .A1(_05337_ ), .A2(_05363_ ), .ZN(_05364_ ) );
INV_X1 _13258_ ( .A(_05349_ ), .ZN(_05365_ ) );
AND2_X1 _13259_ ( .A1(_05352_ ), .A2(_02835_ ), .ZN(_05366_ ) );
NOR2_X1 _13260_ ( .A1(_05352_ ), .A2(_02835_ ), .ZN(_05367_ ) );
OAI211_X1 _13261_ ( .A(_02162_ ), .B(_05357_ ), .C1(_05366_ ), .C2(_05367_ ), .ZN(_05368_ ) );
NAND2_X1 _13262_ ( .A1(_05352_ ), .A2(_02834_ ), .ZN(_05369_ ) );
AOI21_X1 _13263_ ( .A(_05365_ ), .B1(_05368_ ), .B2(_05369_ ), .ZN(_05370_ ) );
INV_X1 _13264_ ( .A(_05344_ ), .ZN(_05371_ ) );
NOR3_X1 _13265_ ( .A1(_05371_ ), .A2(_05341_ ), .A3(_02885_ ), .ZN(_05372_ ) );
AND2_X1 _13266_ ( .A1(_05340_ ), .A2(_02858_ ), .ZN(_05373_ ) );
NOR3_X1 _13267_ ( .A1(_05370_ ), .A2(_05372_ ), .A3(_05373_ ), .ZN(_05374_ ) );
AND2_X2 _13268_ ( .A1(_05364_ ), .A2(_05374_ ), .ZN(_05375_ ) );
XNOR2_X1 _13269_ ( .A(_05141_ ), .B(_02937_ ), .ZN(_05376_ ) );
NOR3_X4 _13270_ ( .A1(_05375_ ), .A2(_05138_ ), .A3(_05376_ ), .ZN(_05377_ ) );
AOI21_X2 _13271_ ( .A(_05160_ ), .B1(_05377_ ), .B2(_05152_ ), .ZN(_05378_ ) );
INV_X1 _13272_ ( .A(\ID_EX_typ [1] ), .ZN(_05379_ ) );
NOR2_X1 _13273_ ( .A1(_05379_ ), .A2(fanout_net_8 ), .ZN(_05380_ ) );
AND2_X1 _13274_ ( .A1(_05380_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05381_ ) );
BUF_X4 _13275_ ( .A(_05381_ ), .Z(_05382_ ) );
INV_X1 _13276_ ( .A(_05382_ ), .ZN(_05383_ ) );
NOR2_X2 _13277_ ( .A1(_05378_ ), .A2(_05383_ ), .ZN(_05384_ ) );
AND2_X1 _13278_ ( .A1(fanout_net_8 ), .A2(\ID_EX_typ [1] ), .ZN(_05385_ ) );
AND2_X2 _13279_ ( .A1(_05385_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ), .ZN(_05386_ ) );
INV_X1 _13280_ ( .A(_05386_ ), .ZN(_05387_ ) );
AND2_X1 _13281_ ( .A1(_02258_ ), .A2(_04866_ ), .ZN(_05388_ ) );
NAND2_X1 _13282_ ( .A1(_02282_ ), .A2(_05099_ ), .ZN(_05389_ ) );
NAND2_X1 _13283_ ( .A1(_05123_ ), .A2(_05389_ ), .ZN(_05390_ ) );
AOI21_X1 _13284_ ( .A(_05388_ ), .B1(_05390_ ), .B2(_04867_ ), .ZN(_05391_ ) );
AOI21_X1 _13285_ ( .A(_05391_ ), .B1(_02315_ ), .B2(_04888_ ), .ZN(_05392_ ) );
NOR2_X1 _13286_ ( .A1(_02315_ ), .A2(_04888_ ), .ZN(_05393_ ) );
OAI21_X1 _13287_ ( .A(_04845_ ), .B1(_05392_ ), .B2(_05393_ ), .ZN(_05394_ ) );
NAND2_X1 _13288_ ( .A1(_02371_ ), .A2(_04778_ ), .ZN(_05395_ ) );
NOR2_X1 _13289_ ( .A1(_04801_ ), .A2(_05395_ ), .ZN(_05396_ ) );
NAND3_X1 _13290_ ( .A1(_04844_ ), .A2(_02319_ ), .A3(_04822_ ), .ZN(_05397_ ) );
OAI21_X1 _13291_ ( .A(_05397_ ), .B1(_02213_ ), .B2(_04843_ ), .ZN(_05398_ ) );
AOI221_X4 _13292_ ( .A(_05396_ ), .B1(_02345_ ), .B2(_04800_ ), .C1(_05398_ ), .C2(_04802_ ), .ZN(_05399_ ) );
AND2_X1 _13293_ ( .A1(_05394_ ), .A2(_05399_ ), .ZN(_05400_ ) );
INV_X1 _13294_ ( .A(_05400_ ), .ZN(_05401_ ) );
NAND2_X1 _13295_ ( .A1(_05401_ ), .A2(_05078_ ), .ZN(_05402_ ) );
NAND3_X1 _13296_ ( .A1(_05028_ ), .A2(_02592_ ), .A3(_05004_ ), .ZN(_05403_ ) );
INV_X1 _13297_ ( .A(_02518_ ), .ZN(_05404_ ) );
INV_X1 _13298_ ( .A(_05077_ ), .ZN(_05405_ ) );
NAND3_X1 _13299_ ( .A1(_04936_ ), .A2(_02422_ ), .A3(_04912_ ), .ZN(_05406_ ) );
OAI21_X1 _13300_ ( .A(_05406_ ), .B1(_02577_ ), .B2(_04935_ ), .ZN(_05407_ ) );
AND2_X1 _13301_ ( .A1(_02448_ ), .A2(_04981_ ), .ZN(_05408_ ) );
NAND2_X1 _13302_ ( .A1(_04960_ ), .A2(_05408_ ), .ZN(_05409_ ) );
INV_X1 _13303_ ( .A(_04958_ ), .ZN(_05410_ ) );
NAND2_X1 _13304_ ( .A1(_05409_ ), .A2(_05410_ ), .ZN(_05411_ ) );
AOI21_X1 _13305_ ( .A(_05407_ ), .B1(_05411_ ), .B2(_04937_ ), .ZN(_05412_ ) );
OAI221_X1 _13306_ ( .A(_05403_ ), .B1(_05404_ ), .B2(_05027_ ), .C1(_05405_ ), .C2(_05412_ ), .ZN(_05413_ ) );
INV_X1 _13307_ ( .A(_05073_ ), .ZN(_05414_ ) );
NAND2_X1 _13308_ ( .A1(_02588_ ), .A2(_05050_ ), .ZN(_05415_ ) );
AOI21_X1 _13309_ ( .A(_05074_ ), .B1(_05414_ ), .B2(_05415_ ), .ZN(_05416_ ) );
AOI21_X1 _13310_ ( .A(_05413_ ), .B1(_05029_ ), .B2(_05416_ ), .ZN(_05417_ ) );
NAND2_X2 _13311_ ( .A1(_05402_ ), .A2(_05417_ ), .ZN(_05418_ ) );
AND2_X2 _13312_ ( .A1(_05418_ ), .A2(_04757_ ), .ZN(_05419_ ) );
NAND3_X1 _13313_ ( .A1(_04709_ ), .A2(_02642_ ), .A3(_04682_ ), .ZN(_05420_ ) );
INV_X1 _13314_ ( .A(_02618_ ), .ZN(_05421_ ) );
OAI21_X1 _13315_ ( .A(_05420_ ), .B1(_05421_ ), .B2(_04708_ ), .ZN(_05422_ ) );
AND2_X1 _13316_ ( .A1(_02666_ ), .A2(_04753_ ), .ZN(_05423_ ) );
AND2_X1 _13317_ ( .A1(_04732_ ), .A2(_05423_ ), .ZN(_05424_ ) );
AOI21_X1 _13318_ ( .A(_05424_ ), .B1(_02688_ ), .B2(_04731_ ), .ZN(_05425_ ) );
INV_X1 _13319_ ( .A(_05425_ ), .ZN(_05426_ ) );
AOI21_X1 _13320_ ( .A(_05422_ ), .B1(_05426_ ), .B2(_04710_ ), .ZN(_05427_ ) );
INV_X1 _13321_ ( .A(_04661_ ), .ZN(_05428_ ) );
NOR2_X1 _13322_ ( .A1(_05427_ ), .A2(_05428_ ), .ZN(_05429_ ) );
INV_X1 _13323_ ( .A(_05429_ ), .ZN(_05430_ ) );
AND2_X1 _13324_ ( .A1(_02770_ ), .A2(_04659_ ), .ZN(_05431_ ) );
NOR2_X1 _13325_ ( .A1(_04635_ ), .A2(_05431_ ), .ZN(_05432_ ) );
NOR2_X1 _13326_ ( .A1(_05432_ ), .A2(_04636_ ), .ZN(_05433_ ) );
AND3_X1 _13327_ ( .A1(_05433_ ), .A2(_04609_ ), .A3(_04586_ ), .ZN(_05434_ ) );
INV_X1 _13328_ ( .A(_05434_ ), .ZN(_05435_ ) );
AND2_X1 _13329_ ( .A1(_02748_ ), .A2(_04585_ ), .ZN(_05436_ ) );
AND2_X1 _13330_ ( .A1(_04609_ ), .A2(_05436_ ), .ZN(_05437_ ) );
AOI21_X1 _13331_ ( .A(_05437_ ), .B1(_02726_ ), .B2(_04608_ ), .ZN(_05438_ ) );
AND3_X1 _13332_ ( .A1(_05430_ ), .A2(_05435_ ), .A3(_05438_ ), .ZN(_05439_ ) );
INV_X1 _13333_ ( .A(_05439_ ), .ZN(_05440_ ) );
OAI21_X1 _13334_ ( .A(_04559_ ), .B1(_05419_ ), .B2(_05440_ ), .ZN(_05441_ ) );
OR3_X1 _13335_ ( .A1(_04480_ ), .A2(_02885_ ), .A3(_04508_ ), .ZN(_05442_ ) );
INV_X1 _13336_ ( .A(_02858_ ), .ZN(_05443_ ) );
OAI21_X1 _13337_ ( .A(_05442_ ), .B1(_05443_ ), .B2(_04478_ ), .ZN(_05444_ ) );
INV_X1 _13338_ ( .A(_04557_ ), .ZN(_05445_ ) );
OR3_X1 _13339_ ( .A1(_05445_ ), .A2(_05358_ ), .A3(_04533_ ), .ZN(_05446_ ) );
AOI21_X1 _13340_ ( .A(_04556_ ), .B1(_02833_ ), .B2(_02812_ ), .ZN(_05447_ ) );
INV_X1 _13341_ ( .A(_05447_ ), .ZN(_05448_ ) );
NAND2_X1 _13342_ ( .A1(_05446_ ), .A2(_05448_ ), .ZN(_05449_ ) );
AOI21_X1 _13343_ ( .A(_05444_ ), .B1(_05449_ ), .B2(_04511_ ), .ZN(_05450_ ) );
INV_X1 _13344_ ( .A(_04456_ ), .ZN(_05451_ ) );
NOR2_X1 _13345_ ( .A1(_05450_ ), .A2(_05451_ ), .ZN(_05452_ ) );
NOR2_X1 _13346_ ( .A1(_02937_ ), .A2(_04408_ ), .ZN(_05453_ ) );
NAND2_X1 _13347_ ( .A1(_04385_ ), .A2(_05453_ ), .ZN(_05454_ ) );
NOR2_X1 _13348_ ( .A1(_05137_ ), .A2(_04384_ ), .ZN(_05455_ ) );
INV_X1 _13349_ ( .A(_05455_ ), .ZN(_05456_ ) );
NAND2_X1 _13350_ ( .A1(_05454_ ), .A2(_05456_ ), .ZN(_05457_ ) );
AND3_X1 _13351_ ( .A1(_05457_ ), .A2(_04433_ ), .A3(_04455_ ), .ZN(_05458_ ) );
NOR2_X1 _13352_ ( .A1(_02962_ ), .A2(_04454_ ), .ZN(_05459_ ) );
NAND2_X1 _13353_ ( .A1(_04433_ ), .A2(_05459_ ), .ZN(_05460_ ) );
INV_X1 _13354_ ( .A(_02987_ ), .ZN(_05461_ ) );
OAI21_X1 _13355_ ( .A(_05460_ ), .B1(_05461_ ), .B2(_04432_ ), .ZN(_05462_ ) );
NOR3_X1 _13356_ ( .A1(_05452_ ), .A2(_05458_ ), .A3(_05462_ ), .ZN(_05463_ ) );
AOI21_X1 _13357_ ( .A(_05387_ ), .B1(_05441_ ), .B2(_05463_ ), .ZN(_05464_ ) );
AND2_X1 _13358_ ( .A1(_05127_ ), .A2(\ID_EX_typ [2] ), .ZN(_05465_ ) );
AND3_X1 _13359_ ( .A1(_05441_ ), .A2(_05463_ ), .A3(_05465_ ), .ZN(_05466_ ) );
OR4_X2 _13360_ ( .A1(_05384_ ), .A2(_05464_ ), .A3(_05128_ ), .A4(_05466_ ), .ZN(_05467_ ) );
INV_X1 _13361_ ( .A(\ID_EX_typ [2] ), .ZN(_05468_ ) );
NOR3_X1 _13362_ ( .A1(_05468_ ), .A2(fanout_net_8 ), .A3(\ID_EX_typ [1] ), .ZN(_05469_ ) );
AND2_X1 _13363_ ( .A1(_05378_ ), .A2(_05469_ ), .ZN(_05470_ ) );
OAI221_X2 _13364_ ( .A(_04324_ ), .B1(_05125_ ), .B2(_05129_ ), .C1(_05467_ ), .C2(_05470_ ), .ZN(_05471_ ) );
NAND4_X1 _13365_ ( .A1(_05078_ ), .A2(_05124_ ), .A3(_04845_ ), .A4(_04890_ ), .ZN(_05472_ ) );
NAND2_X1 _13366_ ( .A1(_04757_ ), .A2(_04559_ ), .ZN(_05473_ ) );
OAI21_X1 _13367_ ( .A(_04323_ ), .B1(_05472_ ), .B2(_05473_ ), .ZN(_05474_ ) );
AND2_X4 _13368_ ( .A1(_05471_ ), .A2(_05474_ ), .ZN(_05475_ ) );
BUF_X4 _13369_ ( .A(_05475_ ), .Z(_05476_ ) );
MUX2_X1 _13370_ ( .A(_04241_ ), .B(_04321_ ), .S(_05476_ ), .Z(_05477_ ) );
BUF_X4 _13371_ ( .A(_04159_ ), .Z(_05478_ ) );
BUF_X4 _13372_ ( .A(_05478_ ), .Z(_05479_ ) );
AOI21_X1 _13373_ ( .A(_04229_ ), .B1(_05477_ ), .B2(_05479_ ), .ZN(_05480_ ) );
INV_X1 _13374_ ( .A(\ID_EX_typ [6] ), .ZN(_05481_ ) );
NAND2_X1 _13375_ ( .A1(_05481_ ), .A2(\ID_EX_typ [5] ), .ZN(_05482_ ) );
NOR2_X2 _13376_ ( .A1(_05482_ ), .A2(_03344_ ), .ZN(_05483_ ) );
INV_X1 _13377_ ( .A(_05483_ ), .ZN(_05484_ ) );
BUF_X4 _13378_ ( .A(_05484_ ), .Z(_05485_ ) );
BUF_X4 _13379_ ( .A(_05485_ ), .Z(_05486_ ) );
BUF_X4 _13380_ ( .A(_05126_ ), .Z(_05487_ ) );
BUF_X2 _13381_ ( .A(_05487_ ), .Z(_05488_ ) );
AOI21_X1 _13382_ ( .A(_05485_ ), .B1(_04321_ ), .B2(_05488_ ), .ZN(_05489_ ) );
OR2_X1 _13383_ ( .A1(_05489_ ), .A2(fanout_net_3 ), .ZN(_05490_ ) );
OR3_X1 _13384_ ( .A1(_03001_ ), .A2(fanout_net_3 ), .A3(_05488_ ), .ZN(_05491_ ) );
AOI22_X1 _13385_ ( .A1(_05480_ ), .A2(_05486_ ), .B1(_05490_ ), .B2(_05491_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_10_D ) );
AND2_X1 _13386_ ( .A1(_04302_ ), .A2(_04309_ ), .ZN(_05492_ ) );
NOR3_X1 _13387_ ( .A1(_05492_ ), .A2(_04306_ ), .A3(_04315_ ), .ZN(_05493_ ) );
NOR2_X1 _13388_ ( .A1(\ID_EX_pc [18] ), .A2(\ID_EX_imm [18] ), .ZN(_05494_ ) );
NOR3_X1 _13389_ ( .A1(_05493_ ), .A2(_05494_ ), .A3(_04311_ ), .ZN(_05495_ ) );
NOR2_X1 _13390_ ( .A1(_05495_ ), .A2(_04311_ ), .ZN(_05496_ ) );
XNOR2_X1 _13391_ ( .A(_05496_ ), .B(_04303_ ), .ZN(_05497_ ) );
MUX2_X1 _13392_ ( .A(_05497_ ), .B(_03006_ ), .S(fanout_net_8 ), .Z(_05498_ ) );
BUF_X4 _13393_ ( .A(_05484_ ), .Z(_05499_ ) );
BUF_X4 _13394_ ( .A(_05499_ ), .Z(_05500_ ) );
NOR2_X1 _13395_ ( .A1(_05498_ ), .A2(_05500_ ), .ZN(_05501_ ) );
INV_X4 _13396_ ( .A(_05475_ ), .ZN(_05502_ ) );
BUF_X4 _13397_ ( .A(_05502_ ), .Z(_05503_ ) );
BUF_X4 _13398_ ( .A(_05503_ ), .Z(_05504_ ) );
AND2_X1 _13399_ ( .A1(_04234_ ), .A2(_04239_ ), .ZN(_05505_ ) );
INV_X1 _13400_ ( .A(_05505_ ), .ZN(_05506_ ) );
NOR2_X1 _13401_ ( .A1(_05506_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_13_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05507_ ) );
XNOR2_X1 _13402_ ( .A(_05507_ ), .B(\ID_EX_pc [19] ), .ZN(_05508_ ) );
AOI21_X1 _13403_ ( .A(fanout_net_10 ), .B1(_05504_ ), .B2(_05508_ ), .ZN(_05509_ ) );
BUF_X4 _13404_ ( .A(_05502_ ), .Z(_05510_ ) );
BUF_X4 _13405_ ( .A(_05510_ ), .Z(_05511_ ) );
OAI21_X1 _13406_ ( .A(_05509_ ), .B1(_05511_ ), .B2(_05497_ ), .ZN(_05512_ ) );
AND4_X1 _13407_ ( .A1(_04167_ ), .A2(_04168_ ), .A3(_04163_ ), .A4(_04175_ ), .ZN(_05513_ ) );
AND4_X1 _13408_ ( .A1(_03823_ ), .A2(_05513_ ), .A3(_04166_ ), .A4(_04178_ ), .ZN(_05514_ ) );
BUF_X2 _13409_ ( .A(_05514_ ), .Z(_05515_ ) );
BUF_X2 _13410_ ( .A(_05515_ ), .Z(_05516_ ) );
INV_X1 _13411_ ( .A(\EX_LS_result_csreg_mem [19] ), .ZN(_05517_ ) );
AND4_X1 _13412_ ( .A1(_04161_ ), .A2(_04165_ ), .A3(_04177_ ), .A4(_04162_ ), .ZN(_05518_ ) );
AND3_X1 _13413_ ( .A1(_05518_ ), .A2(_04173_ ), .A3(_04174_ ), .ZN(_05519_ ) );
BUF_X2 _13414_ ( .A(_05519_ ), .Z(_05520_ ) );
BUF_X2 _13415_ ( .A(_05520_ ), .Z(_05521_ ) );
AND3_X1 _13416_ ( .A1(_05516_ ), .A2(_05517_ ), .A3(_05521_ ), .ZN(_05522_ ) );
AND2_X2 _13417_ ( .A1(_05514_ ), .A2(_05519_ ), .ZN(_05523_ ) );
AND4_X1 _13418_ ( .A1(\ID_EX_csr [10] ), .A2(_04142_ ), .A3(\ID_EX_csr [4] ), .A4(\ID_EX_csr [11] ), .ZN(_05524_ ) );
AND3_X1 _13419_ ( .A1(_05524_ ), .A2(_04185_ ), .A3(_04183_ ), .ZN(_05525_ ) );
AND2_X2 _13420_ ( .A1(_05525_ ), .A2(_04196_ ), .ZN(_05526_ ) );
NOR2_X1 _13421_ ( .A1(_05523_ ), .A2(_05526_ ), .ZN(_05527_ ) );
NAND4_X1 _13422_ ( .A1(_04118_ ), .A2(_04142_ ), .A3(_04145_ ), .A4(_04158_ ), .ZN(_05528_ ) );
INV_X1 _13423_ ( .A(_04183_ ), .ZN(_05529_ ) );
NOR2_X1 _13424_ ( .A1(_05528_ ), .A2(_05529_ ), .ZN(_05530_ ) );
BUF_X4 _13425_ ( .A(_05530_ ), .Z(_05531_ ) );
BUF_X4 _13426_ ( .A(_05531_ ), .Z(_05532_ ) );
BUF_X4 _13427_ ( .A(_05532_ ), .Z(_05533_ ) );
BUF_X4 _13428_ ( .A(_05533_ ), .Z(_05534_ ) );
BUF_X4 _13429_ ( .A(_04196_ ), .Z(_05535_ ) );
BUF_X4 _13430_ ( .A(_04200_ ), .Z(_05536_ ) );
BUF_X4 _13431_ ( .A(_05536_ ), .Z(_05537_ ) );
BUF_X4 _13432_ ( .A(_05537_ ), .Z(_05538_ ) );
NAND4_X1 _13433_ ( .A1(_05534_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][19] ), .A4(_05538_ ), .ZN(_05539_ ) );
BUF_X4 _13434_ ( .A(_04185_ ), .Z(_05540_ ) );
BUF_X4 _13435_ ( .A(_05540_ ), .Z(_05541_ ) );
BUF_X4 _13436_ ( .A(_05541_ ), .Z(_05542_ ) );
BUF_X4 _13437_ ( .A(_05542_ ), .Z(_05543_ ) );
NAND4_X1 _13438_ ( .A1(_05534_ ), .A2(_04218_ ), .A3(\mtvec [19] ), .A4(_05543_ ), .ZN(_05544_ ) );
BUF_X4 _13439_ ( .A(_05533_ ), .Z(_05545_ ) );
BUF_X2 _13440_ ( .A(_04191_ ), .Z(_05546_ ) );
NAND4_X1 _13441_ ( .A1(_05545_ ), .A2(_05546_ ), .A3(\mepc [19] ), .A4(_05538_ ), .ZN(_05547_ ) );
NAND4_X1 _13442_ ( .A1(_05545_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_05543_ ), .A4(_04223_ ), .ZN(_05548_ ) );
AND4_X1 _13443_ ( .A1(_05539_ ), .A2(_05544_ ), .A3(_05547_ ), .A4(_05548_ ), .ZN(_05549_ ) );
AOI211_X1 _13444_ ( .A(_04160_ ), .B(_05522_ ), .C1(_05527_ ), .C2(_05549_ ), .ZN(_05550_ ) );
BUF_X4 _13445_ ( .A(_05483_ ), .Z(_05551_ ) );
BUF_X4 _13446_ ( .A(_05551_ ), .Z(_05552_ ) );
NOR2_X1 _13447_ ( .A1(_05550_ ), .A2(_05552_ ), .ZN(_05553_ ) );
AOI211_X1 _13448_ ( .A(fanout_net_3 ), .B(_05501_ ), .C1(_05512_ ), .C2(_05553_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_11_D ) );
XOR2_X1 _13449_ ( .A(_05505_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_13_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .Z(_05554_ ) );
AOI21_X1 _13450_ ( .A(fanout_net_10 ), .B1(_05511_ ), .B2(_05554_ ), .ZN(_05555_ ) );
XNOR2_X1 _13451_ ( .A(_05493_ ), .B(_04304_ ), .ZN(_05556_ ) );
OAI21_X1 _13452_ ( .A(_05555_ ), .B1(_05511_ ), .B2(_05556_ ), .ZN(_05557_ ) );
AND3_X1 _13453_ ( .A1(_05516_ ), .A2(_03998_ ), .A3(_05521_ ), .ZN(_05558_ ) );
NAND4_X1 _13454_ ( .A1(_05534_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][18] ), .A4(_05538_ ), .ZN(_05559_ ) );
NAND4_X1 _13455_ ( .A1(_05534_ ), .A2(_04218_ ), .A3(\mtvec [18] ), .A4(_05543_ ), .ZN(_05560_ ) );
NAND4_X1 _13456_ ( .A1(_05534_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_05543_ ), .A4(_04223_ ), .ZN(_05561_ ) );
NAND4_X1 _13457_ ( .A1(_05545_ ), .A2(_05546_ ), .A3(\mepc [18] ), .A4(_05538_ ), .ZN(_05562_ ) );
AND4_X1 _13458_ ( .A1(_05559_ ), .A2(_05560_ ), .A3(_05561_ ), .A4(_05562_ ), .ZN(_05563_ ) );
AOI211_X1 _13459_ ( .A(_04160_ ), .B(_05558_ ), .C1(_05527_ ), .C2(_05563_ ), .ZN(_05564_ ) );
NOR2_X1 _13460_ ( .A1(_05564_ ), .A2(_05552_ ), .ZN(_05565_ ) );
AOI21_X1 _13461_ ( .A(_05485_ ), .B1(_05556_ ), .B2(_05488_ ), .ZN(_05566_ ) );
OR2_X1 _13462_ ( .A1(_05566_ ), .A2(fanout_net_3 ), .ZN(_05567_ ) );
OR3_X1 _13463_ ( .A1(_03009_ ), .A2(fanout_net_3 ), .A3(_05488_ ), .ZN(_05568_ ) );
AOI22_X1 _13464_ ( .A1(_05557_ ), .A2(_05565_ ), .B1(_05567_ ), .B2(_05568_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_12_D ) );
CLKBUF_X2 _13465_ ( .A(_05483_ ), .Z(_05569_ ) );
INV_X1 _13466_ ( .A(_04305_ ), .ZN(_05570_ ) );
AOI21_X1 _13467_ ( .A(_05570_ ), .B1(_04284_ ), .B2(_04301_ ), .ZN(_05571_ ) );
OR2_X1 _13468_ ( .A1(_05571_ ), .A2(_04314_ ), .ZN(_05572_ ) );
XNOR2_X1 _13469_ ( .A(_05572_ ), .B(_04308_ ), .ZN(_05573_ ) );
MUX2_X1 _13470_ ( .A(_05573_ ), .B(_03013_ ), .S(fanout_net_8 ), .Z(_05574_ ) );
AND3_X1 _13471_ ( .A1(_05471_ ), .A2(_05474_ ), .A3(_05573_ ), .ZN(_05575_ ) );
INV_X1 _13472_ ( .A(\ID_EX_pc [17] ), .ZN(_05576_ ) );
NAND3_X1 _13473_ ( .A1(_04233_ ), .A2(\ID_EX_pc [9] ), .A3(_04236_ ), .ZN(_05577_ ) );
INV_X1 _13474_ ( .A(\ID_EX_pc [12] ), .ZN(_05578_ ) );
NOR2_X1 _13475_ ( .A1(_05577_ ), .A2(_05578_ ), .ZN(_05579_ ) );
NAND3_X1 _13476_ ( .A1(_05579_ ), .A2(\ID_EX_pc [13] ), .A3(_04238_ ), .ZN(_05580_ ) );
INV_X1 _13477_ ( .A(\ID_EX_pc [16] ), .ZN(_05581_ ) );
OAI21_X1 _13478_ ( .A(_05576_ ), .B1(_05580_ ), .B2(_05581_ ), .ZN(_05582_ ) );
AOI21_X1 _13479_ ( .A(_05475_ ), .B1(_05506_ ), .B2(_05582_ ), .ZN(_05583_ ) );
OR3_X1 _13480_ ( .A1(_05575_ ), .A2(_05583_ ), .A3(fanout_net_10 ), .ZN(_05584_ ) );
OR3_X1 _13481_ ( .A1(_04171_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_04180_ ), .ZN(_05585_ ) );
NOR2_X1 _13482_ ( .A1(_04192_ ), .A2(_04197_ ), .ZN(_05586_ ) );
BUF_X4 _13483_ ( .A(_04205_ ), .Z(_05587_ ) );
NAND3_X1 _13484_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][17] ), .A3(_05587_ ), .ZN(_05588_ ) );
NAND3_X1 _13485_ ( .A1(_04226_ ), .A2(\mepc [17] ), .A3(_05587_ ), .ZN(_05589_ ) );
BUF_X4 _13486_ ( .A(_04221_ ), .Z(_05590_ ) );
NAND3_X1 _13487_ ( .A1(_04213_ ), .A2(\mycsreg.CSReg[0][17] ), .A3(_05590_ ), .ZN(_05591_ ) );
NAND4_X1 _13488_ ( .A1(_05586_ ), .A2(_05588_ ), .A3(_05589_ ), .A4(_05591_ ), .ZN(_05592_ ) );
BUF_X2 _13489_ ( .A(_04212_ ), .Z(_05593_ ) );
BUF_X2 _13490_ ( .A(_04216_ ), .Z(_05594_ ) );
BUF_X2 _13491_ ( .A(_05594_ ), .Z(_05595_ ) );
NAND3_X1 _13492_ ( .A1(_05593_ ), .A2(\mtvec [17] ), .A3(_05595_ ), .ZN(_05596_ ) );
OAI21_X1 _13493_ ( .A(_05596_ ), .B1(_04171_ ), .B2(_04180_ ), .ZN(_05597_ ) );
OAI211_X1 _13494_ ( .A(_05585_ ), .B(fanout_net_10 ), .C1(_05592_ ), .C2(_05597_ ), .ZN(_05598_ ) );
AND2_X1 _13495_ ( .A1(_05598_ ), .A2(_05499_ ), .ZN(_05599_ ) );
AOI221_X1 _13496_ ( .A(fanout_net_3 ), .B1(_05569_ ), .B2(_05574_ ), .C1(_05584_ ), .C2(_05599_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_13_D ) );
BUF_X4 _13497_ ( .A(_05515_ ), .Z(_05600_ ) );
BUF_X4 _13498_ ( .A(_05520_ ), .Z(_05601_ ) );
NAND3_X1 _13499_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [16] ), .A3(_05601_ ), .ZN(_05602_ ) );
BUF_X4 _13500_ ( .A(_05530_ ), .Z(_05603_ ) );
BUF_X2 _13501_ ( .A(_05603_ ), .Z(_05604_ ) );
BUF_X4 _13502_ ( .A(_05541_ ), .Z(_05605_ ) );
NAND4_X1 _13503_ ( .A1(_05604_ ), .A2(_04217_ ), .A3(\mtvec [16] ), .A4(_05605_ ), .ZN(_05606_ ) );
BUF_X4 _13504_ ( .A(_05532_ ), .Z(_05607_ ) );
NAND4_X1 _13505_ ( .A1(_05607_ ), .A2(\mycsreg.CSReg[0][16] ), .A3(_05605_ ), .A4(_05590_ ), .ZN(_05608_ ) );
BUF_X2 _13506_ ( .A(_04195_ ), .Z(_05609_ ) );
BUF_X4 _13507_ ( .A(_05536_ ), .Z(_05610_ ) );
NAND4_X1 _13508_ ( .A1(_05607_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][16] ), .A4(_05610_ ), .ZN(_05611_ ) );
NAND3_X1 _13509_ ( .A1(_05606_ ), .A2(_05608_ ), .A3(_05611_ ), .ZN(_05612_ ) );
AND2_X1 _13510_ ( .A1(_05525_ ), .A2(_04191_ ), .ZN(_05613_ ) );
BUF_X2 _13511_ ( .A(_05531_ ), .Z(_05614_ ) );
AND4_X1 _13512_ ( .A1(\mepc [16] ), .A2(_05614_ ), .A3(_04191_ ), .A4(_05536_ ), .ZN(_05615_ ) );
NOR4_X1 _13513_ ( .A1(_05612_ ), .A2(_05613_ ), .A3(_05526_ ), .A4(_05615_ ), .ZN(_05616_ ) );
BUF_X4 _13514_ ( .A(_05523_ ), .Z(_05617_ ) );
OAI21_X1 _13515_ ( .A(_05602_ ), .B1(_05616_ ), .B2(_05617_ ), .ZN(_05618_ ) );
AOI21_X1 _13516_ ( .A(_05551_ ), .B1(_05618_ ), .B2(fanout_net_10 ), .ZN(_05619_ ) );
AND3_X1 _13517_ ( .A1(_04234_ ), .A2(_04238_ ), .A3(_04237_ ), .ZN(_05620_ ) );
XNOR2_X1 _13518_ ( .A(_05620_ ), .B(_05581_ ), .ZN(_05621_ ) );
AND2_X1 _13519_ ( .A1(_05503_ ), .A2(_05621_ ), .ZN(_05622_ ) );
XNOR2_X1 _13520_ ( .A(_04302_ ), .B(_05570_ ), .ZN(_05623_ ) );
AOI21_X1 _13521_ ( .A(_05622_ ), .B1(_05476_ ), .B2(_05623_ ), .ZN(_05624_ ) );
OAI21_X1 _13522_ ( .A(_05619_ ), .B1(_05624_ ), .B2(fanout_net_10 ), .ZN(_05625_ ) );
AOI21_X1 _13523_ ( .A(_05485_ ), .B1(_05623_ ), .B2(_05488_ ), .ZN(_05626_ ) );
BUF_X4 _13524_ ( .A(_05487_ ), .Z(_05627_ ) );
BUF_X4 _13525_ ( .A(_05627_ ), .Z(_05628_ ) );
OAI21_X1 _13526_ ( .A(_05626_ ), .B1(_03014_ ), .B2(_05628_ ), .ZN(_05629_ ) );
AND3_X1 _13527_ ( .A1(_05625_ ), .A2(_01682_ ), .A3(_05629_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_14_D ) );
OR2_X1 _13528_ ( .A1(_04282_ ), .A2(_04283_ ), .ZN(_05630_ ) );
AND2_X1 _13529_ ( .A1(_05630_ ), .A2(_04251_ ), .ZN(_05631_ ) );
OR2_X1 _13530_ ( .A1(_05631_ ), .A2(_04300_ ), .ZN(_05632_ ) );
AOI21_X1 _13531_ ( .A(_04292_ ), .B1(_05632_ ), .B2(_04257_ ), .ZN(_05633_ ) );
NOR2_X1 _13532_ ( .A1(\ID_EX_pc [14] ), .A2(\ID_EX_imm [14] ), .ZN(_05634_ ) );
NOR3_X1 _13533_ ( .A1(_05633_ ), .A2(_05634_ ), .A3(_04285_ ), .ZN(_05635_ ) );
NOR2_X1 _13534_ ( .A1(_05635_ ), .A2(_04285_ ), .ZN(_05636_ ) );
XNOR2_X1 _13535_ ( .A(_05636_ ), .B(_04252_ ), .ZN(_05637_ ) );
MUX2_X1 _13536_ ( .A(_05637_ ), .B(_03019_ ), .S(fanout_net_8 ), .Z(_05638_ ) );
NOR2_X1 _13537_ ( .A1(_05638_ ), .A2(_05500_ ), .ZN(_05639_ ) );
NAND2_X1 _13538_ ( .A1(_04234_ ), .A2(_04237_ ), .ZN(_05640_ ) );
NOR2_X1 _13539_ ( .A1(_05640_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_17_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05641_ ) );
XNOR2_X1 _13540_ ( .A(_05641_ ), .B(\ID_EX_pc [15] ), .ZN(_05642_ ) );
AOI21_X1 _13541_ ( .A(fanout_net_10 ), .B1(_05504_ ), .B2(_05642_ ), .ZN(_05643_ ) );
OAI21_X1 _13542_ ( .A(_05643_ ), .B1(_05511_ ), .B2(_05637_ ), .ZN(_05644_ ) );
INV_X1 _13543_ ( .A(_05523_ ), .ZN(_05645_ ) );
BUF_X2 _13544_ ( .A(_05645_ ), .Z(_05646_ ) );
INV_X2 _13545_ ( .A(_05526_ ), .ZN(_05647_ ) );
BUF_X2 _13546_ ( .A(_05531_ ), .Z(_05648_ ) );
BUF_X2 _13547_ ( .A(_05540_ ), .Z(_05649_ ) );
AND4_X1 _13548_ ( .A1(\mtvec [15] ), .A2(_05648_ ), .A3(_05594_ ), .A4(_05649_ ), .ZN(_05650_ ) );
NAND4_X1 _13549_ ( .A1(_05604_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][15] ), .A4(_05610_ ), .ZN(_05651_ ) );
NAND4_X1 _13550_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_05605_ ), .A4(_05590_ ), .ZN(_05652_ ) );
NAND2_X1 _13551_ ( .A1(_05651_ ), .A2(_05652_ ), .ZN(_05653_ ) );
AND2_X1 _13552_ ( .A1(_05531_ ), .A2(_04200_ ), .ZN(_05654_ ) );
AND2_X1 _13553_ ( .A1(_05654_ ), .A2(_04191_ ), .ZN(_05655_ ) );
AOI211_X1 _13554_ ( .A(_05650_ ), .B(_05653_ ), .C1(_05655_ ), .C2(\mepc [15] ), .ZN(_05656_ ) );
NAND3_X1 _13555_ ( .A1(_05646_ ), .A2(_05647_ ), .A3(_05656_ ), .ZN(_05657_ ) );
OAI211_X1 _13556_ ( .A(_05657_ ), .B(fanout_net_10 ), .C1(\EX_LS_result_csreg_mem [15] ), .C2(_05646_ ), .ZN(_05658_ ) );
AND2_X1 _13557_ ( .A1(_05658_ ), .A2(_05500_ ), .ZN(_05659_ ) );
AOI211_X1 _13558_ ( .A(fanout_net_3 ), .B(_05639_ ), .C1(_05644_ ), .C2(_05659_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_15_D ) );
XNOR2_X1 _13559_ ( .A(_05633_ ), .B(_04253_ ), .ZN(_05660_ ) );
NAND2_X1 _13560_ ( .A1(_05660_ ), .A2(_05627_ ), .ZN(_05661_ ) );
AOI21_X1 _13561_ ( .A(_05499_ ), .B1(_03020_ ), .B2(fanout_net_8 ), .ZN(_05662_ ) );
XNOR2_X1 _13562_ ( .A(_05640_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_17_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05663_ ) );
NAND2_X1 _13563_ ( .A1(_05510_ ), .A2(_05663_ ), .ZN(_05664_ ) );
OAI211_X1 _13564_ ( .A(_05664_ ), .B(_04160_ ), .C1(_05504_ ), .C2(_05660_ ), .ZN(_05665_ ) );
NAND4_X1 _13565_ ( .A1(_05532_ ), .A2(_04216_ ), .A3(\mtvec [14] ), .A4(_05541_ ), .ZN(_05666_ ) );
NAND4_X1 _13566_ ( .A1(_05603_ ), .A2(\mycsreg.CSReg[0][14] ), .A3(_05540_ ), .A4(_04221_ ), .ZN(_05667_ ) );
NAND4_X1 _13567_ ( .A1(_05603_ ), .A2(_04196_ ), .A3(\mycsreg.CSReg[3][14] ), .A4(_04200_ ), .ZN(_05668_ ) );
AND3_X1 _13568_ ( .A1(_05666_ ), .A2(_05667_ ), .A3(_05668_ ), .ZN(_05669_ ) );
NAND2_X1 _13569_ ( .A1(_05525_ ), .A2(_04191_ ), .ZN(_05670_ ) );
BUF_X2 _13570_ ( .A(_05670_ ), .Z(_05671_ ) );
BUF_X4 _13571_ ( .A(_04191_ ), .Z(_05672_ ) );
NAND4_X1 _13572_ ( .A1(_05607_ ), .A2(_05672_ ), .A3(\mepc [14] ), .A4(_05610_ ), .ZN(_05673_ ) );
NAND4_X1 _13573_ ( .A1(_05669_ ), .A2(_05671_ ), .A3(_05647_ ), .A4(_05673_ ), .ZN(_05674_ ) );
NAND2_X1 _13574_ ( .A1(_05645_ ), .A2(_05674_ ), .ZN(_05675_ ) );
NAND3_X1 _13575_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [14] ), .A3(_05601_ ), .ZN(_05676_ ) );
AOI21_X1 _13576_ ( .A(_05478_ ), .B1(_05675_ ), .B2(_05676_ ), .ZN(_05677_ ) );
BUF_X4 _13577_ ( .A(_05483_ ), .Z(_05678_ ) );
NOR2_X1 _13578_ ( .A1(_05677_ ), .A2(_05678_ ), .ZN(_05679_ ) );
AOI221_X1 _13579_ ( .A(fanout_net_3 ), .B1(_05661_ ), .B2(_05662_ ), .C1(_05665_ ), .C2(_05679_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_16_D ) );
AND2_X1 _13580_ ( .A1(_05632_ ), .A2(_04255_ ), .ZN(_05680_ ) );
OR2_X1 _13581_ ( .A1(_05680_ ), .A2(_04289_ ), .ZN(_05681_ ) );
XOR2_X1 _13582_ ( .A(_05681_ ), .B(_04256_ ), .Z(_05682_ ) );
INV_X1 _13583_ ( .A(_05682_ ), .ZN(_05683_ ) );
MUX2_X1 _13584_ ( .A(_05683_ ), .B(_03023_ ), .S(fanout_net_8 ), .Z(_05684_ ) );
AND2_X1 _13585_ ( .A1(_05684_ ), .A2(_05551_ ), .ZN(_05685_ ) );
BUF_X2 _13586_ ( .A(_04171_ ), .Z(_05686_ ) );
BUF_X2 _13587_ ( .A(_04180_ ), .Z(_05687_ ) );
OR3_X1 _13588_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [13] ), .A3(_05687_ ), .ZN(_05688_ ) );
NAND3_X1 _13589_ ( .A1(_04214_ ), .A2(\mtvec [13] ), .A3(_04218_ ), .ZN(_05689_ ) );
NAND3_X1 _13590_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][13] ), .A3(_04207_ ), .ZN(_05690_ ) );
NAND3_X1 _13591_ ( .A1(_04193_ ), .A2(_05689_ ), .A3(_05690_ ), .ZN(_05691_ ) );
NAND3_X1 _13592_ ( .A1(_04226_ ), .A2(\mepc [13] ), .A3(_04207_ ), .ZN(_05692_ ) );
NAND3_X1 _13593_ ( .A1(_04214_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_04223_ ), .ZN(_05693_ ) );
OAI211_X1 _13594_ ( .A(_05692_ ), .B(_05693_ ), .C1(_04172_ ), .C2(_04181_ ), .ZN(_05694_ ) );
OAI211_X1 _13595_ ( .A(_05688_ ), .B(fanout_net_10 ), .C1(_05691_ ), .C2(_05694_ ), .ZN(_05695_ ) );
INV_X1 _13596_ ( .A(_05695_ ), .ZN(_05696_ ) );
INV_X1 _13597_ ( .A(\ID_EX_pc [13] ), .ZN(_05697_ ) );
XNOR2_X1 _13598_ ( .A(_05579_ ), .B(_05697_ ), .ZN(_05698_ ) );
MUX2_X1 _13599_ ( .A(_05698_ ), .B(_05682_ ), .S(_05476_ ), .Z(_05699_ ) );
AOI21_X1 _13600_ ( .A(_05696_ ), .B1(_05699_ ), .B2(_05479_ ), .ZN(_05700_ ) );
AOI211_X1 _13601_ ( .A(fanout_net_3 ), .B(_05685_ ), .C1(_05700_ ), .C2(_05486_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_17_D ) );
OAI21_X1 _13602_ ( .A(fanout_net_8 ), .B1(_03024_ ), .B2(_03015_ ), .ZN(_05701_ ) );
XOR2_X1 _13603_ ( .A(_05632_ ), .B(_04255_ ), .Z(_05702_ ) );
OAI21_X1 _13604_ ( .A(_05701_ ), .B1(fanout_net_8 ), .B2(_05702_ ), .ZN(_05703_ ) );
XNOR2_X1 _13605_ ( .A(_05577_ ), .B(_05578_ ), .ZN(_05704_ ) );
NAND2_X1 _13606_ ( .A1(_05510_ ), .A2(_05704_ ), .ZN(_05705_ ) );
OAI211_X1 _13607_ ( .A(_05705_ ), .B(_04160_ ), .C1(_05504_ ), .C2(_05702_ ), .ZN(_05706_ ) );
NAND4_X1 _13608_ ( .A1(_05604_ ), .A2(_04217_ ), .A3(\mtvec [12] ), .A4(_05605_ ), .ZN(_05707_ ) );
NAND4_X1 _13609_ ( .A1(_05607_ ), .A2(\mycsreg.CSReg[0][12] ), .A3(_05649_ ), .A4(_05590_ ), .ZN(_05708_ ) );
BUF_X4 _13610_ ( .A(_05603_ ), .Z(_05709_ ) );
NAND4_X1 _13611_ ( .A1(_05709_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][12] ), .A4(_05610_ ), .ZN(_05710_ ) );
NAND3_X1 _13612_ ( .A1(_05707_ ), .A2(_05708_ ), .A3(_05710_ ), .ZN(_05711_ ) );
BUF_X4 _13613_ ( .A(_04200_ ), .Z(_05712_ ) );
NAND4_X1 _13614_ ( .A1(_05709_ ), .A2(_05672_ ), .A3(\mepc [12] ), .A4(_05712_ ), .ZN(_05713_ ) );
NAND3_X1 _13615_ ( .A1(_05647_ ), .A2(_05671_ ), .A3(_05713_ ), .ZN(_05714_ ) );
OAI21_X1 _13616_ ( .A(_05645_ ), .B1(_05711_ ), .B2(_05714_ ), .ZN(_05715_ ) );
NAND3_X1 _13617_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [12] ), .A3(_05601_ ), .ZN(_05716_ ) );
AOI21_X1 _13618_ ( .A(_05478_ ), .B1(_05715_ ), .B2(_05716_ ), .ZN(_05717_ ) );
NOR2_X1 _13619_ ( .A1(_05717_ ), .A2(_05678_ ), .ZN(_05718_ ) );
AOI221_X1 _13620_ ( .A(fanout_net_3 ), .B1(_05569_ ), .B2(_05703_ ), .C1(_05706_ ), .C2(_05718_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_18_D ) );
AND2_X1 _13621_ ( .A1(_05630_ ), .A2(_04242_ ), .ZN(_05719_ ) );
OR2_X1 _13622_ ( .A1(_05719_ ), .A2(_04295_ ), .ZN(_05720_ ) );
AOI21_X1 _13623_ ( .A(_04243_ ), .B1(_05720_ ), .B2(_04294_ ), .ZN(_05721_ ) );
NOR2_X1 _13624_ ( .A1(_05721_ ), .A2(_04293_ ), .ZN(_05722_ ) );
NOR2_X1 _13625_ ( .A1(_05722_ ), .A2(_04298_ ), .ZN(_05723_ ) );
XNOR2_X1 _13626_ ( .A(_05723_ ), .B(_04250_ ), .ZN(_05724_ ) );
MUX2_X1 _13627_ ( .A(_05724_ ), .B(_04156_ ), .S(fanout_net_8 ), .Z(_05725_ ) );
NOR2_X1 _13628_ ( .A1(_05725_ ), .A2(_05500_ ), .ZN(_05726_ ) );
INV_X1 _13629_ ( .A(_04234_ ), .ZN(_05727_ ) );
NOR2_X1 _13630_ ( .A1(_05727_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_21_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05728_ ) );
XNOR2_X1 _13631_ ( .A(_05728_ ), .B(\ID_EX_pc [11] ), .ZN(_05729_ ) );
AOI21_X1 _13632_ ( .A(fanout_net_10 ), .B1(_05504_ ), .B2(_05729_ ), .ZN(_05730_ ) );
OAI21_X1 _13633_ ( .A(_05730_ ), .B1(_05511_ ), .B2(_05724_ ), .ZN(_05731_ ) );
NAND4_X1 _13634_ ( .A1(_05533_ ), .A2(\mycsreg.CSReg[0][11] ), .A3(_05542_ ), .A4(_05590_ ), .ZN(_05732_ ) );
NAND4_X1 _13635_ ( .A1(_05533_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][11] ), .A4(_05537_ ), .ZN(_05733_ ) );
NAND4_X1 _13636_ ( .A1(_05533_ ), .A2(_05546_ ), .A3(\mepc [11] ), .A4(_05537_ ), .ZN(_05734_ ) );
NAND3_X1 _13637_ ( .A1(_05732_ ), .A2(_05733_ ), .A3(_05734_ ), .ZN(_05735_ ) );
NAND4_X1 _13638_ ( .A1(_05533_ ), .A2(_04217_ ), .A3(\mtvec [11] ), .A4(_05605_ ), .ZN(_05736_ ) );
NAND3_X1 _13639_ ( .A1(_05647_ ), .A2(_05671_ ), .A3(_05736_ ), .ZN(_05737_ ) );
OAI21_X1 _13640_ ( .A(_05646_ ), .B1(_05735_ ), .B2(_05737_ ), .ZN(_05738_ ) );
NAND3_X1 _13641_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [11] ), .A3(_05601_ ), .ZN(_05739_ ) );
AOI21_X1 _13642_ ( .A(_05479_ ), .B1(_05738_ ), .B2(_05739_ ), .ZN(_05740_ ) );
NOR2_X1 _13643_ ( .A1(_05740_ ), .A2(_05552_ ), .ZN(_05741_ ) );
AOI211_X1 _13644_ ( .A(fanout_net_3 ), .B(_05726_ ), .C1(_05731_ ), .C2(_05741_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_19_D ) );
AND2_X1 _13645_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_05742_ ) );
INV_X1 _13646_ ( .A(_05742_ ), .ZN(_05743_ ) );
XOR2_X1 _13647_ ( .A(\ID_EX_pc [24] ), .B(\ID_EX_imm [24] ), .Z(_05744_ ) );
XOR2_X1 _13648_ ( .A(\ID_EX_pc [23] ), .B(\ID_EX_imm [23] ), .Z(_05745_ ) );
XOR2_X1 _13649_ ( .A(\ID_EX_pc [22] ), .B(\ID_EX_imm [22] ), .Z(_05746_ ) );
AND2_X1 _13650_ ( .A1(_05745_ ), .A2(_05746_ ), .ZN(_05747_ ) );
AND2_X1 _13651_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_05748_ ) );
NOR2_X1 _13652_ ( .A1(\ID_EX_pc [21] ), .A2(\ID_EX_imm [21] ), .ZN(_05749_ ) );
NOR2_X1 _13653_ ( .A1(_05748_ ), .A2(_05749_ ), .ZN(_05750_ ) );
AND4_X1 _13654_ ( .A1(_04318_ ), .A2(_04319_ ), .A3(_05747_ ), .A4(_05750_ ), .ZN(_05751_ ) );
AND2_X1 _13655_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_05752_ ) );
AND2_X1 _13656_ ( .A1(_05745_ ), .A2(_05752_ ), .ZN(_05753_ ) );
AOI21_X1 _13657_ ( .A(_05753_ ), .B1(\ID_EX_pc [23] ), .B2(\ID_EX_imm [23] ), .ZN(_05754_ ) );
INV_X1 _13658_ ( .A(_05749_ ), .ZN(_05755_ ) );
AND2_X1 _13659_ ( .A1(\ID_EX_pc [20] ), .A2(\ID_EX_imm [20] ), .ZN(_05756_ ) );
AOI21_X1 _13660_ ( .A(_05748_ ), .B1(_05755_ ), .B2(_05756_ ), .ZN(_05757_ ) );
INV_X1 _13661_ ( .A(_05747_ ), .ZN(_05758_ ) );
OAI21_X1 _13662_ ( .A(_05754_ ), .B1(_05757_ ), .B2(_05758_ ), .ZN(_05759_ ) );
OAI21_X1 _13663_ ( .A(_05744_ ), .B1(_05751_ ), .B2(_05759_ ), .ZN(_05760_ ) );
NAND2_X1 _13664_ ( .A1(\ID_EX_pc [24] ), .A2(\ID_EX_imm [24] ), .ZN(_05761_ ) );
AND2_X1 _13665_ ( .A1(_05760_ ), .A2(_05761_ ), .ZN(_05762_ ) );
NOR2_X1 _13666_ ( .A1(\ID_EX_pc [25] ), .A2(\ID_EX_imm [25] ), .ZN(_05763_ ) );
OAI21_X1 _13667_ ( .A(_05743_ ), .B1(_05762_ ), .B2(_05763_ ), .ZN(_05764_ ) );
XOR2_X1 _13668_ ( .A(\ID_EX_pc [27] ), .B(\ID_EX_imm [27] ), .Z(_05765_ ) );
XOR2_X1 _13669_ ( .A(\ID_EX_pc [26] ), .B(\ID_EX_imm [26] ), .Z(_05766_ ) );
NAND3_X1 _13670_ ( .A1(_05764_ ), .A2(_05765_ ), .A3(_05766_ ), .ZN(_05767_ ) );
AND2_X1 _13671_ ( .A1(\ID_EX_pc [26] ), .A2(\ID_EX_imm [26] ), .ZN(_05768_ ) );
AND2_X1 _13672_ ( .A1(_05765_ ), .A2(_05768_ ), .ZN(_05769_ ) );
AOI21_X1 _13673_ ( .A(_05769_ ), .B1(\ID_EX_pc [27] ), .B2(\ID_EX_imm [27] ), .ZN(_05770_ ) );
AND2_X1 _13674_ ( .A1(_05767_ ), .A2(_05770_ ), .ZN(_05771_ ) );
AND2_X1 _13675_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_05772_ ) );
NOR2_X1 _13676_ ( .A1(\ID_EX_pc [28] ), .A2(\ID_EX_imm [28] ), .ZN(_05773_ ) );
NOR3_X1 _13677_ ( .A1(_05771_ ), .A2(_05772_ ), .A3(_05773_ ), .ZN(_05774_ ) );
OR2_X1 _13678_ ( .A1(_05774_ ), .A2(_05772_ ), .ZN(_05775_ ) );
XNOR2_X1 _13679_ ( .A(\ID_EX_pc [29] ), .B(\ID_EX_imm [29] ), .ZN(_05776_ ) );
XNOR2_X1 _13680_ ( .A(_05775_ ), .B(_05776_ ), .ZN(_05777_ ) );
INV_X1 _13681_ ( .A(_05777_ ), .ZN(_05778_ ) );
OAI21_X1 _13682_ ( .A(_05551_ ), .B1(_05778_ ), .B2(fanout_net_8 ), .ZN(_05779_ ) );
AOI21_X1 _13683_ ( .A(_05779_ ), .B1(_03027_ ), .B2(fanout_net_8 ), .ZN(_05780_ ) );
AND2_X1 _13684_ ( .A1(\ID_EX_pc [27] ), .A2(\ID_EX_pc [26] ), .ZN(_05781_ ) );
AND3_X1 _13685_ ( .A1(_04235_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_05782_ ) );
AND2_X1 _13686_ ( .A1(\ID_EX_pc [23] ), .A2(\ID_EX_pc [22] ), .ZN(_05783_ ) );
AND4_X1 _13687_ ( .A1(\ID_EX_pc [25] ), .A2(_05782_ ), .A3(\ID_EX_pc [24] ), .A4(_05783_ ), .ZN(_05784_ ) );
AND3_X1 _13688_ ( .A1(_05505_ ), .A2(_05781_ ), .A3(_05784_ ), .ZN(_05785_ ) );
INV_X1 _13689_ ( .A(_05785_ ), .ZN(_05786_ ) );
NOR2_X1 _13690_ ( .A1(_05786_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05787_ ) );
XNOR2_X1 _13691_ ( .A(_05787_ ), .B(\ID_EX_pc [29] ), .ZN(_05788_ ) );
MUX2_X1 _13692_ ( .A(_05788_ ), .B(_05778_ ), .S(_05476_ ), .Z(_05789_ ) );
OR2_X1 _13693_ ( .A1(_05789_ ), .A2(fanout_net_10 ), .ZN(_05790_ ) );
NAND4_X1 _13694_ ( .A1(_05533_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][29] ), .A4(_05537_ ), .ZN(_05791_ ) );
NAND4_X1 _13695_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[0][29] ), .A3(_05605_ ), .A4(_05590_ ), .ZN(_05792_ ) );
NAND4_X1 _13696_ ( .A1(_05604_ ), .A2(_05546_ ), .A3(\mepc [29] ), .A4(_05610_ ), .ZN(_05793_ ) );
NAND3_X1 _13697_ ( .A1(_05791_ ), .A2(_05792_ ), .A3(_05793_ ), .ZN(_05794_ ) );
NAND4_X1 _13698_ ( .A1(_05604_ ), .A2(_04217_ ), .A3(\mtvec [29] ), .A4(_05605_ ), .ZN(_05795_ ) );
NAND2_X1 _13699_ ( .A1(_05671_ ), .A2(_05795_ ), .ZN(_05796_ ) );
OAI21_X1 _13700_ ( .A(_05645_ ), .B1(_05794_ ), .B2(_05796_ ), .ZN(_05797_ ) );
NAND3_X1 _13701_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [29] ), .A3(_05601_ ), .ZN(_05798_ ) );
AOI21_X1 _13702_ ( .A(_05479_ ), .B1(_05797_ ), .B2(_05798_ ), .ZN(_05799_ ) );
NOR2_X1 _13703_ ( .A1(_05799_ ), .A2(_05552_ ), .ZN(_05800_ ) );
AOI211_X1 _13704_ ( .A(fanout_net_3 ), .B(_05780_ ), .C1(_05790_ ), .C2(_05800_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_1_D ) );
XNOR2_X1 _13705_ ( .A(_05721_ ), .B(_04247_ ), .ZN(_05801_ ) );
NAND2_X1 _13706_ ( .A1(_05801_ ), .A2(_05627_ ), .ZN(_05802_ ) );
AOI21_X1 _13707_ ( .A(_05499_ ), .B1(_04116_ ), .B2(fanout_net_8 ), .ZN(_05803_ ) );
XNOR2_X1 _13708_ ( .A(_04234_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_21_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05804_ ) );
OR2_X1 _13709_ ( .A1(_05476_ ), .A2(_05804_ ), .ZN(_05805_ ) );
OAI211_X1 _13710_ ( .A(_05805_ ), .B(_04160_ ), .C1(_05504_ ), .C2(_05801_ ), .ZN(_05806_ ) );
AND3_X1 _13711_ ( .A1(_05515_ ), .A2(_03999_ ), .A3(_05520_ ), .ZN(_05807_ ) );
NAND4_X1 _13712_ ( .A1(_05531_ ), .A2(_04195_ ), .A3(\mycsreg.CSReg[3][10] ), .A4(_04200_ ), .ZN(_05808_ ) );
NAND4_X1 _13713_ ( .A1(_05531_ ), .A2(_04216_ ), .A3(\mtvec [10] ), .A4(_05540_ ), .ZN(_05809_ ) );
NAND4_X1 _13714_ ( .A1(_05531_ ), .A2(\mycsreg.CSReg[0][10] ), .A3(_04185_ ), .A4(_04221_ ), .ZN(_05810_ ) );
NAND4_X1 _13715_ ( .A1(_05531_ ), .A2(_04190_ ), .A3(\mepc [10] ), .A4(_04200_ ), .ZN(_05811_ ) );
AND4_X1 _13716_ ( .A1(_05808_ ), .A2(_05809_ ), .A3(_05810_ ), .A4(_05811_ ), .ZN(_05812_ ) );
AOI211_X1 _13717_ ( .A(_04159_ ), .B(_05807_ ), .C1(_05527_ ), .C2(_05812_ ), .ZN(_05813_ ) );
NOR2_X1 _13718_ ( .A1(_05813_ ), .A2(_05678_ ), .ZN(_05814_ ) );
AOI221_X1 _13719_ ( .A(fanout_net_3 ), .B1(_05802_ ), .B2(_05803_ ), .C1(_05806_ ), .C2(_05814_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_20_D ) );
NAND2_X1 _13720_ ( .A1(_04121_ ), .A2(fanout_net_8 ), .ZN(_05815_ ) );
XNOR2_X1 _13721_ ( .A(_05720_ ), .B(_04245_ ), .ZN(_05816_ ) );
BUF_X4 _13722_ ( .A(_05627_ ), .Z(_05817_ ) );
NAND2_X1 _13723_ ( .A1(_05816_ ), .A2(_05817_ ), .ZN(_05818_ ) );
AOI21_X1 _13724_ ( .A(_05500_ ), .B1(_05815_ ), .B2(_05818_ ), .ZN(_05819_ ) );
INV_X1 _13725_ ( .A(\ID_EX_pc [9] ), .ZN(_05820_ ) );
XNOR2_X1 _13726_ ( .A(_04233_ ), .B(_05820_ ), .ZN(_05821_ ) );
INV_X1 _13727_ ( .A(_05816_ ), .ZN(_05822_ ) );
MUX2_X1 _13728_ ( .A(_05821_ ), .B(_05822_ ), .S(_05476_ ), .Z(_05823_ ) );
NAND2_X1 _13729_ ( .A1(_05823_ ), .A2(_05479_ ), .ZN(_05824_ ) );
AND4_X1 _13730_ ( .A1(\mycsreg.CSReg[0][9] ), .A2(_05531_ ), .A3(_05540_ ), .A4(_04221_ ), .ZN(_05825_ ) );
AOI21_X1 _13731_ ( .A(_05825_ ), .B1(_05655_ ), .B2(\mepc [9] ), .ZN(_05826_ ) );
NAND4_X1 _13732_ ( .A1(_05532_ ), .A2(_04216_ ), .A3(\mtvec [9] ), .A4(_05541_ ), .ZN(_05827_ ) );
NAND4_X1 _13733_ ( .A1(_05532_ ), .A2(_04196_ ), .A3(\mycsreg.CSReg[3][9] ), .A4(_05536_ ), .ZN(_05828_ ) );
AND2_X1 _13734_ ( .A1(_05827_ ), .A2(_05828_ ), .ZN(_05829_ ) );
NAND4_X1 _13735_ ( .A1(_05645_ ), .A2(_05647_ ), .A3(_05826_ ), .A4(_05829_ ), .ZN(_05830_ ) );
INV_X1 _13736_ ( .A(\EX_LS_result_csreg_mem [9] ), .ZN(_05831_ ) );
NAND3_X1 _13737_ ( .A1(_05515_ ), .A2(_05831_ ), .A3(_05520_ ), .ZN(_05832_ ) );
AND2_X1 _13738_ ( .A1(_05830_ ), .A2(_05832_ ), .ZN(_05833_ ) );
AOI21_X1 _13739_ ( .A(_05552_ ), .B1(_05833_ ), .B2(fanout_net_10 ), .ZN(_05834_ ) );
AOI211_X1 _13740_ ( .A(fanout_net_3 ), .B(_05819_ ), .C1(_05824_ ), .C2(_05834_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_21_D ) );
XOR2_X1 _13741_ ( .A(_05630_ ), .B(_04242_ ), .Z(_05835_ ) );
INV_X1 _13742_ ( .A(_05835_ ), .ZN(_05836_ ) );
OAI21_X1 _13743_ ( .A(_05551_ ), .B1(_05836_ ), .B2(fanout_net_8 ), .ZN(_05837_ ) );
AOI21_X1 _13744_ ( .A(_05837_ ), .B1(_04123_ ), .B2(fanout_net_8 ), .ZN(_05838_ ) );
INV_X1 _13745_ ( .A(\ID_EX_pc [8] ), .ZN(_05839_ ) );
XNOR2_X1 _13746_ ( .A(_04232_ ), .B(_05839_ ), .ZN(_05840_ ) );
AND2_X1 _13747_ ( .A1(_05503_ ), .A2(_05840_ ), .ZN(_05841_ ) );
AOI21_X1 _13748_ ( .A(_05841_ ), .B1(_05476_ ), .B2(_05835_ ), .ZN(_05842_ ) );
OR2_X1 _13749_ ( .A1(_05842_ ), .A2(fanout_net_10 ), .ZN(_05843_ ) );
NAND3_X1 _13750_ ( .A1(_05516_ ), .A2(\EX_LS_result_csreg_mem [8] ), .A3(_05521_ ), .ZN(_05844_ ) );
AND4_X1 _13751_ ( .A1(\mycsreg.CSReg[3][8] ), .A2(_05614_ ), .A3(_05609_ ), .A4(_05536_ ), .ZN(_05845_ ) );
NOR3_X1 _13752_ ( .A1(_05613_ ), .A2(_05526_ ), .A3(_05845_ ), .ZN(_05846_ ) );
BUF_X2 _13753_ ( .A(_05614_ ), .Z(_05847_ ) );
NAND4_X1 _13754_ ( .A1(_05847_ ), .A2(_05595_ ), .A3(\mtvec [8] ), .A4(_05542_ ), .ZN(_05848_ ) );
NAND4_X1 _13755_ ( .A1(_05847_ ), .A2(_05546_ ), .A3(\mepc [8] ), .A4(_05537_ ), .ZN(_05849_ ) );
BUF_X2 _13756_ ( .A(_04222_ ), .Z(_05850_ ) );
NAND4_X1 _13757_ ( .A1(_05847_ ), .A2(\mycsreg.CSReg[0][8] ), .A3(_05542_ ), .A4(_05850_ ), .ZN(_05851_ ) );
AND4_X1 _13758_ ( .A1(_05846_ ), .A2(_05848_ ), .A3(_05849_ ), .A4(_05851_ ), .ZN(_05852_ ) );
OAI21_X1 _13759_ ( .A(_05844_ ), .B1(_05852_ ), .B2(_05617_ ), .ZN(_05853_ ) );
AOI21_X1 _13760_ ( .A(_05552_ ), .B1(_05853_ ), .B2(fanout_net_10 ), .ZN(_05854_ ) );
AOI211_X1 _13761_ ( .A(fanout_net_3 ), .B(_05838_ ), .C1(_05843_ ), .C2(_05854_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_22_D ) );
NAND2_X1 _13762_ ( .A1(_04280_ ), .A2(_04281_ ), .ZN(_05855_ ) );
NOR2_X1 _13763_ ( .A1(_04283_ ), .A2(_04259_ ), .ZN(_05856_ ) );
XNOR2_X1 _13764_ ( .A(_05855_ ), .B(_05856_ ), .ZN(_05857_ ) );
OAI21_X1 _13765_ ( .A(_05551_ ), .B1(_05857_ ), .B2(fanout_net_8 ), .ZN(_05858_ ) );
AOI21_X1 _13766_ ( .A(_05858_ ), .B1(_04130_ ), .B2(fanout_net_8 ), .ZN(_05859_ ) );
NAND3_X1 _13767_ ( .A1(_04213_ ), .A2(\mtvec [7] ), .A3(_04217_ ), .ZN(_05860_ ) );
NAND3_X1 _13768_ ( .A1(_04213_ ), .A2(\mycsreg.CSReg[0][7] ), .A3(_05590_ ), .ZN(_05861_ ) );
AND2_X1 _13769_ ( .A1(_05860_ ), .A2(_05861_ ), .ZN(_05862_ ) );
AND3_X1 _13770_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][7] ), .A3(_04206_ ), .ZN(_05863_ ) );
AND2_X1 _13771_ ( .A1(_04226_ ), .A2(_04206_ ), .ZN(_05864_ ) );
AOI21_X1 _13772_ ( .A(_05863_ ), .B1(\mepc [7] ), .B2(_05864_ ), .ZN(_05865_ ) );
OAI211_X1 _13773_ ( .A(_05862_ ), .B(_05865_ ), .C1(_05686_ ), .C2(_05687_ ), .ZN(_05866_ ) );
OR3_X1 _13774_ ( .A1(_04171_ ), .A2(\EX_LS_result_csreg_mem [7] ), .A3(_04180_ ), .ZN(_05867_ ) );
NAND2_X1 _13775_ ( .A1(_05866_ ), .A2(_05867_ ), .ZN(_05868_ ) );
INV_X1 _13776_ ( .A(_04231_ ), .ZN(_05869_ ) );
NOR2_X1 _13777_ ( .A1(_05869_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05870_ ) );
XNOR2_X1 _13778_ ( .A(_05870_ ), .B(\ID_EX_pc [7] ), .ZN(_05871_ ) );
MUX2_X1 _13779_ ( .A(_05871_ ), .B(_05857_ ), .S(_05476_ ), .Z(_05872_ ) );
MUX2_X1 _13780_ ( .A(_05868_ ), .B(_05872_ ), .S(_05479_ ), .Z(_05873_ ) );
AOI211_X1 _13781_ ( .A(fanout_net_3 ), .B(_05859_ ), .C1(_05873_ ), .C2(_05486_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_23_D ) );
NAND2_X1 _13782_ ( .A1(_04136_ ), .A2(fanout_net_8 ), .ZN(_05874_ ) );
XOR2_X1 _13783_ ( .A(_04278_ ), .B(_04279_ ), .Z(_05875_ ) );
AOI21_X1 _13784_ ( .A(_05499_ ), .B1(_05875_ ), .B2(_05487_ ), .ZN(_05876_ ) );
XNOR2_X1 _13785_ ( .A(_04231_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05877_ ) );
OR2_X1 _13786_ ( .A1(_05475_ ), .A2(_05877_ ), .ZN(_05878_ ) );
OAI211_X1 _13787_ ( .A(_05878_ ), .B(_04160_ ), .C1(_05504_ ), .C2(_05875_ ), .ZN(_05879_ ) );
BUF_X2 _13788_ ( .A(_05483_ ), .Z(_05880_ ) );
NAND3_X1 _13789_ ( .A1(_05515_ ), .A2(\EX_LS_result_csreg_mem [6] ), .A3(_05520_ ), .ZN(_05881_ ) );
NAND4_X1 _13790_ ( .A1(_05603_ ), .A2(_04216_ ), .A3(\mtvec [6] ), .A4(_05540_ ), .ZN(_05882_ ) );
AND2_X1 _13791_ ( .A1(_05670_ ), .A2(_05882_ ), .ZN(_05883_ ) );
NAND4_X1 _13792_ ( .A1(_05648_ ), .A2(\mycsreg.CSReg[0][6] ), .A3(_05541_ ), .A4(_04222_ ), .ZN(_05884_ ) );
NAND4_X1 _13793_ ( .A1(_05648_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][6] ), .A4(_05712_ ), .ZN(_05885_ ) );
NAND4_X1 _13794_ ( .A1(_05614_ ), .A2(_05672_ ), .A3(\mepc [6] ), .A4(_05712_ ), .ZN(_05886_ ) );
AND4_X1 _13795_ ( .A1(_05883_ ), .A2(_05884_ ), .A3(_05885_ ), .A4(_05886_ ), .ZN(_05887_ ) );
OAI21_X1 _13796_ ( .A(_05881_ ), .B1(_05887_ ), .B2(_05523_ ), .ZN(_05888_ ) );
AOI21_X1 _13797_ ( .A(_05880_ ), .B1(_05888_ ), .B2(fanout_net_10 ), .ZN(_05889_ ) );
AOI221_X4 _13798_ ( .A(fanout_net_3 ), .B1(_05874_ ), .B2(_05876_ ), .C1(_05879_ ), .C2(_05889_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_24_D ) );
NOR2_X1 _13799_ ( .A1(_04260_ ), .A2(_04277_ ), .ZN(_05890_ ) );
XOR2_X1 _13800_ ( .A(_04276_ ), .B(_05890_ ), .Z(_05891_ ) );
MUX2_X1 _13801_ ( .A(_05891_ ), .B(_04141_ ), .S(fanout_net_8 ), .Z(_05892_ ) );
XNOR2_X1 _13802_ ( .A(_04230_ ), .B(\ID_EX_pc [5] ), .ZN(_05893_ ) );
AOI21_X1 _13803_ ( .A(fanout_net_10 ), .B1(_05503_ ), .B2(_05893_ ), .ZN(_05894_ ) );
INV_X1 _13804_ ( .A(_05891_ ), .ZN(_05895_ ) );
OAI21_X1 _13805_ ( .A(_05894_ ), .B1(_05504_ ), .B2(_05895_ ), .ZN(_05896_ ) );
NAND3_X1 _13806_ ( .A1(_05515_ ), .A2(\EX_LS_result_csreg_mem [5] ), .A3(_05520_ ), .ZN(_05897_ ) );
NAND4_X1 _13807_ ( .A1(_05648_ ), .A2(\mycsreg.CSReg[0][5] ), .A3(_05649_ ), .A4(_04222_ ), .ZN(_05898_ ) );
NAND4_X1 _13808_ ( .A1(_05648_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][5] ), .A4(_05712_ ), .ZN(_05899_ ) );
NAND4_X1 _13809_ ( .A1(_05648_ ), .A2(_05672_ ), .A3(\mepc [5] ), .A4(_05712_ ), .ZN(_05900_ ) );
NAND3_X1 _13810_ ( .A1(_05898_ ), .A2(_05899_ ), .A3(_05900_ ), .ZN(_05901_ ) );
NAND4_X1 _13811_ ( .A1(_05648_ ), .A2(_05594_ ), .A3(\mtvec [5] ), .A4(_05649_ ), .ZN(_05902_ ) );
NAND2_X1 _13812_ ( .A1(_05670_ ), .A2(_05902_ ), .ZN(_05903_ ) );
NOR2_X1 _13813_ ( .A1(_05901_ ), .A2(_05903_ ), .ZN(_05904_ ) );
OAI21_X1 _13814_ ( .A(_05897_ ), .B1(_05523_ ), .B2(_05904_ ), .ZN(_05905_ ) );
AOI21_X1 _13815_ ( .A(_05880_ ), .B1(_05905_ ), .B2(fanout_net_10 ), .ZN(_05906_ ) );
AOI221_X1 _13816_ ( .A(fanout_net_3 ), .B1(_05569_ ), .B2(_05892_ ), .C1(_05896_ ), .C2(_05906_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_25_D ) );
NAND2_X1 _13817_ ( .A1(_04143_ ), .A2(fanout_net_8 ), .ZN(_05907_ ) );
NAND2_X1 _13818_ ( .A1(_04271_ ), .A2(_04272_ ), .ZN(_05908_ ) );
XNOR2_X1 _13819_ ( .A(_05908_ ), .B(_04273_ ), .ZN(_05909_ ) );
AOI21_X1 _13820_ ( .A(_05499_ ), .B1(_05909_ ), .B2(_05487_ ), .ZN(_05910_ ) );
AND2_X1 _13821_ ( .A1(\ID_EX_pc [3] ), .A2(\ID_EX_pc [2] ), .ZN(_05911_ ) );
XNOR2_X1 _13822_ ( .A(_05911_ ), .B(\ID_EX_pc [4] ), .ZN(_05912_ ) );
NAND2_X1 _13823_ ( .A1(_05503_ ), .A2(_05912_ ), .ZN(_05913_ ) );
OAI211_X1 _13824_ ( .A(_05913_ ), .B(_04160_ ), .C1(_05504_ ), .C2(_05909_ ), .ZN(_05914_ ) );
NAND4_X1 _13825_ ( .A1(_05614_ ), .A2(_05594_ ), .A3(\mtvec [4] ), .A4(_05541_ ), .ZN(_05915_ ) );
NAND4_X1 _13826_ ( .A1(_05532_ ), .A2(_04196_ ), .A3(\mycsreg.CSReg[3][4] ), .A4(_05536_ ), .ZN(_05916_ ) );
AND2_X1 _13827_ ( .A1(_05915_ ), .A2(_05916_ ), .ZN(_05917_ ) );
NAND4_X1 _13828_ ( .A1(_05607_ ), .A2(_05672_ ), .A3(\mepc [4] ), .A4(_05610_ ), .ZN(_05918_ ) );
NAND4_X1 _13829_ ( .A1(_05607_ ), .A2(\mycsreg.CSReg[0][4] ), .A3(_05605_ ), .A4(_05590_ ), .ZN(_05919_ ) );
NAND4_X1 _13830_ ( .A1(_05917_ ), .A2(_05671_ ), .A3(_05918_ ), .A4(_05919_ ), .ZN(_05920_ ) );
NAND2_X1 _13831_ ( .A1(_05645_ ), .A2(_05920_ ), .ZN(_05921_ ) );
NAND3_X1 _13832_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [4] ), .A3(_05601_ ), .ZN(_05922_ ) );
AOI21_X1 _13833_ ( .A(_04159_ ), .B1(_05921_ ), .B2(_05922_ ), .ZN(_05923_ ) );
NOR2_X1 _13834_ ( .A1(_05923_ ), .A2(_05678_ ), .ZN(_05924_ ) );
AOI221_X1 _13835_ ( .A(fanout_net_3 ), .B1(_05907_ ), .B2(_05910_ ), .C1(_05914_ ), .C2(_05924_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_26_D ) );
AND4_X1 _13836_ ( .A1(_04269_ ), .A2(_04268_ ), .A3(_04272_ ), .A4(_04270_ ), .ZN(_05925_ ) );
AOI22_X1 _13837_ ( .A1(_04268_ ), .A2(_04270_ ), .B1(_04269_ ), .B2(_04272_ ), .ZN(_05926_ ) );
OAI21_X1 _13838_ ( .A(_05627_ ), .B1(_05925_ ), .B2(_05926_ ), .ZN(_05927_ ) );
AOI21_X1 _13839_ ( .A(_05499_ ), .B1(_04148_ ), .B2(fanout_net_8 ), .ZN(_05928_ ) );
XNOR2_X1 _13840_ ( .A(\ID_EX_pc [3] ), .B(\ID_EX_pc [2] ), .ZN(_05929_ ) );
NAND2_X1 _13841_ ( .A1(_05503_ ), .A2(_05929_ ), .ZN(_05930_ ) );
OR2_X1 _13842_ ( .A1(_05925_ ), .A2(_05926_ ), .ZN(_05931_ ) );
OAI211_X1 _13843_ ( .A(_05930_ ), .B(_04160_ ), .C1(_05510_ ), .C2(_05931_ ), .ZN(_05932_ ) );
NAND4_X1 _13844_ ( .A1(_05532_ ), .A2(_04216_ ), .A3(\mtvec [3] ), .A4(_05541_ ), .ZN(_05933_ ) );
NAND4_X1 _13845_ ( .A1(_05532_ ), .A2(_04196_ ), .A3(\mycsreg.CSReg[3][3] ), .A4(_05536_ ), .ZN(_05934_ ) );
AND2_X1 _13846_ ( .A1(_05933_ ), .A2(_05934_ ), .ZN(_05935_ ) );
NAND4_X1 _13847_ ( .A1(_05607_ ), .A2(_05672_ ), .A3(\mepc [3] ), .A4(_05610_ ), .ZN(_05936_ ) );
NAND4_X1 _13848_ ( .A1(_05709_ ), .A2(\mycsreg.CSReg[0][3] ), .A3(_05649_ ), .A4(_04222_ ), .ZN(_05937_ ) );
NAND4_X1 _13849_ ( .A1(_05935_ ), .A2(_05671_ ), .A3(_05936_ ), .A4(_05937_ ), .ZN(_05938_ ) );
NAND2_X1 _13850_ ( .A1(_05646_ ), .A2(_05938_ ), .ZN(_05939_ ) );
AND3_X1 _13851_ ( .A1(_05515_ ), .A2(\EX_LS_result_csreg_mem [3] ), .A3(_05520_ ), .ZN(_05940_ ) );
INV_X1 _13852_ ( .A(_05940_ ), .ZN(_05941_ ) );
AOI21_X1 _13853_ ( .A(_04159_ ), .B1(_05939_ ), .B2(_05941_ ), .ZN(_05942_ ) );
NOR2_X1 _13854_ ( .A1(_05942_ ), .A2(_05678_ ), .ZN(_05943_ ) );
AOI221_X1 _13855_ ( .A(fanout_net_3 ), .B1(_05927_ ), .B2(_05928_ ), .C1(_05932_ ), .C2(_05943_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_27_D ) );
NOR3_X1 _13856_ ( .A1(_04151_ ), .A2(_04146_ ), .A3(_05488_ ), .ZN(_05944_ ) );
XOR2_X1 _13857_ ( .A(_04266_ ), .B(_04267_ ), .Z(_05945_ ) );
INV_X1 _13858_ ( .A(_05945_ ), .ZN(_05946_ ) );
OAI21_X1 _13859_ ( .A(_05551_ ), .B1(_05946_ ), .B2(fanout_net_8 ), .ZN(_05947_ ) );
NOR2_X1 _13860_ ( .A1(_05944_ ), .A2(_05947_ ), .ZN(_05948_ ) );
MUX2_X1 _13861_ ( .A(\ID_EX_pc [2] ), .B(_05946_ ), .S(_05476_ ), .Z(_05949_ ) );
OR2_X1 _13862_ ( .A1(_05949_ ), .A2(fanout_net_10 ), .ZN(_05950_ ) );
AND3_X1 _13863_ ( .A1(_05515_ ), .A2(_03977_ ), .A3(_05520_ ), .ZN(_05951_ ) );
NAND4_X1 _13864_ ( .A1(_05603_ ), .A2(_04196_ ), .A3(\mycsreg.CSReg[3][2] ), .A4(_04200_ ), .ZN(_05952_ ) );
NAND4_X1 _13865_ ( .A1(_05603_ ), .A2(_04216_ ), .A3(\mtvec [2] ), .A4(_05540_ ), .ZN(_05953_ ) );
NAND4_X1 _13866_ ( .A1(_05603_ ), .A2(\mycsreg.CSReg[0][2] ), .A3(_05540_ ), .A4(_04221_ ), .ZN(_05954_ ) );
NAND4_X1 _13867_ ( .A1(_05531_ ), .A2(_04191_ ), .A3(\mepc [2] ), .A4(_04200_ ), .ZN(_05955_ ) );
AND4_X1 _13868_ ( .A1(_05952_ ), .A2(_05953_ ), .A3(_05954_ ), .A4(_05955_ ), .ZN(_05956_ ) );
AOI211_X1 _13869_ ( .A(_04160_ ), .B(_05951_ ), .C1(_05527_ ), .C2(_05956_ ), .ZN(_05957_ ) );
NOR2_X1 _13870_ ( .A1(_05957_ ), .A2(_05552_ ), .ZN(_05958_ ) );
AOI211_X1 _13871_ ( .A(fanout_net_3 ), .B(_05948_ ), .C1(_05950_ ), .C2(_05958_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_28_D ) );
NAND2_X1 _13872_ ( .A1(_04101_ ), .A2(fanout_net_8 ), .ZN(_05959_ ) );
XOR2_X1 _13873_ ( .A(_04262_ ), .B(_04263_ ), .Z(_05960_ ) );
AOI21_X1 _13874_ ( .A(_05499_ ), .B1(_05960_ ), .B2(_05487_ ), .ZN(_05961_ ) );
NAND2_X1 _13875_ ( .A1(_05503_ ), .A2(\myexu.pc_jump_$_DFFE_PP0P__Q_29_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05962_ ) );
OAI211_X1 _13876_ ( .A(_05962_ ), .B(_05478_ ), .C1(_05510_ ), .C2(_05960_ ), .ZN(_05963_ ) );
NAND3_X1 _13877_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_05601_ ), .ZN(_05964_ ) );
NAND4_X1 _13878_ ( .A1(_05607_ ), .A2(_05672_ ), .A3(\mepc [1] ), .A4(_05610_ ), .ZN(_05965_ ) );
NAND4_X1 _13879_ ( .A1(_05709_ ), .A2(_04217_ ), .A3(\mtvec [1] ), .A4(_05649_ ), .ZN(_05966_ ) );
NAND4_X1 _13880_ ( .A1(_05709_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_05649_ ), .A4(_04222_ ), .ZN(_05967_ ) );
NAND4_X1 _13881_ ( .A1(_05709_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][1] ), .A4(_05712_ ), .ZN(_05968_ ) );
AND4_X1 _13882_ ( .A1(_05965_ ), .A2(_05966_ ), .A3(_05967_ ), .A4(_05968_ ), .ZN(_05969_ ) );
OAI21_X1 _13883_ ( .A(_05964_ ), .B1(_05617_ ), .B2(_05969_ ), .ZN(_05970_ ) );
AOI21_X1 _13884_ ( .A(_05880_ ), .B1(_05970_ ), .B2(fanout_net_10 ), .ZN(_05971_ ) );
AOI221_X1 _13885_ ( .A(fanout_net_3 ), .B1(_05959_ ), .B2(_05961_ ), .C1(_05963_ ), .C2(_05971_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_29_D ) );
XNOR2_X1 _13886_ ( .A(_05785_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_05972_ ) );
OR2_X1 _13887_ ( .A1(_05475_ ), .A2(_05972_ ), .ZN(_05973_ ) );
XOR2_X1 _13888_ ( .A(\ID_EX_pc [28] ), .B(\ID_EX_imm [28] ), .Z(_05974_ ) );
XNOR2_X1 _13889_ ( .A(_05771_ ), .B(_05974_ ), .ZN(_05975_ ) );
OAI211_X1 _13890_ ( .A(_05973_ ), .B(_05478_ ), .C1(_05510_ ), .C2(_05975_ ), .ZN(_05976_ ) );
NAND4_X1 _13891_ ( .A1(_05614_ ), .A2(\mycsreg.CSReg[0][28] ), .A3(_05541_ ), .A4(_04222_ ), .ZN(_05977_ ) );
NAND4_X1 _13892_ ( .A1(_05614_ ), .A2(_04196_ ), .A3(\mycsreg.CSReg[3][28] ), .A4(_05536_ ), .ZN(_05978_ ) );
NAND4_X1 _13893_ ( .A1(_05614_ ), .A2(_04191_ ), .A3(\mepc [28] ), .A4(_05536_ ), .ZN(_05979_ ) );
NAND3_X1 _13894_ ( .A1(_05977_ ), .A2(_05978_ ), .A3(_05979_ ), .ZN(_05980_ ) );
NAND4_X1 _13895_ ( .A1(_05614_ ), .A2(_05594_ ), .A3(\mtvec [28] ), .A4(_05541_ ), .ZN(_05981_ ) );
NAND2_X1 _13896_ ( .A1(_05670_ ), .A2(_05981_ ), .ZN(_05982_ ) );
OAI21_X1 _13897_ ( .A(_05645_ ), .B1(_05980_ ), .B2(_05982_ ), .ZN(_05983_ ) );
NAND3_X1 _13898_ ( .A1(_05515_ ), .A2(\EX_LS_result_csreg_mem [28] ), .A3(_05520_ ), .ZN(_05984_ ) );
AOI21_X1 _13899_ ( .A(_04159_ ), .B1(_05983_ ), .B2(_05984_ ), .ZN(_05985_ ) );
NOR2_X1 _13900_ ( .A1(_05985_ ), .A2(_05483_ ), .ZN(_05986_ ) );
NAND2_X1 _13901_ ( .A1(_03028_ ), .A2(fanout_net_8 ), .ZN(_05987_ ) );
BUF_X2 _13902_ ( .A(_05487_ ), .Z(_05988_ ) );
AOI21_X1 _13903_ ( .A(_05485_ ), .B1(_05975_ ), .B2(_05988_ ), .ZN(_05989_ ) );
AOI221_X1 _13904_ ( .A(fanout_net_3 ), .B1(_05976_ ), .B2(_05986_ ), .C1(_05987_ ), .C2(_05989_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_2_D ) );
XOR2_X1 _13905_ ( .A(\ID_EX_pc [0] ), .B(\ID_EX_imm [0] ), .Z(_05990_ ) );
AOI21_X1 _13906_ ( .A(_05500_ ), .B1(_05990_ ), .B2(_05628_ ), .ZN(_05991_ ) );
NAND2_X1 _13907_ ( .A1(_05511_ ), .A2(\myexu.pc_jump_$_DFFE_PP0P__Q_30_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_05992_ ) );
OAI211_X1 _13908_ ( .A(_05992_ ), .B(_05479_ ), .C1(_05511_ ), .C2(_05990_ ), .ZN(_05993_ ) );
NOR3_X1 _13909_ ( .A1(_04172_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_04181_ ), .ZN(_05994_ ) );
NAND3_X1 _13910_ ( .A1(_04214_ ), .A2(\mycsreg.CSReg[0][0] ), .A3(_04223_ ), .ZN(_05995_ ) );
NAND3_X1 _13911_ ( .A1(_04226_ ), .A2(\mepc [0] ), .A3(_05587_ ), .ZN(_05996_ ) );
NAND2_X1 _13912_ ( .A1(_05995_ ), .A2(_05996_ ), .ZN(_05997_ ) );
NOR2_X1 _13913_ ( .A1(_04210_ ), .A2(_05997_ ), .ZN(_05998_ ) );
NAND3_X1 _13914_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][0] ), .A3(_04207_ ), .ZN(_05999_ ) );
NAND2_X1 _13915_ ( .A1(_04198_ ), .A2(_05999_ ), .ZN(_06000_ ) );
AND3_X1 _13916_ ( .A1(_05593_ ), .A2(\mtvec [0] ), .A3(_05595_ ), .ZN(_06001_ ) );
NOR2_X1 _13917_ ( .A1(_06000_ ), .A2(_06001_ ), .ZN(_06002_ ) );
AOI21_X1 _13918_ ( .A(_05994_ ), .B1(_05998_ ), .B2(_06002_ ), .ZN(_06003_ ) );
AOI21_X1 _13919_ ( .A(_05552_ ), .B1(_06003_ ), .B2(fanout_net_10 ), .ZN(_06004_ ) );
AOI211_X1 _13920_ ( .A(fanout_net_3 ), .B(_05991_ ), .C1(_05993_ ), .C2(_06004_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_30_D ) );
AND2_X1 _13921_ ( .A1(_05764_ ), .A2(_05766_ ), .ZN(_06005_ ) );
NOR2_X1 _13922_ ( .A1(_06005_ ), .A2(_05768_ ), .ZN(_06006_ ) );
XNOR2_X1 _13923_ ( .A(_06006_ ), .B(_05765_ ), .ZN(_06007_ ) );
MUX2_X1 _13924_ ( .A(_06007_ ), .B(_03031_ ), .S(fanout_net_8 ), .Z(_06008_ ) );
NOR2_X1 _13925_ ( .A1(_06008_ ), .A2(_05500_ ), .ZN(_06009_ ) );
NAND2_X1 _13926_ ( .A1(_05505_ ), .A2(_05784_ ), .ZN(_06010_ ) );
NOR2_X1 _13927_ ( .A1(_06010_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_06011_ ) );
XNOR2_X1 _13928_ ( .A(_06011_ ), .B(\ID_EX_pc [27] ), .ZN(_06012_ ) );
AOI21_X1 _13929_ ( .A(fanout_net_10 ), .B1(_05504_ ), .B2(_06012_ ), .ZN(_06013_ ) );
OAI21_X1 _13930_ ( .A(_06013_ ), .B1(_05511_ ), .B2(_06007_ ), .ZN(_06014_ ) );
BUF_X2 _13931_ ( .A(_05483_ ), .Z(_06015_ ) );
BUF_X4 _13932_ ( .A(_06015_ ), .Z(_06016_ ) );
NAND3_X1 _13933_ ( .A1(_05516_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_05521_ ), .ZN(_06017_ ) );
NAND4_X1 _13934_ ( .A1(_05709_ ), .A2(_05594_ ), .A3(\mtvec [27] ), .A4(_05649_ ), .ZN(_06018_ ) );
AND2_X1 _13935_ ( .A1(_05670_ ), .A2(_06018_ ), .ZN(_06019_ ) );
NAND4_X1 _13936_ ( .A1(_05847_ ), .A2(\mycsreg.CSReg[0][27] ), .A3(_05542_ ), .A4(_05850_ ), .ZN(_06020_ ) );
NAND4_X1 _13937_ ( .A1(_05533_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][27] ), .A4(_05537_ ), .ZN(_06021_ ) );
NAND4_X1 _13938_ ( .A1(_05533_ ), .A2(_05546_ ), .A3(\mepc [27] ), .A4(_05537_ ), .ZN(_06022_ ) );
AND4_X1 _13939_ ( .A1(_06019_ ), .A2(_06020_ ), .A3(_06021_ ), .A4(_06022_ ), .ZN(_06023_ ) );
OAI21_X1 _13940_ ( .A(_06017_ ), .B1(_06023_ ), .B2(_05617_ ), .ZN(_06024_ ) );
AOI21_X1 _13941_ ( .A(_06016_ ), .B1(_06024_ ), .B2(fanout_net_10 ), .ZN(_06025_ ) );
AOI211_X1 _13942_ ( .A(fanout_net_4 ), .B(_06009_ ), .C1(_06014_ ), .C2(_06025_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_3_D ) );
XOR2_X1 _13943_ ( .A(_05764_ ), .B(_05766_ ), .Z(_06026_ ) );
NAND2_X1 _13944_ ( .A1(_06026_ ), .A2(_05627_ ), .ZN(_06027_ ) );
AOI21_X1 _13945_ ( .A(_05484_ ), .B1(_03032_ ), .B2(fanout_net_8 ), .ZN(_06028_ ) );
XNOR2_X1 _13946_ ( .A(_06010_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_06029_ ) );
NAND2_X1 _13947_ ( .A1(_05503_ ), .A2(_06029_ ), .ZN(_06030_ ) );
OAI211_X1 _13948_ ( .A(_06030_ ), .B(_05478_ ), .C1(_05510_ ), .C2(_06026_ ), .ZN(_06031_ ) );
NAND4_X1 _13949_ ( .A1(_05532_ ), .A2(_04191_ ), .A3(\mepc [26] ), .A4(_05536_ ), .ZN(_06032_ ) );
NAND4_X1 _13950_ ( .A1(_05532_ ), .A2(_04216_ ), .A3(\mtvec [26] ), .A4(_05540_ ), .ZN(_06033_ ) );
NAND4_X1 _13951_ ( .A1(_05603_ ), .A2(\mycsreg.CSReg[0][26] ), .A3(_05540_ ), .A4(_04221_ ), .ZN(_06034_ ) );
NAND4_X1 _13952_ ( .A1(_05603_ ), .A2(_04196_ ), .A3(\mycsreg.CSReg[3][26] ), .A4(_04200_ ), .ZN(_06035_ ) );
AND4_X1 _13953_ ( .A1(_06032_ ), .A2(_06033_ ), .A3(_06034_ ), .A4(_06035_ ), .ZN(_06036_ ) );
OR2_X1 _13954_ ( .A1(_05523_ ), .A2(_06036_ ), .ZN(_06037_ ) );
NAND3_X1 _13955_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [26] ), .A3(_05601_ ), .ZN(_06038_ ) );
AOI21_X1 _13956_ ( .A(_04159_ ), .B1(_06037_ ), .B2(_06038_ ), .ZN(_06039_ ) );
NOR2_X1 _13957_ ( .A1(_06039_ ), .A2(_05678_ ), .ZN(_06040_ ) );
AOI221_X1 _13958_ ( .A(fanout_net_4 ), .B1(_06027_ ), .B2(_06028_ ), .C1(_06031_ ), .C2(_06040_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_4_D ) );
OAI21_X1 _13959_ ( .A(_05551_ ), .B1(_03035_ ), .B2(_05988_ ), .ZN(_06041_ ) );
NOR2_X1 _13960_ ( .A1(_05742_ ), .A2(_05763_ ), .ZN(_06042_ ) );
XNOR2_X1 _13961_ ( .A(_05762_ ), .B(_06042_ ), .ZN(_06043_ ) );
AOI21_X1 _13962_ ( .A(_06041_ ), .B1(_05628_ ), .B2(_06043_ ), .ZN(_06044_ ) );
NOR4_X1 _13963_ ( .A1(_05577_ ), .A2(_04287_ ), .A3(_05697_ ), .A4(_05578_ ), .ZN(_06045_ ) );
NAND3_X1 _13964_ ( .A1(_06045_ ), .A2(\ID_EX_pc [16] ), .A3(\ID_EX_pc [14] ), .ZN(_06046_ ) );
NOR2_X1 _13965_ ( .A1(_06046_ ), .A2(_05576_ ), .ZN(_06047_ ) );
NAND4_X1 _13966_ ( .A1(_06047_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [19] ), .A4(\ID_EX_pc [18] ), .ZN(_06048_ ) );
INV_X1 _13967_ ( .A(\ID_EX_pc [20] ), .ZN(_06049_ ) );
INV_X1 _13968_ ( .A(\ID_EX_pc [23] ), .ZN(_06050_ ) );
NOR3_X1 _13969_ ( .A1(_06048_ ), .A2(_06049_ ), .A3(_06050_ ), .ZN(_06051_ ) );
NAND3_X1 _13970_ ( .A1(_06051_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_pc [22] ), .ZN(_06052_ ) );
INV_X1 _13971_ ( .A(\ID_EX_pc [25] ), .ZN(_06053_ ) );
XNOR2_X1 _13972_ ( .A(_06052_ ), .B(_06053_ ), .ZN(_06054_ ) );
NAND2_X1 _13973_ ( .A1(_05511_ ), .A2(_06054_ ), .ZN(_06055_ ) );
OAI211_X1 _13974_ ( .A(_06055_ ), .B(_05479_ ), .C1(_05511_ ), .C2(_06043_ ), .ZN(_06056_ ) );
NAND3_X1 _13975_ ( .A1(_05516_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_05521_ ), .ZN(_06057_ ) );
AND4_X1 _13976_ ( .A1(\mycsreg.CSReg[0][25] ), .A2(_05847_ ), .A3(_05542_ ), .A4(_05850_ ), .ZN(_06058_ ) );
NAND4_X1 _13977_ ( .A1(_05847_ ), .A2(_05595_ ), .A3(\mtvec [25] ), .A4(_05542_ ), .ZN(_06059_ ) );
NAND4_X1 _13978_ ( .A1(_05847_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][25] ), .A4(_05537_ ), .ZN(_06060_ ) );
NAND2_X1 _13979_ ( .A1(_06059_ ), .A2(_06060_ ), .ZN(_06061_ ) );
AOI211_X1 _13980_ ( .A(_06058_ ), .B(_06061_ ), .C1(_05655_ ), .C2(\mepc [25] ), .ZN(_06062_ ) );
OAI21_X1 _13981_ ( .A(_06057_ ), .B1(_06062_ ), .B2(_05617_ ), .ZN(_06063_ ) );
AOI21_X1 _13982_ ( .A(_06016_ ), .B1(_06063_ ), .B2(fanout_net_10 ), .ZN(_06064_ ) );
AOI211_X1 _13983_ ( .A(fanout_net_4 ), .B(_06044_ ), .C1(_06056_ ), .C2(_06064_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_5_D ) );
NAND3_X1 _13984_ ( .A1(_03036_ ), .A2(fanout_net_9 ), .A3(_02809_ ), .ZN(_06065_ ) );
OR3_X1 _13985_ ( .A1(_05751_ ), .A2(_05759_ ), .A3(_05744_ ), .ZN(_06066_ ) );
AND2_X1 _13986_ ( .A1(_06066_ ), .A2(_05760_ ), .ZN(_06067_ ) );
AOI21_X1 _13987_ ( .A(_05484_ ), .B1(_06067_ ), .B2(_05487_ ), .ZN(_06068_ ) );
AND3_X1 _13988_ ( .A1(_04234_ ), .A2(_04239_ ), .A3(_05782_ ), .ZN(_06069_ ) );
AND3_X1 _13989_ ( .A1(_06069_ ), .A2(\ID_EX_pc [24] ), .A3(_05783_ ), .ZN(_06070_ ) );
AOI21_X1 _13990_ ( .A(\ID_EX_pc [24] ), .B1(_06069_ ), .B2(_05783_ ), .ZN(_06071_ ) );
OAI21_X1 _13991_ ( .A(_05503_ ), .B1(_06070_ ), .B2(_06071_ ), .ZN(_06072_ ) );
OAI211_X1 _13992_ ( .A(_06072_ ), .B(_05478_ ), .C1(_05510_ ), .C2(_06067_ ), .ZN(_06073_ ) );
NAND3_X1 _13993_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_05601_ ), .ZN(_06074_ ) );
NAND4_X1 _13994_ ( .A1(_05648_ ), .A2(\mycsreg.CSReg[0][24] ), .A3(_05649_ ), .A4(_04222_ ), .ZN(_06075_ ) );
NAND4_X1 _13995_ ( .A1(_05648_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][24] ), .A4(_05712_ ), .ZN(_06076_ ) );
NAND4_X1 _13996_ ( .A1(_05648_ ), .A2(_05672_ ), .A3(\mepc [24] ), .A4(_05712_ ), .ZN(_06077_ ) );
NAND3_X1 _13997_ ( .A1(_06075_ ), .A2(_06076_ ), .A3(_06077_ ), .ZN(_06078_ ) );
AND4_X1 _13998_ ( .A1(\mtvec [24] ), .A2(_05614_ ), .A3(_05594_ ), .A4(_05541_ ), .ZN(_06079_ ) );
NOR4_X1 _13999_ ( .A1(_06078_ ), .A2(_06079_ ), .A3(_05613_ ), .A4(_05526_ ), .ZN(_06080_ ) );
OAI21_X1 _14000_ ( .A(_06074_ ), .B1(_06080_ ), .B2(_05617_ ), .ZN(_06081_ ) );
AOI21_X1 _14001_ ( .A(_05880_ ), .B1(_06081_ ), .B2(fanout_net_10 ), .ZN(_06082_ ) );
AOI221_X1 _14002_ ( .A(fanout_net_4 ), .B1(_06065_ ), .B2(_06068_ ), .C1(_06073_ ), .C2(_06082_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_6_D ) );
AOI21_X1 _14003_ ( .A(_04320_ ), .B1(_04310_ ), .B2(_04317_ ), .ZN(_06083_ ) );
OR2_X1 _14004_ ( .A1(_06083_ ), .A2(_05756_ ), .ZN(_06084_ ) );
AOI21_X1 _14005_ ( .A(_05748_ ), .B1(_06084_ ), .B2(_05755_ ), .ZN(_06085_ ) );
NOR2_X1 _14006_ ( .A1(\ID_EX_pc [22] ), .A2(\ID_EX_imm [22] ), .ZN(_06086_ ) );
NOR3_X1 _14007_ ( .A1(_06085_ ), .A2(_05752_ ), .A3(_06086_ ), .ZN(_06087_ ) );
NOR2_X1 _14008_ ( .A1(_06087_ ), .A2(_05752_ ), .ZN(_06088_ ) );
XNOR2_X1 _14009_ ( .A(_06088_ ), .B(_05745_ ), .ZN(_06089_ ) );
NAND2_X1 _14010_ ( .A1(_06089_ ), .A2(_05627_ ), .ZN(_06090_ ) );
AOI21_X1 _14011_ ( .A(_05484_ ), .B1(_03040_ ), .B2(fanout_net_9 ), .ZN(_06091_ ) );
INV_X1 _14012_ ( .A(_06069_ ), .ZN(_06092_ ) );
NOR2_X1 _14013_ ( .A1(_06092_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_06093_ ) );
XNOR2_X1 _14014_ ( .A(_06093_ ), .B(\ID_EX_pc [23] ), .ZN(_06094_ ) );
NAND2_X1 _14015_ ( .A1(_05503_ ), .A2(_06094_ ), .ZN(_06095_ ) );
OAI211_X1 _14016_ ( .A(_06095_ ), .B(_05478_ ), .C1(_05510_ ), .C2(_06089_ ), .ZN(_06096_ ) );
NAND3_X1 _14017_ ( .A1(_05600_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_05601_ ), .ZN(_06097_ ) );
NAND4_X1 _14018_ ( .A1(_05607_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_05605_ ), .A4(_05590_ ), .ZN(_06098_ ) );
NAND4_X1 _14019_ ( .A1(_05709_ ), .A2(_05594_ ), .A3(\mtvec [23] ), .A4(_05649_ ), .ZN(_06099_ ) );
NAND4_X1 _14020_ ( .A1(_05709_ ), .A2(_05672_ ), .A3(\mepc [23] ), .A4(_05712_ ), .ZN(_06100_ ) );
NAND4_X1 _14021_ ( .A1(_05709_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][23] ), .A4(_05712_ ), .ZN(_06101_ ) );
AND4_X1 _14022_ ( .A1(_06098_ ), .A2(_06099_ ), .A3(_06100_ ), .A4(_06101_ ), .ZN(_06102_ ) );
OAI21_X1 _14023_ ( .A(_06097_ ), .B1(_05617_ ), .B2(_06102_ ), .ZN(_06103_ ) );
AOI21_X1 _14024_ ( .A(_05880_ ), .B1(_06103_ ), .B2(fanout_net_10 ), .ZN(_06104_ ) );
AOI221_X1 _14025_ ( .A(fanout_net_4 ), .B1(_06090_ ), .B2(_06091_ ), .C1(_06096_ ), .C2(_06104_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_7_D ) );
XNOR2_X1 _14026_ ( .A(_06085_ ), .B(_05746_ ), .ZN(_06105_ ) );
NAND2_X1 _14027_ ( .A1(_06105_ ), .A2(_05627_ ), .ZN(_06106_ ) );
AOI21_X1 _14028_ ( .A(_05484_ ), .B1(_03041_ ), .B2(fanout_net_9 ), .ZN(_06107_ ) );
XNOR2_X1 _14029_ ( .A(_06069_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_06108_ ) );
OR2_X1 _14030_ ( .A1(_05475_ ), .A2(_06108_ ), .ZN(_06109_ ) );
OAI211_X1 _14031_ ( .A(_06109_ ), .B(_05478_ ), .C1(_05510_ ), .C2(_06105_ ), .ZN(_06110_ ) );
OR3_X1 _14032_ ( .A1(_04171_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_04180_ ), .ZN(_06111_ ) );
NAND3_X1 _14033_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_05587_ ), .ZN(_06112_ ) );
NAND3_X1 _14034_ ( .A1(_04226_ ), .A2(\mepc [22] ), .A3(_05587_ ), .ZN(_06113_ ) );
NAND3_X1 _14035_ ( .A1(_04213_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_05850_ ), .ZN(_06114_ ) );
NAND4_X1 _14036_ ( .A1(_05586_ ), .A2(_06112_ ), .A3(_06113_ ), .A4(_06114_ ), .ZN(_06115_ ) );
NAND3_X1 _14037_ ( .A1(_04213_ ), .A2(\mtvec [22] ), .A3(_04217_ ), .ZN(_06116_ ) );
OAI21_X1 _14038_ ( .A(_06116_ ), .B1(_04171_ ), .B2(_04180_ ), .ZN(_06117_ ) );
OAI211_X1 _14039_ ( .A(_06111_ ), .B(fanout_net_10 ), .C1(_06115_ ), .C2(_06117_ ), .ZN(_06118_ ) );
AND2_X1 _14040_ ( .A1(_06118_ ), .A2(_05499_ ), .ZN(_06119_ ) );
AOI221_X4 _14041_ ( .A(fanout_net_4 ), .B1(_06106_ ), .B2(_06107_ ), .C1(_06110_ ), .C2(_06119_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_8_D ) );
INV_X1 _14042_ ( .A(_04210_ ), .ZN(_06120_ ) );
NAND3_X1 _14043_ ( .A1(_05593_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_05850_ ), .ZN(_06121_ ) );
NAND3_X1 _14044_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][21] ), .A3(_05587_ ), .ZN(_06122_ ) );
NAND3_X1 _14045_ ( .A1(_04226_ ), .A2(\mepc [21] ), .A3(_05587_ ), .ZN(_06123_ ) );
AND4_X1 _14046_ ( .A1(_04193_ ), .A2(_06121_ ), .A3(_06122_ ), .A4(_06123_ ), .ZN(_06124_ ) );
AND3_X1 _14047_ ( .A1(_05593_ ), .A2(\mtvec [21] ), .A3(_05595_ ), .ZN(_06125_ ) );
INV_X1 _14048_ ( .A(_06125_ ), .ZN(_06126_ ) );
NAND3_X1 _14049_ ( .A1(_06120_ ), .A2(_06124_ ), .A3(_06126_ ), .ZN(_06127_ ) );
NOR3_X1 _14050_ ( .A1(_04172_ ), .A2(\EX_LS_result_csreg_mem [21] ), .A3(_04181_ ), .ZN(_06128_ ) );
INV_X1 _14051_ ( .A(_06128_ ), .ZN(_06129_ ) );
NAND3_X1 _14052_ ( .A1(_06127_ ), .A2(fanout_net_10 ), .A3(_06129_ ), .ZN(_06130_ ) );
INV_X1 _14053_ ( .A(_06130_ ), .ZN(_06131_ ) );
INV_X1 _14054_ ( .A(_04240_ ), .ZN(_06132_ ) );
NOR2_X1 _14055_ ( .A1(_06132_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_06133_ ) );
INV_X1 _14056_ ( .A(\ID_EX_pc [21] ), .ZN(_06134_ ) );
XNOR2_X1 _14057_ ( .A(_06133_ ), .B(_06134_ ), .ZN(_06135_ ) );
XOR2_X1 _14058_ ( .A(_06084_ ), .B(_05750_ ), .Z(_06136_ ) );
MUX2_X1 _14059_ ( .A(_06135_ ), .B(_06136_ ), .S(_05476_ ), .Z(_06137_ ) );
AOI21_X1 _14060_ ( .A(_06131_ ), .B1(_06137_ ), .B2(_05479_ ), .ZN(_06138_ ) );
AOI21_X1 _14061_ ( .A(_05485_ ), .B1(_06136_ ), .B2(_05488_ ), .ZN(_06139_ ) );
OR2_X1 _14062_ ( .A1(_06139_ ), .A2(fanout_net_4 ), .ZN(_06140_ ) );
OR3_X1 _14063_ ( .A1(_03000_ ), .A2(fanout_net_4 ), .A3(_05488_ ), .ZN(_06141_ ) );
AOI22_X1 _14064_ ( .A1(_06138_ ), .A2(_05486_ ), .B1(_06140_ ), .B2(_06141_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_9_D ) );
OR3_X1 _14065_ ( .A1(_04170_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_04179_ ), .ZN(_06142_ ) );
NAND3_X1 _14066_ ( .A1(_04213_ ), .A2(\mtvec [30] ), .A3(_05594_ ), .ZN(_06143_ ) );
NAND3_X1 _14067_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][30] ), .A3(_04206_ ), .ZN(_06144_ ) );
NAND3_X1 _14068_ ( .A1(_04193_ ), .A2(_06143_ ), .A3(_06144_ ), .ZN(_06145_ ) );
NAND3_X1 _14069_ ( .A1(_04225_ ), .A2(\mepc [30] ), .A3(_04206_ ), .ZN(_06146_ ) );
NAND3_X1 _14070_ ( .A1(_04212_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_04222_ ), .ZN(_06147_ ) );
OAI211_X1 _14071_ ( .A(_06146_ ), .B(_06147_ ), .C1(_04171_ ), .C2(_04180_ ), .ZN(_06148_ ) );
OAI211_X1 _14072_ ( .A(_06142_ ), .B(fanout_net_10 ), .C1(_06145_ ), .C2(_06148_ ), .ZN(_06149_ ) );
INV_X1 _14073_ ( .A(_06149_ ), .ZN(_06150_ ) );
NOR2_X1 _14074_ ( .A1(_05580_ ), .A2(_05581_ ), .ZN(_06151_ ) );
AND3_X1 _14075_ ( .A1(_06151_ ), .A2(\ID_EX_pc [17] ), .A3(_04235_ ), .ZN(_06152_ ) );
AND3_X1 _14076_ ( .A1(_06152_ ), .A2(\ID_EX_pc [21] ), .A3(\ID_EX_pc [20] ), .ZN(_06153_ ) );
AND3_X1 _14077_ ( .A1(_06153_ ), .A2(\ID_EX_pc [24] ), .A3(_05783_ ), .ZN(_06154_ ) );
AND3_X1 _14078_ ( .A1(_06154_ ), .A2(\ID_EX_pc [25] ), .A3(_05781_ ), .ZN(_06155_ ) );
AND3_X1 _14079_ ( .A1(_06155_ ), .A2(\ID_EX_pc [29] ), .A3(\ID_EX_pc [28] ), .ZN(_06156_ ) );
XNOR2_X1 _14080_ ( .A(_06156_ ), .B(\myexu.result_reg_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_06157_ ) );
AND2_X1 _14081_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_06158_ ) );
OR2_X1 _14082_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_imm [29] ), .ZN(_06159_ ) );
AOI21_X1 _14083_ ( .A(_06158_ ), .B1(_05775_ ), .B2(_06159_ ), .ZN(_06160_ ) );
XNOR2_X1 _14084_ ( .A(\ID_EX_pc [30] ), .B(\ID_EX_imm [30] ), .ZN(_06161_ ) );
XOR2_X1 _14085_ ( .A(_06160_ ), .B(_06161_ ), .Z(_06162_ ) );
MUX2_X1 _14086_ ( .A(_06157_ ), .B(_06162_ ), .S(_05475_ ), .Z(_06163_ ) );
AOI21_X1 _14087_ ( .A(_06150_ ), .B1(_06163_ ), .B2(_05478_ ), .ZN(_06164_ ) );
OR2_X1 _14088_ ( .A1(_02994_ ), .A2(_05627_ ), .ZN(_06165_ ) );
AOI21_X1 _14089_ ( .A(_05499_ ), .B1(_06162_ ), .B2(_05988_ ), .ZN(_06166_ ) );
AOI221_X1 _14090_ ( .A(fanout_net_4 ), .B1(_05485_ ), .B2(_06164_ ), .C1(_06165_ ), .C2(_06166_ ), .ZN(\myexu.pc_jump_$_DFFE_PP0P__Q_D ) );
NOR2_X1 _14091_ ( .A1(_06160_ ), .A2(_06161_ ), .ZN(_06167_ ) );
AND2_X1 _14092_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_imm [30] ), .ZN(_06168_ ) );
OR2_X1 _14093_ ( .A1(_06167_ ), .A2(_06168_ ), .ZN(_06169_ ) );
XNOR2_X1 _14094_ ( .A(\ID_EX_pc [31] ), .B(\ID_EX_imm [31] ), .ZN(_06170_ ) );
XNOR2_X1 _14095_ ( .A(_06169_ ), .B(_06170_ ), .ZN(_06171_ ) );
OAI21_X1 _14096_ ( .A(_05678_ ), .B1(_06171_ ), .B2(fanout_net_9 ), .ZN(_06172_ ) );
AOI21_X1 _14097_ ( .A(_06172_ ), .B1(_02990_ ), .B2(fanout_net_9 ), .ZN(_06173_ ) );
OR3_X1 _14098_ ( .A1(_04170_ ), .A2(\EX_LS_result_csreg_mem [31] ), .A3(_04179_ ), .ZN(_06174_ ) );
NAND3_X1 _14099_ ( .A1(_04212_ ), .A2(\mtvec [31] ), .A3(_04216_ ), .ZN(_06175_ ) );
NAND3_X1 _14100_ ( .A1(_04212_ ), .A2(\mycsreg.CSReg[0][31] ), .A3(_04221_ ), .ZN(_06176_ ) );
NAND3_X1 _14101_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][31] ), .A3(_04205_ ), .ZN(_06177_ ) );
NAND3_X1 _14102_ ( .A1(_04225_ ), .A2(\mepc [31] ), .A3(_04205_ ), .ZN(_06178_ ) );
NAND4_X1 _14103_ ( .A1(_06175_ ), .A2(_06176_ ), .A3(_06177_ ), .A4(_06178_ ), .ZN(_06179_ ) );
OAI21_X1 _14104_ ( .A(_06174_ ), .B1(_04210_ ), .B2(_06179_ ), .ZN(_06180_ ) );
INV_X1 _14105_ ( .A(_06180_ ), .ZN(_06181_ ) );
INV_X1 _14106_ ( .A(_06156_ ), .ZN(_06182_ ) );
NOR2_X1 _14107_ ( .A1(_06182_ ), .A2(\myexu.result_reg_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ), .ZN(_06183_ ) );
INV_X1 _14108_ ( .A(\ID_EX_pc [31] ), .ZN(_06184_ ) );
XNOR2_X1 _14109_ ( .A(_06183_ ), .B(_06184_ ), .ZN(_06185_ ) );
MUX2_X1 _14110_ ( .A(_06185_ ), .B(_06171_ ), .S(_05475_ ), .Z(_06186_ ) );
MUX2_X1 _14111_ ( .A(_06181_ ), .B(_06186_ ), .S(_04159_ ), .Z(_06187_ ) );
AND2_X1 _14112_ ( .A1(_06187_ ), .A2(_05485_ ), .ZN(_06188_ ) );
OR3_X1 _14113_ ( .A1(_06173_ ), .A2(fanout_net_4 ), .A3(_06188_ ), .ZN(\myexu.pc_jump_$_DFFE_PP1P__Q_D ) );
NOR2_X1 _14114_ ( .A1(_06134_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_10_D ) );
NOR2_X1 _14115_ ( .A1(_06049_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_11_D ) );
INV_X1 _14116_ ( .A(\ID_EX_pc [19] ), .ZN(_06189_ ) );
NOR2_X1 _14117_ ( .A1(_06189_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_12_D ) );
INV_X1 _14118_ ( .A(\ID_EX_pc [18] ), .ZN(_06190_ ) );
NOR2_X1 _14119_ ( .A1(_06190_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_13_D ) );
NOR2_X1 _14120_ ( .A1(_05576_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_14_D ) );
NOR2_X1 _14121_ ( .A1(_05581_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_15_D ) );
NOR2_X1 _14122_ ( .A1(_04287_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_16_D ) );
INV_X1 _14123_ ( .A(\ID_EX_pc [14] ), .ZN(_06191_ ) );
NOR2_X1 _14124_ ( .A1(_06191_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_17_D ) );
NOR2_X1 _14125_ ( .A1(_05697_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_18_D ) );
NOR2_X1 _14126_ ( .A1(_05578_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_19_D ) );
AND2_X1 _14127_ ( .A1(_01735_ ), .A2(\ID_EX_pc [30] ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_1_D ) );
INV_X1 _14128_ ( .A(\ID_EX_pc [11] ), .ZN(_06192_ ) );
NOR2_X1 _14129_ ( .A1(_06192_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_20_D ) );
AND2_X1 _14130_ ( .A1(_01564_ ), .A2(\ID_EX_pc [10] ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_21_D ) );
NOR2_X1 _14131_ ( .A1(_05820_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_22_D ) );
NOR2_X1 _14132_ ( .A1(_05839_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_23_D ) );
INV_X1 _14133_ ( .A(\ID_EX_pc [7] ), .ZN(_06193_ ) );
NOR2_X1 _14134_ ( .A1(_06193_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_24_D ) );
INV_X1 _14135_ ( .A(\ID_EX_pc [6] ), .ZN(_06194_ ) );
NOR2_X1 _14136_ ( .A1(_06194_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_25_D ) );
AND2_X1 _14137_ ( .A1(_01564_ ), .A2(\ID_EX_pc [5] ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_26_D ) );
INV_X1 _14138_ ( .A(\ID_EX_pc [4] ), .ZN(_06195_ ) );
NOR2_X1 _14139_ ( .A1(_06195_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_27_D ) );
INV_X1 _14140_ ( .A(\ID_EX_pc [3] ), .ZN(_06196_ ) );
NOR2_X1 _14141_ ( .A1(_06196_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_28_D ) );
INV_X1 _14142_ ( .A(\ID_EX_pc [2] ), .ZN(_06197_ ) );
NOR2_X1 _14143_ ( .A1(_06197_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_29_D ) );
AND2_X1 _14144_ ( .A1(_01564_ ), .A2(\ID_EX_pc [29] ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_2_D ) );
NOR2_X1 _14145_ ( .A1(_04265_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_30_D ) );
INV_X1 _14146_ ( .A(\ID_EX_pc [0] ), .ZN(_06198_ ) );
NOR2_X1 _14147_ ( .A1(_06198_ ), .A2(fanout_net_4 ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_31_D ) );
INV_X1 _14148_ ( .A(\ID_EX_pc [28] ), .ZN(_06199_ ) );
NOR2_X1 _14149_ ( .A1(_06199_ ), .A2(reset ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_3_D ) );
AND2_X1 _14150_ ( .A1(_01564_ ), .A2(\ID_EX_pc [27] ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_4_D ) );
INV_X1 _14151_ ( .A(\ID_EX_pc [26] ), .ZN(_06200_ ) );
NOR2_X1 _14152_ ( .A1(_06200_ ), .A2(reset ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_5_D ) );
NOR2_X1 _14153_ ( .A1(_06053_ ), .A2(reset ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_6_D ) );
INV_X1 _14154_ ( .A(\ID_EX_pc [24] ), .ZN(_06201_ ) );
NOR2_X1 _14155_ ( .A1(_06201_ ), .A2(reset ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_7_D ) );
NOR2_X1 _14156_ ( .A1(_06050_ ), .A2(reset ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_8_D ) );
INV_X1 _14157_ ( .A(\ID_EX_pc [22] ), .ZN(_06202_ ) );
NOR2_X1 _14158_ ( .A1(_06202_ ), .A2(reset ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_9_D ) );
NOR2_X1 _14159_ ( .A1(_06184_ ), .A2(reset ), .ZN(\myexu.pc_out_$_DFFE_PP0P__Q_D ) );
OAI211_X1 _14160_ ( .A(_02992_ ), .B(_04097_ ), .C1(_05988_ ), .C2(\ID_EX_imm [21] ), .ZN(_06203_ ) );
INV_X1 _14161_ ( .A(_02793_ ), .ZN(_06204_ ) );
AOI21_X1 _14162_ ( .A(_06203_ ), .B1(_06204_ ), .B2(_05628_ ), .ZN(_06205_ ) );
BUF_X4 _14163_ ( .A(_05468_ ), .Z(_06206_ ) );
BUF_X4 _14164_ ( .A(_06206_ ), .Z(_06207_ ) );
NOR2_X1 _14165_ ( .A1(_04210_ ), .A2(_06125_ ), .ZN(_06208_ ) );
AOI21_X1 _14166_ ( .A(_06128_ ), .B1(_06208_ ), .B2(_06124_ ), .ZN(_06209_ ) );
OAI21_X1 _14167_ ( .A(_06205_ ), .B1(_06207_ ), .B2(_06209_ ), .ZN(_06210_ ) );
NOR2_X1 _14168_ ( .A1(_05379_ ), .A2(\ID_EX_typ [2] ), .ZN(_06211_ ) );
BUF_X4 _14169_ ( .A(_06211_ ), .Z(_06212_ ) );
BUF_X4 _14170_ ( .A(_06212_ ), .Z(_06213_ ) );
NAND4_X1 _14171_ ( .A1(_05534_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][21] ), .A4(_05538_ ), .ZN(_06214_ ) );
AND2_X1 _14172_ ( .A1(_05671_ ), .A2(_06214_ ), .ZN(_06215_ ) );
NAND4_X1 _14173_ ( .A1(_05534_ ), .A2(_04218_ ), .A3(\mtvec [21] ), .A4(_05543_ ), .ZN(_06216_ ) );
NAND4_X1 _14174_ ( .A1(_05534_ ), .A2(_05546_ ), .A3(\mepc [21] ), .A4(_05538_ ), .ZN(_06217_ ) );
NAND4_X1 _14175_ ( .A1(_05534_ ), .A2(\mycsreg.CSReg[0][21] ), .A3(_05543_ ), .A4(_04223_ ), .ZN(_06218_ ) );
AND3_X1 _14176_ ( .A1(_06216_ ), .A2(_06217_ ), .A3(_06218_ ), .ZN(_06219_ ) );
AOI22_X1 _14177_ ( .A1(_06215_ ), .A2(_06219_ ), .B1(_05516_ ), .B2(_05521_ ), .ZN(_06220_ ) );
AND3_X1 _14178_ ( .A1(_05516_ ), .A2(\EX_LS_result_csreg_mem [21] ), .A3(_05521_ ), .ZN(_06221_ ) );
OAI211_X1 _14179_ ( .A(_04126_ ), .B(_06213_ ), .C1(_06220_ ), .C2(_06221_ ), .ZN(_06222_ ) );
MUX2_X1 _14180_ ( .A(_06134_ ), .B(_04634_ ), .S(_04133_ ), .Z(_06223_ ) );
OAI211_X1 _14181_ ( .A(_06210_ ), .B(_06222_ ), .C1(_04127_ ), .C2(_06223_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ) );
BUF_X4 _14182_ ( .A(_04105_ ), .Z(_06224_ ) );
AND3_X1 _14183_ ( .A1(_05515_ ), .A2(\EX_LS_result_csreg_mem [20] ), .A3(_05520_ ), .ZN(_06225_ ) );
NAND4_X1 _14184_ ( .A1(_05604_ ), .A2(\mycsreg.CSReg[0][20] ), .A3(_05605_ ), .A4(_05590_ ), .ZN(_06226_ ) );
NAND4_X1 _14185_ ( .A1(_05604_ ), .A2(_05672_ ), .A3(\mepc [20] ), .A4(_05610_ ), .ZN(_06227_ ) );
NAND4_X1 _14186_ ( .A1(_05607_ ), .A2(_05609_ ), .A3(\mycsreg.CSReg[3][20] ), .A4(_05610_ ), .ZN(_06228_ ) );
AND3_X1 _14187_ ( .A1(_06226_ ), .A2(_06227_ ), .A3(_06228_ ), .ZN(_06229_ ) );
NAND4_X1 _14188_ ( .A1(_05847_ ), .A2(_05595_ ), .A3(\mtvec [20] ), .A4(_05542_ ), .ZN(_06230_ ) );
NAND4_X1 _14189_ ( .A1(_06229_ ), .A2(_06230_ ), .A3(_05671_ ), .A4(_05647_ ), .ZN(_06231_ ) );
AOI211_X1 _14190_ ( .A(_05468_ ), .B(_06225_ ), .C1(_05646_ ), .C2(_06231_ ), .ZN(_06232_ ) );
NAND2_X1 _14191_ ( .A1(_02770_ ), .A2(_05817_ ), .ZN(_06233_ ) );
NAND2_X1 _14192_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [20] ), .ZN(_06234_ ) );
AOI21_X1 _14193_ ( .A(_06232_ ), .B1(_06233_ ), .B2(_06234_ ), .ZN(_06235_ ) );
INV_X1 _14194_ ( .A(_06211_ ), .ZN(_06236_ ) );
BUF_X4 _14195_ ( .A(_06236_ ), .Z(_06237_ ) );
AOI211_X1 _14196_ ( .A(_04182_ ), .B(_06237_ ), .C1(_04211_ ), .C2(_04228_ ), .ZN(_06238_ ) );
OAI21_X1 _14197_ ( .A(_06224_ ), .B1(_06235_ ), .B2(_06238_ ), .ZN(_06239_ ) );
BUF_X4 _14198_ ( .A(_04105_ ), .Z(_06240_ ) );
BUF_X4 _14199_ ( .A(_06240_ ), .Z(_06241_ ) );
BUF_X4 _14200_ ( .A(_04132_ ), .Z(_06242_ ) );
BUF_X4 _14201_ ( .A(_06242_ ), .Z(_06243_ ) );
MUX2_X1 _14202_ ( .A(_06049_ ), .B(_04659_ ), .S(_06243_ ), .Z(_06244_ ) );
OAI21_X1 _14203_ ( .A(_06239_ ), .B1(_06241_ ), .B2(_06244_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _14204_ ( .A1(_05593_ ), .A2(\mycsreg.CSReg[0][19] ), .A3(_05850_ ), .ZN(_06245_ ) );
OAI21_X1 _14205_ ( .A(_06245_ ), .B1(_04171_ ), .B2(_04180_ ), .ZN(_06246_ ) );
NAND3_X1 _14206_ ( .A1(_04213_ ), .A2(\mtvec [19] ), .A3(_04217_ ), .ZN(_06247_ ) );
NAND3_X1 _14207_ ( .A1(_04226_ ), .A2(\mepc [19] ), .A3(_05587_ ), .ZN(_06248_ ) );
NAND3_X1 _14208_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][19] ), .A3(_05587_ ), .ZN(_06249_ ) );
NAND4_X1 _14209_ ( .A1(_04198_ ), .A2(_06247_ ), .A3(_06248_ ), .A4(_06249_ ), .ZN(_06250_ ) );
NOR2_X1 _14210_ ( .A1(_06246_ ), .A2(_06250_ ), .ZN(_06251_ ) );
NOR3_X1 _14211_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_05687_ ), .ZN(_06252_ ) );
NOR2_X1 _14212_ ( .A1(_06251_ ), .A2(_06252_ ), .ZN(_06253_ ) );
BUF_X4 _14213_ ( .A(_05487_ ), .Z(_06254_ ) );
OAI22_X1 _14214_ ( .A1(_06253_ ), .A2(_06206_ ), .B1(_06254_ ), .B2(\ID_EX_imm [19] ), .ZN(_06255_ ) );
AOI21_X1 _14215_ ( .A(_06255_ ), .B1(_05421_ ), .B2(_05628_ ), .ZN(_06256_ ) );
OR3_X1 _14216_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [19] ), .A3(_05687_ ), .ZN(_06257_ ) );
OAI211_X1 _14217_ ( .A(_06257_ ), .B(_06212_ ), .C1(_06250_ ), .C2(_06246_ ), .ZN(_06258_ ) );
INV_X1 _14218_ ( .A(_06258_ ), .ZN(_06259_ ) );
OAI21_X1 _14219_ ( .A(_06224_ ), .B1(_06256_ ), .B2(_06259_ ), .ZN(_06260_ ) );
MUX2_X1 _14220_ ( .A(_06189_ ), .B(_04707_ ), .S(_06243_ ), .Z(_06261_ ) );
OAI21_X1 _14221_ ( .A(_06260_ ), .B1(_06241_ ), .B2(_06261_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _14222_ ( .A1(_04213_ ), .A2(\mycsreg.CSReg[0][18] ), .A3(_05850_ ), .ZN(_06262_ ) );
OAI21_X1 _14223_ ( .A(_06262_ ), .B1(_04171_ ), .B2(_04180_ ), .ZN(_06263_ ) );
NAND3_X1 _14224_ ( .A1(_04213_ ), .A2(\mtvec [18] ), .A3(_04217_ ), .ZN(_06264_ ) );
NAND3_X1 _14225_ ( .A1(_04226_ ), .A2(\mepc [18] ), .A3(_05587_ ), .ZN(_06265_ ) );
NAND3_X1 _14226_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][18] ), .A3(_04206_ ), .ZN(_06266_ ) );
NAND4_X1 _14227_ ( .A1(_04198_ ), .A2(_06264_ ), .A3(_06265_ ), .A4(_06266_ ), .ZN(_06267_ ) );
NOR2_X1 _14228_ ( .A1(_06263_ ), .A2(_06267_ ), .ZN(_06268_ ) );
NOR3_X1 _14229_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [18] ), .A3(_05687_ ), .ZN(_06269_ ) );
NOR2_X1 _14230_ ( .A1(_06268_ ), .A2(_06269_ ), .ZN(_06270_ ) );
OAI22_X1 _14231_ ( .A1(_06270_ ), .A2(_06206_ ), .B1(_06254_ ), .B2(\ID_EX_imm [18] ), .ZN(_06271_ ) );
AOI21_X1 _14232_ ( .A(_06271_ ), .B1(_05210_ ), .B2(_05628_ ), .ZN(_06272_ ) );
INV_X1 _14233_ ( .A(_06269_ ), .ZN(_06273_ ) );
OAI211_X1 _14234_ ( .A(_06273_ ), .B(_06212_ ), .C1(_06267_ ), .C2(_06263_ ), .ZN(_06274_ ) );
INV_X1 _14235_ ( .A(_06274_ ), .ZN(_06275_ ) );
OAI21_X1 _14236_ ( .A(_06224_ ), .B1(_06272_ ), .B2(_06275_ ), .ZN(_06276_ ) );
MUX2_X1 _14237_ ( .A(_06190_ ), .B(_04682_ ), .S(_04133_ ), .Z(_06277_ ) );
OAI21_X1 _14238_ ( .A(_06276_ ), .B1(_06241_ ), .B2(_06277_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ) );
NOR3_X1 _14239_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [17] ), .A3(_05687_ ), .ZN(_06278_ ) );
AND4_X1 _14240_ ( .A1(_05586_ ), .A2(_05588_ ), .A3(_05589_ ), .A4(_05591_ ), .ZN(_06279_ ) );
AND3_X1 _14241_ ( .A1(_05593_ ), .A2(\mtvec [17] ), .A3(_05595_ ), .ZN(_06280_ ) );
NOR2_X1 _14242_ ( .A1(_04210_ ), .A2(_06280_ ), .ZN(_06281_ ) );
AOI21_X1 _14243_ ( .A(_06278_ ), .B1(_06279_ ), .B2(_06281_ ), .ZN(_06282_ ) );
AOI21_X1 _14244_ ( .A(fanout_net_9 ), .B1(_02668_ ), .B2(_02687_ ), .ZN(_06283_ ) );
AND2_X1 _14245_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [17] ), .ZN(_06284_ ) );
OAI221_X1 _14246_ ( .A(_04113_ ), .B1(_06207_ ), .B2(_06282_ ), .C1(_06283_ ), .C2(_06284_ ), .ZN(_06285_ ) );
BUF_X4 _14247_ ( .A(_04105_ ), .Z(_06286_ ) );
NAND3_X1 _14248_ ( .A1(_06282_ ), .A2(_06286_ ), .A3(_06213_ ), .ZN(_06287_ ) );
MUX2_X1 _14249_ ( .A(_05576_ ), .B(_04731_ ), .S(_06242_ ), .Z(_06288_ ) );
OAI211_X1 _14250_ ( .A(_06285_ ), .B(_06287_ ), .C1(_04127_ ), .C2(_06288_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ) );
OAI211_X1 _14251_ ( .A(_02992_ ), .B(_04097_ ), .C1(_05988_ ), .C2(\ID_EX_imm [16] ), .ZN(_06289_ ) );
AOI21_X1 _14252_ ( .A(_06289_ ), .B1(_05200_ ), .B2(_05817_ ), .ZN(_06290_ ) );
OAI21_X1 _14253_ ( .A(_06290_ ), .B1(_06207_ ), .B2(_05618_ ), .ZN(_06291_ ) );
NAND3_X1 _14254_ ( .A1(_05618_ ), .A2(_06286_ ), .A3(_06213_ ), .ZN(_06292_ ) );
MUX2_X1 _14255_ ( .A(_05581_ ), .B(_04753_ ), .S(_06242_ ), .Z(_06293_ ) );
OAI211_X1 _14256_ ( .A(_06291_ ), .B(_06292_ ), .C1(_04127_ ), .C2(_06293_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ) );
NAND3_X1 _14257_ ( .A1(_04212_ ), .A2(\mtvec [15] ), .A3(_05594_ ), .ZN(_06294_ ) );
NAND3_X1 _14258_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][15] ), .A3(_04206_ ), .ZN(_06295_ ) );
NAND3_X1 _14259_ ( .A1(_04198_ ), .A2(_06294_ ), .A3(_06295_ ), .ZN(_06296_ ) );
AND3_X1 _14260_ ( .A1(_04225_ ), .A2(\mepc [15] ), .A3(_04206_ ), .ZN(_06297_ ) );
AND3_X1 _14261_ ( .A1(_04212_ ), .A2(\mycsreg.CSReg[0][15] ), .A3(_04222_ ), .ZN(_06298_ ) );
NOR4_X1 _14262_ ( .A1(_04210_ ), .A2(_06296_ ), .A3(_06297_ ), .A4(_06298_ ), .ZN(_06299_ ) );
NOR3_X1 _14263_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [15] ), .A3(_05687_ ), .ZN(_06300_ ) );
NOR2_X1 _14264_ ( .A1(_06299_ ), .A2(_06300_ ), .ZN(_06301_ ) );
OAI22_X1 _14265_ ( .A1(_06301_ ), .A2(_06206_ ), .B1(_06254_ ), .B2(\ID_EX_imm [15] ), .ZN(_06302_ ) );
AOI21_X1 _14266_ ( .A(_06302_ ), .B1(_05628_ ), .B2(_05404_ ), .ZN(_06303_ ) );
OR3_X1 _14267_ ( .A1(_06299_ ), .A2(_06300_ ), .A3(_06236_ ), .ZN(_06304_ ) );
INV_X1 _14268_ ( .A(_06304_ ), .ZN(_06305_ ) );
OAI21_X1 _14269_ ( .A(_06224_ ), .B1(_06303_ ), .B2(_06305_ ), .ZN(_06306_ ) );
MUX2_X1 _14270_ ( .A(_04287_ ), .B(_05026_ ), .S(_04133_ ), .Z(_06307_ ) );
OAI21_X1 _14271_ ( .A(_06306_ ), .B1(_06241_ ), .B2(_06307_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ) );
NAND3_X1 _14272_ ( .A1(_02476_ ), .A2(_02495_ ), .A3(_06254_ ), .ZN(_06308_ ) );
OR2_X1 _14273_ ( .A1(_05487_ ), .A2(\ID_EX_imm [14] ), .ZN(_06309_ ) );
NAND3_X1 _14274_ ( .A1(_05675_ ), .A2(\ID_EX_typ [2] ), .A3(_05676_ ), .ZN(_06310_ ) );
AND3_X1 _14275_ ( .A1(_06308_ ), .A2(_06309_ ), .A3(_06310_ ), .ZN(_06311_ ) );
AOI21_X1 _14276_ ( .A(_06237_ ), .B1(_05675_ ), .B2(_05676_ ), .ZN(_06312_ ) );
OAI21_X1 _14277_ ( .A(_06224_ ), .B1(_06311_ ), .B2(_06312_ ), .ZN(_06313_ ) );
MUX2_X1 _14278_ ( .A(_06191_ ), .B(_05004_ ), .S(_04133_ ), .Z(_06314_ ) );
OAI21_X1 _14279_ ( .A(_06313_ ), .B1(_06241_ ), .B2(_06314_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ) );
OAI211_X1 _14280_ ( .A(_02992_ ), .B(_04097_ ), .C1(_05988_ ), .C2(\ID_EX_imm [13] ), .ZN(_06315_ ) );
INV_X1 _14281_ ( .A(_02565_ ), .ZN(_06316_ ) );
AOI21_X1 _14282_ ( .A(_06315_ ), .B1(_06316_ ), .B2(_05817_ ), .ZN(_06317_ ) );
NAND3_X1 _14283_ ( .A1(_05516_ ), .A2(\EX_LS_result_csreg_mem [13] ), .A3(_05521_ ), .ZN(_06318_ ) );
NAND4_X1 _14284_ ( .A1(_05534_ ), .A2(\mycsreg.CSReg[0][13] ), .A3(_05543_ ), .A4(_04223_ ), .ZN(_06319_ ) );
NAND4_X1 _14285_ ( .A1(_05545_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][13] ), .A4(_05538_ ), .ZN(_06320_ ) );
NAND4_X1 _14286_ ( .A1(_05545_ ), .A2(_05546_ ), .A3(\mepc [13] ), .A4(_05538_ ), .ZN(_06321_ ) );
NAND3_X1 _14287_ ( .A1(_06319_ ), .A2(_06320_ ), .A3(_06321_ ), .ZN(_06322_ ) );
NAND4_X1 _14288_ ( .A1(_05545_ ), .A2(_04218_ ), .A3(\mtvec [13] ), .A4(_05543_ ), .ZN(_06323_ ) );
NAND2_X1 _14289_ ( .A1(_05671_ ), .A2(_06323_ ), .ZN(_06324_ ) );
NOR2_X1 _14290_ ( .A1(_06322_ ), .A2(_06324_ ), .ZN(_06325_ ) );
OAI21_X1 _14291_ ( .A(_06318_ ), .B1(_05617_ ), .B2(_06325_ ), .ZN(_06326_ ) );
OAI21_X1 _14292_ ( .A(_06317_ ), .B1(_06207_ ), .B2(_06326_ ), .ZN(_06327_ ) );
NAND3_X1 _14293_ ( .A1(_06326_ ), .A2(_06286_ ), .A3(_06213_ ), .ZN(_06328_ ) );
MUX2_X1 _14294_ ( .A(_05697_ ), .B(_05072_ ), .S(_06242_ ), .Z(_06329_ ) );
OAI211_X1 _14295_ ( .A(_06327_ ), .B(_06328_ ), .C1(_04127_ ), .C2(_06329_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ) );
AND3_X1 _14296_ ( .A1(_05715_ ), .A2(\ID_EX_typ [2] ), .A3(_05716_ ), .ZN(_06330_ ) );
NAND2_X1 _14297_ ( .A1(_02588_ ), .A2(_05817_ ), .ZN(_06331_ ) );
NAND2_X1 _14298_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [12] ), .ZN(_06332_ ) );
AOI21_X1 _14299_ ( .A(_06330_ ), .B1(_06331_ ), .B2(_06332_ ), .ZN(_06333_ ) );
AOI21_X1 _14300_ ( .A(_06237_ ), .B1(_05715_ ), .B2(_05716_ ), .ZN(_06334_ ) );
OAI21_X1 _14301_ ( .A(_06224_ ), .B1(_06333_ ), .B2(_06334_ ), .ZN(_06335_ ) );
MUX2_X1 _14302_ ( .A(_05578_ ), .B(_05050_ ), .S(_04133_ ), .Z(_06336_ ) );
OAI21_X1 _14303_ ( .A(_06335_ ), .B1(_06241_ ), .B2(_06336_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ) );
OAI211_X1 _14304_ ( .A(_02992_ ), .B(_04097_ ), .C1(_05988_ ), .C2(\ID_EX_imm [30] ), .ZN(_06337_ ) );
AOI21_X1 _14305_ ( .A(_06337_ ), .B1(_02962_ ), .B2(_05817_ ), .ZN(_06338_ ) );
NAND3_X1 _14306_ ( .A1(_05516_ ), .A2(\EX_LS_result_csreg_mem [30] ), .A3(_05521_ ), .ZN(_06339_ ) );
NAND4_X1 _14307_ ( .A1(_05545_ ), .A2(\mycsreg.CSReg[0][30] ), .A3(_05543_ ), .A4(_04223_ ), .ZN(_06340_ ) );
NAND4_X1 _14308_ ( .A1(_05545_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][30] ), .A4(_05538_ ), .ZN(_06341_ ) );
NAND4_X1 _14309_ ( .A1(_05545_ ), .A2(_05546_ ), .A3(\mepc [30] ), .A4(_05538_ ), .ZN(_06342_ ) );
NAND3_X1 _14310_ ( .A1(_06340_ ), .A2(_06341_ ), .A3(_06342_ ), .ZN(_06343_ ) );
NAND4_X1 _14311_ ( .A1(_05545_ ), .A2(_04218_ ), .A3(\mtvec [30] ), .A4(_05543_ ), .ZN(_06344_ ) );
NAND2_X1 _14312_ ( .A1(_05671_ ), .A2(_06344_ ), .ZN(_06345_ ) );
NOR2_X1 _14313_ ( .A1(_06343_ ), .A2(_06345_ ), .ZN(_06346_ ) );
OAI21_X1 _14314_ ( .A(_06339_ ), .B1(_05617_ ), .B2(_06346_ ), .ZN(_06347_ ) );
OAI21_X1 _14315_ ( .A(_06338_ ), .B1(_06207_ ), .B2(_06347_ ), .ZN(_06348_ ) );
NAND3_X1 _14316_ ( .A1(_06347_ ), .A2(_06286_ ), .A3(_06213_ ), .ZN(_06349_ ) );
AND4_X1 _14317_ ( .A1(\ID_EX_pc [30] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06350_ ) );
AOI21_X1 _14318_ ( .A(_06350_ ), .B1(_04454_ ), .B2(_06243_ ), .ZN(_06351_ ) );
OAI211_X1 _14319_ ( .A(_06348_ ), .B(_06349_ ), .C1(_04127_ ), .C2(_06351_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ) );
NAND3_X1 _14320_ ( .A1(_05738_ ), .A2(\ID_EX_typ [2] ), .A3(_05739_ ), .ZN(_06352_ ) );
NAND3_X1 _14321_ ( .A1(_02379_ ), .A2(_02398_ ), .A3(_05627_ ), .ZN(_06353_ ) );
NAND2_X1 _14322_ ( .A1(_02576_ ), .A2(fanout_net_9 ), .ZN(_06354_ ) );
AND3_X1 _14323_ ( .A1(_06352_ ), .A2(_06353_ ), .A3(_06354_ ), .ZN(_06355_ ) );
AOI21_X1 _14324_ ( .A(_06237_ ), .B1(_05738_ ), .B2(_05739_ ), .ZN(_06356_ ) );
OAI21_X1 _14325_ ( .A(_06224_ ), .B1(_06355_ ), .B2(_06356_ ), .ZN(_06357_ ) );
MUX2_X1 _14326_ ( .A(_06192_ ), .B(_04934_ ), .S(_04133_ ), .Z(_06358_ ) );
OAI21_X1 _14327_ ( .A(_06357_ ), .B1(_06241_ ), .B2(_06358_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ) );
NAND3_X1 _14328_ ( .A1(_05645_ ), .A2(_05647_ ), .A3(_05812_ ), .ZN(_06359_ ) );
INV_X1 _14329_ ( .A(_05807_ ), .ZN(_06360_ ) );
AND2_X1 _14330_ ( .A1(_06359_ ), .A2(_06360_ ), .ZN(_06361_ ) );
OAI22_X1 _14331_ ( .A1(_06361_ ), .A2(_05468_ ), .B1(_05487_ ), .B2(\ID_EX_imm [10] ), .ZN(_06362_ ) );
AOI21_X1 _14332_ ( .A(_06362_ ), .B1(_05988_ ), .B2(_02574_ ), .ZN(_06363_ ) );
AOI211_X1 _14333_ ( .A(_05807_ ), .B(_06236_ ), .C1(_05527_ ), .C2(_05812_ ), .ZN(_06364_ ) );
OR3_X1 _14334_ ( .A1(_06363_ ), .A2(_04106_ ), .A3(_06364_ ), .ZN(_06365_ ) );
NAND4_X1 _14335_ ( .A1(\ID_EX_pc [10] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06366_ ) );
OAI211_X1 _14336_ ( .A(_04107_ ), .B(_06366_ ), .C1(_04912_ ), .C2(_04131_ ), .ZN(_06367_ ) );
AND2_X1 _14337_ ( .A1(_06365_ ), .A2(_06367_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ) );
OAI22_X1 _14338_ ( .A1(_05833_ ), .A2(_06206_ ), .B1(_06254_ ), .B2(\ID_EX_imm [9] ), .ZN(_06368_ ) );
AOI21_X1 _14339_ ( .A(_06368_ ), .B1(_05628_ ), .B2(_02582_ ), .ZN(_06369_ ) );
AND3_X1 _14340_ ( .A1(_05830_ ), .A2(_05832_ ), .A3(_06211_ ), .ZN(_06370_ ) );
OAI21_X1 _14341_ ( .A(_06224_ ), .B1(_06369_ ), .B2(_06370_ ), .ZN(_06371_ ) );
MUX2_X1 _14342_ ( .A(_05820_ ), .B(_04957_ ), .S(_04133_ ), .Z(_06372_ ) );
OAI21_X1 _14343_ ( .A(_06371_ ), .B1(_06241_ ), .B2(_06372_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ) );
OAI211_X1 _14344_ ( .A(_02992_ ), .B(_04097_ ), .C1(_06254_ ), .C2(\ID_EX_imm [8] ), .ZN(_06373_ ) );
AOI21_X1 _14345_ ( .A(_06373_ ), .B1(_05323_ ), .B2(_05817_ ), .ZN(_06374_ ) );
OAI21_X1 _14346_ ( .A(_06374_ ), .B1(_06207_ ), .B2(_05853_ ), .ZN(_06375_ ) );
NAND3_X1 _14347_ ( .A1(_05853_ ), .A2(_06286_ ), .A3(_06213_ ), .ZN(_06376_ ) );
MUX2_X1 _14348_ ( .A(_05839_ ), .B(_04981_ ), .S(_06242_ ), .Z(_06377_ ) );
OAI211_X1 _14349_ ( .A(_06375_ ), .B(_06376_ ), .C1(_04127_ ), .C2(_06377_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ) );
AOI22_X1 _14350_ ( .A1(_05868_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_06378_ ) );
OAI211_X1 _14351_ ( .A(_06378_ ), .B(_04126_ ), .C1(fanout_net_9 ), .C2(_02345_ ), .ZN(_06379_ ) );
NAND4_X1 _14352_ ( .A1(_05866_ ), .A2(_06240_ ), .A3(_05867_ ), .A4(_06213_ ), .ZN(_06380_ ) );
MUX2_X1 _14353_ ( .A(_06193_ ), .B(_04800_ ), .S(_06242_ ), .Z(_06381_ ) );
OAI211_X1 _14354_ ( .A(_06379_ ), .B(_06380_ ), .C1(_04127_ ), .C2(_06381_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ) );
OAI211_X1 _14355_ ( .A(_02992_ ), .B(_04097_ ), .C1(_06254_ ), .C2(\ID_EX_imm [6] ), .ZN(_06382_ ) );
INV_X1 _14356_ ( .A(_02371_ ), .ZN(_06383_ ) );
AOI21_X1 _14357_ ( .A(_06382_ ), .B1(_06383_ ), .B2(_05817_ ), .ZN(_06384_ ) );
OAI21_X1 _14358_ ( .A(_06384_ ), .B1(_06207_ ), .B2(_05888_ ), .ZN(_06385_ ) );
NAND3_X1 _14359_ ( .A1(_05888_ ), .A2(_06240_ ), .A3(_06213_ ), .ZN(_06386_ ) );
BUF_X4 _14360_ ( .A(_04113_ ), .Z(_06387_ ) );
MUX2_X1 _14361_ ( .A(_06194_ ), .B(_04778_ ), .S(_06242_ ), .Z(_06388_ ) );
OAI211_X1 _14362_ ( .A(_06385_ ), .B(_06386_ ), .C1(_06387_ ), .C2(_06388_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ) );
OAI211_X1 _14363_ ( .A(_02991_ ), .B(_04097_ ), .C1(_06254_ ), .C2(\ID_EX_imm [5] ), .ZN(_06389_ ) );
AOI21_X1 _14364_ ( .A(_06389_ ), .B1(_02213_ ), .B2(_05817_ ), .ZN(_06390_ ) );
OAI21_X1 _14365_ ( .A(_06390_ ), .B1(_06207_ ), .B2(_05905_ ), .ZN(_06391_ ) );
NAND3_X1 _14366_ ( .A1(_05905_ ), .A2(_06240_ ), .A3(_06213_ ), .ZN(_06392_ ) );
AND4_X1 _14367_ ( .A1(\ID_EX_pc [5] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06393_ ) );
AOI21_X1 _14368_ ( .A(_06393_ ), .B1(_04843_ ), .B2(_06243_ ), .ZN(_06394_ ) );
OAI211_X1 _14369_ ( .A(_06391_ ), .B(_06392_ ), .C1(_06387_ ), .C2(_06394_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ) );
NAND3_X1 _14370_ ( .A1(_02190_ ), .A2(_02209_ ), .A3(_06254_ ), .ZN(_06395_ ) );
NAND2_X1 _14371_ ( .A1(_02320_ ), .A2(fanout_net_9 ), .ZN(_06396_ ) );
NAND3_X1 _14372_ ( .A1(_05921_ ), .A2(\ID_EX_typ [2] ), .A3(_05922_ ), .ZN(_06397_ ) );
AND3_X1 _14373_ ( .A1(_06395_ ), .A2(_06396_ ), .A3(_06397_ ), .ZN(_06398_ ) );
AOI21_X1 _14374_ ( .A(_06237_ ), .B1(_05921_ ), .B2(_05922_ ), .ZN(_06399_ ) );
OAI21_X1 _14375_ ( .A(_06286_ ), .B1(_06398_ ), .B2(_06399_ ), .ZN(_06400_ ) );
MUX2_X1 _14376_ ( .A(_06195_ ), .B(_04822_ ), .S(_04133_ ), .Z(_06401_ ) );
OAI21_X1 _14377_ ( .A(_06400_ ), .B1(_06241_ ), .B2(_06401_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ) );
BUF_X4 _14378_ ( .A(_04105_ ), .Z(_06402_ ) );
AOI211_X1 _14379_ ( .A(_05468_ ), .B(_05940_ ), .C1(_05646_ ), .C2(_05938_ ), .ZN(_06403_ ) );
NAND2_X1 _14380_ ( .A1(_02235_ ), .A2(_05817_ ), .ZN(_06404_ ) );
NAND2_X1 _14381_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [3] ), .ZN(_06405_ ) );
AOI21_X1 _14382_ ( .A(_06403_ ), .B1(_06404_ ), .B2(_06405_ ), .ZN(_06406_ ) );
AOI21_X1 _14383_ ( .A(_06237_ ), .B1(_05939_ ), .B2(_05941_ ), .ZN(_06407_ ) );
OAI21_X1 _14384_ ( .A(_06402_ ), .B1(_06406_ ), .B2(_06407_ ), .ZN(_06408_ ) );
BUF_X4 _14385_ ( .A(_04106_ ), .Z(_06409_ ) );
NAND3_X1 _14386_ ( .A1(_03343_ ), .A2(_06196_ ), .A3(\ID_EX_typ [7] ), .ZN(_06410_ ) );
OAI211_X1 _14387_ ( .A(_06409_ ), .B(_06410_ ), .C1(_04888_ ), .C2(_04131_ ), .ZN(_06411_ ) );
NAND2_X1 _14388_ ( .A1(_06408_ ), .A2(_06411_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ) );
NAND3_X1 _14389_ ( .A1(_05645_ ), .A2(_05647_ ), .A3(_05956_ ), .ZN(_06412_ ) );
INV_X1 _14390_ ( .A(_05951_ ), .ZN(_06413_ ) );
AND2_X1 _14391_ ( .A1(_06412_ ), .A2(_06413_ ), .ZN(_06414_ ) );
OAI22_X1 _14392_ ( .A1(_06414_ ), .A2(_06206_ ), .B1(_06254_ ), .B2(\ID_EX_imm [2] ), .ZN(_06415_ ) );
AOI21_X1 _14393_ ( .A(_06415_ ), .B1(_05628_ ), .B2(_05281_ ), .ZN(_06416_ ) );
AOI211_X1 _14394_ ( .A(_05951_ ), .B(_06237_ ), .C1(_05527_ ), .C2(_05956_ ), .ZN(_06417_ ) );
OAI21_X1 _14395_ ( .A(_06286_ ), .B1(_06416_ ), .B2(_06417_ ), .ZN(_06418_ ) );
MUX2_X1 _14396_ ( .A(_06197_ ), .B(_04866_ ), .S(_04133_ ), .Z(_06419_ ) );
OAI21_X1 _14397_ ( .A(_06418_ ), .B1(_06241_ ), .B2(_06419_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ) );
AND3_X1 _14398_ ( .A1(_05797_ ), .A2(\ID_EX_typ [2] ), .A3(_05798_ ), .ZN(_06420_ ) );
NAND2_X1 _14399_ ( .A1(_02909_ ), .A2(_05488_ ), .ZN(_06421_ ) );
NAND2_X1 _14400_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [29] ), .ZN(_06422_ ) );
AOI21_X1 _14401_ ( .A(_06420_ ), .B1(_06421_ ), .B2(_06422_ ), .ZN(_06423_ ) );
AOI21_X1 _14402_ ( .A(_06237_ ), .B1(_05797_ ), .B2(_05798_ ), .ZN(_06424_ ) );
OAI21_X1 _14403_ ( .A(_06286_ ), .B1(_06423_ ), .B2(_06424_ ), .ZN(_06425_ ) );
AND4_X1 _14404_ ( .A1(\ID_EX_pc [29] ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06426_ ) );
AOI21_X1 _14405_ ( .A(_06426_ ), .B1(_04384_ ), .B2(_06243_ ), .ZN(_06427_ ) );
OAI21_X1 _14406_ ( .A(_06425_ ), .B1(_04127_ ), .B2(_06427_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ) );
OR3_X1 _14407_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [1] ), .A3(_05687_ ), .ZN(_06428_ ) );
NAND3_X1 _14408_ ( .A1(_04214_ ), .A2(\mtvec [1] ), .A3(_04218_ ), .ZN(_06429_ ) );
NAND3_X1 _14409_ ( .A1(_04214_ ), .A2(\mycsreg.CSReg[0][1] ), .A3(_04223_ ), .ZN(_06430_ ) );
NAND3_X1 _14410_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][1] ), .A3(_04207_ ), .ZN(_06431_ ) );
NAND3_X1 _14411_ ( .A1(_04226_ ), .A2(\mepc [1] ), .A3(_04207_ ), .ZN(_06432_ ) );
NAND4_X1 _14412_ ( .A1(_06429_ ), .A2(_06430_ ), .A3(_06431_ ), .A4(_06432_ ), .ZN(_06433_ ) );
OAI21_X1 _14413_ ( .A(_06428_ ), .B1(_04210_ ), .B2(_06433_ ), .ZN(_06434_ ) );
AOI22_X1 _14414_ ( .A1(_06434_ ), .A2(\ID_EX_typ [2] ), .B1(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .B2(fanout_net_9 ), .ZN(_06435_ ) );
OAI211_X1 _14415_ ( .A(_06240_ ), .B(_06435_ ), .C1(_02282_ ), .C2(fanout_net_9 ), .ZN(_06436_ ) );
AND2_X1 _14416_ ( .A1(_06429_ ), .A2(_06430_ ), .ZN(_06437_ ) );
AND2_X1 _14417_ ( .A1(_06431_ ), .A2(_06432_ ), .ZN(_06438_ ) );
OAI211_X1 _14418_ ( .A(_06437_ ), .B(_06438_ ), .C1(_04172_ ), .C2(_04181_ ), .ZN(_06439_ ) );
NAND4_X1 _14419_ ( .A1(_06439_ ), .A2(_06240_ ), .A3(_06428_ ), .A4(_06212_ ), .ZN(_06440_ ) );
MUX2_X1 _14420_ ( .A(_04265_ ), .B(_05099_ ), .S(_06243_ ), .Z(_06441_ ) );
OAI211_X1 _14421_ ( .A(_06436_ ), .B(_06440_ ), .C1(_06441_ ), .C2(_04114_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ) );
AND3_X1 _14422_ ( .A1(_02306_ ), .A2(_05988_ ), .A3(_02308_ ), .ZN(_06442_ ) );
AND2_X1 _14423_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [0] ), .ZN(_06443_ ) );
OAI221_X1 _14424_ ( .A(_04113_ ), .B1(_06206_ ), .B2(_06003_ ), .C1(_06442_ ), .C2(_06443_ ), .ZN(_06444_ ) );
NAND2_X1 _14425_ ( .A1(_05998_ ), .A2(_06002_ ), .ZN(_06445_ ) );
OR3_X1 _14426_ ( .A1(_04172_ ), .A2(\EX_LS_result_csreg_mem [0] ), .A3(_04181_ ), .ZN(_06446_ ) );
NAND4_X1 _14427_ ( .A1(_06445_ ), .A2(_06240_ ), .A3(_06446_ ), .A4(_06212_ ), .ZN(_06447_ ) );
MUX2_X1 _14428_ ( .A(_06198_ ), .B(_05121_ ), .S(_06242_ ), .Z(_06448_ ) );
OAI211_X1 _14429_ ( .A(_06444_ ), .B(_06447_ ), .C1(_06387_ ), .C2(_06448_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ) );
AND3_X1 _14430_ ( .A1(_05983_ ), .A2(\ID_EX_typ [2] ), .A3(_05984_ ), .ZN(_06449_ ) );
NOR2_X1 _14431_ ( .A1(_05488_ ), .A2(\ID_EX_imm [28] ), .ZN(_06450_ ) );
AOI21_X1 _14432_ ( .A(fanout_net_9 ), .B1(_02931_ ), .B2(_02932_ ), .ZN(_06451_ ) );
NOR3_X1 _14433_ ( .A1(_06449_ ), .A2(_06450_ ), .A3(_06451_ ), .ZN(_06452_ ) );
AOI21_X1 _14434_ ( .A(_06237_ ), .B1(_05983_ ), .B2(_05984_ ), .ZN(_06453_ ) );
OAI21_X1 _14435_ ( .A(_06402_ ), .B1(_06452_ ), .B2(_06453_ ), .ZN(_06454_ ) );
NAND3_X1 _14436_ ( .A1(_03343_ ), .A2(_06199_ ), .A3(\ID_EX_typ [7] ), .ZN(_06455_ ) );
OAI211_X1 _14437_ ( .A(_06409_ ), .B(_06455_ ), .C1(_04408_ ), .C2(_04131_ ), .ZN(_06456_ ) );
NAND2_X1 _14438_ ( .A1(_06454_ ), .A2(_06456_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _14439_ ( .A(fanout_net_9 ), .B1(_02838_ ), .B2(_02857_ ), .ZN(_06457_ ) );
AND2_X1 _14440_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [27] ), .ZN(_06458_ ) );
OAI221_X1 _14441_ ( .A(_04113_ ), .B1(_06206_ ), .B2(_06024_ ), .C1(_06457_ ), .C2(_06458_ ), .ZN(_06459_ ) );
NAND3_X1 _14442_ ( .A1(_04214_ ), .A2(\mtvec [27] ), .A3(_04218_ ), .ZN(_06460_ ) );
NAND3_X1 _14443_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][27] ), .A3(_04207_ ), .ZN(_06461_ ) );
AND3_X1 _14444_ ( .A1(_04193_ ), .A2(_06460_ ), .A3(_06461_ ), .ZN(_06462_ ) );
AND2_X1 _14445_ ( .A1(_04214_ ), .A2(_04223_ ), .ZN(_06463_ ) );
AOI22_X1 _14446_ ( .A1(_06463_ ), .A2(\mycsreg.CSReg[0][27] ), .B1(\mepc [27] ), .B2(_05864_ ), .ZN(_06464_ ) );
NAND3_X1 _14447_ ( .A1(_06120_ ), .A2(_06462_ ), .A3(_06464_ ), .ZN(_06465_ ) );
OR3_X1 _14448_ ( .A1(_04172_ ), .A2(\EX_LS_result_csreg_mem [27] ), .A3(_04181_ ), .ZN(_06466_ ) );
NAND4_X1 _14449_ ( .A1(_06465_ ), .A2(_06240_ ), .A3(_06466_ ), .A4(_06212_ ), .ZN(_06467_ ) );
AND3_X1 _14450_ ( .A1(_03343_ ), .A2(\ID_EX_pc [27] ), .A3(\ID_EX_typ [7] ), .ZN(_06468_ ) );
AOI21_X1 _14451_ ( .A(_06468_ ), .B1(_04478_ ), .B2(_06243_ ), .ZN(_06469_ ) );
OAI211_X1 _14452_ ( .A(_06459_ ), .B(_06467_ ), .C1(_06469_ ), .C2(_04114_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ) );
AND2_X1 _14453_ ( .A1(_06037_ ), .A2(_06038_ ), .ZN(_06470_ ) );
INV_X1 _14454_ ( .A(_06470_ ), .ZN(_06471_ ) );
NAND3_X1 _14455_ ( .A1(_02860_ ), .A2(_05988_ ), .A3(_02879_ ), .ZN(_06472_ ) );
NAND2_X1 _14456_ ( .A1(fanout_net_9 ), .A2(\myexu.src1_plus_imm_$_NOT__Y_3_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ), .ZN(_06473_ ) );
AND2_X1 _14457_ ( .A1(_06472_ ), .A2(_06473_ ), .ZN(_06474_ ) );
AOI21_X1 _14458_ ( .A(_06237_ ), .B1(_06037_ ), .B2(_06038_ ), .ZN(_06475_ ) );
OAI221_X1 _14459_ ( .A(_06224_ ), .B1(_06471_ ), .B2(_06207_ ), .C1(_06474_ ), .C2(_06475_ ), .ZN(_06476_ ) );
NAND4_X1 _14460_ ( .A1(_06200_ ), .A2(\ID_EX_typ [7] ), .A3(\ID_EX_typ [6] ), .A4(\ID_EX_typ [5] ), .ZN(_06477_ ) );
OAI211_X1 _14461_ ( .A(_06409_ ), .B(_06477_ ), .C1(_04508_ ), .C2(_04131_ ), .ZN(_06478_ ) );
NAND2_X1 _14462_ ( .A1(_06476_ ), .A2(_06478_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ) );
NAND3_X1 _14463_ ( .A1(_05593_ ), .A2(\mtvec [25] ), .A3(_05595_ ), .ZN(_06479_ ) );
NAND3_X1 _14464_ ( .A1(_05593_ ), .A2(\mycsreg.CSReg[0][25] ), .A3(_05850_ ), .ZN(_06480_ ) );
AND2_X1 _14465_ ( .A1(_06479_ ), .A2(_06480_ ), .ZN(_06481_ ) );
AND3_X1 _14466_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][25] ), .A3(_04206_ ), .ZN(_06482_ ) );
AOI21_X1 _14467_ ( .A(_06482_ ), .B1(\mepc [25] ), .B2(_05864_ ), .ZN(_06483_ ) );
OAI211_X1 _14468_ ( .A(_06481_ ), .B(_06483_ ), .C1(_04172_ ), .C2(_04181_ ), .ZN(_06484_ ) );
OR3_X1 _14469_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [25] ), .A3(_05687_ ), .ZN(_06485_ ) );
NAND2_X1 _14470_ ( .A1(_06484_ ), .A2(_06485_ ), .ZN(_06486_ ) );
AOI22_X1 _14471_ ( .A1(_06486_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(_02811_ ), .ZN(_06487_ ) );
OAI211_X1 _14472_ ( .A(_06487_ ), .B(_04126_ ), .C1(fanout_net_9 ), .C2(_02834_ ), .ZN(_06488_ ) );
NAND4_X1 _14473_ ( .A1(_06484_ ), .A2(_04126_ ), .A3(_06485_ ), .A4(_06212_ ), .ZN(_06489_ ) );
AND3_X1 _14474_ ( .A1(_03343_ ), .A2(\ID_EX_pc [25] ), .A3(\ID_EX_typ [7] ), .ZN(_06490_ ) );
AOI21_X1 _14475_ ( .A(_06490_ ), .B1(_04556_ ), .B2(_06243_ ), .ZN(_06491_ ) );
OAI211_X1 _14476_ ( .A(_06488_ ), .B(_06489_ ), .C1(_06387_ ), .C2(_06491_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ) );
AOI21_X1 _14477_ ( .A(fanout_net_9 ), .B1(_02160_ ), .B2(_02161_ ), .ZN(_06492_ ) );
AND2_X1 _14478_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [24] ), .ZN(_06493_ ) );
OAI221_X1 _14479_ ( .A(_04113_ ), .B1(_06206_ ), .B2(_06081_ ), .C1(_06492_ ), .C2(_06493_ ), .ZN(_06494_ ) );
NAND3_X1 _14480_ ( .A1(_04214_ ), .A2(\mtvec [24] ), .A3(_04218_ ), .ZN(_06495_ ) );
NAND3_X1 _14481_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][24] ), .A3(_04207_ ), .ZN(_06496_ ) );
AND4_X1 _14482_ ( .A1(_04193_ ), .A2(_04198_ ), .A3(_06495_ ), .A4(_06496_ ), .ZN(_06497_ ) );
AOI22_X1 _14483_ ( .A1(_06463_ ), .A2(\mycsreg.CSReg[0][24] ), .B1(\mepc [24] ), .B2(_05864_ ), .ZN(_06498_ ) );
NAND3_X1 _14484_ ( .A1(_06497_ ), .A2(_06120_ ), .A3(_06498_ ), .ZN(_06499_ ) );
OR3_X1 _14485_ ( .A1(_04172_ ), .A2(\EX_LS_result_csreg_mem [24] ), .A3(_04181_ ), .ZN(_06500_ ) );
NAND4_X1 _14486_ ( .A1(_06499_ ), .A2(_04126_ ), .A3(_06500_ ), .A4(_06212_ ), .ZN(_06501_ ) );
AND3_X1 _14487_ ( .A1(_03343_ ), .A2(\ID_EX_pc [24] ), .A3(\ID_EX_typ [7] ), .ZN(_06502_ ) );
AOI21_X1 _14488_ ( .A(_06502_ ), .B1(_04533_ ), .B2(_06243_ ), .ZN(_06503_ ) );
OAI211_X1 _14489_ ( .A(_06494_ ), .B(_06501_ ), .C1(_06387_ ), .C2(_06503_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ) );
NAND3_X1 _14490_ ( .A1(_05593_ ), .A2(\mtvec [23] ), .A3(_05595_ ), .ZN(_06504_ ) );
NAND3_X1 _14491_ ( .A1(_05593_ ), .A2(\mycsreg.CSReg[0][23] ), .A3(_05850_ ), .ZN(_06505_ ) );
AND2_X1 _14492_ ( .A1(_06504_ ), .A2(_06505_ ), .ZN(_06506_ ) );
AND3_X1 _14493_ ( .A1(_04202_ ), .A2(\mycsreg.CSReg[3][23] ), .A3(_04206_ ), .ZN(_06507_ ) );
AOI21_X1 _14494_ ( .A(_06507_ ), .B1(\mepc [23] ), .B2(_05864_ ), .ZN(_06508_ ) );
OAI211_X1 _14495_ ( .A(_06506_ ), .B(_06508_ ), .C1(_04172_ ), .C2(_04181_ ), .ZN(_06509_ ) );
OR3_X1 _14496_ ( .A1(_05686_ ), .A2(\EX_LS_result_csreg_mem [23] ), .A3(_05687_ ), .ZN(_06510_ ) );
NAND2_X1 _14497_ ( .A1(_06509_ ), .A2(_06510_ ), .ZN(_06511_ ) );
AOI22_X1 _14498_ ( .A1(_06511_ ), .A2(\ID_EX_typ [2] ), .B1(fanout_net_9 ), .B2(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ), .ZN(_06512_ ) );
OAI211_X1 _14499_ ( .A(_06512_ ), .B(_04126_ ), .C1(_02726_ ), .C2(fanout_net_9 ), .ZN(_06513_ ) );
NAND4_X1 _14500_ ( .A1(_06509_ ), .A2(_04126_ ), .A3(_06510_ ), .A4(_06212_ ), .ZN(_06514_ ) );
MUX2_X1 _14501_ ( .A(_06050_ ), .B(_04608_ ), .S(_06242_ ), .Z(_06515_ ) );
OAI211_X1 _14502_ ( .A(_06513_ ), .B(_06514_ ), .C1(_06387_ ), .C2(_06515_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ) );
NAND3_X1 _14503_ ( .A1(_05516_ ), .A2(\EX_LS_result_csreg_mem [22] ), .A3(_05521_ ), .ZN(_06516_ ) );
NAND4_X1 _14504_ ( .A1(_05847_ ), .A2(_05595_ ), .A3(\mtvec [22] ), .A4(_05542_ ), .ZN(_06517_ ) );
NAND4_X1 _14505_ ( .A1(_05847_ ), .A2(\mycsreg.CSReg[0][22] ), .A3(_05542_ ), .A4(_05850_ ), .ZN(_06518_ ) );
NAND4_X1 _14506_ ( .A1(_05533_ ), .A2(_05535_ ), .A3(\mycsreg.CSReg[3][22] ), .A4(_05537_ ), .ZN(_06519_ ) );
NAND3_X1 _14507_ ( .A1(_06517_ ), .A2(_06518_ ), .A3(_06519_ ), .ZN(_06520_ ) );
AND4_X1 _14508_ ( .A1(\mepc [22] ), .A2(_05604_ ), .A3(_05546_ ), .A4(_05537_ ), .ZN(_06521_ ) );
NOR4_X1 _14509_ ( .A1(_06520_ ), .A2(_05613_ ), .A3(_06521_ ), .A4(_05526_ ), .ZN(_06522_ ) );
OAI21_X1 _14510_ ( .A(_06516_ ), .B1(_06522_ ), .B2(_05617_ ), .ZN(_06523_ ) );
AOI21_X1 _14511_ ( .A(fanout_net_9 ), .B1(_02728_ ), .B2(_02747_ ), .ZN(_06524_ ) );
AND2_X1 _14512_ ( .A1(fanout_net_9 ), .A2(\ID_EX_imm [22] ), .ZN(_06525_ ) );
OAI221_X1 _14513_ ( .A(_04113_ ), .B1(_06206_ ), .B2(_06523_ ), .C1(_06524_ ), .C2(_06525_ ), .ZN(_06526_ ) );
AND3_X1 _14514_ ( .A1(_04203_ ), .A2(\mycsreg.CSReg[3][22] ), .A3(_04207_ ), .ZN(_06527_ ) );
NOR3_X1 _14515_ ( .A1(_06527_ ), .A2(_04192_ ), .A3(_04197_ ), .ZN(_06528_ ) );
AND2_X1 _14516_ ( .A1(_06114_ ), .A2(_06113_ ), .ZN(_06529_ ) );
NAND4_X1 _14517_ ( .A1(_06120_ ), .A2(_06528_ ), .A3(_06529_ ), .A4(_06116_ ), .ZN(_06530_ ) );
NAND4_X1 _14518_ ( .A1(_06530_ ), .A2(_04126_ ), .A3(_06111_ ), .A4(_06212_ ), .ZN(_06531_ ) );
MUX2_X1 _14519_ ( .A(_06202_ ), .B(_04585_ ), .S(_06242_ ), .Z(_06532_ ) );
OAI211_X1 _14520_ ( .A(_06526_ ), .B(_06531_ ), .C1(_06387_ ), .C2(_06532_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ) );
AOI22_X1 _14521_ ( .A1(_06180_ ), .A2(\ID_EX_typ [2] ), .B1(\ID_EX_typ [0] ), .B2(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ), .ZN(_06533_ ) );
OAI211_X1 _14522_ ( .A(_06533_ ), .B(_04126_ ), .C1(_02988_ ), .C2(\ID_EX_typ [0] ), .ZN(_06534_ ) );
NAND3_X1 _14523_ ( .A1(_06181_ ), .A2(_06240_ ), .A3(_06213_ ), .ZN(_06535_ ) );
AND3_X1 _14524_ ( .A1(_03343_ ), .A2(\ID_EX_pc [31] ), .A3(\ID_EX_typ [7] ), .ZN(_06536_ ) );
AOI21_X1 _14525_ ( .A(_06536_ ), .B1(_04432_ ), .B2(_06243_ ), .ZN(_06537_ ) );
OAI211_X1 _14526_ ( .A(_06534_ ), .B(_06535_ ), .C1(_06537_ ), .C2(_04114_ ), .ZN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ) );
OAI21_X1 _14527_ ( .A(_06286_ ), .B1(_06220_ ), .B2(_06221_ ), .ZN(_06538_ ) );
AND2_X2 _14528_ ( .A1(fanout_net_10 ), .A2(\ID_EX_typ [2] ), .ZN(_06539_ ) );
NOR3_X1 _14529_ ( .A1(_05133_ ), .A2(\ID_EX_typ [0] ), .A3(\ID_EX_typ [1] ), .ZN(_06540_ ) );
NOR3_X1 _14530_ ( .A1(_05379_ ), .A2(\ID_EX_typ [0] ), .A3(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__B_A_$_OR__A_Y_$_OR__A_B ), .ZN(_06541_ ) );
OAI21_X1 _14531_ ( .A(_06539_ ), .B1(_06540_ ), .B2(_06541_ ), .ZN(_06542_ ) );
NOR2_X1 _14532_ ( .A1(_04159_ ), .A2(\ID_EX_typ [2] ), .ZN(_06543_ ) );
OAI211_X1 _14533_ ( .A(_06543_ ), .B(_05379_ ), .C1(_05126_ ), .C2(_05133_ ), .ZN(_06544_ ) );
AND2_X1 _14534_ ( .A1(_06542_ ), .A2(_06544_ ), .ZN(_06545_ ) );
NOR2_X1 _14535_ ( .A1(_05482_ ), .A2(\ID_EX_typ [7] ), .ZN(_06546_ ) );
INV_X1 _14536_ ( .A(_06546_ ), .ZN(_06547_ ) );
NOR2_X1 _14537_ ( .A1(_06545_ ), .A2(_06547_ ), .ZN(_06548_ ) );
BUF_X4 _14538_ ( .A(_06548_ ), .Z(_06549_ ) );
AND2_X2 _14539_ ( .A1(_05385_ ), .A2(\ID_EX_typ [2] ), .ZN(_06550_ ) );
BUF_X4 _14540_ ( .A(_06550_ ), .Z(_06551_ ) );
AND2_X4 _14541_ ( .A1(_05271_ ), .A2(_05275_ ), .ZN(_06552_ ) );
AND2_X4 _14542_ ( .A1(_06552_ ), .A2(_05267_ ), .ZN(_06553_ ) );
INV_X1 _14543_ ( .A(_05262_ ), .ZN(_06554_ ) );
AND2_X4 _14544_ ( .A1(_06553_ ), .A2(_06554_ ), .ZN(_06555_ ) );
AND2_X4 _14545_ ( .A1(_06555_ ), .A2(_05287_ ), .ZN(_06556_ ) );
INV_X1 _14546_ ( .A(_05291_ ), .ZN(_06557_ ) );
OAI21_X4 _14547_ ( .A(_05299_ ), .B1(_06556_ ), .B2(_06557_ ), .ZN(_06558_ ) );
OR3_X4 _14548_ ( .A1(_06558_ ), .A2(_05324_ ), .A3(_05311_ ), .ZN(_06559_ ) );
INV_X1 _14549_ ( .A(_05251_ ), .ZN(_06560_ ) );
NOR3_X4 _14550_ ( .A1(_06559_ ), .A2(_05330_ ), .A3(_06560_ ), .ZN(_06561_ ) );
NAND4_X1 _14551_ ( .A1(_05223_ ), .A2(_05219_ ), .A3(_05224_ ), .A4(_05220_ ), .ZN(_06562_ ) );
NOR3_X1 _14552_ ( .A1(_05315_ ), .A2(_05231_ ), .A3(_06562_ ), .ZN(_06563_ ) );
AND3_X2 _14553_ ( .A1(_06561_ ), .A2(_05246_ ), .A3(_06563_ ), .ZN(_06564_ ) );
AND2_X1 _14554_ ( .A1(_05178_ ), .A2(_05183_ ), .ZN(_06565_ ) );
AND3_X1 _14555_ ( .A1(_05203_ ), .A2(_05193_ ), .A3(_05189_ ), .ZN(_06566_ ) );
AND2_X1 _14556_ ( .A1(_06566_ ), .A2(_05198_ ), .ZN(_06567_ ) );
AND3_X4 _14557_ ( .A1(_06564_ ), .A2(_06565_ ), .A3(_06567_ ), .ZN(_06568_ ) );
NOR4_X1 _14558_ ( .A1(_05344_ ), .A2(_05164_ ), .A3(_05340_ ), .A4(_05352_ ), .ZN(_06569_ ) );
AND4_X1 _14559_ ( .A1(_05355_ ), .A2(_06569_ ), .A3(_05356_ ), .A4(_05158_ ), .ZN(_06570_ ) );
NAND4_X1 _14560_ ( .A1(_06570_ ), .A2(_05172_ ), .A3(_05141_ ), .A4(_05146_ ), .ZN(_06571_ ) );
NOR2_X2 _14561_ ( .A1(_06568_ ), .A2(_06571_ ), .ZN(_06572_ ) );
AOI21_X4 _14562_ ( .A(_06572_ ), .B1(_05134_ ), .B2(_05135_ ), .ZN(_06573_ ) );
AND4_X1 _14563_ ( .A1(_05164_ ), .A2(_05344_ ), .A3(_05340_ ), .A4(_05352_ ), .ZN(_06574_ ) );
NAND4_X1 _14564_ ( .A1(_06574_ ), .A2(_05357_ ), .A3(_05159_ ), .A4(_06565_ ), .ZN(_06575_ ) );
NOR4_X1 _14565_ ( .A1(_06575_ ), .A2(_05172_ ), .A3(_05141_ ), .A4(_05146_ ), .ZN(_06576_ ) );
AND3_X1 _14566_ ( .A1(_06564_ ), .A2(_06567_ ), .A3(_06576_ ), .ZN(_06577_ ) );
NOR2_X1 _14567_ ( .A1(_06577_ ), .A2(_05136_ ), .ZN(_06578_ ) );
AND2_X1 _14568_ ( .A1(_06561_ ), .A2(_05246_ ), .ZN(_06579_ ) );
INV_X1 _14569_ ( .A(_06579_ ), .ZN(_06580_ ) );
AOI211_X1 _14570_ ( .A(_05225_ ), .B(_05221_ ), .C1(_05230_ ), .C2(_05229_ ), .ZN(_06581_ ) );
NAND3_X1 _14571_ ( .A1(_06580_ ), .A2(_05315_ ), .A3(_06581_ ), .ZN(_06582_ ) );
INV_X1 _14572_ ( .A(_06564_ ), .ZN(_06583_ ) );
AND2_X1 _14573_ ( .A1(_06582_ ), .A2(_06583_ ), .ZN(_06584_ ) );
OAI211_X1 _14574_ ( .A(_06560_ ), .B(_05324_ ), .C1(_06558_ ), .C2(_05311_ ), .ZN(_06585_ ) );
OAI21_X1 _14575_ ( .A(_06585_ ), .B1(_06559_ ), .B2(_06560_ ), .ZN(_06586_ ) );
OR4_X1 _14576_ ( .A1(_05295_ ), .A2(_06556_ ), .A3(_05299_ ), .A4(_06557_ ), .ZN(_06587_ ) );
OAI21_X1 _14577_ ( .A(_06587_ ), .B1(_05311_ ), .B2(_06558_ ), .ZN(_06588_ ) );
NAND3_X1 _14578_ ( .A1(_06586_ ), .A2(_02988_ ), .A3(_06588_ ), .ZN(_06589_ ) );
NOR4_X2 _14579_ ( .A1(_06573_ ), .A2(_06578_ ), .A3(_06584_ ), .A4(_06589_ ), .ZN(_06590_ ) );
OR4_X1 _14580_ ( .A1(_05178_ ), .A2(_05183_ ), .A3(_05198_ ), .A4(_05189_ ), .ZN(_06591_ ) );
NOR4_X1 _14581_ ( .A1(_06564_ ), .A2(_05203_ ), .A3(_05193_ ), .A4(_06591_ ), .ZN(_06592_ ) );
NOR2_X1 _14582_ ( .A1(_06592_ ), .A2(_06568_ ), .ZN(_06593_ ) );
NOR2_X1 _14583_ ( .A1(_06559_ ), .A2(_06560_ ), .ZN(_06594_ ) );
NOR3_X1 _14584_ ( .A1(_06594_ ), .A2(_05246_ ), .A3(_05242_ ), .ZN(_06595_ ) );
NOR2_X1 _14585_ ( .A1(_06579_ ), .A2(_06595_ ), .ZN(_06596_ ) );
NOR2_X1 _14586_ ( .A1(_06593_ ), .A2(_06596_ ), .ZN(_06597_ ) );
AND2_X4 _14587_ ( .A1(_06590_ ), .A2(_06597_ ), .ZN(_06598_ ) );
XNOR2_X1 _14588_ ( .A(_06556_ ), .B(_05291_ ), .ZN(_06599_ ) );
NAND2_X1 _14589_ ( .A1(_06598_ ), .A2(_06599_ ), .ZN(_06600_ ) );
XNOR2_X1 _14590_ ( .A(_06555_ ), .B(_05287_ ), .ZN(_06601_ ) );
NOR2_X1 _14591_ ( .A1(_06601_ ), .A2(_05291_ ), .ZN(_06602_ ) );
INV_X1 _14592_ ( .A(_06602_ ), .ZN(_06603_ ) );
INV_X1 _14593_ ( .A(_06601_ ), .ZN(_06604_ ) );
AOI211_X1 _14594_ ( .A(_06596_ ), .B(_06589_ ), .C1(_06582_ ), .C2(_06583_ ), .ZN(_06605_ ) );
OAI221_X1 _14595_ ( .A(_06605_ ), .B1(_05136_ ), .B2(_06577_ ), .C1(_06568_ ), .C2(_06592_ ), .ZN(_06606_ ) );
NOR2_X2 _14596_ ( .A1(_06606_ ), .A2(_06573_ ), .ZN(_06607_ ) );
BUF_X2 _14597_ ( .A(_06607_ ), .Z(_06608_ ) );
BUF_X2 _14598_ ( .A(_05271_ ), .Z(_06609_ ) );
BUF_X4 _14599_ ( .A(_06609_ ), .Z(_06610_ ) );
BUF_X4 _14600_ ( .A(_06610_ ), .Z(_06611_ ) );
BUF_X4 _14601_ ( .A(_06611_ ), .Z(_06612_ ) );
BUF_X4 _14602_ ( .A(_05275_ ), .Z(_06613_ ) );
BUF_X4 _14603_ ( .A(_06613_ ), .Z(_06614_ ) );
BUF_X4 _14604_ ( .A(_06614_ ), .Z(_06615_ ) );
XNOR2_X1 _14605_ ( .A(_06612_ ), .B(_06615_ ), .ZN(_06616_ ) );
BUF_X4 _14606_ ( .A(_05282_ ), .Z(_06617_ ) );
BUF_X4 _14607_ ( .A(_06617_ ), .Z(_06618_ ) );
BUF_X4 _14608_ ( .A(_06618_ ), .Z(_06619_ ) );
BUF_X2 _14609_ ( .A(_06619_ ), .Z(_06620_ ) );
NOR2_X1 _14610_ ( .A1(_06616_ ), .A2(_06620_ ), .ZN(_06621_ ) );
INV_X1 _14611_ ( .A(_06621_ ), .ZN(_06622_ ) );
BUF_X4 _14612_ ( .A(_05262_ ), .Z(_06623_ ) );
XNOR2_X1 _14613_ ( .A(_06553_ ), .B(_06623_ ), .ZN(_06624_ ) );
INV_X1 _14614_ ( .A(_06624_ ), .ZN(_06625_ ) );
BUF_X2 _14615_ ( .A(_06625_ ), .Z(_06626_ ) );
NAND3_X1 _14616_ ( .A1(_06608_ ), .A2(_06622_ ), .A3(_06626_ ), .ZN(_06627_ ) );
AOI22_X1 _14617_ ( .A1(_06600_ ), .A2(_06603_ ), .B1(_06604_ ), .B2(_06627_ ), .ZN(_06628_ ) );
BUF_X4 _14618_ ( .A(_05267_ ), .Z(_06629_ ) );
BUF_X4 _14619_ ( .A(_06629_ ), .Z(_06630_ ) );
BUF_X2 _14620_ ( .A(_06630_ ), .Z(_06631_ ) );
BUF_X4 _14621_ ( .A(_06613_ ), .Z(_06632_ ) );
NOR2_X1 _14622_ ( .A1(_06632_ ), .A2(_02748_ ), .ZN(_06633_ ) );
INV_X1 _14623_ ( .A(_05271_ ), .ZN(_06634_ ) );
BUF_X4 _14624_ ( .A(_06634_ ), .Z(_06635_ ) );
BUF_X4 _14625_ ( .A(_05273_ ), .Z(_06636_ ) );
BUF_X4 _14626_ ( .A(_05274_ ), .Z(_06637_ ) );
AOI21_X1 _14627_ ( .A(_02793_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06638_ ) );
NOR3_X1 _14628_ ( .A1(_06633_ ), .A2(_06635_ ), .A3(_06638_ ), .ZN(_06639_ ) );
NOR2_X1 _14629_ ( .A1(_06632_ ), .A2(_02162_ ), .ZN(_06640_ ) );
BUF_X4 _14630_ ( .A(_06636_ ), .Z(_06641_ ) );
BUF_X4 _14631_ ( .A(_06637_ ), .Z(_06642_ ) );
AOI21_X1 _14632_ ( .A(_02726_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06643_ ) );
NOR3_X1 _14633_ ( .A1(_06640_ ), .A2(_06643_ ), .A3(_06610_ ), .ZN(_06644_ ) );
OAI21_X1 _14634_ ( .A(_06631_ ), .B1(_06639_ ), .B2(_06644_ ), .ZN(_06645_ ) );
NOR2_X1 _14635_ ( .A1(_06613_ ), .A2(_02880_ ), .ZN(_06646_ ) );
AOI21_X1 _14636_ ( .A(_02834_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06647_ ) );
OAI21_X1 _14637_ ( .A(_06611_ ), .B1(_06646_ ), .B2(_06647_ ), .ZN(_06648_ ) );
BUF_X2 _14638_ ( .A(_06635_ ), .Z(_06649_ ) );
NOR2_X1 _14639_ ( .A1(_06613_ ), .A2(_02933_ ), .ZN(_06650_ ) );
AOI21_X1 _14640_ ( .A(_02858_ ), .B1(_05273_ ), .B2(_05274_ ), .ZN(_06651_ ) );
OAI21_X1 _14641_ ( .A(_06649_ ), .B1(_06650_ ), .B2(_06651_ ), .ZN(_06652_ ) );
NAND3_X1 _14642_ ( .A1(_06648_ ), .A2(_06652_ ), .A3(_06619_ ), .ZN(_06653_ ) );
NAND2_X1 _14643_ ( .A1(_06645_ ), .A2(_06653_ ), .ZN(_06654_ ) );
NAND2_X1 _14644_ ( .A1(_06613_ ), .A2(_05137_ ), .ZN(_06655_ ) );
BUF_X2 _14645_ ( .A(_05271_ ), .Z(_06656_ ) );
BUF_X4 _14646_ ( .A(_06636_ ), .Z(_06657_ ) );
BUF_X4 _14647_ ( .A(_06637_ ), .Z(_06658_ ) );
NAND3_X1 _14648_ ( .A1(_02962_ ), .A2(_06657_ ), .A3(_06658_ ), .ZN(_06659_ ) );
AND3_X1 _14649_ ( .A1(_06655_ ), .A2(_06656_ ), .A3(_06659_ ), .ZN(_06660_ ) );
AND2_X1 _14650_ ( .A1(_06614_ ), .A2(_02988_ ), .ZN(_06661_ ) );
AOI21_X1 _14651_ ( .A(_06660_ ), .B1(_06649_ ), .B2(_06661_ ), .ZN(_06662_ ) );
BUF_X4 _14652_ ( .A(_06618_ ), .Z(_06663_ ) );
NOR2_X1 _14653_ ( .A1(_06662_ ), .A2(_06663_ ), .ZN(_06664_ ) );
BUF_X2 _14654_ ( .A(_06623_ ), .Z(_06665_ ) );
MUX2_X1 _14655_ ( .A(_06654_ ), .B(_06664_ ), .S(_06665_ ), .Z(_06666_ ) );
BUF_X2 _14656_ ( .A(_05287_ ), .Z(_06667_ ) );
BUF_X2 _14657_ ( .A(_06667_ ), .Z(_06668_ ) );
BUF_X2 _14658_ ( .A(_06668_ ), .Z(_06669_ ) );
AND2_X1 _14659_ ( .A1(_06666_ ), .A2(_06669_ ), .ZN(_06670_ ) );
OAI21_X1 _14660_ ( .A(_06551_ ), .B1(_06628_ ), .B2(_06670_ ), .ZN(_06671_ ) );
NOR2_X1 _14661_ ( .A1(_05237_ ), .A2(_05314_ ), .ZN(_06672_ ) );
INV_X1 _14662_ ( .A(_06672_ ), .ZN(_06673_ ) );
NAND3_X1 _14663_ ( .A1(_05314_ ), .A2(_05236_ ), .A3(_05235_ ), .ZN(_06674_ ) );
AND3_X1 _14664_ ( .A1(_05234_ ), .A2(_06673_ ), .A3(_06674_ ), .ZN(_06675_ ) );
AND3_X1 _14665_ ( .A1(_06675_ ), .A2(_05226_ ), .A3(_05222_ ), .ZN(_06676_ ) );
INV_X1 _14666_ ( .A(_06676_ ), .ZN(_06677_ ) );
AND2_X1 _14667_ ( .A1(_05247_ ), .A2(_05243_ ), .ZN(_06678_ ) );
AND3_X1 _14668_ ( .A1(_06678_ ), .A2(_05252_ ), .A3(_05257_ ), .ZN(_06679_ ) );
INV_X1 _14669_ ( .A(_06679_ ), .ZN(_06680_ ) );
AND3_X1 _14670_ ( .A1(_05269_ ), .A2(_02282_ ), .A3(_05270_ ), .ZN(_06681_ ) );
INV_X1 _14671_ ( .A(_06681_ ), .ZN(_06682_ ) );
NAND2_X1 _14672_ ( .A1(_05271_ ), .A2(_02283_ ), .ZN(_06683_ ) );
INV_X1 _14673_ ( .A(_04110_ ), .ZN(_06684_ ) );
NOR2_X1 _14674_ ( .A1(_05275_ ), .A2(_06684_ ), .ZN(_06685_ ) );
AND3_X1 _14675_ ( .A1(_06682_ ), .A2(_06683_ ), .A3(_06685_ ), .ZN(_06686_ ) );
NOR2_X1 _14676_ ( .A1(_06686_ ), .A2(_06681_ ), .ZN(_06687_ ) );
INV_X1 _14677_ ( .A(_05268_ ), .ZN(_06688_ ) );
NOR2_X1 _14678_ ( .A1(_06687_ ), .A2(_06688_ ), .ZN(_06689_ ) );
NOR2_X1 _14679_ ( .A1(_05267_ ), .A2(_05281_ ), .ZN(_06690_ ) );
NOR2_X1 _14680_ ( .A1(_06689_ ), .A2(_06690_ ), .ZN(_06691_ ) );
OAI21_X1 _14681_ ( .A(_06691_ ), .B1(_02315_ ), .B2(_06554_ ), .ZN(_06692_ ) );
NOR2_X1 _14682_ ( .A1(_05262_ ), .A2(_02235_ ), .ZN(_06693_ ) );
INV_X1 _14683_ ( .A(_06693_ ), .ZN(_06694_ ) );
AND4_X1 _14684_ ( .A1(_05296_ ), .A2(_05288_ ), .A3(_05300_ ), .A4(_05292_ ), .ZN(_06695_ ) );
NAND3_X1 _14685_ ( .A1(_06692_ ), .A2(_06694_ ), .A3(_06695_ ), .ZN(_06696_ ) );
AND2_X1 _14686_ ( .A1(_05291_ ), .A2(_02188_ ), .ZN(_06697_ ) );
INV_X1 _14687_ ( .A(_06697_ ), .ZN(_06698_ ) );
NOR2_X1 _14688_ ( .A1(_05287_ ), .A2(_05305_ ), .ZN(_06699_ ) );
NAND2_X1 _14689_ ( .A1(_05292_ ), .A2(_06699_ ), .ZN(_06700_ ) );
AOI211_X1 _14690_ ( .A(_05303_ ), .B(_05304_ ), .C1(_06698_ ), .C2(_06700_ ), .ZN(_06701_ ) );
NOR2_X1 _14691_ ( .A1(_05295_ ), .A2(_02376_ ), .ZN(_06702_ ) );
OR2_X1 _14692_ ( .A1(_05299_ ), .A2(_06383_ ), .ZN(_06703_ ) );
AND3_X1 _14693_ ( .A1(_02376_ ), .A2(_05294_ ), .A3(_05293_ ), .ZN(_06704_ ) );
NOR3_X1 _14694_ ( .A1(_06703_ ), .A2(_06704_ ), .A3(_06702_ ), .ZN(_06705_ ) );
NOR3_X1 _14695_ ( .A1(_06701_ ), .A2(_06702_ ), .A3(_06705_ ), .ZN(_06706_ ) );
AOI211_X1 _14696_ ( .A(_06677_ ), .B(_06680_ ), .C1(_06696_ ), .C2(_06706_ ), .ZN(_06707_ ) );
NOR2_X1 _14697_ ( .A1(_05225_ ), .A2(_05404_ ), .ZN(_06708_ ) );
NOR2_X1 _14698_ ( .A1(_05251_ ), .A2(_02582_ ), .ZN(_06709_ ) );
NAND3_X1 _14699_ ( .A1(_02582_ ), .A2(_05250_ ), .A3(_05249_ ), .ZN(_06710_ ) );
NOR2_X1 _14700_ ( .A1(_05256_ ), .A2(_05323_ ), .ZN(_06711_ ) );
AOI21_X1 _14701_ ( .A(_06709_ ), .B1(_06710_ ), .B2(_06711_ ), .ZN(_06712_ ) );
INV_X1 _14702_ ( .A(_06712_ ), .ZN(_06713_ ) );
AND2_X1 _14703_ ( .A1(_06713_ ), .A2(_06678_ ), .ZN(_06714_ ) );
NOR2_X1 _14704_ ( .A1(_05246_ ), .A2(_02577_ ), .ZN(_06715_ ) );
NOR2_X1 _14705_ ( .A1(_05242_ ), .A2(_02574_ ), .ZN(_06716_ ) );
AND2_X1 _14706_ ( .A1(_05247_ ), .A2(_06716_ ), .ZN(_06717_ ) );
NOR3_X4 _14707_ ( .A1(_06714_ ), .A2(_06715_ ), .A3(_06717_ ), .ZN(_06718_ ) );
NOR2_X1 _14708_ ( .A1(_06718_ ), .A2(_06677_ ), .ZN(_06719_ ) );
INV_X1 _14709_ ( .A(_05222_ ), .ZN(_06720_ ) );
INV_X1 _14710_ ( .A(_05233_ ), .ZN(_06721_ ) );
AOI21_X1 _14711_ ( .A(_05232_ ), .B1(_06721_ ), .B2(_06672_ ), .ZN(_06722_ ) );
NOR3_X1 _14712_ ( .A1(_05319_ ), .A2(_06720_ ), .A3(_06722_ ), .ZN(_06723_ ) );
INV_X1 _14713_ ( .A(_02592_ ), .ZN(_06724_ ) );
NOR2_X1 _14714_ ( .A1(_05221_ ), .A2(_06724_ ), .ZN(_06725_ ) );
AND2_X1 _14715_ ( .A1(_05226_ ), .A2(_06725_ ), .ZN(_06726_ ) );
OR4_X4 _14716_ ( .A1(_06708_ ), .A2(_06719_ ), .A3(_06723_ ), .A4(_06726_ ), .ZN(_06727_ ) );
NOR2_X1 _14717_ ( .A1(_06707_ ), .A2(_06727_ ), .ZN(_06728_ ) );
INV_X1 _14718_ ( .A(_06728_ ), .ZN(_06729_ ) );
AND2_X1 _14719_ ( .A1(_05199_ ), .A2(_05335_ ), .ZN(_06730_ ) );
AND3_X1 _14720_ ( .A1(_06730_ ), .A2(_05194_ ), .A3(_05190_ ), .ZN(_06731_ ) );
AND2_X1 _14721_ ( .A1(_06729_ ), .A2(_06731_ ), .ZN(_06732_ ) );
INV_X1 _14722_ ( .A(_06732_ ), .ZN(_06733_ ) );
INV_X1 _14723_ ( .A(_02688_ ), .ZN(_06734_ ) );
NOR2_X1 _14724_ ( .A1(_05198_ ), .A2(_06734_ ), .ZN(_06735_ ) );
NOR2_X1 _14725_ ( .A1(_05203_ ), .A2(_05200_ ), .ZN(_06736_ ) );
AOI21_X1 _14726_ ( .A(_06735_ ), .B1(_05199_ ), .B2(_06736_ ), .ZN(_06737_ ) );
INV_X1 _14727_ ( .A(_05190_ ), .ZN(_06738_ ) );
INV_X1 _14728_ ( .A(_05194_ ), .ZN(_06739_ ) );
NOR3_X1 _14729_ ( .A1(_06737_ ), .A2(_06738_ ), .A3(_06739_ ), .ZN(_06740_ ) );
NOR2_X1 _14730_ ( .A1(_05193_ ), .A2(_05421_ ), .ZN(_06741_ ) );
NAND2_X1 _14731_ ( .A1(_05211_ ), .A2(_02642_ ), .ZN(_06742_ ) );
AND3_X1 _14732_ ( .A1(_05421_ ), .A2(_05192_ ), .A3(_05191_ ), .ZN(_06743_ ) );
NOR3_X1 _14733_ ( .A1(_06742_ ), .A2(_06743_ ), .A3(_06741_ ), .ZN(_06744_ ) );
NOR3_X1 _14734_ ( .A1(_06740_ ), .A2(_06741_ ), .A3(_06744_ ), .ZN(_06745_ ) );
AOI21_X1 _14735_ ( .A(_05180_ ), .B1(_06733_ ), .B2(_06745_ ), .ZN(_06746_ ) );
NOR2_X1 _14736_ ( .A1(_05178_ ), .A2(_02799_ ), .ZN(_06747_ ) );
OR3_X1 _14737_ ( .A1(_06746_ ), .A2(_06747_ ), .A3(_05184_ ), .ZN(_06748_ ) );
OAI21_X1 _14738_ ( .A(_05184_ ), .B1(_06746_ ), .B2(_06747_ ), .ZN(_06749_ ) );
NOR2_X1 _14739_ ( .A1(\ID_EX_typ [1] ), .A2(\ID_EX_typ [2] ), .ZN(_06750_ ) );
INV_X1 _14740_ ( .A(_06750_ ), .ZN(_06751_ ) );
NOR2_X1 _14741_ ( .A1(_05128_ ), .A2(_06751_ ), .ZN(_06752_ ) );
AND3_X1 _14742_ ( .A1(_06748_ ), .A2(_06749_ ), .A3(_06752_ ), .ZN(_06753_ ) );
BUF_X2 _14743_ ( .A(_05465_ ), .Z(_06754_ ) );
NOR2_X1 _14744_ ( .A1(_06614_ ), .A2(_02258_ ), .ZN(_06755_ ) );
AOI21_X1 _14745_ ( .A(_02235_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06756_ ) );
OR3_X1 _14746_ ( .A1(_06755_ ), .A2(_06756_ ), .A3(_06611_ ), .ZN(_06757_ ) );
BUF_X2 _14747_ ( .A(_06613_ ), .Z(_06758_ ) );
NOR2_X1 _14748_ ( .A1(_06758_ ), .A2(_02319_ ), .ZN(_06759_ ) );
AOI21_X1 _14749_ ( .A(_02188_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06760_ ) );
OR3_X1 _14750_ ( .A1(_06759_ ), .A2(_06649_ ), .A3(_06760_ ), .ZN(_06761_ ) );
NAND3_X1 _14751_ ( .A1(_06757_ ), .A2(_06761_ ), .A3(_06631_ ), .ZN(_06762_ ) );
BUF_X4 _14752_ ( .A(_06630_ ), .Z(_06763_ ) );
BUF_X4 _14753_ ( .A(_06763_ ), .Z(_06764_ ) );
BUF_X4 _14754_ ( .A(_06649_ ), .Z(_06765_ ) );
AOI21_X1 _14755_ ( .A(_02282_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06766_ ) );
NOR3_X1 _14756_ ( .A1(_05276_ ), .A2(_06765_ ), .A3(_06766_ ), .ZN(_06767_ ) );
OAI21_X1 _14757_ ( .A(_06762_ ), .B1(_06764_ ), .B2(_06767_ ), .ZN(_06768_ ) );
BUF_X4 _14758_ ( .A(_06623_ ), .Z(_06769_ ) );
BUF_X2 _14759_ ( .A(_06769_ ), .Z(_06770_ ) );
NOR2_X1 _14760_ ( .A1(_06768_ ), .A2(_06770_ ), .ZN(_06771_ ) );
BUF_X2 _14761_ ( .A(_06667_ ), .Z(_06772_ ) );
BUF_X2 _14762_ ( .A(_06772_ ), .Z(_06773_ ) );
OAI21_X1 _14763_ ( .A(_06754_ ), .B1(_06771_ ), .B2(_06773_ ), .ZN(_06774_ ) );
AOI21_X1 _14764_ ( .A(_02399_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06775_ ) );
INV_X1 _14765_ ( .A(_06775_ ), .ZN(_06776_ ) );
BUF_X2 _14766_ ( .A(_06635_ ), .Z(_06777_ ) );
OAI211_X1 _14767_ ( .A(_06776_ ), .B(_06777_ ), .C1(_02422_ ), .C2(_06615_ ), .ZN(_06778_ ) );
AOI21_X1 _14768_ ( .A(_02565_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06779_ ) );
INV_X1 _14769_ ( .A(_06779_ ), .ZN(_06780_ ) );
BUF_X4 _14770_ ( .A(_06610_ ), .Z(_06781_ ) );
OAI211_X1 _14771_ ( .A(_06780_ ), .B(_06781_ ), .C1(_02588_ ), .C2(_06615_ ), .ZN(_06782_ ) );
BUF_X2 _14772_ ( .A(_06630_ ), .Z(_06783_ ) );
AND3_X1 _14773_ ( .A1(_06778_ ), .A2(_06782_ ), .A3(_06783_ ), .ZN(_06784_ ) );
BUF_X4 _14774_ ( .A(_06554_ ), .Z(_06785_ ) );
BUF_X2 _14775_ ( .A(_06785_ ), .Z(_06786_ ) );
BUF_X2 _14776_ ( .A(_06786_ ), .Z(_06787_ ) );
NOR2_X1 _14777_ ( .A1(_06758_ ), .A2(_02448_ ), .ZN(_06788_ ) );
AOI21_X1 _14778_ ( .A(_02472_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06789_ ) );
OAI21_X1 _14779_ ( .A(_06781_ ), .B1(_06788_ ), .B2(_06789_ ), .ZN(_06790_ ) );
NOR2_X1 _14780_ ( .A1(_06758_ ), .A2(_02371_ ), .ZN(_06791_ ) );
AOI21_X1 _14781_ ( .A(_02345_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06792_ ) );
OAI21_X1 _14782_ ( .A(_06765_ ), .B1(_06791_ ), .B2(_06792_ ), .ZN(_06793_ ) );
AOI21_X1 _14783_ ( .A(_06783_ ), .B1(_06790_ ), .B2(_06793_ ), .ZN(_06794_ ) );
OR3_X1 _14784_ ( .A1(_06784_ ), .A2(_06787_ ), .A3(_06794_ ), .ZN(_06795_ ) );
NOR2_X1 _14785_ ( .A1(_06615_ ), .A2(_02592_ ), .ZN(_06796_ ) );
AOI21_X1 _14786_ ( .A(_02518_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06797_ ) );
OR3_X1 _14787_ ( .A1(_06796_ ), .A2(_06612_ ), .A3(_06797_ ), .ZN(_06798_ ) );
AOI21_X1 _14788_ ( .A(_02688_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06799_ ) );
INV_X1 _14789_ ( .A(_06799_ ), .ZN(_06800_ ) );
BUF_X4 _14790_ ( .A(_06781_ ), .Z(_06801_ ) );
OAI211_X1 _14791_ ( .A(_06800_ ), .B(_06801_ ), .C1(_02666_ ), .C2(_06615_ ), .ZN(_06802_ ) );
AOI21_X1 _14792_ ( .A(_06764_ ), .B1(_06798_ ), .B2(_06802_ ), .ZN(_06803_ ) );
NOR2_X1 _14793_ ( .A1(_06758_ ), .A2(_02770_ ), .ZN(_06804_ ) );
OAI21_X1 _14794_ ( .A(_06612_ ), .B1(_06804_ ), .B2(_06638_ ), .ZN(_06805_ ) );
BUF_X4 _14795_ ( .A(_06777_ ), .Z(_06806_ ) );
NOR2_X1 _14796_ ( .A1(_06614_ ), .A2(_02642_ ), .ZN(_06807_ ) );
AOI21_X1 _14797_ ( .A(_02618_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06808_ ) );
OAI21_X1 _14798_ ( .A(_06806_ ), .B1(_06807_ ), .B2(_06808_ ), .ZN(_06809_ ) );
AND3_X1 _14799_ ( .A1(_06805_ ), .A2(_06809_ ), .A3(_06631_ ), .ZN(_06810_ ) );
OAI21_X1 _14800_ ( .A(_06787_ ), .B1(_06803_ ), .B2(_06810_ ), .ZN(_06811_ ) );
AND2_X1 _14801_ ( .A1(_06811_ ), .A2(_06773_ ), .ZN(_06812_ ) );
AOI21_X1 _14802_ ( .A(_06774_ ), .B1(_06795_ ), .B2(_06812_ ), .ZN(_06813_ ) );
AND2_X1 _14803_ ( .A1(_05184_ ), .A2(_05386_ ), .ZN(_06814_ ) );
BUF_X4 _14804_ ( .A(_05383_ ), .Z(_06815_ ) );
AOI21_X1 _14805_ ( .A(_06815_ ), .B1(_05183_ ), .B2(_06204_ ), .ZN(_06816_ ) );
OR2_X1 _14806_ ( .A1(_06814_ ), .A2(_06816_ ), .ZN(_06817_ ) );
BUF_X2 _14807_ ( .A(_06668_ ), .Z(_06818_ ) );
AND2_X1 _14808_ ( .A1(_05380_ ), .A2(\ID_EX_typ [2] ), .ZN(_06819_ ) );
BUF_X2 _14809_ ( .A(_06819_ ), .Z(_06820_ ) );
NAND3_X1 _14810_ ( .A1(_06666_ ), .A2(_06818_ ), .A3(_06820_ ), .ZN(_06821_ ) );
OR3_X1 _14811_ ( .A1(_05183_ ), .A2(_06204_ ), .A3(_05129_ ), .ZN(_06822_ ) );
NAND2_X1 _14812_ ( .A1(_06821_ ), .A2(_06822_ ), .ZN(_06823_ ) );
NOR4_X1 _14813_ ( .A1(_06753_ ), .A2(_06813_ ), .A3(_06817_ ), .A4(_06823_ ), .ZN(_06824_ ) );
AOI21_X1 _14814_ ( .A(_06549_ ), .B1(_06671_ ), .B2(_06824_ ), .ZN(_06825_ ) );
BUF_X4 _14815_ ( .A(_06547_ ), .Z(_06826_ ) );
NAND2_X1 _14816_ ( .A1(_05418_ ), .A2(_04756_ ), .ZN(_06827_ ) );
AND2_X1 _14817_ ( .A1(_06827_ ), .A2(_05427_ ), .ZN(_06828_ ) );
INV_X1 _14818_ ( .A(_04660_ ), .ZN(_06829_ ) );
NOR2_X1 _14819_ ( .A1(_06828_ ), .A2(_06829_ ), .ZN(_06830_ ) );
OR3_X1 _14820_ ( .A1(_06830_ ), .A2(_04637_ ), .A3(_05431_ ), .ZN(_06831_ ) );
AND3_X1 _14821_ ( .A1(_04322_ ), .A2(\ID_EX_typ [3] ), .A3(_05468_ ), .ZN(_06832_ ) );
AND2_X1 _14822_ ( .A1(_06832_ ), .A2(_05133_ ), .ZN(_06833_ ) );
BUF_X4 _14823_ ( .A(_06833_ ), .Z(_06834_ ) );
BUF_X4 _14824_ ( .A(_06834_ ), .Z(_06835_ ) );
OAI21_X1 _14825_ ( .A(_04637_ ), .B1(_06830_ ), .B2(_05431_ ), .ZN(_06836_ ) );
NAND3_X1 _14826_ ( .A1(_06831_ ), .A2(_06835_ ), .A3(_06836_ ), .ZN(_06837_ ) );
AND2_X2 _14827_ ( .A1(_06540_ ), .A2(_06539_ ), .ZN(_06838_ ) );
BUF_X2 _14828_ ( .A(_06838_ ), .Z(_06839_ ) );
AND2_X2 _14829_ ( .A1(_06541_ ), .A2(_06539_ ), .ZN(_06840_ ) );
BUF_X4 _14830_ ( .A(_06840_ ), .Z(_06841_ ) );
AOI22_X1 _14831_ ( .A1(_06136_ ), .A2(_06839_ ), .B1(\ID_EX_imm [21] ), .B2(_06841_ ), .ZN(_06842_ ) );
AOI21_X1 _14832_ ( .A(_06826_ ), .B1(_06837_ ), .B2(_06842_ ), .ZN(_06843_ ) );
OR2_X1 _14833_ ( .A1(_06843_ ), .A2(_05569_ ), .ZN(_06844_ ) );
BUF_X4 _14834_ ( .A(_05485_ ), .Z(_06845_ ) );
OAI22_X1 _14835_ ( .A1(_06825_ ), .A2(_06844_ ), .B1(_06845_ ), .B2(_06135_ ), .ZN(_06846_ ) );
OAI21_X1 _14836_ ( .A(_06538_ ), .B1(_06846_ ), .B2(_06387_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_10_D ) );
AND2_X1 _14837_ ( .A1(_05646_ ), .A2(_06231_ ), .ZN(_06847_ ) );
OAI21_X1 _14838_ ( .A(_06286_ ), .B1(_06847_ ), .B2(_06225_ ), .ZN(_06848_ ) );
OAI21_X1 _14839_ ( .A(_06834_ ), .B1(_06828_ ), .B2(_06829_ ), .ZN(_06849_ ) );
AOI21_X1 _14840_ ( .A(_06849_ ), .B1(_06829_ ), .B2(_06828_ ), .ZN(_06850_ ) );
BUF_X2 _14841_ ( .A(_06838_ ), .Z(_06851_ ) );
AND2_X1 _14842_ ( .A1(_04321_ ), .A2(_06851_ ), .ZN(_06852_ ) );
AND3_X1 _14843_ ( .A1(_06541_ ), .A2(\ID_EX_imm [20] ), .A3(_06539_ ), .ZN(_06853_ ) );
NOR3_X1 _14844_ ( .A1(_06850_ ), .A2(_06852_ ), .A3(_06853_ ), .ZN(_06854_ ) );
AOI21_X1 _14845_ ( .A(_05482_ ), .B1(_06854_ ), .B2(_03344_ ), .ZN(_06855_ ) );
INV_X1 _14846_ ( .A(_06550_ ), .ZN(_06856_ ) );
INV_X1 _14847_ ( .A(_06632_ ), .ZN(_06857_ ) );
OAI21_X1 _14848_ ( .A(_06631_ ), .B1(_06806_ ), .B2(_06857_ ), .ZN(_06858_ ) );
AND3_X1 _14849_ ( .A1(_06607_ ), .A2(_06625_ ), .A3(_06858_ ), .ZN(_06859_ ) );
AND2_X1 _14850_ ( .A1(_06607_ ), .A2(_06599_ ), .ZN(_06860_ ) );
OAI22_X1 _14851_ ( .A1(_06859_ ), .A2(_06601_ ), .B1(_06860_ ), .B2(_06602_ ), .ZN(_06861_ ) );
NOR2_X1 _14852_ ( .A1(_06613_ ), .A2(_02834_ ), .ZN(_06862_ ) );
AOI21_X1 _14853_ ( .A(_02162_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06863_ ) );
NOR2_X1 _14854_ ( .A1(_06862_ ), .A2(_06863_ ), .ZN(_06864_ ) );
BUF_X2 _14855_ ( .A(_06634_ ), .Z(_06865_ ) );
NOR2_X1 _14856_ ( .A1(_06864_ ), .A2(_06865_ ), .ZN(_06866_ ) );
AOI21_X1 _14857_ ( .A(_02880_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06867_ ) );
INV_X1 _14858_ ( .A(_06867_ ), .ZN(_06868_ ) );
NAND3_X1 _14859_ ( .A1(_05443_ ), .A2(_06657_ ), .A3(_06658_ ), .ZN(_06869_ ) );
AOI21_X1 _14860_ ( .A(_06609_ ), .B1(_06868_ ), .B2(_06869_ ), .ZN(_06870_ ) );
OR3_X1 _14861_ ( .A1(_06866_ ), .A2(_06629_ ), .A3(_06870_ ), .ZN(_06871_ ) );
NOR2_X1 _14862_ ( .A1(_06632_ ), .A2(_02793_ ), .ZN(_06872_ ) );
AOI21_X1 _14863_ ( .A(_02770_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06873_ ) );
OAI21_X1 _14864_ ( .A(_06656_ ), .B1(_06872_ ), .B2(_06873_ ), .ZN(_06874_ ) );
NOR2_X1 _14865_ ( .A1(_06613_ ), .A2(_02726_ ), .ZN(_06875_ ) );
AOI21_X1 _14866_ ( .A(_02748_ ), .B1(_05273_ ), .B2(_05274_ ), .ZN(_06876_ ) );
OAI21_X1 _14867_ ( .A(_06635_ ), .B1(_06875_ ), .B2(_06876_ ), .ZN(_06877_ ) );
NAND3_X1 _14868_ ( .A1(_06874_ ), .A2(_06877_ ), .A3(_06630_ ), .ZN(_06878_ ) );
NAND2_X1 _14869_ ( .A1(_06871_ ), .A2(_06878_ ), .ZN(_06879_ ) );
NOR2_X1 _14870_ ( .A1(_06613_ ), .A2(_02909_ ), .ZN(_06880_ ) );
AOI21_X1 _14871_ ( .A(_02933_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06881_ ) );
NOR2_X1 _14872_ ( .A1(_06880_ ), .A2(_06881_ ), .ZN(_06882_ ) );
INV_X1 _14873_ ( .A(_02962_ ), .ZN(_06883_ ) );
MUX2_X1 _14874_ ( .A(_02988_ ), .B(_06883_ ), .S(_06613_ ), .Z(_06884_ ) );
MUX2_X1 _14875_ ( .A(_06882_ ), .B(_06884_ ), .S(_06634_ ), .Z(_06885_ ) );
AND2_X1 _14876_ ( .A1(_06885_ ), .A2(_06763_ ), .ZN(_06886_ ) );
MUX2_X1 _14877_ ( .A(_06879_ ), .B(_06886_ ), .S(_06769_ ), .Z(_06887_ ) );
CLKBUF_X2 _14878_ ( .A(_06772_ ), .Z(_06888_ ) );
NAND2_X1 _14879_ ( .A1(_06887_ ), .A2(_06888_ ), .ZN(_06889_ ) );
AOI21_X1 _14880_ ( .A(_06856_ ), .B1(_06861_ ), .B2(_06889_ ), .ZN(_06890_ ) );
INV_X1 _14881_ ( .A(_06754_ ), .ZN(_06891_ ) );
NOR2_X1 _14882_ ( .A1(_06758_ ), .A2(_02345_ ), .ZN(_06892_ ) );
AOI21_X1 _14883_ ( .A(_02448_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06893_ ) );
NOR3_X1 _14884_ ( .A1(_06892_ ), .A2(_06777_ ), .A3(_06893_ ), .ZN(_06894_ ) );
NOR2_X1 _14885_ ( .A1(_06632_ ), .A2(_02188_ ), .ZN(_06895_ ) );
AOI21_X1 _14886_ ( .A(_02371_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06896_ ) );
NOR3_X1 _14887_ ( .A1(_06895_ ), .A2(_06896_ ), .A3(_06611_ ), .ZN(_06897_ ) );
NOR2_X1 _14888_ ( .A1(_06894_ ), .A2(_06897_ ), .ZN(_06898_ ) );
NOR2_X1 _14889_ ( .A1(_06898_ ), .A2(_06783_ ), .ZN(_06899_ ) );
BUF_X4 _14890_ ( .A(_06785_ ), .Z(_06900_ ) );
NOR2_X1 _14891_ ( .A1(_06632_ ), .A2(_02399_ ), .ZN(_06901_ ) );
AOI21_X1 _14892_ ( .A(_02588_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06902_ ) );
OR3_X1 _14893_ ( .A1(_06901_ ), .A2(_06649_ ), .A3(_06902_ ), .ZN(_06903_ ) );
NOR2_X1 _14894_ ( .A1(_06758_ ), .A2(_02472_ ), .ZN(_06904_ ) );
AOI21_X1 _14895_ ( .A(_02422_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06905_ ) );
OR3_X1 _14896_ ( .A1(_06904_ ), .A2(_06905_ ), .A3(_06610_ ), .ZN(_06906_ ) );
AOI21_X1 _14897_ ( .A(_06619_ ), .B1(_06903_ ), .B2(_06906_ ), .ZN(_06907_ ) );
OR3_X1 _14898_ ( .A1(_06899_ ), .A2(_06900_ ), .A3(_06907_ ), .ZN(_06908_ ) );
NOR2_X1 _14899_ ( .A1(_06758_ ), .A2(_02518_ ), .ZN(_06909_ ) );
AOI21_X1 _14900_ ( .A(_02666_ ), .B1(_06641_ ), .B2(_06642_ ), .ZN(_06910_ ) );
OR3_X1 _14901_ ( .A1(_06909_ ), .A2(_06649_ ), .A3(_06910_ ), .ZN(_06911_ ) );
NOR2_X1 _14902_ ( .A1(_06632_ ), .A2(_02565_ ), .ZN(_06912_ ) );
AOI21_X1 _14903_ ( .A(_02592_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06913_ ) );
OR3_X1 _14904_ ( .A1(_06912_ ), .A2(_06913_ ), .A3(_06610_ ), .ZN(_06914_ ) );
AOI21_X1 _14905_ ( .A(_06763_ ), .B1(_06911_ ), .B2(_06914_ ), .ZN(_06915_ ) );
NOR2_X1 _14906_ ( .A1(_06632_ ), .A2(_02618_ ), .ZN(_06916_ ) );
OAI21_X1 _14907_ ( .A(_06611_ ), .B1(_06916_ ), .B2(_06873_ ), .ZN(_06917_ ) );
NOR2_X1 _14908_ ( .A1(_06758_ ), .A2(_02688_ ), .ZN(_06918_ ) );
AOI21_X1 _14909_ ( .A(_02642_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06919_ ) );
OAI21_X1 _14910_ ( .A(_06777_ ), .B1(_06918_ ), .B2(_06919_ ), .ZN(_06920_ ) );
AND3_X1 _14911_ ( .A1(_06917_ ), .A2(_06920_ ), .A3(_06763_ ), .ZN(_06921_ ) );
OR3_X1 _14912_ ( .A1(_06915_ ), .A2(_06921_ ), .A3(_06769_ ), .ZN(_06922_ ) );
NAND3_X1 _14913_ ( .A1(_06908_ ), .A2(_06888_ ), .A3(_06922_ ), .ZN(_06923_ ) );
NOR2_X1 _14914_ ( .A1(_06632_ ), .A2(_02235_ ), .ZN(_06924_ ) );
AOI21_X1 _14915_ ( .A(_02319_ ), .B1(_06657_ ), .B2(_06658_ ), .ZN(_06925_ ) );
OAI21_X1 _14916_ ( .A(_06610_ ), .B1(_06924_ ), .B2(_06925_ ), .ZN(_06926_ ) );
NOR2_X1 _14917_ ( .A1(_06632_ ), .A2(_02282_ ), .ZN(_06927_ ) );
AOI21_X1 _14918_ ( .A(_02258_ ), .B1(_06636_ ), .B2(_06637_ ), .ZN(_06928_ ) );
OAI21_X1 _14919_ ( .A(_06649_ ), .B1(_06927_ ), .B2(_06928_ ), .ZN(_06929_ ) );
NAND3_X1 _14920_ ( .A1(_06926_ ), .A2(_06929_ ), .A3(_06630_ ), .ZN(_06930_ ) );
NAND4_X1 _14921_ ( .A1(_06618_ ), .A2(_04110_ ), .A3(_06611_ ), .A4(_06615_ ), .ZN(_06931_ ) );
AND2_X1 _14922_ ( .A1(_06930_ ), .A2(_06931_ ), .ZN(_06932_ ) );
OR3_X1 _14923_ ( .A1(_06932_ ), .A2(_06772_ ), .A3(_06665_ ), .ZN(_06933_ ) );
AOI21_X1 _14924_ ( .A(_06891_ ), .B1(_06923_ ), .B2(_06933_ ), .ZN(_06934_ ) );
AND3_X1 _14925_ ( .A1(_06887_ ), .A2(_06888_ ), .A3(_06820_ ), .ZN(_06935_ ) );
OR3_X1 _14926_ ( .A1(_06890_ ), .A2(_06934_ ), .A3(_06935_ ), .ZN(_06936_ ) );
AND2_X1 _14927_ ( .A1(_06733_ ), .A2(_06745_ ), .ZN(_06937_ ) );
OAI21_X1 _14928_ ( .A(_06752_ ), .B1(_06937_ ), .B2(_05180_ ), .ZN(_06938_ ) );
AOI21_X1 _14929_ ( .A(_06938_ ), .B1(_05180_ ), .B2(_06937_ ), .ZN(_06939_ ) );
BUF_X2 _14930_ ( .A(_05386_ ), .Z(_06940_ ) );
AND2_X1 _14931_ ( .A1(_05179_ ), .A2(_06940_ ), .ZN(_06941_ ) );
NOR3_X1 _14932_ ( .A1(_05178_ ), .A2(_02799_ ), .A3(_05129_ ), .ZN(_06942_ ) );
AOI21_X1 _14933_ ( .A(_06815_ ), .B1(_05178_ ), .B2(_02799_ ), .ZN(_06943_ ) );
OR3_X1 _14934_ ( .A1(_06941_ ), .A2(_06942_ ), .A3(_06943_ ), .ZN(_06944_ ) );
OR3_X1 _14935_ ( .A1(_06936_ ), .A2(_06939_ ), .A3(_06944_ ), .ZN(_06945_ ) );
INV_X1 _14936_ ( .A(_06548_ ), .ZN(_06946_ ) );
BUF_X4 _14937_ ( .A(_06946_ ), .Z(_06947_ ) );
BUF_X4 _14938_ ( .A(_06947_ ), .Z(_06948_ ) );
AOI21_X1 _14939_ ( .A(_06855_ ), .B1(_06945_ ), .B2(_06948_ ), .ZN(_06949_ ) );
OAI21_X1 _14940_ ( .A(_06409_ ), .B1(_04241_ ), .B2(_05486_ ), .ZN(_06950_ ) );
OAI21_X1 _14941_ ( .A(_06848_ ), .B1(_06949_ ), .B2(_06950_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _14942_ ( .A1(_05646_ ), .A2(_05647_ ), .A3(_05549_ ), .ZN(_06951_ ) );
BUF_X4 _14943_ ( .A(_04105_ ), .Z(_06952_ ) );
INV_X1 _14944_ ( .A(_05522_ ), .ZN(_06953_ ) );
NAND3_X1 _14945_ ( .A1(_06951_ ), .A2(_06952_ ), .A3(_06953_ ), .ZN(_06954_ ) );
INV_X1 _14946_ ( .A(_06834_ ), .ZN(_06955_ ) );
BUF_X4 _14947_ ( .A(_06955_ ), .Z(_06956_ ) );
NAND2_X1 _14948_ ( .A1(_02642_ ), .A2(_04682_ ), .ZN(_06957_ ) );
AOI21_X1 _14949_ ( .A(_05426_ ), .B1(_05418_ ), .B2(_04755_ ), .ZN(_06958_ ) );
INV_X1 _14950_ ( .A(_04683_ ), .ZN(_06959_ ) );
OAI21_X1 _14951_ ( .A(_06957_ ), .B1(_06958_ ), .B2(_06959_ ), .ZN(_06960_ ) );
AOI21_X1 _14952_ ( .A(_06956_ ), .B1(_06960_ ), .B2(_04709_ ), .ZN(_06961_ ) );
OAI21_X1 _14953_ ( .A(_06961_ ), .B1(_04709_ ), .B2(_06960_ ), .ZN(_06962_ ) );
AOI22_X1 _14954_ ( .A1(_05497_ ), .A2(_06851_ ), .B1(\ID_EX_imm [19] ), .B2(_06841_ ), .ZN(_06963_ ) );
AOI21_X1 _14955_ ( .A(_06826_ ), .B1(_06962_ ), .B2(_06963_ ), .ZN(_06964_ ) );
OR2_X1 _14956_ ( .A1(_06964_ ), .A2(_05569_ ), .ZN(_06965_ ) );
BUF_X4 _14957_ ( .A(_06856_ ), .Z(_06966_ ) );
AND2_X2 _14958_ ( .A1(_06599_ ), .A2(_06601_ ), .ZN(_06967_ ) );
AND2_X1 _14959_ ( .A1(_06598_ ), .A2(_06967_ ), .ZN(_06968_ ) );
NOR3_X1 _14960_ ( .A1(_06804_ ), .A2(_06865_ ), .A3(_06808_ ), .ZN(_06969_ ) );
NOR3_X1 _14961_ ( .A1(_06633_ ), .A2(_06638_ ), .A3(_06609_ ), .ZN(_06970_ ) );
NOR3_X1 _14962_ ( .A1(_06969_ ), .A2(_06970_ ), .A3(_06617_ ), .ZN(_06971_ ) );
OAI21_X1 _14963_ ( .A(_06656_ ), .B1(_06640_ ), .B2(_06643_ ), .ZN(_06972_ ) );
OAI21_X1 _14964_ ( .A(_06865_ ), .B1(_06646_ ), .B2(_06647_ ), .ZN(_06973_ ) );
AOI21_X1 _14965_ ( .A(_05267_ ), .B1(_06972_ ), .B2(_06973_ ), .ZN(_06974_ ) );
NOR2_X1 _14966_ ( .A1(_06971_ ), .A2(_06974_ ), .ZN(_06975_ ) );
OR3_X1 _14967_ ( .A1(_06650_ ), .A2(_06634_ ), .A3(_06651_ ), .ZN(_06976_ ) );
NAND3_X1 _14968_ ( .A1(_06655_ ), .A2(_06634_ ), .A3(_06659_ ), .ZN(_06977_ ) );
AOI21_X1 _14969_ ( .A(_06617_ ), .B1(_06976_ ), .B2(_06977_ ), .ZN(_06978_ ) );
AND4_X1 _14970_ ( .A1(_02988_ ), .A2(_06617_ ), .A3(_06609_ ), .A4(_06758_ ), .ZN(_06979_ ) );
OR2_X1 _14971_ ( .A1(_06978_ ), .A2(_06979_ ), .ZN(_06980_ ) );
MUX2_X1 _14972_ ( .A(_06975_ ), .B(_06980_ ), .S(_06623_ ), .Z(_06981_ ) );
AOI21_X1 _14973_ ( .A(_06968_ ), .B1(_06669_ ), .B2(_06981_ ), .ZN(_06982_ ) );
XNOR2_X1 _14974_ ( .A(_06552_ ), .B(_06630_ ), .ZN(_06983_ ) );
NAND4_X1 _14975_ ( .A1(_06608_ ), .A2(_06626_ ), .A3(_06983_ ), .A4(_06599_ ), .ZN(_06984_ ) );
AOI21_X1 _14976_ ( .A(_06966_ ), .B1(_06982_ ), .B2(_06984_ ), .ZN(_06985_ ) );
BUF_X2 _14977_ ( .A(_06820_ ), .Z(_06986_ ) );
NAND3_X1 _14978_ ( .A1(_06981_ ), .A2(_06669_ ), .A3(_06986_ ), .ZN(_06987_ ) );
BUF_X4 _14979_ ( .A(_05306_ ), .Z(_06988_ ) );
BUF_X4 _14980_ ( .A(_06988_ ), .Z(_06989_ ) );
NOR3_X1 _14981_ ( .A1(_06796_ ), .A2(_06765_ ), .A3(_06797_ ), .ZN(_06990_ ) );
NOR2_X1 _14982_ ( .A1(_06615_ ), .A2(_02588_ ), .ZN(_06991_ ) );
NOR3_X1 _14983_ ( .A1(_06991_ ), .A2(_06779_ ), .A3(_06781_ ), .ZN(_06992_ ) );
NOR2_X1 _14984_ ( .A1(_06990_ ), .A2(_06992_ ), .ZN(_06993_ ) );
NOR2_X1 _14985_ ( .A1(_06993_ ), .A2(_06764_ ), .ZN(_06994_ ) );
BUF_X4 _14986_ ( .A(_06769_ ), .Z(_06995_ ) );
OR3_X1 _14987_ ( .A1(_06807_ ), .A2(_06777_ ), .A3(_06808_ ), .ZN(_06996_ ) );
OAI211_X1 _14988_ ( .A(_06800_ ), .B(_06765_ ), .C1(_02666_ ), .C2(_06615_ ), .ZN(_06997_ ) );
AOI21_X1 _14989_ ( .A(_06663_ ), .B1(_06996_ ), .B2(_06997_ ), .ZN(_06998_ ) );
OR3_X1 _14990_ ( .A1(_06994_ ), .A2(_06995_ ), .A3(_06998_ ), .ZN(_06999_ ) );
BUF_X4 _14991_ ( .A(_06995_ ), .Z(_07000_ ) );
NOR2_X1 _14992_ ( .A1(_06758_ ), .A2(_02422_ ), .ZN(_07001_ ) );
OAI21_X1 _14993_ ( .A(_06612_ ), .B1(_07001_ ), .B2(_06775_ ), .ZN(_07002_ ) );
OAI21_X1 _14994_ ( .A(_06765_ ), .B1(_06788_ ), .B2(_06789_ ), .ZN(_07003_ ) );
AOI21_X1 _14995_ ( .A(_06663_ ), .B1(_07002_ ), .B2(_07003_ ), .ZN(_07004_ ) );
OAI21_X1 _14996_ ( .A(_06612_ ), .B1(_06791_ ), .B2(_06792_ ), .ZN(_07005_ ) );
OAI21_X1 _14997_ ( .A(_06765_ ), .B1(_06759_ ), .B2(_06760_ ), .ZN(_07006_ ) );
AOI21_X1 _14998_ ( .A(_06783_ ), .B1(_07005_ ), .B2(_07006_ ), .ZN(_07007_ ) );
OAI21_X1 _14999_ ( .A(_07000_ ), .B1(_07004_ ), .B2(_07007_ ), .ZN(_07008_ ) );
AOI21_X1 _15000_ ( .A(_06989_ ), .B1(_06999_ ), .B2(_07008_ ), .ZN(_07009_ ) );
OR3_X1 _15001_ ( .A1(_06755_ ), .A2(_06777_ ), .A3(_06756_ ), .ZN(_07010_ ) );
OR3_X1 _15002_ ( .A1(_05276_ ), .A2(_06766_ ), .A3(_06781_ ), .ZN(_07011_ ) );
AOI21_X1 _15003_ ( .A(_06620_ ), .B1(_07010_ ), .B2(_07011_ ), .ZN(_07012_ ) );
AND2_X1 _15004_ ( .A1(_07012_ ), .A2(_06787_ ), .ZN(_07013_ ) );
OAI21_X1 _15005_ ( .A(_06754_ ), .B1(_07013_ ), .B2(_06818_ ), .ZN(_07014_ ) );
OAI221_X1 _15006_ ( .A(_06987_ ), .B1(_06743_ ), .B2(_06815_ ), .C1(_07009_ ), .C2(_07014_ ), .ZN(_07015_ ) );
BUF_X4 _15007_ ( .A(_05128_ ), .Z(_07016_ ) );
BUF_X4 _15008_ ( .A(_07016_ ), .Z(_07017_ ) );
NAND2_X1 _15009_ ( .A1(_06741_ ), .A2(_07017_ ), .ZN(_07018_ ) );
OAI21_X1 _15010_ ( .A(_06730_ ), .B1(_06707_ ), .B2(_06727_ ), .ZN(_07019_ ) );
AND2_X1 _15011_ ( .A1(_07019_ ), .A2(_06737_ ), .ZN(_07020_ ) );
OAI21_X1 _15012_ ( .A(_06742_ ), .B1(_07020_ ), .B2(_06738_ ), .ZN(_07021_ ) );
XNOR2_X1 _15013_ ( .A(_07021_ ), .B(_05194_ ), .ZN(_07022_ ) );
INV_X1 _15014_ ( .A(_06752_ ), .ZN(_07023_ ) );
BUF_X4 _15015_ ( .A(_07023_ ), .Z(_07024_ ) );
OAI221_X1 _15016_ ( .A(_07018_ ), .B1(_06739_ ), .B2(_05387_ ), .C1(_07022_ ), .C2(_07024_ ), .ZN(_07025_ ) );
OR3_X1 _15017_ ( .A1(_06985_ ), .A2(_07015_ ), .A3(_07025_ ), .ZN(_07026_ ) );
AOI21_X1 _15018_ ( .A(_06965_ ), .B1(_07026_ ), .B2(_06948_ ), .ZN(_07027_ ) );
NAND2_X1 _15019_ ( .A1(_05508_ ), .A2(_06016_ ), .ZN(_07028_ ) );
NAND2_X1 _15020_ ( .A1(_07028_ ), .A2(_04108_ ), .ZN(_07029_ ) );
OAI21_X1 _15021_ ( .A(_06954_ ), .B1(_07027_ ), .B2(_07029_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_12_D ) );
NAND3_X1 _15022_ ( .A1(_05646_ ), .A2(_05647_ ), .A3(_05563_ ), .ZN(_07030_ ) );
INV_X1 _15023_ ( .A(_05558_ ), .ZN(_07031_ ) );
NAND3_X1 _15024_ ( .A1(_07030_ ), .A2(_06952_ ), .A3(_07031_ ), .ZN(_07032_ ) );
OAI21_X1 _15025_ ( .A(_06834_ ), .B1(_06958_ ), .B2(_06959_ ), .ZN(_07033_ ) );
AOI21_X1 _15026_ ( .A(_07033_ ), .B1(_06959_ ), .B2(_06958_ ), .ZN(_07034_ ) );
AND2_X1 _15027_ ( .A1(_05556_ ), .A2(_06851_ ), .ZN(_07035_ ) );
AND3_X1 _15028_ ( .A1(_06541_ ), .A2(\ID_EX_imm [18] ), .A3(_06539_ ), .ZN(_07036_ ) );
NOR3_X1 _15029_ ( .A1(_07034_ ), .A2(_07035_ ), .A3(_07036_ ), .ZN(_07037_ ) );
AOI21_X1 _15030_ ( .A(_05482_ ), .B1(_07037_ ), .B2(_03344_ ), .ZN(_07038_ ) );
NOR2_X1 _15031_ ( .A1(_06635_ ), .A2(_06614_ ), .ZN(_07039_ ) );
INV_X1 _15032_ ( .A(_07039_ ), .ZN(_07040_ ) );
NAND4_X1 _15033_ ( .A1(_06598_ ), .A2(_07040_ ), .A3(_06626_ ), .A4(_06983_ ), .ZN(_07041_ ) );
AOI22_X1 _15034_ ( .A1(_07041_ ), .A2(_06604_ ), .B1(_06600_ ), .B2(_06603_ ), .ZN(_07042_ ) );
OR3_X1 _15035_ ( .A1(_06916_ ), .A2(_06865_ ), .A3(_06919_ ), .ZN(_07043_ ) );
OR3_X1 _15036_ ( .A1(_06872_ ), .A2(_06873_ ), .A3(_06609_ ), .ZN(_07044_ ) );
NAND3_X1 _15037_ ( .A1(_07043_ ), .A2(_07044_ ), .A3(_06763_ ), .ZN(_07045_ ) );
OR3_X1 _15038_ ( .A1(_06862_ ), .A2(_06863_ ), .A3(_06609_ ), .ZN(_07046_ ) );
OR3_X1 _15039_ ( .A1(_06875_ ), .A2(_06634_ ), .A3(_06876_ ), .ZN(_07047_ ) );
NAND3_X1 _15040_ ( .A1(_07046_ ), .A2(_07047_ ), .A3(_06618_ ), .ZN(_07048_ ) );
AND2_X1 _15041_ ( .A1(_07045_ ), .A2(_07048_ ), .ZN(_07049_ ) );
AND3_X1 _15042_ ( .A1(_06868_ ), .A2(_06609_ ), .A3(_06869_ ), .ZN(_07050_ ) );
NOR3_X1 _15043_ ( .A1(_06880_ ), .A2(_06881_ ), .A3(_06609_ ), .ZN(_07051_ ) );
OR3_X1 _15044_ ( .A1(_07050_ ), .A2(_07051_ ), .A3(_06618_ ), .ZN(_07052_ ) );
AND2_X1 _15045_ ( .A1(_06884_ ), .A2(_06781_ ), .ZN(_07053_ ) );
OAI21_X1 _15046_ ( .A(_07052_ ), .B1(_06631_ ), .B2(_07053_ ), .ZN(_07054_ ) );
INV_X1 _15047_ ( .A(_07054_ ), .ZN(_07055_ ) );
MUX2_X1 _15048_ ( .A(_07049_ ), .B(_07055_ ), .S(_06665_ ), .Z(_07056_ ) );
AND2_X1 _15049_ ( .A1(_07056_ ), .A2(_06669_ ), .ZN(_07057_ ) );
OAI21_X1 _15050_ ( .A(_06551_ ), .B1(_07042_ ), .B2(_07057_ ), .ZN(_07058_ ) );
XNOR2_X1 _15051_ ( .A(_07020_ ), .B(_05190_ ), .ZN(_07059_ ) );
BUF_X4 _15052_ ( .A(_06752_ ), .Z(_07060_ ) );
NAND2_X1 _15053_ ( .A1(_07059_ ), .A2(_07060_ ), .ZN(_07061_ ) );
OAI21_X1 _15054_ ( .A(_06656_ ), .B1(_06927_ ), .B2(_06928_ ), .ZN(_07062_ ) );
OAI21_X1 _15055_ ( .A(_06865_ ), .B1(_06857_ ), .B2(_06684_ ), .ZN(_07063_ ) );
NAND2_X1 _15056_ ( .A1(_07062_ ), .A2(_07063_ ), .ZN(_07064_ ) );
BUF_X4 _15057_ ( .A(_06663_ ), .Z(_07065_ ) );
NOR3_X1 _15058_ ( .A1(_07064_ ), .A2(_06770_ ), .A3(_07065_ ), .ZN(_07066_ ) );
OAI21_X1 _15059_ ( .A(_06754_ ), .B1(_07066_ ), .B2(_06818_ ), .ZN(_07067_ ) );
OR3_X1 _15060_ ( .A1(_06909_ ), .A2(_06910_ ), .A3(_06781_ ), .ZN(_07068_ ) );
OR3_X1 _15061_ ( .A1(_06918_ ), .A2(_06777_ ), .A3(_06919_ ), .ZN(_07069_ ) );
BUF_X4 _15062_ ( .A(_06764_ ), .Z(_07070_ ) );
NAND3_X1 _15063_ ( .A1(_07068_ ), .A2(_07069_ ), .A3(_07070_ ), .ZN(_07071_ ) );
OR3_X1 _15064_ ( .A1(_06901_ ), .A2(_06902_ ), .A3(_06609_ ), .ZN(_07072_ ) );
OR3_X1 _15065_ ( .A1(_06912_ ), .A2(_06634_ ), .A3(_06913_ ), .ZN(_07073_ ) );
NAND3_X1 _15066_ ( .A1(_07072_ ), .A2(_07073_ ), .A3(_07065_ ), .ZN(_07074_ ) );
BUF_X4 _15067_ ( .A(_06900_ ), .Z(_07075_ ) );
BUF_X4 _15068_ ( .A(_07075_ ), .Z(_07076_ ) );
NAND3_X1 _15069_ ( .A1(_07071_ ), .A2(_07074_ ), .A3(_07076_ ), .ZN(_07077_ ) );
AND2_X1 _15070_ ( .A1(_07077_ ), .A2(_06818_ ), .ZN(_07078_ ) );
NOR3_X1 _15071_ ( .A1(_06904_ ), .A2(_06865_ ), .A3(_06905_ ), .ZN(_07079_ ) );
NOR3_X1 _15072_ ( .A1(_06892_ ), .A2(_06893_ ), .A3(_06656_ ), .ZN(_07080_ ) );
NOR2_X1 _15073_ ( .A1(_07079_ ), .A2(_07080_ ), .ZN(_07081_ ) );
NAND2_X1 _15074_ ( .A1(_07081_ ), .A2(_06763_ ), .ZN(_07082_ ) );
OAI21_X1 _15075_ ( .A(_06656_ ), .B1(_06895_ ), .B2(_06896_ ), .ZN(_07083_ ) );
OAI21_X1 _15076_ ( .A(_06865_ ), .B1(_06924_ ), .B2(_06925_ ), .ZN(_07084_ ) );
NAND2_X1 _15077_ ( .A1(_07083_ ), .A2(_07084_ ), .ZN(_07085_ ) );
NAND2_X1 _15078_ ( .A1(_07085_ ), .A2(_06618_ ), .ZN(_07086_ ) );
NAND3_X1 _15079_ ( .A1(_07082_ ), .A2(_07000_ ), .A3(_07086_ ), .ZN(_07087_ ) );
AOI21_X1 _15080_ ( .A(_07067_ ), .B1(_07078_ ), .B2(_07087_ ), .ZN(_07088_ ) );
NAND3_X1 _15081_ ( .A1(_07056_ ), .A2(_06669_ ), .A3(_06820_ ), .ZN(_07089_ ) );
OAI21_X1 _15082_ ( .A(_07089_ ), .B1(_06742_ ), .B2(_05129_ ), .ZN(_07090_ ) );
BUF_X2 _15083_ ( .A(_05386_ ), .Z(_07091_ ) );
AND2_X1 _15084_ ( .A1(_05190_ ), .A2(_07091_ ), .ZN(_07092_ ) );
AOI21_X1 _15085_ ( .A(_06815_ ), .B1(_05189_ ), .B2(_05210_ ), .ZN(_07093_ ) );
NOR4_X1 _15086_ ( .A1(_07088_ ), .A2(_07090_ ), .A3(_07092_ ), .A4(_07093_ ), .ZN(_07094_ ) );
NAND3_X1 _15087_ ( .A1(_07058_ ), .A2(_07061_ ), .A3(_07094_ ), .ZN(_07095_ ) );
AOI21_X1 _15088_ ( .A(_07038_ ), .B1(_07095_ ), .B2(_06948_ ), .ZN(_07096_ ) );
NAND2_X1 _15089_ ( .A1(_05554_ ), .A2(_06016_ ), .ZN(_07097_ ) );
NAND2_X1 _15090_ ( .A1(_07097_ ), .A2(_04108_ ), .ZN(_07098_ ) );
OAI21_X1 _15091_ ( .A(_07032_ ), .B1(_07096_ ), .B2(_07098_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_13_D ) );
NAND2_X1 _15092_ ( .A1(_06282_ ), .A2(_06402_ ), .ZN(_07099_ ) );
AND2_X1 _15093_ ( .A1(_05418_ ), .A2(_04754_ ), .ZN(_07100_ ) );
OR2_X1 _15094_ ( .A1(_07100_ ), .A2(_05423_ ), .ZN(_07101_ ) );
AOI21_X1 _15095_ ( .A(_06956_ ), .B1(_07101_ ), .B2(_04732_ ), .ZN(_07102_ ) );
OAI21_X1 _15096_ ( .A(_07102_ ), .B1(_04732_ ), .B2(_07101_ ), .ZN(_07103_ ) );
INV_X1 _15097_ ( .A(_06838_ ), .ZN(_07104_ ) );
NOR2_X1 _15098_ ( .A1(_05573_ ), .A2(_07104_ ), .ZN(_07105_ ) );
AOI21_X1 _15099_ ( .A(_07105_ ), .B1(\ID_EX_imm [17] ), .B2(_06841_ ), .ZN(_07106_ ) );
AOI21_X1 _15100_ ( .A(_06826_ ), .B1(_07103_ ), .B2(_07106_ ), .ZN(_07107_ ) );
OR2_X1 _15101_ ( .A1(_07107_ ), .A2(_05569_ ), .ZN(_07108_ ) );
AND3_X1 _15102_ ( .A1(_06608_ ), .A2(_06626_ ), .A3(_06983_ ), .ZN(_07109_ ) );
NAND2_X1 _15103_ ( .A1(_07109_ ), .A2(_06616_ ), .ZN(_07110_ ) );
AOI22_X1 _15104_ ( .A1(_07110_ ), .A2(_06604_ ), .B1(_06603_ ), .B2(_06600_ ), .ZN(_07111_ ) );
OAI21_X1 _15105_ ( .A(_06618_ ), .B1(_06639_ ), .B2(_06644_ ), .ZN(_07112_ ) );
OAI21_X1 _15106_ ( .A(_06611_ ), .B1(_06807_ ), .B2(_06799_ ), .ZN(_07113_ ) );
OAI21_X1 _15107_ ( .A(_06649_ ), .B1(_06804_ ), .B2(_06808_ ), .ZN(_07114_ ) );
NAND3_X1 _15108_ ( .A1(_07113_ ), .A2(_07114_ ), .A3(_06630_ ), .ZN(_07115_ ) );
AND2_X1 _15109_ ( .A1(_07112_ ), .A2(_07115_ ), .ZN(_07116_ ) );
NAND2_X1 _15110_ ( .A1(_06662_ ), .A2(_06618_ ), .ZN(_07117_ ) );
NAND2_X1 _15111_ ( .A1(_06648_ ), .A2(_06652_ ), .ZN(_07118_ ) );
NAND2_X1 _15112_ ( .A1(_07118_ ), .A2(_06763_ ), .ZN(_07119_ ) );
NAND2_X1 _15113_ ( .A1(_07117_ ), .A2(_07119_ ), .ZN(_07120_ ) );
MUX2_X1 _15114_ ( .A(_07116_ ), .B(_07120_ ), .S(_06769_ ), .Z(_07121_ ) );
NOR2_X1 _15115_ ( .A1(_07121_ ), .A2(_06989_ ), .ZN(_07122_ ) );
OAI21_X1 _15116_ ( .A(_06551_ ), .B1(_07111_ ), .B2(_07122_ ), .ZN(_07123_ ) );
INV_X1 _15117_ ( .A(_05335_ ), .ZN(_07124_ ) );
NOR2_X1 _15118_ ( .A1(_06728_ ), .A2(_07124_ ), .ZN(_07125_ ) );
NOR3_X1 _15119_ ( .A1(_07125_ ), .A2(_05199_ ), .A3(_06736_ ), .ZN(_07126_ ) );
NOR2_X1 _15120_ ( .A1(_07126_ ), .A2(_07024_ ), .ZN(_07127_ ) );
OAI21_X1 _15121_ ( .A(_05199_ ), .B1(_07125_ ), .B2(_06736_ ), .ZN(_07128_ ) );
NAND2_X1 _15122_ ( .A1(_07127_ ), .A2(_07128_ ), .ZN(_07129_ ) );
INV_X2 _15123_ ( .A(_06819_ ), .ZN(_07130_ ) );
NOR3_X1 _15124_ ( .A1(_07121_ ), .A2(_06989_ ), .A3(_07130_ ), .ZN(_07131_ ) );
BUF_X2 _15125_ ( .A(_06900_ ), .Z(_07132_ ) );
BUF_X2 _15126_ ( .A(_06783_ ), .Z(_07133_ ) );
AND3_X1 _15127_ ( .A1(_06767_ ), .A2(_07132_ ), .A3(_07133_ ), .ZN(_07134_ ) );
OAI21_X1 _15128_ ( .A(_06754_ ), .B1(_07134_ ), .B2(_06818_ ), .ZN(_07135_ ) );
NAND3_X1 _15129_ ( .A1(_06798_ ), .A2(_06802_ ), .A3(_07133_ ), .ZN(_07136_ ) );
NAND3_X1 _15130_ ( .A1(_06778_ ), .A2(_06782_ ), .A3(_07065_ ), .ZN(_07137_ ) );
NAND3_X1 _15131_ ( .A1(_07136_ ), .A2(_07137_ ), .A3(_07076_ ), .ZN(_07138_ ) );
AND2_X1 _15132_ ( .A1(_07138_ ), .A2(_06818_ ), .ZN(_07139_ ) );
NAND2_X1 _15133_ ( .A1(_06790_ ), .A2(_06793_ ), .ZN(_07140_ ) );
NAND2_X1 _15134_ ( .A1(_07140_ ), .A2(_06631_ ), .ZN(_07141_ ) );
NAND3_X1 _15135_ ( .A1(_06757_ ), .A2(_06761_ ), .A3(_06663_ ), .ZN(_07142_ ) );
NAND3_X1 _15136_ ( .A1(_07141_ ), .A2(_07142_ ), .A3(_07000_ ), .ZN(_07143_ ) );
AOI21_X1 _15137_ ( .A(_07135_ ), .B1(_07139_ ), .B2(_07143_ ), .ZN(_07144_ ) );
AND2_X1 _15138_ ( .A1(_05198_ ), .A2(_06734_ ), .ZN(_07145_ ) );
NOR3_X1 _15139_ ( .A1(_07145_ ), .A2(_06735_ ), .A3(_05387_ ), .ZN(_07146_ ) );
NAND2_X1 _15140_ ( .A1(_06735_ ), .A2(_07016_ ), .ZN(_07147_ ) );
OAI21_X1 _15141_ ( .A(_07147_ ), .B1(_07145_ ), .B2(_06815_ ), .ZN(_07148_ ) );
NOR4_X1 _15142_ ( .A1(_07131_ ), .A2(_07144_ ), .A3(_07146_ ), .A4(_07148_ ), .ZN(_07149_ ) );
NAND3_X1 _15143_ ( .A1(_07123_ ), .A2(_07129_ ), .A3(_07149_ ), .ZN(_07150_ ) );
AOI21_X1 _15144_ ( .A(_07108_ ), .B1(_07150_ ), .B2(_06948_ ), .ZN(_07151_ ) );
AOI21_X1 _15145_ ( .A(_05485_ ), .B1(_05582_ ), .B2(_05506_ ), .ZN(_07152_ ) );
OR2_X1 _15146_ ( .A1(_07152_ ), .A2(_04113_ ), .ZN(_07153_ ) );
OAI21_X1 _15147_ ( .A(_07099_ ), .B1(_07151_ ), .B2(_07153_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_14_D ) );
NAND2_X1 _15148_ ( .A1(_05618_ ), .A2(_06402_ ), .ZN(_07154_ ) );
AOI21_X1 _15149_ ( .A(_06956_ ), .B1(_05418_ ), .B2(_04754_ ), .ZN(_07155_ ) );
OAI21_X1 _15150_ ( .A(_07155_ ), .B1(_04754_ ), .B2(_05418_ ), .ZN(_07156_ ) );
BUF_X4 _15151_ ( .A(_06840_ ), .Z(_07157_ ) );
AOI22_X1 _15152_ ( .A1(_05623_ ), .A2(_06851_ ), .B1(\ID_EX_imm [16] ), .B2(_07157_ ), .ZN(_07158_ ) );
AOI21_X1 _15153_ ( .A(_06826_ ), .B1(_07156_ ), .B2(_07158_ ), .ZN(_07159_ ) );
OR2_X1 _15154_ ( .A1(_07159_ ), .A2(_05569_ ), .ZN(_07160_ ) );
OAI211_X1 _15155_ ( .A(_06608_ ), .B(_06599_ ), .C1(_06989_ ), .C2(_06555_ ), .ZN(_07161_ ) );
NOR3_X1 _15156_ ( .A1(_06918_ ), .A2(_06865_ ), .A3(_06910_ ), .ZN(_07162_ ) );
NOR3_X1 _15157_ ( .A1(_06916_ ), .A2(_06919_ ), .A3(_06656_ ), .ZN(_07163_ ) );
OAI21_X1 _15158_ ( .A(_06629_ ), .B1(_07162_ ), .B2(_07163_ ), .ZN(_07164_ ) );
NAND3_X1 _15159_ ( .A1(_06874_ ), .A2(_06877_ ), .A3(_06617_ ), .ZN(_07165_ ) );
NAND2_X1 _15160_ ( .A1(_07164_ ), .A2(_07165_ ), .ZN(_07166_ ) );
OAI21_X1 _15161_ ( .A(_05267_ ), .B1(_06866_ ), .B2(_06870_ ), .ZN(_07167_ ) );
OAI21_X1 _15162_ ( .A(_07167_ ), .B1(_06885_ ), .B2(_06629_ ), .ZN(_07168_ ) );
INV_X1 _15163_ ( .A(_07168_ ), .ZN(_07169_ ) );
MUX2_X1 _15164_ ( .A(_07166_ ), .B(_07169_ ), .S(_06623_ ), .Z(_07170_ ) );
NAND2_X1 _15165_ ( .A1(_07170_ ), .A2(_06669_ ), .ZN(_07171_ ) );
AOI21_X1 _15166_ ( .A(_06966_ ), .B1(_07161_ ), .B2(_07171_ ), .ZN(_07172_ ) );
OAI21_X1 _15167_ ( .A(_07060_ ), .B1(_06729_ ), .B2(_05335_ ), .ZN(_07173_ ) );
NOR2_X1 _15168_ ( .A1(_07173_ ), .A2(_07125_ ), .ZN(_07174_ ) );
NAND3_X1 _15169_ ( .A1(_07170_ ), .A2(_06669_ ), .A3(_06986_ ), .ZN(_07175_ ) );
NOR3_X1 _15170_ ( .A1(_06894_ ), .A2(_06897_ ), .A3(_06619_ ), .ZN(_07176_ ) );
AOI21_X1 _15171_ ( .A(_06763_ ), .B1(_06926_ ), .B2(_06929_ ), .ZN(_07177_ ) );
OR3_X1 _15172_ ( .A1(_07176_ ), .A2(_07075_ ), .A3(_07177_ ), .ZN(_07178_ ) );
NAND3_X1 _15173_ ( .A1(_06911_ ), .A2(_06914_ ), .A3(_06631_ ), .ZN(_07179_ ) );
NAND3_X1 _15174_ ( .A1(_06903_ ), .A2(_06906_ ), .A3(_06663_ ), .ZN(_07180_ ) );
NAND3_X1 _15175_ ( .A1(_07179_ ), .A2(_07180_ ), .A3(_06787_ ), .ZN(_07181_ ) );
NAND3_X1 _15176_ ( .A1(_07178_ ), .A2(_06818_ ), .A3(_07181_ ), .ZN(_07182_ ) );
AND2_X1 _15177_ ( .A1(_06615_ ), .A2(_04110_ ), .ZN(_07183_ ) );
AND3_X1 _15178_ ( .A1(_07183_ ), .A2(_06631_ ), .A3(_06801_ ), .ZN(_07184_ ) );
NAND2_X1 _15179_ ( .A1(_07184_ ), .A2(_06787_ ), .ZN(_07185_ ) );
BUF_X2 _15180_ ( .A(_06988_ ), .Z(_07186_ ) );
AOI21_X1 _15181_ ( .A(_06891_ ), .B1(_07185_ ), .B2(_07186_ ), .ZN(_07187_ ) );
NAND2_X1 _15182_ ( .A1(_07182_ ), .A2(_07187_ ), .ZN(_07188_ ) );
NAND3_X1 _15183_ ( .A1(_05204_ ), .A2(_02666_ ), .A3(_07016_ ), .ZN(_07189_ ) );
AOI21_X1 _15184_ ( .A(_06815_ ), .B1(_05203_ ), .B2(_05200_ ), .ZN(_07190_ ) );
AOI21_X1 _15185_ ( .A(_07190_ ), .B1(_05335_ ), .B2(_07091_ ), .ZN(_07191_ ) );
NAND4_X1 _15186_ ( .A1(_07175_ ), .A2(_07188_ ), .A3(_07189_ ), .A4(_07191_ ), .ZN(_07192_ ) );
OR3_X1 _15187_ ( .A1(_07172_ ), .A2(_07174_ ), .A3(_07192_ ), .ZN(_07193_ ) );
AOI21_X1 _15188_ ( .A(_07160_ ), .B1(_07193_ ), .B2(_06948_ ), .ZN(_07194_ ) );
OAI21_X1 _15189_ ( .A(_06409_ ), .B1(_05621_ ), .B2(_05486_ ), .ZN(_07195_ ) );
OAI21_X1 _15190_ ( .A(_07154_ ), .B1(_07194_ ), .B2(_07195_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_15_D ) );
OAI211_X1 _15191_ ( .A(_05657_ ), .B(_06240_ ), .C1(\EX_LS_result_csreg_mem [15] ), .C2(_05646_ ), .ZN(_07196_ ) );
BUF_X4 _15192_ ( .A(_06547_ ), .Z(_07197_ ) );
AND2_X1 _15193_ ( .A1(_02592_ ), .A2(_05004_ ), .ZN(_07198_ ) );
NAND2_X1 _15194_ ( .A1(_05401_ ), .A2(_04983_ ), .ZN(_07199_ ) );
AND2_X1 _15195_ ( .A1(_07199_ ), .A2(_05412_ ), .ZN(_07200_ ) );
INV_X1 _15196_ ( .A(_05051_ ), .ZN(_07201_ ) );
NOR2_X1 _15197_ ( .A1(_07200_ ), .A2(_07201_ ), .ZN(_07202_ ) );
AOI21_X1 _15198_ ( .A(_07202_ ), .B1(_02588_ ), .B2(_05050_ ), .ZN(_07203_ ) );
OAI21_X1 _15199_ ( .A(_05414_ ), .B1(_07203_ ), .B2(_05074_ ), .ZN(_07204_ ) );
AOI21_X1 _15200_ ( .A(_07198_ ), .B1(_07204_ ), .B2(_05005_ ), .ZN(_07205_ ) );
XNOR2_X1 _15201_ ( .A(_07205_ ), .B(_05028_ ), .ZN(_07206_ ) );
NAND2_X1 _15202_ ( .A1(_07206_ ), .A2(_06835_ ), .ZN(_07207_ ) );
AOI22_X1 _15203_ ( .A1(_05637_ ), .A2(_06851_ ), .B1(\ID_EX_imm [15] ), .B2(_07157_ ), .ZN(_07208_ ) );
AOI21_X1 _15204_ ( .A(_07197_ ), .B1(_07207_ ), .B2(_07208_ ), .ZN(_07209_ ) );
OR2_X1 _15205_ ( .A1(_07209_ ), .A2(_05569_ ), .ZN(_07210_ ) );
INV_X1 _15206_ ( .A(_06968_ ), .ZN(_07211_ ) );
AND3_X1 _15207_ ( .A1(_06976_ ), .A2(_06617_ ), .A3(_06977_ ), .ZN(_07212_ ) );
AOI21_X1 _15208_ ( .A(_06617_ ), .B1(_06972_ ), .B2(_06973_ ), .ZN(_07213_ ) );
OR3_X1 _15209_ ( .A1(_07212_ ), .A2(_07075_ ), .A3(_07213_ ), .ZN(_07214_ ) );
OR3_X1 _15210_ ( .A1(_06969_ ), .A2(_06970_ ), .A3(_06783_ ), .ZN(_07215_ ) );
NOR2_X1 _15211_ ( .A1(_06614_ ), .A2(_02666_ ), .ZN(_07216_ ) );
OAI21_X1 _15212_ ( .A(_06610_ ), .B1(_07216_ ), .B2(_06797_ ), .ZN(_07217_ ) );
OAI21_X1 _15213_ ( .A(_06635_ ), .B1(_06807_ ), .B2(_06799_ ), .ZN(_07218_ ) );
NAND2_X1 _15214_ ( .A1(_07217_ ), .A2(_07218_ ), .ZN(_07219_ ) );
NAND2_X1 _15215_ ( .A1(_07219_ ), .A2(_07133_ ), .ZN(_07220_ ) );
NAND3_X1 _15216_ ( .A1(_07215_ ), .A2(_07132_ ), .A3(_07220_ ), .ZN(_07221_ ) );
NAND3_X1 _15217_ ( .A1(_07214_ ), .A2(_06773_ ), .A3(_07221_ ), .ZN(_07222_ ) );
NAND3_X1 _15218_ ( .A1(_06661_ ), .A2(_06783_ ), .A3(_06612_ ), .ZN(_07223_ ) );
OAI21_X1 _15219_ ( .A(_07186_ ), .B1(_07223_ ), .B2(_06770_ ), .ZN(_07224_ ) );
NAND2_X1 _15220_ ( .A1(_07222_ ), .A2(_07224_ ), .ZN(_07225_ ) );
AOI21_X1 _15221_ ( .A(_06966_ ), .B1(_07211_ ), .B2(_07225_ ), .ZN(_07226_ ) );
AND2_X1 _15222_ ( .A1(_06696_ ), .A2(_06706_ ), .ZN(_07227_ ) );
OR2_X1 _15223_ ( .A1(_07227_ ), .A2(_06680_ ), .ZN(_07228_ ) );
AND2_X1 _15224_ ( .A1(_07228_ ), .A2(_06718_ ), .ZN(_07229_ ) );
INV_X1 _15225_ ( .A(_05238_ ), .ZN(_07230_ ) );
OR4_X1 _15226_ ( .A1(_05232_ ), .A2(_07229_ ), .A3(_05233_ ), .A4(_07230_ ), .ZN(_07231_ ) );
AOI21_X1 _15227_ ( .A(_06720_ ), .B1(_07231_ ), .B2(_06722_ ), .ZN(_07232_ ) );
OR3_X1 _15228_ ( .A1(_07232_ ), .A2(_05226_ ), .A3(_06725_ ), .ZN(_07233_ ) );
OAI21_X1 _15229_ ( .A(_05226_ ), .B1(_07232_ ), .B2(_06725_ ), .ZN(_07234_ ) );
AND3_X1 _15230_ ( .A1(_07233_ ), .A2(_06752_ ), .A3(_07234_ ), .ZN(_07235_ ) );
NAND3_X1 _15231_ ( .A1(_07222_ ), .A2(_06986_ ), .A3(_07224_ ), .ZN(_07236_ ) );
NAND2_X1 _15232_ ( .A1(_06993_ ), .A2(_07070_ ), .ZN(_07237_ ) );
NAND2_X1 _15233_ ( .A1(_07002_ ), .A2(_07003_ ), .ZN(_07238_ ) );
NAND2_X1 _15234_ ( .A1(_07238_ ), .A2(_07065_ ), .ZN(_07239_ ) );
NAND2_X1 _15235_ ( .A1(_07237_ ), .A2(_07239_ ), .ZN(_07240_ ) );
NAND2_X1 _15236_ ( .A1(_07240_ ), .A2(_07076_ ), .ZN(_07241_ ) );
NAND2_X1 _15237_ ( .A1(_07005_ ), .A2(_07006_ ), .ZN(_07242_ ) );
NAND2_X1 _15238_ ( .A1(_07242_ ), .A2(_07133_ ), .ZN(_07243_ ) );
NAND3_X1 _15239_ ( .A1(_07010_ ), .A2(_07011_ ), .A3(_07065_ ), .ZN(_07244_ ) );
NAND2_X1 _15240_ ( .A1(_07243_ ), .A2(_07244_ ), .ZN(_07245_ ) );
NAND2_X1 _15241_ ( .A1(_07245_ ), .A2(_07000_ ), .ZN(_07246_ ) );
AND2_X1 _15242_ ( .A1(_06667_ ), .A2(_05465_ ), .ZN(_07247_ ) );
BUF_X4 _15243_ ( .A(_07247_ ), .Z(_07248_ ) );
NAND3_X1 _15244_ ( .A1(_07241_ ), .A2(_07246_ ), .A3(_07248_ ), .ZN(_07249_ ) );
NAND2_X1 _15245_ ( .A1(_06708_ ), .A2(_07017_ ), .ZN(_07250_ ) );
AOI21_X1 _15246_ ( .A(_05383_ ), .B1(_05225_ ), .B2(_05404_ ), .ZN(_07251_ ) );
AOI21_X1 _15247_ ( .A(_07251_ ), .B1(_05226_ ), .B2(_06940_ ), .ZN(_07252_ ) );
NAND4_X1 _15248_ ( .A1(_07236_ ), .A2(_07249_ ), .A3(_07250_ ), .A4(_07252_ ), .ZN(_07253_ ) );
OR3_X1 _15249_ ( .A1(_07226_ ), .A2(_07235_ ), .A3(_07253_ ), .ZN(_07254_ ) );
AOI21_X1 _15250_ ( .A(_07210_ ), .B1(_07254_ ), .B2(_06948_ ), .ZN(_07255_ ) );
NAND2_X1 _15251_ ( .A1(_05642_ ), .A2(_06016_ ), .ZN(_07256_ ) );
NAND2_X1 _15252_ ( .A1(_07256_ ), .A2(_04108_ ), .ZN(_07257_ ) );
OAI21_X1 _15253_ ( .A(_07196_ ), .B1(_07255_ ), .B2(_07257_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_16_D ) );
AND2_X1 _15254_ ( .A1(_05675_ ), .A2(_05676_ ), .ZN(_07258_ ) );
INV_X1 _15255_ ( .A(_07258_ ), .ZN(_07259_ ) );
AND2_X1 _15256_ ( .A1(_05663_ ), .A2(_05880_ ), .ZN(_07260_ ) );
AND2_X1 _15257_ ( .A1(_05222_ ), .A2(_06940_ ), .ZN(_07261_ ) );
AND2_X1 _15258_ ( .A1(_07039_ ), .A2(_06630_ ), .ZN(_07262_ ) );
INV_X1 _15259_ ( .A(_07262_ ), .ZN(_07263_ ) );
OAI211_X1 _15260_ ( .A(_06598_ ), .B(_06967_ ), .C1(_06625_ ), .C2(_07263_ ), .ZN(_07264_ ) );
AND3_X1 _15261_ ( .A1(_07046_ ), .A2(_07047_ ), .A3(_05267_ ), .ZN(_07265_ ) );
NOR3_X1 _15262_ ( .A1(_07050_ ), .A2(_07051_ ), .A3(_05267_ ), .ZN(_07266_ ) );
OR3_X1 _15263_ ( .A1(_07265_ ), .A2(_07266_ ), .A3(_06554_ ), .ZN(_07267_ ) );
OR3_X1 _15264_ ( .A1(_06909_ ), .A2(_06865_ ), .A3(_06913_ ), .ZN(_07268_ ) );
OR3_X1 _15265_ ( .A1(_06918_ ), .A2(_06910_ ), .A3(_06656_ ), .ZN(_07269_ ) );
NAND3_X1 _15266_ ( .A1(_07268_ ), .A2(_07269_ ), .A3(_06629_ ), .ZN(_07270_ ) );
NAND3_X1 _15267_ ( .A1(_07043_ ), .A2(_07044_ ), .A3(_06617_ ), .ZN(_07271_ ) );
NAND3_X1 _15268_ ( .A1(_07270_ ), .A2(_07271_ ), .A3(_06785_ ), .ZN(_07272_ ) );
NAND3_X1 _15269_ ( .A1(_07267_ ), .A2(_06667_ ), .A3(_07272_ ), .ZN(_07273_ ) );
AND3_X1 _15270_ ( .A1(_06884_ ), .A2(_05267_ ), .A3(_06656_ ), .ZN(_07274_ ) );
AND2_X1 _15271_ ( .A1(_07274_ ), .A2(_06554_ ), .ZN(_07275_ ) );
OR2_X1 _15272_ ( .A1(_07275_ ), .A2(_06667_ ), .ZN(_07276_ ) );
NAND2_X1 _15273_ ( .A1(_07273_ ), .A2(_07276_ ), .ZN(_07277_ ) );
AOI21_X1 _15274_ ( .A(_06856_ ), .B1(_07264_ ), .B2(_07277_ ), .ZN(_07278_ ) );
AND3_X1 _15275_ ( .A1(_07273_ ), .A2(_06819_ ), .A3(_07276_ ), .ZN(_07279_ ) );
NOR2_X1 _15276_ ( .A1(_07081_ ), .A2(_06629_ ), .ZN(_07280_ ) );
AOI21_X1 _15277_ ( .A(_06617_ ), .B1(_07073_ ), .B2(_07072_ ), .ZN(_07281_ ) );
OAI21_X1 _15278_ ( .A(_06785_ ), .B1(_07280_ ), .B2(_07281_ ), .ZN(_07282_ ) );
MUX2_X1 _15279_ ( .A(_07064_ ), .B(_07085_ ), .S(_06629_ ), .Z(_07283_ ) );
OAI21_X1 _15280_ ( .A(_07282_ ), .B1(_06785_ ), .B2(_07283_ ), .ZN(_07284_ ) );
AND2_X1 _15281_ ( .A1(_07284_ ), .A2(_07247_ ), .ZN(_07285_ ) );
OR3_X2 _15282_ ( .A1(_07278_ ), .A2(_07279_ ), .A3(_07285_ ), .ZN(_07286_ ) );
AOI21_X1 _15283_ ( .A(_05383_ ), .B1(_05221_ ), .B2(_06724_ ), .ZN(_07287_ ) );
NOR3_X1 _15284_ ( .A1(_05221_ ), .A2(_06724_ ), .A3(_05129_ ), .ZN(_07288_ ) );
OR4_X2 _15285_ ( .A1(_07261_ ), .A2(_07286_ ), .A3(_07287_ ), .A4(_07288_ ), .ZN(_07289_ ) );
AND3_X1 _15286_ ( .A1(_07231_ ), .A2(_06720_ ), .A3(_06722_ ), .ZN(_07290_ ) );
NOR3_X1 _15287_ ( .A1(_07290_ ), .A2(_07232_ ), .A3(_07024_ ), .ZN(_07291_ ) );
OAI21_X1 _15288_ ( .A(_06947_ ), .B1(_07289_ ), .B2(_07291_ ), .ZN(_07292_ ) );
AOI21_X1 _15289_ ( .A(_06955_ ), .B1(_07204_ ), .B2(_05005_ ), .ZN(_07293_ ) );
OAI21_X1 _15290_ ( .A(_07293_ ), .B1(_05005_ ), .B2(_07204_ ), .ZN(_07294_ ) );
AOI22_X1 _15291_ ( .A1(_05660_ ), .A2(_06838_ ), .B1(\ID_EX_imm [14] ), .B2(_07157_ ), .ZN(_07295_ ) );
AOI21_X1 _15292_ ( .A(_07197_ ), .B1(_07294_ ), .B2(_07295_ ), .ZN(_07296_ ) );
NOR2_X1 _15293_ ( .A1(_07296_ ), .A2(_06015_ ), .ZN(_07297_ ) );
AOI21_X1 _15294_ ( .A(_07260_ ), .B1(_07292_ ), .B2(_07297_ ), .ZN(_07298_ ) );
MUX2_X1 _15295_ ( .A(_07259_ ), .B(_07298_ ), .S(_04107_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_17_D ) );
NAND2_X1 _15296_ ( .A1(_06326_ ), .A2(_06402_ ), .ZN(_07299_ ) );
NOR2_X1 _15297_ ( .A1(_06768_ ), .A2(_07075_ ), .ZN(_07300_ ) );
NOR3_X1 _15298_ ( .A1(_06784_ ), .A2(_06665_ ), .A3(_06794_ ), .ZN(_07301_ ) );
OAI21_X1 _15299_ ( .A(_07248_ ), .B1(_07300_ ), .B2(_07301_ ), .ZN(_07302_ ) );
AOI22_X1 _15300_ ( .A1(_05234_ ), .A2(_06940_ ), .B1(_05232_ ), .B2(_07016_ ), .ZN(_07303_ ) );
NAND3_X1 _15301_ ( .A1(_07113_ ), .A2(_07114_ ), .A3(_06619_ ), .ZN(_07304_ ) );
OAI21_X1 _15302_ ( .A(_06781_ ), .B1(_06796_ ), .B2(_06779_ ), .ZN(_07305_ ) );
OAI21_X1 _15303_ ( .A(_06765_ ), .B1(_07216_ ), .B2(_06797_ ), .ZN(_07306_ ) );
NAND2_X1 _15304_ ( .A1(_07305_ ), .A2(_07306_ ), .ZN(_07307_ ) );
OAI211_X1 _15305_ ( .A(_07304_ ), .B(_06786_ ), .C1(_07307_ ), .C2(_06620_ ), .ZN(_07308_ ) );
OAI211_X1 _15306_ ( .A(_07308_ ), .B(_06668_ ), .C1(_06654_ ), .C2(_07132_ ), .ZN(_07309_ ) );
NAND3_X1 _15307_ ( .A1(_06664_ ), .A2(_06988_ ), .A3(_07132_ ), .ZN(_07310_ ) );
AND2_X1 _15308_ ( .A1(_07309_ ), .A2(_07310_ ), .ZN(_07311_ ) );
OAI211_X1 _15309_ ( .A(_07302_ ), .B(_07303_ ), .C1(_07311_ ), .C2(_07130_ ), .ZN(_07312_ ) );
BUF_X2 _15310_ ( .A(_06967_ ), .Z(_07313_ ) );
OAI211_X1 _15311_ ( .A(_06598_ ), .B(_07313_ ), .C1(_06622_ ), .C2(_06626_ ), .ZN(_07314_ ) );
AOI21_X1 _15312_ ( .A(_06966_ ), .B1(_07314_ ), .B2(_07311_ ), .ZN(_07315_ ) );
BUF_X4 _15313_ ( .A(_05382_ ), .Z(_07316_ ) );
AOI211_X1 _15314_ ( .A(_07312_ ), .B(_07315_ ), .C1(_06721_ ), .C2(_07316_ ), .ZN(_07317_ ) );
AOI21_X1 _15315_ ( .A(_07230_ ), .B1(_07228_ ), .B2(_06718_ ), .ZN(_07318_ ) );
OR2_X1 _15316_ ( .A1(_07318_ ), .A2(_06672_ ), .ZN(_07319_ ) );
AOI21_X1 _15317_ ( .A(_07024_ ), .B1(_07319_ ), .B2(_05234_ ), .ZN(_07320_ ) );
OAI21_X1 _15318_ ( .A(_07320_ ), .B1(_05234_ ), .B2(_07319_ ), .ZN(_07321_ ) );
AOI21_X1 _15319_ ( .A(_06549_ ), .B1(_07317_ ), .B2(_07321_ ), .ZN(_07322_ ) );
INV_X1 _15320_ ( .A(_06840_ ), .ZN(_07323_ ) );
OAI22_X1 _15321_ ( .A1(_05683_ ), .A2(_07104_ ), .B1(_02567_ ), .B2(_07323_ ), .ZN(_07324_ ) );
XNOR2_X1 _15322_ ( .A(_07203_ ), .B(_05075_ ), .ZN(_07325_ ) );
AOI21_X1 _15323_ ( .A(_07324_ ), .B1(_07325_ ), .B2(_06835_ ), .ZN(_07326_ ) );
AOI21_X1 _15324_ ( .A(_05482_ ), .B1(_07326_ ), .B2(_03344_ ), .ZN(_07327_ ) );
OAI22_X1 _15325_ ( .A1(_07322_ ), .A2(_07327_ ), .B1(_06845_ ), .B2(_05698_ ), .ZN(_07328_ ) );
OAI21_X1 _15326_ ( .A(_07299_ ), .B1(_07328_ ), .B2(_06387_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_18_D ) );
AND2_X1 _15327_ ( .A1(_05715_ ), .A2(_05716_ ), .ZN(_07329_ ) );
INV_X1 _15328_ ( .A(_07329_ ), .ZN(_07330_ ) );
AND2_X1 _15329_ ( .A1(_05704_ ), .A2(_05880_ ), .ZN(_07331_ ) );
NOR3_X1 _15330_ ( .A1(_06552_ ), .A2(_06623_ ), .A3(_06618_ ), .ZN(_07332_ ) );
INV_X1 _15331_ ( .A(_07332_ ), .ZN(_07333_ ) );
NAND4_X1 _15332_ ( .A1(_06607_ ), .A2(_06601_ ), .A3(_06599_ ), .A4(_07333_ ), .ZN(_07334_ ) );
NOR3_X1 _15333_ ( .A1(_07162_ ), .A2(_07163_ ), .A3(_06629_ ), .ZN(_07335_ ) );
OAI21_X1 _15334_ ( .A(_06610_ ), .B1(_06912_ ), .B2(_06902_ ), .ZN(_07336_ ) );
OAI21_X1 _15335_ ( .A(_06635_ ), .B1(_06909_ ), .B2(_06913_ ), .ZN(_07337_ ) );
AOI21_X1 _15336_ ( .A(_06617_ ), .B1(_07336_ ), .B2(_07337_ ), .ZN(_07338_ ) );
OAI21_X1 _15337_ ( .A(_06785_ ), .B1(_07335_ ), .B2(_07338_ ), .ZN(_07339_ ) );
OAI211_X1 _15338_ ( .A(_06667_ ), .B(_07339_ ), .C1(_06879_ ), .C2(_06785_ ), .ZN(_07340_ ) );
NAND4_X1 _15339_ ( .A1(_06885_ ), .A2(_05306_ ), .A3(_06785_ ), .A4(_06783_ ), .ZN(_07341_ ) );
AND2_X1 _15340_ ( .A1(_07340_ ), .A2(_07341_ ), .ZN(_07342_ ) );
AOI21_X1 _15341_ ( .A(_06856_ ), .B1(_07334_ ), .B2(_07342_ ), .ZN(_07343_ ) );
AOI21_X1 _15342_ ( .A(_07130_ ), .B1(_07340_ ), .B2(_07341_ ), .ZN(_07344_ ) );
INV_X1 _15343_ ( .A(_07247_ ), .ZN(_07345_ ) );
OR2_X1 _15344_ ( .A1(_06932_ ), .A2(_06900_ ), .ZN(_07346_ ) );
OAI21_X1 _15345_ ( .A(_06900_ ), .B1(_06899_ ), .B2(_06907_ ), .ZN(_07347_ ) );
AOI21_X1 _15346_ ( .A(_07345_ ), .B1(_07346_ ), .B2(_07347_ ), .ZN(_07348_ ) );
OR3_X1 _15347_ ( .A1(_07343_ ), .A2(_07344_ ), .A3(_07348_ ), .ZN(_07349_ ) );
OAI21_X1 _15348_ ( .A(_06752_ ), .B1(_07229_ ), .B2(_07230_ ), .ZN(_07350_ ) );
AOI21_X1 _15349_ ( .A(_07350_ ), .B1(_07230_ ), .B2(_07229_ ), .ZN(_07351_ ) );
AOI22_X1 _15350_ ( .A1(_06672_ ), .A2(_07016_ ), .B1(_06674_ ), .B2(_05382_ ), .ZN(_07352_ ) );
OAI21_X1 _15351_ ( .A(_07352_ ), .B1(_07230_ ), .B2(_05387_ ), .ZN(_07353_ ) );
NOR3_X1 _15352_ ( .A1(_07349_ ), .A2(_07351_ ), .A3(_07353_ ), .ZN(_07354_ ) );
OR2_X1 _15353_ ( .A1(_07354_ ), .A2(_06548_ ), .ZN(_07355_ ) );
AOI22_X1 _15354_ ( .A1(_05702_ ), .A2(_06838_ ), .B1(\ID_EX_imm [12] ), .B2(_07157_ ), .ZN(_07356_ ) );
OAI21_X1 _15355_ ( .A(_06834_ ), .B1(_07200_ ), .B2(_07201_ ), .ZN(_07357_ ) );
AND3_X1 _15356_ ( .A1(_07199_ ), .A2(_07201_ ), .A3(_05412_ ), .ZN(_07358_ ) );
OAI21_X1 _15357_ ( .A(_07356_ ), .B1(_07357_ ), .B2(_07358_ ), .ZN(_07359_ ) );
AOI21_X1 _15358_ ( .A(_05678_ ), .B1(_07359_ ), .B2(_06546_ ), .ZN(_07360_ ) );
AOI21_X1 _15359_ ( .A(_07331_ ), .B1(_07355_ ), .B2(_07360_ ), .ZN(_07361_ ) );
MUX2_X1 _15360_ ( .A(_07330_ ), .B(_07361_ ), .S(_04107_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_19_D ) );
NAND2_X1 _15361_ ( .A1(_06347_ ), .A2(_06402_ ), .ZN(_07362_ ) );
OAI211_X1 _15362_ ( .A(_06598_ ), .B(_06602_ ), .C1(_06625_ ), .C2(_07263_ ), .ZN(_07363_ ) );
INV_X1 _15363_ ( .A(_07363_ ), .ZN(_07364_ ) );
AND2_X1 _15364_ ( .A1(_07275_ ), .A2(_06772_ ), .ZN(_07365_ ) );
OR3_X1 _15365_ ( .A1(_07364_ ), .A2(_06968_ ), .A3(_07365_ ), .ZN(_07366_ ) );
NAND2_X1 _15366_ ( .A1(_07366_ ), .A2(_06551_ ), .ZN(_07367_ ) );
AOI211_X1 _15367_ ( .A(_06777_ ), .B(_06880_ ), .C1(_02962_ ), .C2(_06615_ ), .ZN(_07368_ ) );
NOR2_X1 _15368_ ( .A1(_06614_ ), .A2(_02858_ ), .ZN(_07369_ ) );
NOR3_X1 _15369_ ( .A1(_07369_ ), .A2(_06781_ ), .A3(_06881_ ), .ZN(_07370_ ) );
OR3_X1 _15370_ ( .A1(_07368_ ), .A2(_06619_ ), .A3(_07370_ ), .ZN(_07371_ ) );
NOR2_X1 _15371_ ( .A1(_06862_ ), .A2(_06867_ ), .ZN(_07372_ ) );
NOR2_X1 _15372_ ( .A1(_06875_ ), .A2(_06863_ ), .ZN(_07373_ ) );
MUX2_X1 _15373_ ( .A(_07372_ ), .B(_07373_ ), .S(_06765_ ), .Z(_07374_ ) );
OAI211_X1 _15374_ ( .A(_07371_ ), .B(_07075_ ), .C1(_07374_ ), .C2(_07133_ ), .ZN(_07375_ ) );
OAI21_X1 _15375_ ( .A(_06612_ ), .B1(_06872_ ), .B2(_06876_ ), .ZN(_07376_ ) );
OAI21_X1 _15376_ ( .A(_06765_ ), .B1(_06916_ ), .B2(_06873_ ), .ZN(_07377_ ) );
NAND2_X1 _15377_ ( .A1(_07376_ ), .A2(_07377_ ), .ZN(_07378_ ) );
NAND2_X1 _15378_ ( .A1(_07378_ ), .A2(_06764_ ), .ZN(_07379_ ) );
NAND3_X1 _15379_ ( .A1(_07068_ ), .A2(_07069_ ), .A3(_06663_ ), .ZN(_07380_ ) );
NAND3_X1 _15380_ ( .A1(_07379_ ), .A2(_07380_ ), .A3(_06665_ ), .ZN(_07381_ ) );
NAND3_X1 _15381_ ( .A1(_07375_ ), .A2(_06668_ ), .A3(_07381_ ), .ZN(_07382_ ) );
AND2_X1 _15382_ ( .A1(_07382_ ), .A2(_06754_ ), .ZN(_07383_ ) );
OAI21_X1 _15383_ ( .A(_07383_ ), .B1(_06669_ ), .B2(_07284_ ), .ZN(_07384_ ) );
OAI21_X1 _15384_ ( .A(_07316_ ), .B1(_06883_ ), .B2(_05146_ ), .ZN(_07385_ ) );
AND3_X1 _15385_ ( .A1(_07275_ ), .A2(_06667_ ), .A3(_06819_ ), .ZN(_07386_ ) );
INV_X1 _15386_ ( .A(_05146_ ), .ZN(_07387_ ) );
NOR2_X1 _15387_ ( .A1(_07387_ ), .A2(_02962_ ), .ZN(_07388_ ) );
AOI221_X4 _15388_ ( .A(_07386_ ), .B1(_07388_ ), .B2(_05128_ ), .C1(_05147_ ), .C2(_05386_ ), .ZN(_07389_ ) );
AND4_X1 _15389_ ( .A1(_07367_ ), .A2(_07384_ ), .A3(_07385_ ), .A4(_07389_ ), .ZN(_07390_ ) );
NOR2_X1 _15390_ ( .A1(_05345_ ), .A2(_05347_ ), .ZN(_07391_ ) );
AND4_X1 _15391_ ( .A1(_05341_ ), .A2(_07391_ ), .A3(_05361_ ), .A4(_05353_ ), .ZN(_07392_ ) );
AND2_X1 _15392_ ( .A1(_05179_ ), .A2(_05184_ ), .ZN(_07393_ ) );
AND2_X1 _15393_ ( .A1(_05167_ ), .A2(_05174_ ), .ZN(_07394_ ) );
AND2_X1 _15394_ ( .A1(_07393_ ), .A2(_07394_ ), .ZN(_07395_ ) );
AND3_X1 _15395_ ( .A1(_06729_ ), .A2(_06731_ ), .A3(_07395_ ), .ZN(_07396_ ) );
INV_X1 _15396_ ( .A(_07395_ ), .ZN(_07397_ ) );
NOR2_X1 _15397_ ( .A1(_06745_ ), .A2(_07397_ ), .ZN(_07398_ ) );
NAND2_X1 _15398_ ( .A1(_05184_ ), .A2(_06747_ ), .ZN(_07399_ ) );
OAI21_X1 _15399_ ( .A(_07399_ ), .B1(_06204_ ), .B2(_05183_ ), .ZN(_07400_ ) );
AND2_X1 _15400_ ( .A1(_07400_ ), .A2(_07394_ ), .ZN(_07401_ ) );
NOR4_X1 _15401_ ( .A1(_05165_ ), .A2(_05166_ ), .A3(_05168_ ), .A4(_05171_ ), .ZN(_07402_ ) );
NOR4_X1 _15402_ ( .A1(_07398_ ), .A2(_05165_ ), .A3(_07401_ ), .A4(_07402_ ), .ZN(_07403_ ) );
INV_X1 _15403_ ( .A(_07403_ ), .ZN(_07404_ ) );
OAI21_X1 _15404_ ( .A(_07392_ ), .B1(_07396_ ), .B2(_07404_ ), .ZN(_07405_ ) );
NOR2_X1 _15405_ ( .A1(_05443_ ), .A2(_05340_ ), .ZN(_07406_ ) );
AOI21_X1 _15406_ ( .A(_05367_ ), .B1(_05359_ ), .B2(_05353_ ), .ZN(_07407_ ) );
INV_X1 _15407_ ( .A(_05341_ ), .ZN(_07408_ ) );
NOR4_X1 _15408_ ( .A1(_07407_ ), .A2(_07408_ ), .A3(_05345_ ), .A4(_05347_ ), .ZN(_07409_ ) );
AOI211_X1 _15409_ ( .A(_07406_ ), .B(_07409_ ), .C1(_05341_ ), .C2(_05345_ ), .ZN(_07410_ ) );
NAND2_X1 _15410_ ( .A1(_07405_ ), .A2(_07410_ ), .ZN(_07411_ ) );
NAND3_X1 _15411_ ( .A1(_07411_ ), .A2(_05138_ ), .A3(_05376_ ), .ZN(_07412_ ) );
INV_X1 _15412_ ( .A(_05147_ ), .ZN(_07413_ ) );
AND2_X1 _15413_ ( .A1(_05136_ ), .A2(_02909_ ), .ZN(_07414_ ) );
AND2_X1 _15414_ ( .A1(_05141_ ), .A2(_02933_ ), .ZN(_07415_ ) );
AOI21_X1 _15415_ ( .A(_07414_ ), .B1(_05138_ ), .B2(_07415_ ), .ZN(_07416_ ) );
AND3_X1 _15416_ ( .A1(_07412_ ), .A2(_07413_ ), .A3(_07416_ ), .ZN(_07417_ ) );
AOI21_X1 _15417_ ( .A(_07413_ ), .B1(_07412_ ), .B2(_07416_ ), .ZN(_07418_ ) );
OR3_X1 _15418_ ( .A1(_07417_ ), .A2(_07418_ ), .A3(_07024_ ), .ZN(_07419_ ) );
AOI21_X1 _15419_ ( .A(_06549_ ), .B1(_07390_ ), .B2(_07419_ ), .ZN(_07420_ ) );
AOI22_X1 _15420_ ( .A1(_06162_ ), .A2(_06839_ ), .B1(\ID_EX_imm [30] ), .B2(_06841_ ), .ZN(_07421_ ) );
OAI211_X1 _15421_ ( .A(_04511_ ), .B(_04558_ ), .C1(_05419_ ), .C2(_05440_ ), .ZN(_07422_ ) );
NAND2_X1 _15422_ ( .A1(_07422_ ), .A2(_05450_ ), .ZN(_07423_ ) );
NAND2_X1 _15423_ ( .A1(_07423_ ), .A2(_04410_ ), .ZN(_07424_ ) );
NAND3_X1 _15424_ ( .A1(_07424_ ), .A2(_05456_ ), .A3(_05454_ ), .ZN(_07425_ ) );
AOI21_X1 _15425_ ( .A(_06955_ ), .B1(_07425_ ), .B2(_04455_ ), .ZN(_07426_ ) );
OAI21_X1 _15426_ ( .A(_07426_ ), .B1(_04455_ ), .B2(_07425_ ), .ZN(_07427_ ) );
AOI21_X1 _15427_ ( .A(_06826_ ), .B1(_07421_ ), .B2(_07427_ ), .ZN(_07428_ ) );
OR2_X1 _15428_ ( .A1(_07428_ ), .A2(_05569_ ), .ZN(_07429_ ) );
OAI22_X1 _15429_ ( .A1(_07420_ ), .A2(_07429_ ), .B1(_06845_ ), .B2(_06157_ ), .ZN(_07430_ ) );
OAI21_X1 _15430_ ( .A(_07362_ ), .B1(_07430_ ), .B2(_06387_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_1_D ) );
NAND2_X1 _15431_ ( .A1(_05724_ ), .A2(_06838_ ), .ZN(_07431_ ) );
OAI21_X1 _15432_ ( .A(_07431_ ), .B1(_02576_ ), .B2(_07323_ ), .ZN(_07432_ ) );
NAND3_X1 _15433_ ( .A1(_05401_ ), .A2(_04960_ ), .A3(_04982_ ), .ZN(_07433_ ) );
NAND3_X1 _15434_ ( .A1(_07433_ ), .A2(_05410_ ), .A3(_05409_ ), .ZN(_07434_ ) );
AND2_X1 _15435_ ( .A1(_07434_ ), .A2(_04913_ ), .ZN(_07435_ ) );
AOI21_X1 _15436_ ( .A(_07435_ ), .B1(_02422_ ), .B2(_04912_ ), .ZN(_07436_ ) );
XNOR2_X1 _15437_ ( .A(_07436_ ), .B(_04936_ ), .ZN(_07437_ ) );
AOI21_X1 _15438_ ( .A(_07432_ ), .B1(_07437_ ), .B2(_06835_ ), .ZN(_07438_ ) );
OAI211_X1 _15439_ ( .A(_06608_ ), .B(_06967_ ), .C1(_06625_ ), .C2(_06983_ ), .ZN(_07439_ ) );
OAI211_X1 _15440_ ( .A(_06780_ ), .B(_06635_ ), .C1(_02592_ ), .C2(_06614_ ), .ZN(_07440_ ) );
OAI211_X1 _15441_ ( .A(_06776_ ), .B(_06656_ ), .C1(_02588_ ), .C2(_06614_ ), .ZN(_07441_ ) );
AND3_X1 _15442_ ( .A1(_07440_ ), .A2(_07441_ ), .A3(_06629_ ), .ZN(_07442_ ) );
AOI21_X1 _15443_ ( .A(_06629_ ), .B1(_07217_ ), .B2(_07218_ ), .ZN(_07443_ ) );
OAI21_X1 _15444_ ( .A(_06900_ ), .B1(_07442_ ), .B2(_07443_ ), .ZN(_07444_ ) );
OAI211_X1 _15445_ ( .A(_07444_ ), .B(_06772_ ), .C1(_06975_ ), .C2(_06786_ ), .ZN(_07445_ ) );
OAI211_X1 _15446_ ( .A(_06988_ ), .B(_06786_ ), .C1(_06978_ ), .C2(_06979_ ), .ZN(_07446_ ) );
AND2_X1 _15447_ ( .A1(_07445_ ), .A2(_07446_ ), .ZN(_07447_ ) );
AOI21_X1 _15448_ ( .A(_06966_ ), .B1(_07439_ ), .B2(_07447_ ), .ZN(_07448_ ) );
AOI21_X1 _15449_ ( .A(_07130_ ), .B1(_07445_ ), .B2(_07446_ ), .ZN(_07449_ ) );
NOR3_X1 _15450_ ( .A1(_07004_ ), .A2(_07007_ ), .A3(_06769_ ), .ZN(_07450_ ) );
AOI211_X1 _15451_ ( .A(_06900_ ), .B(_06663_ ), .C1(_07010_ ), .C2(_07011_ ), .ZN(_07451_ ) );
NOR2_X1 _15452_ ( .A1(_07450_ ), .A2(_07451_ ), .ZN(_07452_ ) );
NOR2_X1 _15453_ ( .A1(_07452_ ), .A2(_07345_ ), .ZN(_07453_ ) );
NOR3_X1 _15454_ ( .A1(_07448_ ), .A2(_07449_ ), .A3(_07453_ ), .ZN(_07454_ ) );
AOI211_X1 _15455_ ( .A(_05253_ ), .B(_05258_ ), .C1(_06696_ ), .C2(_06706_ ), .ZN(_07455_ ) );
OR2_X1 _15456_ ( .A1(_07455_ ), .A2(_06713_ ), .ZN(_07456_ ) );
NAND3_X1 _15457_ ( .A1(_02574_ ), .A2(_05241_ ), .A3(_05240_ ), .ZN(_07457_ ) );
AOI21_X1 _15458_ ( .A(_06716_ ), .B1(_07456_ ), .B2(_07457_ ), .ZN(_07458_ ) );
XNOR2_X1 _15459_ ( .A(_07458_ ), .B(_05247_ ), .ZN(_07459_ ) );
NAND2_X1 _15460_ ( .A1(_07459_ ), .A2(_07060_ ), .ZN(_07460_ ) );
NAND2_X1 _15461_ ( .A1(_05247_ ), .A2(_06940_ ), .ZN(_07461_ ) );
AOI21_X1 _15462_ ( .A(_05383_ ), .B1(_05246_ ), .B2(_02577_ ), .ZN(_07462_ ) );
AOI21_X1 _15463_ ( .A(_07462_ ), .B1(_06715_ ), .B2(_07016_ ), .ZN(_07463_ ) );
AND2_X1 _15464_ ( .A1(_07461_ ), .A2(_07463_ ), .ZN(_07464_ ) );
AND3_X1 _15465_ ( .A1(_07454_ ), .A2(_07460_ ), .A3(_07464_ ), .ZN(_07465_ ) );
OAI221_X1 _15466_ ( .A(_05500_ ), .B1(_06826_ ), .B2(_07438_ ), .C1(_07465_ ), .C2(_06549_ ), .ZN(_07466_ ) );
NAND2_X1 _15467_ ( .A1(_05729_ ), .A2(_05551_ ), .ZN(_07467_ ) );
NAND3_X1 _15468_ ( .A1(_07466_ ), .A2(_06409_ ), .A3(_07467_ ), .ZN(_07468_ ) );
AND2_X1 _15469_ ( .A1(_05738_ ), .A2(_05739_ ), .ZN(_07469_ ) );
OAI21_X1 _15470_ ( .A(_07468_ ), .B1(_04108_ ), .B2(_07469_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_20_D ) );
NAND3_X1 _15471_ ( .A1(_06359_ ), .A2(_06952_ ), .A3(_06360_ ), .ZN(_07470_ ) );
AOI21_X1 _15472_ ( .A(_06956_ ), .B1(_07434_ ), .B2(_04913_ ), .ZN(_07471_ ) );
OAI21_X1 _15473_ ( .A(_07471_ ), .B1(_04913_ ), .B2(_07434_ ), .ZN(_07472_ ) );
AOI22_X1 _15474_ ( .A1(_05801_ ), .A2(_06851_ ), .B1(\ID_EX_imm [10] ), .B2(_07157_ ), .ZN(_07473_ ) );
AOI21_X1 _15475_ ( .A(_07197_ ), .B1(_07472_ ), .B2(_07473_ ), .ZN(_07474_ ) );
OR2_X1 _15476_ ( .A1(_07474_ ), .A2(_06015_ ), .ZN(_07475_ ) );
AND3_X1 _15477_ ( .A1(_06607_ ), .A2(_07040_ ), .A3(_06983_ ), .ZN(_07476_ ) );
AND2_X1 _15478_ ( .A1(_06607_ ), .A2(_06625_ ), .ZN(_07477_ ) );
OAI21_X1 _15479_ ( .A(_07313_ ), .B1(_07476_ ), .B2(_07477_ ), .ZN(_07478_ ) );
OR2_X1 _15480_ ( .A1(_07049_ ), .A2(_06786_ ), .ZN(_07479_ ) );
AOI21_X1 _15481_ ( .A(_06631_ ), .B1(_07268_ ), .B2(_07269_ ), .ZN(_07480_ ) );
OR3_X1 _15482_ ( .A1(_06901_ ), .A2(_06649_ ), .A3(_06905_ ), .ZN(_07481_ ) );
OR3_X1 _15483_ ( .A1(_06912_ ), .A2(_06902_ ), .A3(_06611_ ), .ZN(_07482_ ) );
AOI21_X1 _15484_ ( .A(_06619_ ), .B1(_07481_ ), .B2(_07482_ ), .ZN(_07483_ ) );
OR2_X1 _15485_ ( .A1(_07480_ ), .A2(_07483_ ), .ZN(_07484_ ) );
OAI211_X1 _15486_ ( .A(_07479_ ), .B(_06888_ ), .C1(_06770_ ), .C2(_07484_ ), .ZN(_07485_ ) );
NAND3_X1 _15487_ ( .A1(_07055_ ), .A2(_07186_ ), .A3(_06787_ ), .ZN(_07486_ ) );
AND2_X1 _15488_ ( .A1(_07485_ ), .A2(_07486_ ), .ZN(_07487_ ) );
AOI21_X1 _15489_ ( .A(_06966_ ), .B1(_07478_ ), .B2(_07487_ ), .ZN(_07488_ ) );
XNOR2_X1 _15490_ ( .A(_07456_ ), .B(_05243_ ), .ZN(_07489_ ) );
NOR2_X1 _15491_ ( .A1(_07489_ ), .A2(_07024_ ), .ZN(_07490_ ) );
NAND2_X1 _15492_ ( .A1(_07457_ ), .A2(_07316_ ), .ZN(_07491_ ) );
NAND3_X1 _15493_ ( .A1(_07082_ ), .A2(_06900_ ), .A3(_07086_ ), .ZN(_07492_ ) );
NAND4_X1 _15494_ ( .A1(_07062_ ), .A2(_07063_ ), .A3(_06623_ ), .A4(_06763_ ), .ZN(_07493_ ) );
AOI21_X1 _15495_ ( .A(_07345_ ), .B1(_07492_ ), .B2(_07493_ ), .ZN(_07494_ ) );
AOI221_X4 _15496_ ( .A(_07494_ ), .B1(_06716_ ), .B2(_05128_ ), .C1(_05243_ ), .C2(_05386_ ), .ZN(_07495_ ) );
OAI211_X1 _15497_ ( .A(_07491_ ), .B(_07495_ ), .C1(_07487_ ), .C2(_07130_ ), .ZN(_07496_ ) );
OR3_X1 _15498_ ( .A1(_07488_ ), .A2(_07490_ ), .A3(_07496_ ), .ZN(_07497_ ) );
AOI21_X1 _15499_ ( .A(_07475_ ), .B1(_07497_ ), .B2(_06948_ ), .ZN(_07498_ ) );
OAI21_X1 _15500_ ( .A(_04135_ ), .B1(_05804_ ), .B2(_06845_ ), .ZN(_07499_ ) );
OAI21_X1 _15501_ ( .A(_07470_ ), .B1(_07498_ ), .B2(_07499_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_21_D ) );
NAND3_X1 _15502_ ( .A1(_05830_ ), .A2(_06952_ ), .A3(_05832_ ), .ZN(_07500_ ) );
INV_X1 _15503_ ( .A(_04982_ ), .ZN(_07501_ ) );
AOI21_X1 _15504_ ( .A(_07501_ ), .B1(_05394_ ), .B2(_05399_ ), .ZN(_07502_ ) );
OR3_X1 _15505_ ( .A1(_07502_ ), .A2(_04960_ ), .A3(_05408_ ), .ZN(_07503_ ) );
OAI21_X1 _15506_ ( .A(_04960_ ), .B1(_07502_ ), .B2(_05408_ ), .ZN(_07504_ ) );
NAND3_X1 _15507_ ( .A1(_07503_ ), .A2(_06835_ ), .A3(_07504_ ), .ZN(_07505_ ) );
AOI22_X1 _15508_ ( .A1(_05822_ ), .A2(_06851_ ), .B1(\ID_EX_imm [9] ), .B2(_07157_ ), .ZN(_07506_ ) );
AOI21_X1 _15509_ ( .A(_07197_ ), .B1(_07505_ ), .B2(_07506_ ), .ZN(_07507_ ) );
OR2_X1 _15510_ ( .A1(_07507_ ), .A2(_06015_ ), .ZN(_07508_ ) );
INV_X1 _15511_ ( .A(_07313_ ), .ZN(_07509_ ) );
AND3_X1 _15512_ ( .A1(_06607_ ), .A2(_06616_ ), .A3(_06983_ ), .ZN(_07510_ ) );
INV_X1 _15513_ ( .A(_07510_ ), .ZN(_07511_ ) );
INV_X1 _15514_ ( .A(_07477_ ), .ZN(_07512_ ) );
AOI21_X1 _15515_ ( .A(_07509_ ), .B1(_07511_ ), .B2(_07512_ ), .ZN(_07513_ ) );
OAI21_X1 _15516_ ( .A(_06988_ ), .B1(_07120_ ), .B2(_06995_ ), .ZN(_07514_ ) );
NAND3_X1 _15517_ ( .A1(_07305_ ), .A2(_07306_ ), .A3(_06619_ ), .ZN(_07515_ ) );
OAI21_X1 _15518_ ( .A(_06781_ ), .B1(_07001_ ), .B2(_06789_ ), .ZN(_07516_ ) );
OAI21_X1 _15519_ ( .A(_06777_ ), .B1(_06991_ ), .B2(_06775_ ), .ZN(_07517_ ) );
NAND3_X1 _15520_ ( .A1(_07516_ ), .A2(_07517_ ), .A3(_06783_ ), .ZN(_07518_ ) );
NAND2_X1 _15521_ ( .A1(_07515_ ), .A2(_07518_ ), .ZN(_07519_ ) );
NAND2_X1 _15522_ ( .A1(_07519_ ), .A2(_07075_ ), .ZN(_07520_ ) );
OAI211_X1 _15523_ ( .A(_07520_ ), .B(_06668_ ), .C1(_07116_ ), .C2(_07075_ ), .ZN(_07521_ ) );
AND2_X1 _15524_ ( .A1(_07514_ ), .A2(_07521_ ), .ZN(_07522_ ) );
OAI21_X1 _15525_ ( .A(_06550_ ), .B1(_07513_ ), .B2(_07522_ ), .ZN(_07523_ ) );
NAND3_X1 _15526_ ( .A1(_07514_ ), .A2(_07521_ ), .A3(_06986_ ), .ZN(_07524_ ) );
NAND3_X1 _15527_ ( .A1(_07141_ ), .A2(_07142_ ), .A3(_06786_ ), .ZN(_07525_ ) );
NAND3_X1 _15528_ ( .A1(_06767_ ), .A2(_06665_ ), .A3(_07133_ ), .ZN(_07526_ ) );
NAND2_X1 _15529_ ( .A1(_07525_ ), .A2(_07526_ ), .ZN(_07527_ ) );
NAND2_X1 _15530_ ( .A1(_07527_ ), .A2(_07248_ ), .ZN(_07528_ ) );
NAND3_X1 _15531_ ( .A1(_07523_ ), .A2(_07524_ ), .A3(_07528_ ), .ZN(_07529_ ) );
OR2_X1 _15532_ ( .A1(_07227_ ), .A2(_05258_ ), .ZN(_07530_ ) );
INV_X1 _15533_ ( .A(_06711_ ), .ZN(_07531_ ) );
AND3_X1 _15534_ ( .A1(_07530_ ), .A2(_05253_ ), .A3(_07531_ ), .ZN(_07532_ ) );
AOI21_X1 _15535_ ( .A(_05253_ ), .B1(_07530_ ), .B2(_07531_ ), .ZN(_07533_ ) );
NOR3_X1 _15536_ ( .A1(_07532_ ), .A2(_07533_ ), .A3(_07024_ ), .ZN(_07534_ ) );
AOI22_X1 _15537_ ( .A1(_06709_ ), .A2(_07017_ ), .B1(_06710_ ), .B2(_05382_ ), .ZN(_07535_ ) );
OAI21_X1 _15538_ ( .A(_07535_ ), .B1(_05253_ ), .B2(_05387_ ), .ZN(_07536_ ) );
OR3_X1 _15539_ ( .A1(_07529_ ), .A2(_07534_ ), .A3(_07536_ ), .ZN(_07537_ ) );
AOI21_X1 _15540_ ( .A(_07508_ ), .B1(_07537_ ), .B2(_06948_ ), .ZN(_07538_ ) );
OAI21_X1 _15541_ ( .A(_04135_ ), .B1(_05821_ ), .B2(_06845_ ), .ZN(_07539_ ) );
OAI21_X1 _15542_ ( .A(_07500_ ), .B1(_07538_ ), .B2(_07539_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_22_D ) );
NAND2_X1 _15543_ ( .A1(_05853_ ), .A2(_06402_ ), .ZN(_07540_ ) );
OAI22_X1 _15544_ ( .A1(_05836_ ), .A2(_07104_ ), .B1(_02449_ ), .B2(_07323_ ), .ZN(_07541_ ) );
NOR2_X1 _15545_ ( .A1(_07502_ ), .A2(_06956_ ), .ZN(_07542_ ) );
NAND3_X1 _15546_ ( .A1(_05394_ ), .A2(_07501_ ), .A3(_05399_ ), .ZN(_07543_ ) );
AOI21_X1 _15547_ ( .A(_07541_ ), .B1(_07542_ ), .B2(_07543_ ), .ZN(_07544_ ) );
AOI21_X1 _15548_ ( .A(_05482_ ), .B1(_07544_ ), .B2(_03344_ ), .ZN(_07545_ ) );
NAND3_X1 _15549_ ( .A1(_07169_ ), .A2(_06988_ ), .A3(_07132_ ), .ZN(_07546_ ) );
NOR3_X1 _15550_ ( .A1(_06904_ ), .A2(_06635_ ), .A3(_06893_ ), .ZN(_07547_ ) );
NOR3_X1 _15551_ ( .A1(_06901_ ), .A2(_06905_ ), .A3(_06610_ ), .ZN(_07548_ ) );
NOR3_X1 _15552_ ( .A1(_07547_ ), .A2(_07548_ ), .A3(_06618_ ), .ZN(_07549_ ) );
AOI21_X1 _15553_ ( .A(_06630_ ), .B1(_07336_ ), .B2(_07337_ ), .ZN(_07550_ ) );
OAI21_X1 _15554_ ( .A(_06786_ ), .B1(_07549_ ), .B2(_07550_ ), .ZN(_07551_ ) );
OAI211_X1 _15555_ ( .A(_07551_ ), .B(_06668_ ), .C1(_07132_ ), .C2(_07166_ ), .ZN(_07552_ ) );
AOI21_X1 _15556_ ( .A(_07130_ ), .B1(_07546_ ), .B2(_07552_ ), .ZN(_07553_ ) );
OR3_X1 _15557_ ( .A1(_07176_ ), .A2(_06769_ ), .A3(_07177_ ), .ZN(_07554_ ) );
NAND4_X1 _15558_ ( .A1(_07183_ ), .A2(_06665_ ), .A3(_07133_ ), .A4(_06801_ ), .ZN(_07555_ ) );
NAND2_X1 _15559_ ( .A1(_07554_ ), .A2(_07555_ ), .ZN(_07556_ ) );
NOR2_X1 _15560_ ( .A1(_06553_ ), .A2(_06623_ ), .ZN(_07557_ ) );
OAI211_X1 _15561_ ( .A(_07552_ ), .B(_07546_ ), .C1(_07211_ ), .C2(_07557_ ), .ZN(_07558_ ) );
AOI221_X4 _15562_ ( .A(_07553_ ), .B1(_07248_ ), .B2(_07556_ ), .C1(_07558_ ), .C2(_06550_ ), .ZN(_07559_ ) );
NAND3_X1 _15563_ ( .A1(_06696_ ), .A2(_05258_ ), .A3(_06706_ ), .ZN(_07560_ ) );
NAND3_X1 _15564_ ( .A1(_07530_ ), .A2(_07060_ ), .A3(_07560_ ), .ZN(_07561_ ) );
NAND2_X1 _15565_ ( .A1(_05257_ ), .A2(_07091_ ), .ZN(_07562_ ) );
NAND3_X1 _15566_ ( .A1(_05324_ ), .A2(_02448_ ), .A3(_07017_ ), .ZN(_07563_ ) );
OAI21_X1 _15567_ ( .A(_07316_ ), .B1(_05324_ ), .B2(_02448_ ), .ZN(_07564_ ) );
AND3_X1 _15568_ ( .A1(_07562_ ), .A2(_07563_ ), .A3(_07564_ ), .ZN(_07565_ ) );
NAND3_X1 _15569_ ( .A1(_07559_ ), .A2(_07561_ ), .A3(_07565_ ), .ZN(_07566_ ) );
AOI21_X1 _15570_ ( .A(_07545_ ), .B1(_07566_ ), .B2(_06948_ ), .ZN(_07567_ ) );
OAI21_X1 _15571_ ( .A(_04135_ ), .B1(_05840_ ), .B2(_06845_ ), .ZN(_07568_ ) );
OAI21_X1 _15572_ ( .A(_07540_ ), .B1(_07567_ ), .B2(_07568_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_23_D ) );
NAND3_X1 _15573_ ( .A1(_05866_ ), .A2(_06952_ ), .A3(_05867_ ), .ZN(_07569_ ) );
NAND3_X1 _15574_ ( .A1(_06541_ ), .A2(\ID_EX_imm [7] ), .A3(_06539_ ), .ZN(_07570_ ) );
OAI21_X1 _15575_ ( .A(_07570_ ), .B1(_05857_ ), .B2(_07104_ ), .ZN(_07571_ ) );
NOR2_X1 _15576_ ( .A1(_05392_ ), .A2(_05393_ ), .ZN(_07572_ ) );
INV_X1 _15577_ ( .A(_07572_ ), .ZN(_07573_ ) );
AND3_X1 _15578_ ( .A1(_07573_ ), .A2(_04823_ ), .A3(_04844_ ), .ZN(_07574_ ) );
NOR2_X1 _15579_ ( .A1(_07574_ ), .A2(_05398_ ), .ZN(_07575_ ) );
OR2_X1 _15580_ ( .A1(_07575_ ), .A2(_04779_ ), .ZN(_07576_ ) );
AOI21_X1 _15581_ ( .A(_04801_ ), .B1(_07576_ ), .B2(_05395_ ), .ZN(_07577_ ) );
NOR2_X1 _15582_ ( .A1(_07577_ ), .A2(_06956_ ), .ZN(_07578_ ) );
NAND3_X1 _15583_ ( .A1(_07576_ ), .A2(_04801_ ), .A3(_05395_ ), .ZN(_07579_ ) );
AOI21_X1 _15584_ ( .A(_07571_ ), .B1(_07578_ ), .B2(_07579_ ), .ZN(_07580_ ) );
AOI21_X1 _15585_ ( .A(_05482_ ), .B1(_07580_ ), .B2(_03344_ ), .ZN(_07581_ ) );
AND4_X1 _15586_ ( .A1(_06626_ ), .A2(_06590_ ), .A3(_06597_ ), .A4(_07313_ ), .ZN(_07582_ ) );
AOI21_X1 _15587_ ( .A(_06764_ ), .B1(_07440_ ), .B2(_07441_ ), .ZN(_07583_ ) );
OR3_X1 _15588_ ( .A1(_06788_ ), .A2(_06865_ ), .A3(_06792_ ), .ZN(_07584_ ) );
OR3_X1 _15589_ ( .A1(_07001_ ), .A2(_06789_ ), .A3(_06609_ ), .ZN(_07585_ ) );
NAND2_X1 _15590_ ( .A1(_07584_ ), .A2(_07585_ ), .ZN(_07586_ ) );
AOI211_X1 _15591_ ( .A(_06995_ ), .B(_07583_ ), .C1(_07070_ ), .C2(_07586_ ), .ZN(_07587_ ) );
AOI21_X1 _15592_ ( .A(_07132_ ), .B1(_07215_ ), .B2(_07220_ ), .ZN(_07588_ ) );
OR3_X1 _15593_ ( .A1(_07587_ ), .A2(_07186_ ), .A3(_07588_ ), .ZN(_07589_ ) );
OR3_X1 _15594_ ( .A1(_07212_ ), .A2(_06623_ ), .A3(_07213_ ), .ZN(_07590_ ) );
OAI21_X1 _15595_ ( .A(_07590_ ), .B1(_06900_ ), .B2(_07223_ ), .ZN(_07591_ ) );
NAND2_X1 _15596_ ( .A1(_07591_ ), .A2(_06989_ ), .ZN(_07592_ ) );
NAND2_X1 _15597_ ( .A1(_07589_ ), .A2(_07592_ ), .ZN(_07593_ ) );
OAI21_X1 _15598_ ( .A(_06551_ ), .B1(_07582_ ), .B2(_07593_ ), .ZN(_07594_ ) );
OAI21_X1 _15599_ ( .A(_07316_ ), .B1(_05311_ ), .B2(_02345_ ), .ZN(_07595_ ) );
NAND2_X1 _15600_ ( .A1(_05296_ ), .A2(_06940_ ), .ZN(_07596_ ) );
NAND3_X1 _15601_ ( .A1(_05311_ ), .A2(_02345_ ), .A3(_07016_ ), .ZN(_07597_ ) );
NAND3_X1 _15602_ ( .A1(_07243_ ), .A2(_07244_ ), .A3(_07076_ ), .ZN(_07598_ ) );
OAI211_X1 _15603_ ( .A(_07596_ ), .B(_07597_ ), .C1(_07598_ ), .C2(_07345_ ), .ZN(_07599_ ) );
AND3_X1 _15604_ ( .A1(_06692_ ), .A2(_06694_ ), .A3(_05288_ ), .ZN(_07600_ ) );
NOR2_X1 _15605_ ( .A1(_07600_ ), .A2(_06699_ ), .ZN(_07601_ ) );
INV_X1 _15606_ ( .A(_05292_ ), .ZN(_07602_ ) );
NOR2_X1 _15607_ ( .A1(_07601_ ), .A2(_07602_ ), .ZN(_07603_ ) );
OAI21_X1 _15608_ ( .A(_05300_ ), .B1(_07603_ ), .B2(_06697_ ), .ZN(_07604_ ) );
NAND2_X1 _15609_ ( .A1(_07604_ ), .A2(_06703_ ), .ZN(_07605_ ) );
OAI21_X1 _15610_ ( .A(_06752_ ), .B1(_07605_ ), .B2(_05296_ ), .ZN(_07606_ ) );
AOI21_X1 _15611_ ( .A(_07606_ ), .B1(_05296_ ), .B2(_07605_ ), .ZN(_07607_ ) );
AOI211_X1 _15612_ ( .A(_07599_ ), .B(_07607_ ), .C1(_06986_ ), .C2(_07593_ ), .ZN(_07608_ ) );
NAND3_X1 _15613_ ( .A1(_07594_ ), .A2(_07595_ ), .A3(_07608_ ), .ZN(_07609_ ) );
AOI21_X1 _15614_ ( .A(_07581_ ), .B1(_07609_ ), .B2(_06948_ ), .ZN(_07610_ ) );
NAND2_X1 _15615_ ( .A1(_05871_ ), .A2(_06016_ ), .ZN(_07611_ ) );
NAND2_X1 _15616_ ( .A1(_07611_ ), .A2(_06409_ ), .ZN(_07612_ ) );
OAI21_X1 _15617_ ( .A(_07569_ ), .B1(_07610_ ), .B2(_07612_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _15618_ ( .A1(_05888_ ), .A2(_06402_ ), .ZN(_07613_ ) );
NAND2_X1 _15619_ ( .A1(_07575_ ), .A2(_04779_ ), .ZN(_07614_ ) );
NAND3_X1 _15620_ ( .A1(_07576_ ), .A2(_06835_ ), .A3(_07614_ ), .ZN(_07615_ ) );
AOI22_X1 _15621_ ( .A1(_05875_ ), .A2(_06851_ ), .B1(\ID_EX_imm [6] ), .B2(_07157_ ), .ZN(_07616_ ) );
AOI21_X1 _15622_ ( .A(_07197_ ), .B1(_07615_ ), .B2(_07616_ ), .ZN(_07617_ ) );
OR2_X1 _15623_ ( .A1(_07617_ ), .A2(_06015_ ), .ZN(_07618_ ) );
NAND4_X1 _15624_ ( .A1(_06608_ ), .A2(_06626_ ), .A3(_07313_ ), .A4(_07263_ ), .ZN(_07619_ ) );
AOI21_X1 _15625_ ( .A(_06764_ ), .B1(_07481_ ), .B2(_07482_ ), .ZN(_07620_ ) );
NOR3_X1 _15626_ ( .A1(_06904_ ), .A2(_06893_ ), .A3(_06801_ ), .ZN(_07621_ ) );
NOR3_X1 _15627_ ( .A1(_06892_ ), .A2(_06806_ ), .A3(_06896_ ), .ZN(_07622_ ) );
NOR2_X1 _15628_ ( .A1(_07621_ ), .A2(_07622_ ), .ZN(_07623_ ) );
INV_X1 _15629_ ( .A(_07623_ ), .ZN(_07624_ ) );
AOI211_X1 _15630_ ( .A(_06995_ ), .B(_07620_ ), .C1(_07624_ ), .C2(_07070_ ), .ZN(_07625_ ) );
AOI21_X1 _15631_ ( .A(_06787_ ), .B1(_07270_ ), .B2(_07271_ ), .ZN(_07626_ ) );
OAI21_X1 _15632_ ( .A(_06818_ ), .B1(_07625_ ), .B2(_07626_ ), .ZN(_07627_ ) );
OR3_X1 _15633_ ( .A1(_07265_ ), .A2(_07266_ ), .A3(_06769_ ), .ZN(_07628_ ) );
NAND4_X1 _15634_ ( .A1(_06884_ ), .A2(_06665_ ), .A3(_06764_ ), .A4(_06801_ ), .ZN(_07629_ ) );
NAND3_X1 _15635_ ( .A1(_07628_ ), .A2(_07186_ ), .A3(_07629_ ), .ZN(_07630_ ) );
NAND2_X1 _15636_ ( .A1(_07627_ ), .A2(_07630_ ), .ZN(_07631_ ) );
AOI21_X1 _15637_ ( .A(_06966_ ), .B1(_07619_ ), .B2(_07631_ ), .ZN(_07632_ ) );
AND3_X1 _15638_ ( .A1(_07627_ ), .A2(_06986_ ), .A3(_07630_ ), .ZN(_07633_ ) );
NOR4_X1 _15639_ ( .A1(_07283_ ), .A2(_06989_ ), .A3(_07000_ ), .A4(_06891_ ), .ZN(_07634_ ) );
NOR3_X1 _15640_ ( .A1(_07632_ ), .A2(_07633_ ), .A3(_07634_ ), .ZN(_07635_ ) );
OAI211_X1 _15641_ ( .A(_05304_ ), .B(_06698_ ), .C1(_07601_ ), .C2(_07602_ ), .ZN(_07636_ ) );
NAND3_X1 _15642_ ( .A1(_07604_ ), .A2(_07060_ ), .A3(_07636_ ), .ZN(_07637_ ) );
NAND3_X1 _15643_ ( .A1(_06383_ ), .A2(_05298_ ), .A3(_05297_ ), .ZN(_07638_ ) );
NAND3_X1 _15644_ ( .A1(_06703_ ), .A2(_07638_ ), .A3(_07091_ ), .ZN(_07639_ ) );
OR3_X1 _15645_ ( .A1(_05299_ ), .A2(_06383_ ), .A3(_05129_ ), .ZN(_07640_ ) );
NAND2_X1 _15646_ ( .A1(_07638_ ), .A2(_07316_ ), .ZN(_07641_ ) );
AND3_X1 _15647_ ( .A1(_07639_ ), .A2(_07640_ ), .A3(_07641_ ), .ZN(_07642_ ) );
NAND3_X1 _15648_ ( .A1(_07635_ ), .A2(_07637_ ), .A3(_07642_ ), .ZN(_07643_ ) );
AOI21_X1 _15649_ ( .A(_07618_ ), .B1(_07643_ ), .B2(_06947_ ), .ZN(_07644_ ) );
OAI21_X1 _15650_ ( .A(_04135_ ), .B1(_05877_ ), .B2(_06845_ ), .ZN(_07645_ ) );
OAI21_X1 _15651_ ( .A(_07613_ ), .B1(_07644_ ), .B2(_07645_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _15652_ ( .A1(_05905_ ), .A2(_06402_ ), .ZN(_07646_ ) );
AND4_X1 _15653_ ( .A1(_06622_ ), .A2(_06608_ ), .A3(_06626_ ), .A4(_07313_ ), .ZN(_07647_ ) );
NAND2_X1 _15654_ ( .A1(_06666_ ), .A2(_07186_ ), .ZN(_07648_ ) );
NAND3_X1 _15655_ ( .A1(_07516_ ), .A2(_07517_ ), .A3(_06620_ ), .ZN(_07649_ ) );
NOR3_X1 _15656_ ( .A1(_06788_ ), .A2(_06792_ ), .A3(_06612_ ), .ZN(_07650_ ) );
NOR3_X1 _15657_ ( .A1(_06791_ ), .A2(_06806_ ), .A3(_06760_ ), .ZN(_07651_ ) );
NOR2_X1 _15658_ ( .A1(_07650_ ), .A2(_07651_ ), .ZN(_07652_ ) );
OAI211_X1 _15659_ ( .A(_07649_ ), .B(_07132_ ), .C1(_07652_ ), .C2(_07065_ ), .ZN(_07653_ ) );
OAI211_X1 _15660_ ( .A(_07304_ ), .B(_06995_ ), .C1(_07307_ ), .C2(_07065_ ), .ZN(_07654_ ) );
NAND3_X1 _15661_ ( .A1(_07653_ ), .A2(_07654_ ), .A3(_06773_ ), .ZN(_07655_ ) );
NAND2_X1 _15662_ ( .A1(_07648_ ), .A2(_07655_ ), .ZN(_07656_ ) );
OAI21_X1 _15663_ ( .A(_06551_ ), .B1(_07647_ ), .B2(_07656_ ), .ZN(_07657_ ) );
OAI21_X1 _15664_ ( .A(_06752_ ), .B1(_07601_ ), .B2(_07602_ ), .ZN(_07658_ ) );
AOI21_X1 _15665_ ( .A(_07658_ ), .B1(_07602_ ), .B2(_07601_ ), .ZN(_07659_ ) );
OR3_X1 _15666_ ( .A1(_06768_ ), .A2(_06770_ ), .A3(_07345_ ), .ZN(_07660_ ) );
OAI21_X1 _15667_ ( .A(_05382_ ), .B1(_05291_ ), .B2(_02188_ ), .ZN(_07661_ ) );
OAI211_X1 _15668_ ( .A(_07660_ ), .B(_07661_ ), .C1(_07602_ ), .C2(_05387_ ), .ZN(_07662_ ) );
AOI21_X1 _15669_ ( .A(_07130_ ), .B1(_07648_ ), .B2(_07655_ ), .ZN(_07663_ ) );
AND3_X1 _15670_ ( .A1(_05291_ ), .A2(_02188_ ), .A3(_07016_ ), .ZN(_07664_ ) );
NOR4_X1 _15671_ ( .A1(_07659_ ), .A2(_07662_ ), .A3(_07663_ ), .A4(_07664_ ), .ZN(_07665_ ) );
AOI21_X1 _15672_ ( .A(_06549_ ), .B1(_07657_ ), .B2(_07665_ ), .ZN(_07666_ ) );
OAI21_X1 _15673_ ( .A(_04823_ ), .B1(_05392_ ), .B2(_05393_ ), .ZN(_07667_ ) );
NAND2_X1 _15674_ ( .A1(_02319_ ), .A2(_04822_ ), .ZN(_07668_ ) );
NAND2_X1 _15675_ ( .A1(_07667_ ), .A2(_07668_ ), .ZN(_07669_ ) );
XNOR2_X1 _15676_ ( .A(_07669_ ), .B(_04844_ ), .ZN(_07670_ ) );
OR2_X1 _15677_ ( .A1(_07670_ ), .A2(_06956_ ), .ZN(_07671_ ) );
AOI22_X1 _15678_ ( .A1(_05895_ ), .A2(_06839_ ), .B1(\ID_EX_imm [5] ), .B2(_06841_ ), .ZN(_07672_ ) );
AOI21_X1 _15679_ ( .A(_06826_ ), .B1(_07671_ ), .B2(_07672_ ), .ZN(_07673_ ) );
NOR3_X1 _15680_ ( .A1(_07666_ ), .A2(_05552_ ), .A3(_07673_ ), .ZN(_07674_ ) );
NAND2_X1 _15681_ ( .A1(_05893_ ), .A2(_06016_ ), .ZN(_07675_ ) );
NAND2_X1 _15682_ ( .A1(_07675_ ), .A2(_06409_ ), .ZN(_07676_ ) );
OAI21_X1 _15683_ ( .A(_07646_ ), .B1(_07674_ ), .B2(_07676_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_26_D ) );
AND2_X1 _15684_ ( .A1(_05921_ ), .A2(_05922_ ), .ZN(_07677_ ) );
INV_X1 _15685_ ( .A(_07677_ ), .ZN(_07678_ ) );
AND2_X1 _15686_ ( .A1(_05912_ ), .A2(_05483_ ), .ZN(_07679_ ) );
NAND4_X1 _15687_ ( .A1(_06608_ ), .A2(_06626_ ), .A3(_06858_ ), .A4(_07313_ ), .ZN(_07680_ ) );
OR2_X1 _15688_ ( .A1(_06887_ ), .A2(_06888_ ), .ZN(_07681_ ) );
OR3_X1 _15689_ ( .A1(_06895_ ), .A2(_06649_ ), .A3(_06925_ ), .ZN(_07682_ ) );
OR3_X1 _15690_ ( .A1(_06892_ ), .A2(_06896_ ), .A3(_06610_ ), .ZN(_07683_ ) );
AND3_X1 _15691_ ( .A1(_07682_ ), .A2(_07683_ ), .A3(_06783_ ), .ZN(_07684_ ) );
NOR3_X1 _15692_ ( .A1(_07547_ ), .A2(_07548_ ), .A3(_06631_ ), .ZN(_07685_ ) );
NOR3_X1 _15693_ ( .A1(_07684_ ), .A2(_07685_ ), .A3(_06665_ ), .ZN(_07686_ ) );
NOR3_X1 _15694_ ( .A1(_07335_ ), .A2(_06786_ ), .A3(_07338_ ), .ZN(_07687_ ) );
OR3_X1 _15695_ ( .A1(_07686_ ), .A2(_07687_ ), .A3(_06988_ ), .ZN(_07688_ ) );
NAND2_X1 _15696_ ( .A1(_07681_ ), .A2(_07688_ ), .ZN(_07689_ ) );
AOI21_X1 _15697_ ( .A(_06966_ ), .B1(_07680_ ), .B2(_07689_ ), .ZN(_07690_ ) );
NAND3_X1 _15698_ ( .A1(_07681_ ), .A2(_06986_ ), .A3(_07688_ ), .ZN(_07691_ ) );
AOI21_X1 _15699_ ( .A(_05288_ ), .B1(_06692_ ), .B2(_06694_ ), .ZN(_07692_ ) );
OR3_X1 _15700_ ( .A1(_07600_ ), .A2(_07692_ ), .A3(_07023_ ), .ZN(_07693_ ) );
NAND2_X1 _15701_ ( .A1(_05288_ ), .A2(_06940_ ), .ZN(_07694_ ) );
NAND3_X1 _15702_ ( .A1(_06988_ ), .A2(_02319_ ), .A3(_05128_ ), .ZN(_07695_ ) );
OAI21_X1 _15703_ ( .A(_05382_ ), .B1(_06988_ ), .B2(_02319_ ), .ZN(_07696_ ) );
AND3_X1 _15704_ ( .A1(_07694_ ), .A2(_07695_ ), .A3(_07696_ ), .ZN(_07697_ ) );
OR3_X1 _15705_ ( .A1(_06932_ ), .A2(_06770_ ), .A3(_07345_ ), .ZN(_07698_ ) );
NAND4_X1 _15706_ ( .A1(_07691_ ), .A2(_07693_ ), .A3(_07697_ ), .A4(_07698_ ), .ZN(_07699_ ) );
OAI21_X1 _15707_ ( .A(_06947_ ), .B1(_07690_ ), .B2(_07699_ ), .ZN(_07700_ ) );
AND2_X1 _15708_ ( .A1(_07667_ ), .A2(_06834_ ), .ZN(_07701_ ) );
OAI21_X1 _15709_ ( .A(_07701_ ), .B1(_04823_ ), .B2(_07573_ ), .ZN(_07702_ ) );
AOI22_X1 _15710_ ( .A1(_05909_ ), .A2(_06838_ ), .B1(\ID_EX_imm [4] ), .B2(_07157_ ), .ZN(_07703_ ) );
AOI21_X1 _15711_ ( .A(_07197_ ), .B1(_07702_ ), .B2(_07703_ ), .ZN(_07704_ ) );
NOR2_X1 _15712_ ( .A1(_07704_ ), .A2(_06015_ ), .ZN(_07705_ ) );
AOI21_X1 _15713_ ( .A(_07679_ ), .B1(_07700_ ), .B2(_07705_ ), .ZN(_07706_ ) );
MUX2_X1 _15714_ ( .A(_07678_ ), .B(_07706_ ), .S(_04107_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_27_D ) );
AND2_X1 _15715_ ( .A1(_05939_ ), .A2(_05941_ ), .ZN(_07707_ ) );
INV_X1 _15716_ ( .A(_07707_ ), .ZN(_07708_ ) );
AND2_X1 _15717_ ( .A1(_05880_ ), .A2(_05929_ ), .ZN(_07709_ ) );
NOR2_X1 _15718_ ( .A1(_06981_ ), .A2(_06667_ ), .ZN(_07710_ ) );
NOR3_X1 _15719_ ( .A1(_07442_ ), .A2(_06554_ ), .A3(_07443_ ), .ZN(_07711_ ) );
NOR2_X1 _15720_ ( .A1(_06759_ ), .A2(_06756_ ), .ZN(_07712_ ) );
NOR2_X1 _15721_ ( .A1(_06791_ ), .A2(_06760_ ), .ZN(_07713_ ) );
MUX2_X1 _15722_ ( .A(_07712_ ), .B(_07713_ ), .S(_06635_ ), .Z(_07714_ ) );
MUX2_X1 _15723_ ( .A(_07586_ ), .B(_07714_ ), .S(_06630_ ), .Z(_07715_ ) );
AOI211_X1 _15724_ ( .A(_05306_ ), .B(_07711_ ), .C1(_07715_ ), .C2(_06900_ ), .ZN(_07716_ ) );
NOR3_X1 _15725_ ( .A1(_07710_ ), .A2(_07716_ ), .A3(_07130_ ), .ZN(_07717_ ) );
NAND4_X1 _15726_ ( .A1(_06607_ ), .A2(_06625_ ), .A3(_06983_ ), .A4(_06967_ ), .ZN(_07718_ ) );
OR2_X1 _15727_ ( .A1(_07710_ ), .A2(_07716_ ), .ZN(_07719_ ) );
AOI21_X1 _15728_ ( .A(_06856_ ), .B1(_07718_ ), .B2(_07719_ ), .ZN(_07720_ ) );
AOI211_X1 _15729_ ( .A(_07717_ ), .B(_07720_ ), .C1(_07013_ ), .C2(_07248_ ), .ZN(_07721_ ) );
NAND2_X1 _15730_ ( .A1(_05263_ ), .A2(_07091_ ), .ZN(_07722_ ) );
NAND3_X1 _15731_ ( .A1(_07000_ ), .A2(_02235_ ), .A3(_07017_ ), .ZN(_07723_ ) );
OAI21_X1 _15732_ ( .A(_07316_ ), .B1(_07000_ ), .B2(_02235_ ), .ZN(_07724_ ) );
NAND4_X1 _15733_ ( .A1(_07721_ ), .A2(_07722_ ), .A3(_07723_ ), .A4(_07724_ ), .ZN(_07725_ ) );
XNOR2_X1 _15734_ ( .A(_06691_ ), .B(_05263_ ), .ZN(_07726_ ) );
AND2_X1 _15735_ ( .A1(_07726_ ), .A2(_07060_ ), .ZN(_07727_ ) );
OAI21_X1 _15736_ ( .A(_06947_ ), .B1(_07725_ ), .B2(_07727_ ), .ZN(_07728_ ) );
XNOR2_X1 _15737_ ( .A(_05391_ ), .B(_04889_ ), .ZN(_07729_ ) );
NAND2_X1 _15738_ ( .A1(_07729_ ), .A2(_06835_ ), .ZN(_07730_ ) );
OAI21_X1 _15739_ ( .A(_06838_ ), .B1(_05925_ ), .B2(_05926_ ), .ZN(_07731_ ) );
NAND3_X1 _15740_ ( .A1(_06541_ ), .A2(\ID_EX_imm [3] ), .A3(_06539_ ), .ZN(_07732_ ) );
NAND3_X1 _15741_ ( .A1(_07730_ ), .A2(_07731_ ), .A3(_07732_ ), .ZN(_07733_ ) );
AOI21_X1 _15742_ ( .A(_05678_ ), .B1(_07733_ ), .B2(_06546_ ), .ZN(_07734_ ) );
AOI21_X1 _15743_ ( .A(_07709_ ), .B1(_07728_ ), .B2(_07734_ ), .ZN(_07735_ ) );
MUX2_X1 _15744_ ( .A(_07708_ ), .B(_07735_ ), .S(_04107_ ), .Z(\myexu.result_reg_$_DFFE_PP__Q_28_D ) );
NAND3_X1 _15745_ ( .A1(_06412_ ), .A2(_06224_ ), .A3(_06413_ ), .ZN(_07736_ ) );
OAI22_X1 _15746_ ( .A1(_05946_ ), .A2(_07104_ ), .B1(_02259_ ), .B2(_07323_ ), .ZN(_07737_ ) );
OR2_X1 _15747_ ( .A1(_05390_ ), .A2(_04867_ ), .ZN(_07738_ ) );
AOI21_X1 _15748_ ( .A(_06956_ ), .B1(_05390_ ), .B2(_04867_ ), .ZN(_07739_ ) );
AOI21_X1 _15749_ ( .A(_07737_ ), .B1(_07738_ ), .B2(_07739_ ), .ZN(_07740_ ) );
AOI21_X1 _15750_ ( .A(_05482_ ), .B1(_07740_ ), .B2(_03344_ ), .ZN(_07741_ ) );
AND3_X1 _15751_ ( .A1(_07476_ ), .A2(_06626_ ), .A3(_07313_ ), .ZN(_07742_ ) );
NAND2_X1 _15752_ ( .A1(_07056_ ), .A2(_06989_ ), .ZN(_07743_ ) );
NOR2_X1 _15753_ ( .A1(_06924_ ), .A2(_06928_ ), .ZN(_07744_ ) );
NOR2_X1 _15754_ ( .A1(_06895_ ), .A2(_06925_ ), .ZN(_07745_ ) );
MUX2_X1 _15755_ ( .A(_07744_ ), .B(_07745_ ), .S(_06806_ ), .Z(_07746_ ) );
NAND2_X1 _15756_ ( .A1(_07746_ ), .A2(_07070_ ), .ZN(_07747_ ) );
OAI211_X1 _15757_ ( .A(_07747_ ), .B(_07076_ ), .C1(_07070_ ), .C2(_07623_ ), .ZN(_07748_ ) );
OAI211_X1 _15758_ ( .A(_07748_ ), .B(_06669_ ), .C1(_07076_ ), .C2(_07484_ ), .ZN(_07749_ ) );
NAND2_X1 _15759_ ( .A1(_07743_ ), .A2(_07749_ ), .ZN(_07750_ ) );
OAI21_X1 _15760_ ( .A(_06551_ ), .B1(_07742_ ), .B2(_07750_ ), .ZN(_07751_ ) );
NAND2_X1 _15761_ ( .A1(_07750_ ), .A2(_06986_ ), .ZN(_07752_ ) );
NAND2_X1 _15762_ ( .A1(_07066_ ), .A2(_07248_ ), .ZN(_07753_ ) );
AOI21_X1 _15763_ ( .A(_07023_ ), .B1(_06687_ ), .B2(_06688_ ), .ZN(_07754_ ) );
OAI21_X1 _15764_ ( .A(_07754_ ), .B1(_06688_ ), .B2(_06687_ ), .ZN(_07755_ ) );
NAND3_X1 _15765_ ( .A1(_07065_ ), .A2(_02258_ ), .A3(_07017_ ), .ZN(_07756_ ) );
AOI21_X1 _15766_ ( .A(_06815_ ), .B1(_07070_ ), .B2(_05281_ ), .ZN(_07757_ ) );
AOI21_X1 _15767_ ( .A(_07757_ ), .B1(_05268_ ), .B2(_07091_ ), .ZN(_07758_ ) );
AND4_X1 _15768_ ( .A1(_07753_ ), .A2(_07755_ ), .A3(_07756_ ), .A4(_07758_ ), .ZN(_07759_ ) );
NAND3_X1 _15769_ ( .A1(_07751_ ), .A2(_07752_ ), .A3(_07759_ ), .ZN(_07760_ ) );
AOI21_X1 _15770_ ( .A(_07741_ ), .B1(_07760_ ), .B2(_06947_ ), .ZN(_07761_ ) );
OAI21_X1 _15771_ ( .A(_04135_ ), .B1(_05486_ ), .B2(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ), .ZN(_07762_ ) );
OAI21_X1 _15772_ ( .A(_07736_ ), .B1(_07761_ ), .B2(_07762_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_29_D ) );
AND2_X1 _15773_ ( .A1(_05797_ ), .A2(_05798_ ), .ZN(_07763_ ) );
OR2_X1 _15774_ ( .A1(_07763_ ), .A2(_04107_ ), .ZN(_07764_ ) );
AOI21_X1 _15775_ ( .A(_05453_ ), .B1(_07423_ ), .B2(_04409_ ), .ZN(_07765_ ) );
XNOR2_X1 _15776_ ( .A(_07765_ ), .B(_04385_ ), .ZN(_07766_ ) );
AOI22_X1 _15777_ ( .A1(_07766_ ), .A2(_06834_ ), .B1(\ID_EX_imm [29] ), .B2(_06841_ ), .ZN(_07767_ ) );
NAND2_X1 _15778_ ( .A1(_05777_ ), .A2(_06839_ ), .ZN(_07768_ ) );
AOI21_X1 _15779_ ( .A(_07197_ ), .B1(_07767_ ), .B2(_07768_ ), .ZN(_07769_ ) );
OR2_X1 _15780_ ( .A1(_07769_ ), .A2(_06015_ ), .ZN(_07770_ ) );
NOR3_X1 _15781_ ( .A1(_06601_ ), .A2(_06622_ ), .A3(_06625_ ), .ZN(_07771_ ) );
NOR2_X1 _15782_ ( .A1(_06600_ ), .A2(_07771_ ), .ZN(_07772_ ) );
NOR3_X1 _15783_ ( .A1(_06662_ ), .A2(_06623_ ), .A3(_06619_ ), .ZN(_07773_ ) );
AND2_X1 _15784_ ( .A1(_07773_ ), .A2(_06773_ ), .ZN(_07774_ ) );
OAI21_X1 _15785_ ( .A(_06550_ ), .B1(_07772_ ), .B2(_07774_ ), .ZN(_07775_ ) );
OAI21_X1 _15786_ ( .A(_06612_ ), .B1(_06640_ ), .B2(_06647_ ), .ZN(_07776_ ) );
OAI21_X1 _15787_ ( .A(_06806_ ), .B1(_06633_ ), .B2(_06643_ ), .ZN(_07777_ ) );
AND3_X1 _15788_ ( .A1(_07776_ ), .A2(_07777_ ), .A3(_06663_ ), .ZN(_07778_ ) );
NOR2_X1 _15789_ ( .A1(_06646_ ), .A2(_06651_ ), .ZN(_07779_ ) );
INV_X1 _15790_ ( .A(_06650_ ), .ZN(_07780_ ) );
AND2_X1 _15791_ ( .A1(_07780_ ), .A2(_06655_ ), .ZN(_07781_ ) );
MUX2_X1 _15792_ ( .A(_07779_ ), .B(_07781_ ), .S(_06801_ ), .Z(_07782_ ) );
AOI211_X1 _15793_ ( .A(_06995_ ), .B(_07778_ ), .C1(_07782_ ), .C2(_07070_ ), .ZN(_07783_ ) );
NOR3_X1 _15794_ ( .A1(_06803_ ), .A2(_06810_ ), .A3(_06787_ ), .ZN(_07784_ ) );
OAI21_X1 _15795_ ( .A(_06818_ ), .B1(_07783_ ), .B2(_07784_ ), .ZN(_07785_ ) );
OR3_X1 _15796_ ( .A1(_07300_ ), .A2(_06668_ ), .A3(_07301_ ), .ZN(_07786_ ) );
NAND3_X1 _15797_ ( .A1(_07785_ ), .A2(_07786_ ), .A3(_06754_ ), .ZN(_07787_ ) );
OAI21_X1 _15798_ ( .A(_07316_ ), .B1(_05136_ ), .B2(_02909_ ), .ZN(_07788_ ) );
AND3_X1 _15799_ ( .A1(_07773_ ), .A2(_06667_ ), .A3(_06819_ ), .ZN(_07789_ ) );
AOI221_X4 _15800_ ( .A(_07789_ ), .B1(_07414_ ), .B2(_05128_ ), .C1(_05138_ ), .C2(_05386_ ), .ZN(_07790_ ) );
AND4_X1 _15801_ ( .A1(_07775_ ), .A2(_07787_ ), .A3(_07788_ ), .A4(_07790_ ), .ZN(_07791_ ) );
OR2_X1 _15802_ ( .A1(_05141_ ), .A2(_02933_ ), .ZN(_07792_ ) );
AOI21_X1 _15803_ ( .A(_07415_ ), .B1(_07411_ ), .B2(_07792_ ), .ZN(_07793_ ) );
XOR2_X1 _15804_ ( .A(_07793_ ), .B(_05138_ ), .Z(_07794_ ) );
OAI21_X1 _15805_ ( .A(_07791_ ), .B1(_07024_ ), .B2(_07794_ ), .ZN(_07795_ ) );
AOI21_X1 _15806_ ( .A(_07770_ ), .B1(_07795_ ), .B2(_06947_ ), .ZN(_07796_ ) );
NAND2_X1 _15807_ ( .A1(_05788_ ), .A2(_06016_ ), .ZN(_07797_ ) );
NAND2_X1 _15808_ ( .A1(_07797_ ), .A2(_06409_ ), .ZN(_07798_ ) );
OAI21_X1 _15809_ ( .A(_07764_ ), .B1(_07796_ ), .B2(_07798_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_2_D ) );
NAND2_X1 _15810_ ( .A1(_05970_ ), .A2(_06952_ ), .ZN(_07799_ ) );
AOI21_X1 _15811_ ( .A(_06956_ ), .B1(_05100_ ), .B2(_05122_ ), .ZN(_07800_ ) );
OAI21_X1 _15812_ ( .A(_07800_ ), .B1(_05100_ ), .B2(_05122_ ), .ZN(_07801_ ) );
AOI22_X1 _15813_ ( .A1(_05960_ ), .A2(_06851_ ), .B1(\ID_EX_imm [1] ), .B2(_07157_ ), .ZN(_07802_ ) );
AOI21_X1 _15814_ ( .A(_07197_ ), .B1(_07801_ ), .B2(_07802_ ), .ZN(_07803_ ) );
OR2_X1 _15815_ ( .A1(_07803_ ), .A2(_06015_ ), .ZN(_07804_ ) );
AND3_X1 _15816_ ( .A1(_07109_ ), .A2(_06616_ ), .A3(_07313_ ), .ZN(_07805_ ) );
OR2_X1 _15817_ ( .A1(_07121_ ), .A2(_06888_ ), .ZN(_07806_ ) );
OAI21_X1 _15818_ ( .A(_06801_ ), .B1(_06755_ ), .B2(_06766_ ), .ZN(_07807_ ) );
OAI211_X1 _15819_ ( .A(_07807_ ), .B(_06764_ ), .C1(_07712_ ), .C2(_06801_ ), .ZN(_07808_ ) );
OAI211_X1 _15820_ ( .A(_07808_ ), .B(_07132_ ), .C1(_07652_ ), .C2(_07133_ ), .ZN(_07809_ ) );
OAI211_X1 _15821_ ( .A(_07809_ ), .B(_06773_ ), .C1(_07076_ ), .C2(_07519_ ), .ZN(_07810_ ) );
NAND2_X1 _15822_ ( .A1(_07806_ ), .A2(_07810_ ), .ZN(_07811_ ) );
OAI21_X1 _15823_ ( .A(_06551_ ), .B1(_07805_ ), .B2(_07811_ ), .ZN(_07812_ ) );
AOI21_X1 _15824_ ( .A(_07024_ ), .B1(_05272_ ), .B2(_06685_ ), .ZN(_07813_ ) );
OAI21_X1 _15825_ ( .A(_07813_ ), .B1(_05272_ ), .B2(_06685_ ), .ZN(_07814_ ) );
NAND2_X1 _15826_ ( .A1(_07811_ ), .A2(_06986_ ), .ZN(_07815_ ) );
NAND2_X1 _15827_ ( .A1(_07134_ ), .A2(_07248_ ), .ZN(_07816_ ) );
NAND2_X1 _15828_ ( .A1(_06681_ ), .A2(_07017_ ), .ZN(_07817_ ) );
AOI22_X1 _15829_ ( .A1(_05272_ ), .A2(_07091_ ), .B1(_06683_ ), .B2(_07316_ ), .ZN(_07818_ ) );
AND4_X1 _15830_ ( .A1(_07815_ ), .A2(_07816_ ), .A3(_07817_ ), .A4(_07818_ ), .ZN(_07819_ ) );
NAND3_X1 _15831_ ( .A1(_07812_ ), .A2(_07814_ ), .A3(_07819_ ), .ZN(_07820_ ) );
AOI21_X1 _15832_ ( .A(_07804_ ), .B1(_07820_ ), .B2(_06947_ ), .ZN(_07821_ ) );
OAI21_X1 _15833_ ( .A(_04135_ ), .B1(_05486_ ), .B2(\ID_EX_pc [1] ), .ZN(_07822_ ) );
OAI21_X1 _15834_ ( .A(_07799_ ), .B1(_07821_ ), .B2(_07822_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_30_D ) );
AND3_X1 _15835_ ( .A1(_05127_ ), .A2(_06543_ ), .A3(_05133_ ), .ZN(_07823_ ) );
AND4_X1 _15836_ ( .A1(\ID_EX_typ [4] ), .A2(_04322_ ), .A3(\ID_EX_typ [3] ), .A4(_05468_ ), .ZN(_07824_ ) );
OAI21_X1 _15837_ ( .A(_05378_ ), .B1(_07823_ ), .B2(_07824_ ), .ZN(_07825_ ) );
AND3_X1 _15838_ ( .A1(_05990_ ), .A2(_06540_ ), .A3(_06539_ ), .ZN(_07826_ ) );
XNOR2_X1 _15839_ ( .A(_04110_ ), .B(_05121_ ), .ZN(_07827_ ) );
AOI221_X4 _15840_ ( .A(_07826_ ), .B1(\ID_EX_imm [0] ), .B2(_06840_ ), .C1(_07827_ ), .C2(_06834_ ), .ZN(_07828_ ) );
AOI21_X1 _15841_ ( .A(_06547_ ), .B1(_07825_ ), .B2(_07828_ ), .ZN(_07829_ ) );
AND2_X1 _15842_ ( .A1(_05377_ ), .A2(_05152_ ), .ZN(_07830_ ) );
OAI211_X1 _15843_ ( .A(_05157_ ), .B(_05469_ ), .C1(_05461_ ), .C2(_05158_ ), .ZN(_07831_ ) );
NOR3_X1 _15844_ ( .A1(_07830_ ), .A2(_05153_ ), .A3(_07831_ ), .ZN(_07832_ ) );
NAND4_X1 _15845_ ( .A1(_06590_ ), .A2(_05291_ ), .A3(_06556_ ), .A4(_06597_ ), .ZN(_07833_ ) );
OR2_X1 _15846_ ( .A1(_07170_ ), .A2(_06772_ ), .ZN(_07834_ ) );
OR3_X1 _15847_ ( .A1(_07549_ ), .A2(_06785_ ), .A3(_07550_ ), .ZN(_07835_ ) );
NAND3_X1 _15848_ ( .A1(_07682_ ), .A2(_07683_ ), .A3(_06619_ ), .ZN(_07836_ ) );
AOI21_X1 _15849_ ( .A(_06927_ ), .B1(_06684_ ), .B2(_06614_ ), .ZN(_07837_ ) );
MUX2_X1 _15850_ ( .A(_07744_ ), .B(_07837_ ), .S(_06611_ ), .Z(_07838_ ) );
OAI21_X1 _15851_ ( .A(_07836_ ), .B1(_07838_ ), .B2(_06663_ ), .ZN(_07839_ ) );
OAI211_X1 _15852_ ( .A(_07835_ ), .B(_06772_ ), .C1(_07839_ ), .C2(_06769_ ), .ZN(_07840_ ) );
NAND2_X1 _15853_ ( .A1(_07834_ ), .A2(_07840_ ), .ZN(_07841_ ) );
AOI21_X1 _15854_ ( .A(_06856_ ), .B1(_07833_ ), .B2(_07841_ ), .ZN(_07842_ ) );
AND3_X1 _15855_ ( .A1(_07834_ ), .A2(_06820_ ), .A3(_07840_ ), .ZN(_07843_ ) );
AND4_X1 _15856_ ( .A1(_06668_ ), .A2(_07184_ ), .A3(_07075_ ), .A4(_06754_ ), .ZN(_07844_ ) );
NOR4_X1 _15857_ ( .A1(_07832_ ), .A2(_07842_ ), .A3(_07843_ ), .A4(_07844_ ), .ZN(_07845_ ) );
OAI21_X1 _15858_ ( .A(_07060_ ), .B1(_07183_ ), .B2(_05276_ ), .ZN(_07846_ ) );
OAI21_X1 _15859_ ( .A(_06940_ ), .B1(_07183_ ), .B2(_05276_ ), .ZN(_07847_ ) );
NAND3_X1 _15860_ ( .A1(_06857_ ), .A2(_04110_ ), .A3(_07016_ ), .ZN(_07848_ ) );
OAI21_X1 _15861_ ( .A(_05382_ ), .B1(_06857_ ), .B2(_04110_ ), .ZN(_07849_ ) );
AND3_X1 _15862_ ( .A1(_07847_ ), .A2(_07848_ ), .A3(_07849_ ), .ZN(_07850_ ) );
NAND3_X1 _15863_ ( .A1(_07845_ ), .A2(_07846_ ), .A3(_07850_ ), .ZN(_07851_ ) );
AOI211_X1 _15864_ ( .A(_05678_ ), .B(_07829_ ), .C1(_07851_ ), .C2(_06946_ ), .ZN(_07852_ ) );
AND4_X1 _15865_ ( .A1(_06198_ ), .A2(_05481_ ), .A3(\ID_EX_typ [7] ), .A4(\ID_EX_typ [5] ), .ZN(_07853_ ) );
OR3_X1 _15866_ ( .A1(_07852_ ), .A2(_04113_ ), .A3(_07853_ ), .ZN(_07854_ ) );
NAND3_X1 _15867_ ( .A1(_06445_ ), .A2(_06402_ ), .A3(_06446_ ), .ZN(_07855_ ) );
NAND2_X1 _15868_ ( .A1(_07854_ ), .A2(_07855_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_31_D ) );
AND2_X1 _15869_ ( .A1(_05983_ ), .A2(_05984_ ), .ZN(_07856_ ) );
OR2_X1 _15870_ ( .A1(_07856_ ), .A2(_04107_ ), .ZN(_07857_ ) );
AOI22_X1 _15871_ ( .A1(_05975_ ), .A2(_06839_ ), .B1(\ID_EX_imm [28] ), .B2(_06841_ ), .ZN(_07858_ ) );
AOI21_X1 _15872_ ( .A(_06955_ ), .B1(_07423_ ), .B2(_04409_ ), .ZN(_07859_ ) );
OAI21_X1 _15873_ ( .A(_07859_ ), .B1(_04409_ ), .B2(_07423_ ), .ZN(_07860_ ) );
AOI21_X1 _15874_ ( .A(_07197_ ), .B1(_07858_ ), .B2(_07860_ ), .ZN(_07861_ ) );
OR2_X1 _15875_ ( .A1(_07861_ ), .A2(_06015_ ), .ZN(_07862_ ) );
AND2_X1 _15876_ ( .A1(_06860_ ), .A2(_06601_ ), .ZN(_07863_ ) );
NAND3_X1 _15877_ ( .A1(_06608_ ), .A2(_06602_ ), .A3(_07333_ ), .ZN(_07864_ ) );
AND3_X1 _15878_ ( .A1(_06885_ ), .A2(_06785_ ), .A3(_06763_ ), .ZN(_07865_ ) );
NAND2_X1 _15879_ ( .A1(_07865_ ), .A2(_06818_ ), .ZN(_07866_ ) );
NAND2_X1 _15880_ ( .A1(_07864_ ), .A2(_07866_ ), .ZN(_07867_ ) );
OAI21_X1 _15881_ ( .A(_06551_ ), .B1(_07863_ ), .B2(_07867_ ), .ZN(_07868_ ) );
NAND3_X1 _15882_ ( .A1(_05141_ ), .A2(_02933_ ), .A3(_07017_ ), .ZN(_07869_ ) );
AND3_X1 _15883_ ( .A1(_07865_ ), .A2(_06772_ ), .A3(_06820_ ), .ZN(_07870_ ) );
AOI221_X4 _15884_ ( .A(_07870_ ), .B1(_07792_ ), .B2(_05382_ ), .C1(_05376_ ), .C2(_06940_ ), .ZN(_07871_ ) );
AND3_X1 _15885_ ( .A1(_07868_ ), .A2(_07869_ ), .A3(_07871_ ), .ZN(_07872_ ) );
AOI21_X1 _15886_ ( .A(_07024_ ), .B1(_07411_ ), .B2(_05376_ ), .ZN(_07873_ ) );
OAI21_X1 _15887_ ( .A(_07873_ ), .B1(_05376_ ), .B2(_07411_ ), .ZN(_07874_ ) );
AOI21_X1 _15888_ ( .A(_06669_ ), .B1(_07346_ ), .B2(_07347_ ), .ZN(_07875_ ) );
OAI21_X1 _15889_ ( .A(_06801_ ), .B1(_06875_ ), .B2(_06863_ ), .ZN(_07876_ ) );
OAI21_X1 _15890_ ( .A(_06806_ ), .B1(_06872_ ), .B2(_06876_ ), .ZN(_07877_ ) );
AOI21_X1 _15891_ ( .A(_07070_ ), .B1(_07876_ ), .B2(_07877_ ), .ZN(_07878_ ) );
OR3_X1 _15892_ ( .A1(_07369_ ), .A2(_06806_ ), .A3(_06881_ ), .ZN(_07879_ ) );
AOI21_X1 _15893_ ( .A(_07065_ ), .B1(_07372_ ), .B2(_06806_ ), .ZN(_07880_ ) );
AOI21_X1 _15894_ ( .A(_07878_ ), .B1(_07879_ ), .B2(_07880_ ), .ZN(_07881_ ) );
NAND2_X1 _15895_ ( .A1(_07881_ ), .A2(_07076_ ), .ZN(_07882_ ) );
OAI21_X1 _15896_ ( .A(_07000_ ), .B1(_06915_ ), .B2(_06921_ ), .ZN(_07883_ ) );
AOI21_X1 _15897_ ( .A(_06989_ ), .B1(_07882_ ), .B2(_07883_ ), .ZN(_07884_ ) );
OAI21_X1 _15898_ ( .A(_06754_ ), .B1(_07875_ ), .B2(_07884_ ), .ZN(_07885_ ) );
NAND3_X1 _15899_ ( .A1(_07872_ ), .A2(_07874_ ), .A3(_07885_ ), .ZN(_07886_ ) );
AOI21_X1 _15900_ ( .A(_07862_ ), .B1(_07886_ ), .B2(_06947_ ), .ZN(_07887_ ) );
OAI21_X1 _15901_ ( .A(_04135_ ), .B1(_05972_ ), .B2(_06845_ ), .ZN(_07888_ ) );
OAI21_X1 _15902_ ( .A(_07857_ ), .B1(_07887_ ), .B2(_07888_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_3_D ) );
NAND2_X1 _15903_ ( .A1(_06024_ ), .A2(_06952_ ), .ZN(_07889_ ) );
NOR2_X1 _15904_ ( .A1(_06012_ ), .A2(_05500_ ), .ZN(_07890_ ) );
OAI21_X1 _15905_ ( .A(_04558_ ), .B1(_05419_ ), .B2(_05440_ ), .ZN(_07891_ ) );
NAND3_X1 _15906_ ( .A1(_07891_ ), .A2(_05448_ ), .A3(_05446_ ), .ZN(_07892_ ) );
XNOR2_X1 _15907_ ( .A(_02880_ ), .B(_04508_ ), .ZN(_07893_ ) );
AOI21_X1 _15908_ ( .A(_04509_ ), .B1(_07892_ ), .B2(_07893_ ), .ZN(_07894_ ) );
AOI21_X1 _15909_ ( .A(_06955_ ), .B1(_07894_ ), .B2(_04480_ ), .ZN(_07895_ ) );
OAI21_X1 _15910_ ( .A(_07895_ ), .B1(_04480_ ), .B2(_07894_ ), .ZN(_07896_ ) );
OAI21_X1 _15911_ ( .A(_07896_ ), .B1(_02883_ ), .B2(_07323_ ), .ZN(_07897_ ) );
AND2_X1 _15912_ ( .A1(_06007_ ), .A2(_06839_ ), .ZN(_07898_ ) );
OAI21_X1 _15913_ ( .A(_06546_ ), .B1(_07897_ ), .B2(_07898_ ), .ZN(_07899_ ) );
OAI21_X1 _15914_ ( .A(_06786_ ), .B1(_06978_ ), .B2(_06979_ ), .ZN(_07900_ ) );
NOR2_X1 _15915_ ( .A1(_07900_ ), .A2(_06988_ ), .ZN(_07901_ ) );
AOI21_X1 _15916_ ( .A(_07901_ ), .B1(_06598_ ), .B2(_06967_ ), .ZN(_07902_ ) );
OAI211_X1 _15917_ ( .A(_06608_ ), .B(_06602_ ), .C1(_06625_ ), .C2(_06983_ ), .ZN(_07903_ ) );
AOI21_X1 _15918_ ( .A(_06966_ ), .B1(_07902_ ), .B2(_07903_ ), .ZN(_07904_ ) );
NOR3_X1 _15919_ ( .A1(_06994_ ), .A2(_07075_ ), .A3(_06998_ ), .ZN(_07905_ ) );
NOR3_X1 _15920_ ( .A1(_06640_ ), .A2(_06647_ ), .A3(_06612_ ), .ZN(_07906_ ) );
NOR3_X1 _15921_ ( .A1(_06646_ ), .A2(_06765_ ), .A3(_06651_ ), .ZN(_07907_ ) );
NOR2_X1 _15922_ ( .A1(_07906_ ), .A2(_07907_ ), .ZN(_07908_ ) );
OR3_X1 _15923_ ( .A1(_06633_ ), .A2(_06777_ ), .A3(_06643_ ), .ZN(_07909_ ) );
OR3_X1 _15924_ ( .A1(_06804_ ), .A2(_06638_ ), .A3(_06611_ ), .ZN(_07910_ ) );
AND2_X1 _15925_ ( .A1(_07909_ ), .A2(_07910_ ), .ZN(_07911_ ) );
MUX2_X1 _15926_ ( .A(_07908_ ), .B(_07911_ ), .S(_06620_ ), .Z(_07912_ ) );
AOI211_X1 _15927_ ( .A(_07345_ ), .B(_07905_ ), .C1(_07912_ ), .C2(_07076_ ), .ZN(_07913_ ) );
NOR3_X1 _15928_ ( .A1(_07452_ ), .A2(_06773_ ), .A3(_06891_ ), .ZN(_07914_ ) );
NOR3_X1 _15929_ ( .A1(_07900_ ), .A2(_07186_ ), .A3(_07130_ ), .ZN(_07915_ ) );
NOR4_X1 _15930_ ( .A1(_07904_ ), .A2(_07913_ ), .A3(_07914_ ), .A4(_07915_ ), .ZN(_07916_ ) );
NOR2_X2 _15931_ ( .A1(_07396_ ), .A2(_07404_ ), .ZN(_07917_ ) );
OR3_X1 _15932_ ( .A1(_07917_ ), .A2(_05354_ ), .A3(_05362_ ), .ZN(_07918_ ) );
AND2_X1 _15933_ ( .A1(_07918_ ), .A2(_07407_ ), .ZN(_07919_ ) );
INV_X1 _15934_ ( .A(_07391_ ), .ZN(_07920_ ) );
OR2_X2 _15935_ ( .A1(_07919_ ), .A2(_07920_ ), .ZN(_00226_ ) );
AND3_X1 _15936_ ( .A1(_00226_ ), .A2(_07408_ ), .A3(_05346_ ), .ZN(_00227_ ) );
AOI21_X1 _15937_ ( .A(_07408_ ), .B1(_00226_ ), .B2(_05346_ ), .ZN(_00228_ ) );
OR3_X1 _15938_ ( .A1(_00227_ ), .A2(_00228_ ), .A3(_07023_ ), .ZN(_00229_ ) );
AOI21_X1 _15939_ ( .A(_05383_ ), .B1(_05443_ ), .B2(_05340_ ), .ZN(_00230_ ) );
AOI21_X1 _15940_ ( .A(_00230_ ), .B1(_05341_ ), .B2(_06940_ ), .ZN(_00231_ ) );
OR3_X1 _15941_ ( .A1(_05443_ ), .A2(_05340_ ), .A3(_05129_ ), .ZN(_00232_ ) );
AND2_X1 _15942_ ( .A1(_00231_ ), .A2(_00232_ ), .ZN(_00233_ ) );
AND3_X1 _15943_ ( .A1(_07916_ ), .A2(_00229_ ), .A3(_00233_ ), .ZN(_00234_ ) );
OAI21_X1 _15944_ ( .A(_07899_ ), .B1(_00234_ ), .B2(_06549_ ), .ZN(_00235_ ) );
AOI21_X1 _15945_ ( .A(_07890_ ), .B1(_00235_ ), .B2(_05486_ ), .ZN(_00236_ ) );
OAI21_X1 _15946_ ( .A(_07889_ ), .B1(_00236_ ), .B2(_04114_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_4_D ) );
OR2_X1 _15947_ ( .A1(_06470_ ), .A2(_04107_ ), .ZN(_00237_ ) );
AOI21_X1 _15948_ ( .A(_06955_ ), .B1(_07892_ ), .B2(_07893_ ), .ZN(_00238_ ) );
OAI21_X1 _15949_ ( .A(_00238_ ), .B1(_07893_ ), .B2(_07892_ ), .ZN(_00239_ ) );
AOI22_X1 _15950_ ( .A1(_06026_ ), .A2(_06851_ ), .B1(\ID_EX_imm [26] ), .B2(_07157_ ), .ZN(_00240_ ) );
AOI21_X1 _15951_ ( .A(_07197_ ), .B1(_00239_ ), .B2(_00240_ ), .ZN(_00241_ ) );
OR2_X1 _15952_ ( .A1(_00241_ ), .A2(_06015_ ), .ZN(_00242_ ) );
OAI21_X1 _15953_ ( .A(_06602_ ), .B1(_07476_ ), .B2(_07477_ ), .ZN(_00243_ ) );
NOR2_X1 _15954_ ( .A1(_07054_ ), .A2(_06995_ ), .ZN(_00244_ ) );
AND2_X1 _15955_ ( .A1(_00244_ ), .A2(_06888_ ), .ZN(_00245_ ) );
AOI21_X1 _15956_ ( .A(_00245_ ), .B1(_06598_ ), .B2(_07313_ ), .ZN(_00246_ ) );
AOI21_X1 _15957_ ( .A(_06966_ ), .B1(_00243_ ), .B2(_00246_ ), .ZN(_00247_ ) );
NAND2_X1 _15958_ ( .A1(_07492_ ), .A2(_07493_ ), .ZN(_00248_ ) );
NOR2_X1 _15959_ ( .A1(_06772_ ), .A2(_06891_ ), .ZN(_00249_ ) );
AND2_X1 _15960_ ( .A1(_00248_ ), .A2(_00249_ ), .ZN(_00250_ ) );
NOR3_X1 _15961_ ( .A1(_05344_ ), .A2(_02885_ ), .A3(_05129_ ), .ZN(_00251_ ) );
AND3_X1 _15962_ ( .A1(_07376_ ), .A2(_07377_ ), .A3(_06620_ ), .ZN(_00252_ ) );
AOI211_X1 _15963_ ( .A(_06770_ ), .B(_00252_ ), .C1(_07070_ ), .C2(_07374_ ), .ZN(_00253_ ) );
AOI21_X1 _15964_ ( .A(_07076_ ), .B1(_07071_ ), .B2(_07074_ ), .ZN(_00254_ ) );
NOR3_X1 _15965_ ( .A1(_00253_ ), .A2(_07345_ ), .A3(_00254_ ), .ZN(_00255_ ) );
NOR4_X1 _15966_ ( .A1(_00247_ ), .A2(_00250_ ), .A3(_00251_ ), .A4(_00255_ ), .ZN(_00256_ ) );
NAND3_X1 _15967_ ( .A1(_07918_ ), .A2(_07920_ ), .A3(_07407_ ), .ZN(_00257_ ) );
NAND3_X1 _15968_ ( .A1(_00226_ ), .A2(_07060_ ), .A3(_00257_ ), .ZN(_00258_ ) );
AND3_X1 _15969_ ( .A1(_00244_ ), .A2(_06668_ ), .A3(_06820_ ), .ZN(_00259_ ) );
AOI221_X4 _15970_ ( .A(_00259_ ), .B1(_05348_ ), .B2(_07316_ ), .C1(_07391_ ), .C2(_07091_ ), .ZN(_00260_ ) );
NAND3_X1 _15971_ ( .A1(_00256_ ), .A2(_00258_ ), .A3(_00260_ ), .ZN(_00261_ ) );
AOI21_X1 _15972_ ( .A(_00242_ ), .B1(_00261_ ), .B2(_06947_ ), .ZN(_00262_ ) );
NAND2_X1 _15973_ ( .A1(_06029_ ), .A2(_06016_ ), .ZN(_00263_ ) );
NAND2_X1 _15974_ ( .A1(_00263_ ), .A2(_06409_ ), .ZN(_00264_ ) );
OAI21_X1 _15975_ ( .A(_00237_ ), .B1(_00262_ ), .B2(_00264_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_5_D ) );
NOR2_X1 _15976_ ( .A1(_05419_ ), .A2(_05440_ ), .ZN(_00265_ ) );
INV_X1 _15977_ ( .A(_04534_ ), .ZN(_00266_ ) );
OR2_X1 _15978_ ( .A1(_00265_ ), .A2(_00266_ ), .ZN(_00267_ ) );
OAI21_X1 _15979_ ( .A(_00267_ ), .B1(_05358_ ), .B2(_04533_ ), .ZN(_00268_ ) );
AND2_X1 _15980_ ( .A1(_00268_ ), .A2(_04557_ ), .ZN(_00269_ ) );
OAI21_X1 _15981_ ( .A(_06834_ ), .B1(_00268_ ), .B2(_04557_ ), .ZN(_00270_ ) );
OR2_X1 _15982_ ( .A1(_00269_ ), .A2(_00270_ ), .ZN(_00271_ ) );
AOI22_X1 _15983_ ( .A1(_06043_ ), .A2(_06838_ ), .B1(\ID_EX_imm [25] ), .B2(_06840_ ), .ZN(_00272_ ) );
AOI21_X1 _15984_ ( .A(_06547_ ), .B1(_00271_ ), .B2(_00272_ ), .ZN(_00273_ ) );
AND3_X1 _15985_ ( .A1(_07117_ ), .A2(_06786_ ), .A3(_07119_ ), .ZN(_00274_ ) );
AOI21_X1 _15986_ ( .A(_06968_ ), .B1(_06888_ ), .B2(_00274_ ), .ZN(_00275_ ) );
OAI21_X1 _15987_ ( .A(_06602_ ), .B1(_07510_ ), .B2(_07477_ ), .ZN(_00276_ ) );
AOI21_X1 _15988_ ( .A(_06856_ ), .B1(_00275_ ), .B2(_00276_ ), .ZN(_00277_ ) );
NAND2_X1 _15989_ ( .A1(_07527_ ), .A2(_00249_ ), .ZN(_00278_ ) );
AOI21_X1 _15990_ ( .A(_06787_ ), .B1(_07136_ ), .B2(_07137_ ), .ZN(_00279_ ) );
NAND3_X1 _15991_ ( .A1(_07776_ ), .A2(_07777_ ), .A3(_06764_ ), .ZN(_00280_ ) );
NAND3_X1 _15992_ ( .A1(_06805_ ), .A2(_06809_ ), .A3(_06620_ ), .ZN(_00281_ ) );
NAND3_X1 _15993_ ( .A1(_00280_ ), .A2(_00281_ ), .A3(_07075_ ), .ZN(_00282_ ) );
NAND2_X1 _15994_ ( .A1(_00282_ ), .A2(_07248_ ), .ZN(_00283_ ) );
OAI21_X1 _15995_ ( .A(_00278_ ), .B1(_00279_ ), .B2(_00283_ ), .ZN(_00284_ ) );
AND3_X1 _15996_ ( .A1(_00274_ ), .A2(_06888_ ), .A3(_06820_ ), .ZN(_00285_ ) );
NOR3_X1 _15997_ ( .A1(_00277_ ), .A2(_00284_ ), .A3(_00285_ ), .ZN(_00286_ ) );
NOR2_X1 _15998_ ( .A1(_07917_ ), .A2(_05362_ ), .ZN(_00287_ ) );
NOR2_X1 _15999_ ( .A1(_00287_ ), .A2(_05359_ ), .ZN(_00288_ ) );
AOI21_X1 _16000_ ( .A(_07023_ ), .B1(_00288_ ), .B2(_05354_ ), .ZN(_00289_ ) );
OAI21_X1 _16001_ ( .A(_00289_ ), .B1(_05354_ ), .B2(_00288_ ), .ZN(_00290_ ) );
OAI22_X1 _16002_ ( .A1(_05354_ ), .A2(_05387_ ), .B1(_05366_ ), .B2(_06815_ ), .ZN(_00291_ ) );
AOI21_X1 _16003_ ( .A(_00291_ ), .B1(_05367_ ), .B2(_07017_ ), .ZN(_00292_ ) );
NAND3_X1 _16004_ ( .A1(_00286_ ), .A2(_00290_ ), .A3(_00292_ ), .ZN(_00293_ ) );
AOI211_X1 _16005_ ( .A(_05880_ ), .B(_00273_ ), .C1(_00293_ ), .C2(_06946_ ), .ZN(_00294_ ) );
AND2_X1 _16006_ ( .A1(_06054_ ), .A2(_05880_ ), .ZN(_00295_ ) );
OR3_X2 _16007_ ( .A1(_00294_ ), .A2(_04113_ ), .A3(_00295_ ), .ZN(_00296_ ) );
NAND2_X1 _16008_ ( .A1(_06063_ ), .A2(_04114_ ), .ZN(_00297_ ) );
NAND2_X1 _16009_ ( .A1(_00296_ ), .A2(_00297_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_6_D ) );
NAND2_X1 _16010_ ( .A1(_06081_ ), .A2(_06952_ ), .ZN(_00298_ ) );
NOR3_X1 _16011_ ( .A1(_06070_ ), .A2(_06071_ ), .A3(_05500_ ), .ZN(_00299_ ) );
OR3_X1 _16012_ ( .A1(_05419_ ), .A2(_04534_ ), .A3(_05440_ ), .ZN(_00300_ ) );
NAND3_X1 _16013_ ( .A1(_00267_ ), .A2(_06835_ ), .A3(_00300_ ), .ZN(_00301_ ) );
OAI21_X1 _16014_ ( .A(_00301_ ), .B1(_02163_ ), .B2(_07323_ ), .ZN(_00302_ ) );
AND3_X1 _16015_ ( .A1(_06066_ ), .A2(_05760_ ), .A3(_06839_ ), .ZN(_00303_ ) );
OAI21_X1 _16016_ ( .A(_06546_ ), .B1(_00302_ ), .B2(_00303_ ), .ZN(_00304_ ) );
NOR4_X1 _16017_ ( .A1(_06606_ ), .A2(_07557_ ), .A3(_06573_ ), .A4(_06603_ ), .ZN(_00305_ ) );
NOR2_X1 _16018_ ( .A1(_07168_ ), .A2(_06769_ ), .ZN(_00306_ ) );
AND2_X1 _16019_ ( .A1(_00306_ ), .A2(_06667_ ), .ZN(_00307_ ) );
OR2_X1 _16020_ ( .A1(_00305_ ), .A2(_00307_ ), .ZN(_00308_ ) );
OAI21_X1 _16021_ ( .A(_06550_ ), .B1(_00308_ ), .B2(_06968_ ), .ZN(_00309_ ) );
NAND3_X1 _16022_ ( .A1(_00306_ ), .A2(_06773_ ), .A3(_06820_ ), .ZN(_00310_ ) );
AND3_X1 _16023_ ( .A1(_07179_ ), .A2(_07180_ ), .A3(_06665_ ), .ZN(_00311_ ) );
NAND3_X1 _16024_ ( .A1(_07876_ ), .A2(_07877_ ), .A3(_07133_ ), .ZN(_00312_ ) );
NAND3_X1 _16025_ ( .A1(_06917_ ), .A2(_06920_ ), .A3(_06620_ ), .ZN(_00313_ ) );
AOI21_X1 _16026_ ( .A(_06995_ ), .B1(_00312_ ), .B2(_00313_ ), .ZN(_00314_ ) );
OAI21_X1 _16027_ ( .A(_07248_ ), .B1(_00311_ ), .B2(_00314_ ), .ZN(_00315_ ) );
NAND2_X1 _16028_ ( .A1(_07556_ ), .A2(_00249_ ), .ZN(_00316_ ) );
AND4_X1 _16029_ ( .A1(_00309_ ), .A2(_00310_ ), .A3(_00315_ ), .A4(_00316_ ), .ZN(_00317_ ) );
AOI21_X1 _16030_ ( .A(_07023_ ), .B1(_07917_ ), .B2(_05362_ ), .ZN(_00318_ ) );
OAI21_X1 _16031_ ( .A(_00318_ ), .B1(_05362_ ), .B2(_07917_ ), .ZN(_00319_ ) );
OR3_X1 _16032_ ( .A1(_05359_ ), .A2(_05360_ ), .A3(_05387_ ), .ZN(_00320_ ) );
OR3_X1 _16033_ ( .A1(_05357_ ), .A2(_05358_ ), .A3(_05129_ ), .ZN(_00321_ ) );
OR2_X1 _16034_ ( .A1(_05360_ ), .A2(_05383_ ), .ZN(_00322_ ) );
AND3_X1 _16035_ ( .A1(_00320_ ), .A2(_00321_ ), .A3(_00322_ ), .ZN(_00323_ ) );
AND3_X1 _16036_ ( .A1(_00317_ ), .A2(_00319_ ), .A3(_00323_ ), .ZN(_00324_ ) );
OAI21_X1 _16037_ ( .A(_00304_ ), .B1(_00324_ ), .B2(_06549_ ), .ZN(_00325_ ) );
AOI21_X1 _16038_ ( .A(_00299_ ), .B1(_00325_ ), .B2(_05486_ ), .ZN(_00326_ ) );
OAI21_X1 _16039_ ( .A(_00298_ ), .B1(_00326_ ), .B2(_04114_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_7_D ) );
NAND2_X1 _16040_ ( .A1(_06103_ ), .A2(_06952_ ), .ZN(_00327_ ) );
NAND2_X1 _16041_ ( .A1(_06094_ ), .A2(_06016_ ), .ZN(_00328_ ) );
AOI21_X1 _16042_ ( .A(_06891_ ), .B1(_07598_ ), .B2(_06989_ ), .ZN(_00329_ ) );
NAND3_X1 _16043_ ( .A1(_07910_ ), .A2(_07909_ ), .A3(_07133_ ), .ZN(_00330_ ) );
NAND3_X1 _16044_ ( .A1(_06996_ ), .A2(_06620_ ), .A3(_06997_ ), .ZN(_00331_ ) );
AOI21_X1 _16045_ ( .A(_06770_ ), .B1(_00330_ ), .B2(_00331_ ), .ZN(_00332_ ) );
AOI21_X1 _16046_ ( .A(_00332_ ), .B1(_07000_ ), .B2(_07240_ ), .ZN(_00333_ ) );
OAI21_X1 _16047_ ( .A(_00329_ ), .B1(_00333_ ), .B2(_06989_ ), .ZN(_00334_ ) );
AOI21_X1 _16048_ ( .A(_06600_ ), .B1(_06668_ ), .B2(_06624_ ), .ZN(_00335_ ) );
AND2_X1 _16049_ ( .A1(_07591_ ), .A2(_06772_ ), .ZN(_00336_ ) );
OAI21_X1 _16050_ ( .A(_06550_ ), .B1(_00335_ ), .B2(_00336_ ), .ZN(_00337_ ) );
NAND3_X1 _16051_ ( .A1(_07591_ ), .A2(_06773_ ), .A3(_06820_ ), .ZN(_00338_ ) );
AND2_X1 _16052_ ( .A1(_00337_ ), .A2(_00338_ ), .ZN(_00339_ ) );
NAND3_X1 _16053_ ( .A1(_05217_ ), .A2(_02726_ ), .A3(_07017_ ), .ZN(_00340_ ) );
AOI21_X1 _16054_ ( .A(_06815_ ), .B1(_05164_ ), .B2(_02806_ ), .ZN(_00341_ ) );
AOI21_X1 _16055_ ( .A(_00341_ ), .B1(_05167_ ), .B2(_07091_ ), .ZN(_00342_ ) );
AND4_X1 _16056_ ( .A1(_00334_ ), .A2(_00339_ ), .A3(_00340_ ), .A4(_00342_ ), .ZN(_00343_ ) );
INV_X1 _16057_ ( .A(_05174_ ), .ZN(_00344_ ) );
OR3_X1 _16058_ ( .A1(_06937_ ), .A2(_05180_ ), .A3(_05185_ ), .ZN(_00345_ ) );
INV_X1 _16059_ ( .A(_07400_ ), .ZN(_00346_ ) );
AOI21_X1 _16060_ ( .A(_00344_ ), .B1(_00345_ ), .B2(_00346_ ), .ZN(_00347_ ) );
NOR2_X1 _16061_ ( .A1(_05171_ ), .A2(_05168_ ), .ZN(_00348_ ) );
OR3_X1 _16062_ ( .A1(_00347_ ), .A2(_05167_ ), .A3(_00348_ ), .ZN(_00349_ ) );
OAI21_X1 _16063_ ( .A(_05167_ ), .B1(_00347_ ), .B2(_00348_ ), .ZN(_00350_ ) );
NAND3_X1 _16064_ ( .A1(_00349_ ), .A2(_07060_ ), .A3(_00350_ ), .ZN(_00351_ ) );
AOI21_X1 _16065_ ( .A(_06549_ ), .B1(_00343_ ), .B2(_00351_ ), .ZN(_00352_ ) );
NOR4_X1 _16066_ ( .A1(_06828_ ), .A2(_04635_ ), .A3(_04636_ ), .A4(_06829_ ), .ZN(_00353_ ) );
OR2_X1 _16067_ ( .A1(_00353_ ), .A2(_05433_ ), .ZN(_00354_ ) );
AND2_X1 _16068_ ( .A1(_00354_ ), .A2(_04586_ ), .ZN(_00355_ ) );
OR3_X1 _16069_ ( .A1(_00355_ ), .A2(_04609_ ), .A3(_05436_ ), .ZN(_00356_ ) );
OAI21_X1 _16070_ ( .A(_04609_ ), .B1(_00355_ ), .B2(_05436_ ), .ZN(_00357_ ) );
NAND3_X1 _16071_ ( .A1(_00356_ ), .A2(_06835_ ), .A3(_00357_ ), .ZN(_00358_ ) );
AOI22_X1 _16072_ ( .A1(_06089_ ), .A2(_06839_ ), .B1(\ID_EX_imm [23] ), .B2(_06841_ ), .ZN(_00359_ ) );
AOI21_X1 _16073_ ( .A(_06826_ ), .B1(_00358_ ), .B2(_00359_ ), .ZN(_00360_ ) );
OR2_X1 _16074_ ( .A1(_00360_ ), .A2(_05551_ ), .ZN(_00361_ ) );
OAI21_X1 _16075_ ( .A(_00328_ ), .B1(_00352_ ), .B2(_00361_ ), .ZN(_00362_ ) );
OAI21_X1 _16076_ ( .A(_00327_ ), .B1(_00362_ ), .B2(_04114_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_8_D ) );
NAND2_X1 _16077_ ( .A1(_06523_ ), .A2(_06952_ ), .ZN(_00363_ ) );
AND4_X1 _16078_ ( .A1(_06625_ ), .A2(_06607_ ), .A3(_06602_ ), .A4(_07263_ ), .ZN(_00364_ ) );
NAND2_X1 _16079_ ( .A1(_07628_ ), .A2(_07629_ ), .ZN(_00365_ ) );
AND2_X1 _16080_ ( .A1(_00365_ ), .A2(_06888_ ), .ZN(_00366_ ) );
OR3_X1 _16081_ ( .A1(_07863_ ), .A2(_00364_ ), .A3(_00366_ ), .ZN(_00367_ ) );
NAND2_X1 _16082_ ( .A1(_00367_ ), .A2(_06551_ ), .ZN(_00368_ ) );
AND3_X1 _16083_ ( .A1(_00345_ ), .A2(_00344_ ), .A3(_00346_ ), .ZN(_00369_ ) );
OR3_X1 _16084_ ( .A1(_00369_ ), .A2(_00347_ ), .A3(_07023_ ), .ZN(_00370_ ) );
OAI21_X1 _16085_ ( .A(_06770_ ), .B1(_07280_ ), .B2(_07281_ ), .ZN(_00371_ ) );
NAND3_X1 _16086_ ( .A1(_07379_ ), .A2(_07380_ ), .A3(_06787_ ), .ZN(_00372_ ) );
AOI21_X1 _16087_ ( .A(_07186_ ), .B1(_00371_ ), .B2(_00372_ ), .ZN(_00373_ ) );
NOR3_X1 _16088_ ( .A1(_07283_ ), .A2(_06773_ ), .A3(_06770_ ), .ZN(_00374_ ) );
OAI21_X1 _16089_ ( .A(_06754_ ), .B1(_00373_ ), .B2(_00374_ ), .ZN(_00375_ ) );
AOI22_X1 _16090_ ( .A1(_05174_ ), .A2(_07091_ ), .B1(_00348_ ), .B2(_07016_ ), .ZN(_00376_ ) );
AOI21_X1 _16091_ ( .A(_06815_ ), .B1(_05171_ ), .B2(_05168_ ), .ZN(_00377_ ) );
AOI21_X1 _16092_ ( .A(_00377_ ), .B1(_00366_ ), .B2(_06986_ ), .ZN(_00378_ ) );
AND4_X1 _16093_ ( .A1(_00370_ ), .A2(_00375_ ), .A3(_00376_ ), .A4(_00378_ ), .ZN(_00379_ ) );
AOI21_X1 _16094_ ( .A(_06549_ ), .B1(_00368_ ), .B2(_00379_ ), .ZN(_00380_ ) );
AOI21_X1 _16095_ ( .A(_06956_ ), .B1(_00354_ ), .B2(_04586_ ), .ZN(_00381_ ) );
OAI21_X1 _16096_ ( .A(_00381_ ), .B1(_04586_ ), .B2(_00354_ ), .ZN(_00382_ ) );
AOI22_X1 _16097_ ( .A1(_06105_ ), .A2(_06839_ ), .B1(\ID_EX_imm [22] ), .B2(_06841_ ), .ZN(_00383_ ) );
AOI21_X1 _16098_ ( .A(_06826_ ), .B1(_00382_ ), .B2(_00383_ ), .ZN(_00384_ ) );
OR2_X1 _16099_ ( .A1(_00384_ ), .A2(_05569_ ), .ZN(_00385_ ) );
OAI22_X1 _16100_ ( .A1(_00380_ ), .A2(_00385_ ), .B1(_06845_ ), .B2(_06108_ ), .ZN(_00386_ ) );
OAI21_X1 _16101_ ( .A(_00363_ ), .B1(_00386_ ), .B2(_04114_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_9_D ) );
OR2_X1 _16102_ ( .A1(_06180_ ), .A2(_04107_ ), .ZN(_00387_ ) );
NAND2_X1 _16103_ ( .A1(_06171_ ), .A2(_06839_ ), .ZN(_00388_ ) );
AOI21_X1 _16104_ ( .A(_05459_ ), .B1(_07425_ ), .B2(_04455_ ), .ZN(_00389_ ) );
XNOR2_X1 _16105_ ( .A(_00389_ ), .B(_04433_ ), .ZN(_00390_ ) );
AOI22_X1 _16106_ ( .A1(_00390_ ), .A2(_06835_ ), .B1(\ID_EX_imm [31] ), .B2(_06841_ ), .ZN(_00391_ ) );
AOI21_X1 _16107_ ( .A(_06826_ ), .B1(_00388_ ), .B2(_00391_ ), .ZN(_00392_ ) );
NAND3_X1 _16108_ ( .A1(_06553_ ), .A2(_02988_ ), .A3(_07132_ ), .ZN(_00393_ ) );
NOR2_X1 _16109_ ( .A1(_00393_ ), .A2(_07186_ ), .ZN(_00394_ ) );
OAI21_X1 _16110_ ( .A(_06550_ ), .B1(_06860_ ), .B2(_00394_ ), .ZN(_00395_ ) );
NAND3_X1 _16111_ ( .A1(_07241_ ), .A2(_07246_ ), .A3(_00249_ ), .ZN(_00396_ ) );
AOI211_X1 _16112_ ( .A(_06806_ ), .B(_06661_ ), .C1(_06883_ ), .C2(_06857_ ), .ZN(_00397_ ) );
AOI21_X1 _16113_ ( .A(_06801_ ), .B1(_07780_ ), .B2(_06655_ ), .ZN(_00398_ ) );
OR3_X1 _16114_ ( .A1(_00397_ ), .A2(_06620_ ), .A3(_00398_ ), .ZN(_00399_ ) );
OAI21_X1 _16115_ ( .A(_07065_ ), .B1(_07906_ ), .B2(_07907_ ), .ZN(_00400_ ) );
AOI21_X1 _16116_ ( .A(_07000_ ), .B1(_00399_ ), .B2(_00400_ ), .ZN(_00401_ ) );
AND3_X1 _16117_ ( .A1(_00330_ ), .A2(_00331_ ), .A3(_06995_ ), .ZN(_00402_ ) );
OAI21_X1 _16118_ ( .A(_07248_ ), .B1(_00401_ ), .B2(_00402_ ), .ZN(_00403_ ) );
NOR3_X1 _16119_ ( .A1(_00393_ ), .A2(_07186_ ), .A3(_07130_ ), .ZN(_00404_ ) );
AND3_X1 _16120_ ( .A1(_05158_ ), .A2(_02988_ ), .A3(_05128_ ), .ZN(_00405_ ) );
OAI21_X1 _16121_ ( .A(_05382_ ), .B1(_05158_ ), .B2(_02988_ ), .ZN(_00406_ ) );
OAI21_X1 _16122_ ( .A(_00406_ ), .B1(_05155_ ), .B2(_05387_ ), .ZN(_00407_ ) );
NOR3_X1 _16123_ ( .A1(_00404_ ), .A2(_00405_ ), .A3(_00407_ ), .ZN(_00408_ ) );
AND4_X1 _16124_ ( .A1(_00395_ ), .A2(_00396_ ), .A3(_00403_ ), .A4(_00408_ ), .ZN(_00409_ ) );
INV_X1 _16125_ ( .A(_05155_ ), .ZN(_00410_ ) );
OR3_X1 _16126_ ( .A1(_07418_ ), .A2(_00410_ ), .A3(_07388_ ), .ZN(_00411_ ) );
OAI21_X1 _16127_ ( .A(_00410_ ), .B1(_07418_ ), .B2(_07388_ ), .ZN(_00412_ ) );
NAND3_X1 _16128_ ( .A1(_00411_ ), .A2(_07060_ ), .A3(_00412_ ), .ZN(_00413_ ) );
AOI21_X1 _16129_ ( .A(_06549_ ), .B1(_00409_ ), .B2(_00413_ ), .ZN(_00414_ ) );
NOR3_X1 _16130_ ( .A1(_00392_ ), .A2(_05552_ ), .A3(_00414_ ), .ZN(_00415_ ) );
OAI21_X1 _16131_ ( .A(_04135_ ), .B1(_06185_ ), .B2(_06845_ ), .ZN(_00416_ ) );
OAI21_X1 _16132_ ( .A(_00387_ ), .B1(_00415_ ), .B2(_00416_ ), .ZN(\myexu.result_reg_$_DFFE_PP__Q_D ) );
OAI21_X1 _16133_ ( .A(_02017_ ), .B1(_03872_ ), .B2(_03897_ ), .ZN(_00417_ ) );
INV_X1 _16134_ ( .A(\mylsu.state [0] ), .ZN(_00418_ ) );
AOI221_X4 _16135_ ( .A(_01941_ ), .B1(_03954_ ), .B2(_00418_ ), .C1(_02036_ ), .C2(_04016_ ), .ZN(_00419_ ) );
AOI221_X4 _16136_ ( .A(reset ), .B1(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ), .B2(_01941_ ), .C1(_00417_ ), .C2(_00419_ ), .ZN(\myexu.state_$_DFF_PP0__Q_D ) );
NOR2_X1 _16137_ ( .A1(_05481_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_1_D ) );
NOR2_X1 _16138_ ( .A1(_04097_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_2_D ) );
NOR2_X1 _16139_ ( .A1(_05133_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_3_D ) );
NOR2_X1 _16140_ ( .A1(_05479_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_4_D ) );
NOR2_X1 _16141_ ( .A1(_06207_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_5_D ) );
NOR2_X1 _16142_ ( .A1(_05379_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_6_D ) );
NOR2_X1 _16143_ ( .A1(_05628_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_7_D ) );
NOR2_X1 _16144_ ( .A1(_03344_ ), .A2(reset ), .ZN(\myexu.typ_out_$_DFFE_PP0P__Q_D ) );
INV_X1 _16145_ ( .A(IDU_ready_IFU ), .ZN(_00420_ ) );
NAND2_X1 _16146_ ( .A1(_00420_ ), .A2(IDU_valid_EXU ), .ZN(_00421_ ) );
OAI21_X1 _16147_ ( .A(_00421_ ), .B1(_03283_ ), .B2(_03281_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ) );
NOR2_X1 _16148_ ( .A1(_03281_ ), .A2(_03287_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR2_X1 _16149_ ( .A1(_03281_ ), .A2(_03287_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
INV_X1 _16150_ ( .A(_03278_ ), .ZN(_00422_ ) );
NOR4_X1 _16151_ ( .A1(_03287_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03074_ ), .A4(_00422_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ) );
NOR4_X1 _16152_ ( .A1(_03608_ ), .A2(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .A3(_03074_ ), .A4(_03277_ ), .ZN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ) );
AOI21_X1 _16153_ ( .A(_03807_ ), .B1(EXU_valid_LSU ), .B2(IDU_valid_EXU ), .ZN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ) );
OAI21_X1 _16154_ ( .A(_00421_ ), .B1(_00422_ ), .B2(_00420_ ), .ZN(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ) );
OAI22_X1 _16155_ ( .A1(_03278_ ), .A2(_00420_ ), .B1(_01941_ ), .B2(_03328_ ), .ZN(_00423_ ) );
INV_X1 _16156_ ( .A(loaduse_clear ), .ZN(_00424_ ) );
AOI221_X4 _16157_ ( .A(_00423_ ), .B1(\myidu.state [2] ), .B2(_00424_ ), .C1(_03287_ ), .C2(_03807_ ), .ZN(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ) );
NAND3_X1 _16158_ ( .A1(_03077_ ), .A2(\myidu.state [2] ), .A3(loaduse_clear ), .ZN(_00425_ ) );
NAND3_X1 _16159_ ( .A1(_03059_ ), .A2(IDU_valid_EXU ), .A3(_03856_ ), .ZN(_00426_ ) );
AND4_X1 _16160_ ( .A1(_03124_ ), .A2(_03394_ ), .A3(_03198_ ), .A4(_03368_ ), .ZN(_00427_ ) );
AND2_X1 _16161_ ( .A1(_03227_ ), .A2(_00427_ ), .ZN(_00428_ ) );
AOI21_X1 _16162_ ( .A(_00428_ ), .B1(_03353_ ), .B2(_03361_ ), .ZN(_00429_ ) );
INV_X1 _16163_ ( .A(_00429_ ), .ZN(_00430_ ) );
AOI21_X1 _16164_ ( .A(_03364_ ), .B1(_00430_ ), .B2(_03341_ ), .ZN(_00431_ ) );
NAND2_X1 _16165_ ( .A1(_03279_ ), .A2(_03077_ ), .ZN(_00432_ ) );
OAI211_X1 _16166_ ( .A(_00425_ ), .B(_00426_ ), .C1(_00431_ ), .C2(_00432_ ), .ZN(\myidu.state_$_DFF_P__Q_1_D ) );
OAI211_X1 _16167_ ( .A(_03077_ ), .B(_04091_ ), .C1(_03278_ ), .C2(_00420_ ), .ZN(\myidu.state_$_DFF_P__Q_2_D ) );
NAND3_X1 _16168_ ( .A1(_03077_ ), .A2(\myidu.state [2] ), .A3(_00424_ ), .ZN(_00433_ ) );
AOI21_X1 _16169_ ( .A(_03353_ ), .B1(_03340_ ), .B2(_03055_ ), .ZN(_00434_ ) );
NAND4_X1 _16170_ ( .A1(_03278_ ), .A2(IDU_ready_IFU ), .A3(_03059_ ), .A4(_00434_ ), .ZN(_00435_ ) );
AOI21_X1 _16171_ ( .A(_03060_ ), .B1(_03361_ ), .B2(_03353_ ), .ZN(_00436_ ) );
AND2_X1 _16172_ ( .A1(_03124_ ), .A2(_03368_ ), .ZN(_00437_ ) );
BUF_X4 _16173_ ( .A(_00437_ ), .Z(_00438_ ) );
INV_X1 _16174_ ( .A(_00438_ ), .ZN(_00439_ ) );
NOR2_X1 _16175_ ( .A1(_03224_ ), .A2(_03225_ ), .ZN(_00440_ ) );
AND4_X1 _16176_ ( .A1(_03053_ ), .A2(_03166_ ), .A3(_03192_ ), .A4(_03222_ ), .ZN(_00441_ ) );
NOR3_X1 _16177_ ( .A1(_00440_ ), .A2(_03209_ ), .A3(_00441_ ), .ZN(_00442_ ) );
NOR3_X1 _16178_ ( .A1(_03379_ ), .A2(_03294_ ), .A3(_03378_ ), .ZN(_00443_ ) );
NOR3_X1 _16179_ ( .A1(_03225_ ), .A2(_03294_ ), .A3(_03378_ ), .ZN(_00444_ ) );
NOR2_X1 _16180_ ( .A1(_00443_ ), .A2(_00444_ ), .ZN(_00445_ ) );
AOI21_X1 _16181_ ( .A(_03406_ ), .B1(_03208_ ), .B2(_03389_ ), .ZN(_00446_ ) );
NAND4_X1 _16182_ ( .A1(_00442_ ), .A2(_03221_ ), .A3(_00445_ ), .A4(_00446_ ), .ZN(_00447_ ) );
OAI211_X1 _16183_ ( .A(_03278_ ), .B(_00436_ ), .C1(_00439_ ), .C2(_00447_ ), .ZN(_00448_ ) );
OAI211_X1 _16184_ ( .A(_00433_ ), .B(_00435_ ), .C1(_00448_ ), .C2(_00420_ ), .ZN(\myidu.state_$_DFF_P__Q_D ) );
NOR2_X1 _16185_ ( .A1(_03275_ ), .A2(IDU_ready_IFU ), .ZN(_00449_ ) );
NOR2_X1 _16186_ ( .A1(_03275_ ), .A2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(_00450_ ) );
NOR2_X1 _16187_ ( .A1(\myifu.state [0] ), .A2(\myifu.state [1] ), .ZN(_00451_ ) );
NOR4_X1 _16188_ ( .A1(_00449_ ), .A2(_00450_ ), .A3(reset ), .A4(_00451_ ), .ZN(\myifu.check_assert_$_DFFE_PP__Q_E ) );
OAI21_X1 _16189_ ( .A(_01735_ ), .B1(_04095_ ), .B2(_04091_ ), .ZN(\myifu.check_assert_$_ORNOT__A_Y_$_MUX__A_S_$_OR__A_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
CLKBUF_X2 _16190_ ( .A(_03942_ ), .Z(_00452_ ) );
OR3_X1 _16191_ ( .A1(_01964_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00453_ ) );
OAI21_X1 _16192_ ( .A(_00453_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03943_ ), .ZN(_00454_ ) );
MUX2_X1 _16193_ ( .A(\io_master_rdata [31] ), .B(_00454_ ), .S(_02060_ ), .Z(_00455_ ) );
AND2_X1 _16194_ ( .A1(_00455_ ), .A2(_02012_ ), .ZN(\myifu.data_in [31] ) );
OR3_X1 _16195_ ( .A1(_01964_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00456_ ) );
OAI21_X1 _16196_ ( .A(_00456_ ), .B1(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ), .B2(_03943_ ), .ZN(_00457_ ) );
MUX2_X1 _16197_ ( .A(\io_master_rdata [30] ), .B(_00457_ ), .S(_02060_ ), .Z(_00458_ ) );
AND2_X1 _16198_ ( .A1(_00458_ ), .A2(_02012_ ), .ZN(\myifu.data_in [30] ) );
OR3_X1 _16199_ ( .A1(_01964_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00459_ ) );
OAI211_X1 _16200_ ( .A(_02006_ ), .B(_00459_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03944_ ), .ZN(_00460_ ) );
BUF_X8 _16201_ ( .A(_02006_ ), .Z(_00461_ ) );
OAI21_X1 _16202_ ( .A(_00460_ ), .B1(\io_master_rdata [21] ), .B2(_00461_ ), .ZN(_00462_ ) );
NOR2_X1 _16203_ ( .A1(_00462_ ), .A2(_03911_ ), .ZN(\myifu.data_in [21] ) );
OR2_X1 _16204_ ( .A1(_02008_ ), .A2(\io_master_rdata [20] ), .ZN(_00463_ ) );
CLKBUF_X2 _16205_ ( .A(_00452_ ), .Z(_00464_ ) );
CLKBUF_X2 _16206_ ( .A(_00464_ ), .Z(_00465_ ) );
OR3_X1 _16207_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00466_ ) );
OAI211_X1 _16208_ ( .A(_02008_ ), .B(_00466_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00467_ ) );
AND3_X1 _16209_ ( .A1(_00463_ ), .A2(_00467_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [20] ) );
OR2_X1 _16210_ ( .A1(_02008_ ), .A2(\io_master_rdata [19] ), .ZN(_00468_ ) );
OR3_X1 _16211_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00469_ ) );
OAI211_X1 _16212_ ( .A(_02008_ ), .B(_00469_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00470_ ) );
AND3_X1 _16213_ ( .A1(_00468_ ), .A2(_00470_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [19] ) );
MUX2_X1 _16214_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03944_ ), .Z(_00471_ ) );
OR2_X1 _16215_ ( .A1(_02062_ ), .A2(_00471_ ), .ZN(_00472_ ) );
INV_X1 _16216_ ( .A(\io_master_rdata [18] ), .ZN(_00473_ ) );
OR2_X1 _16217_ ( .A1(_02060_ ), .A2(_00473_ ), .ZN(_00474_ ) );
AOI21_X1 _16218_ ( .A(_03796_ ), .B1(_00472_ ), .B2(_00474_ ), .ZN(\myifu.data_in [18] ) );
BUF_X2 _16219_ ( .A(_02007_ ), .Z(_00475_ ) );
OR2_X1 _16220_ ( .A1(_00475_ ), .A2(\io_master_rdata [17] ), .ZN(_00476_ ) );
OR3_X1 _16221_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00477_ ) );
OAI211_X1 _16222_ ( .A(_00475_ ), .B(_00477_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00478_ ) );
AND3_X1 _16223_ ( .A1(_00476_ ), .A2(_00478_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [17] ) );
OR2_X1 _16224_ ( .A1(_00475_ ), .A2(\io_master_rdata [16] ), .ZN(_00479_ ) );
OR3_X1 _16225_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00480_ ) );
OAI211_X1 _16226_ ( .A(_00475_ ), .B(_00480_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03945_ ), .ZN(_00481_ ) );
AND3_X1 _16227_ ( .A1(_00479_ ), .A2(_00481_ ), .A3(\io_master_arburst [0] ), .ZN(\myifu.data_in [16] ) );
OR3_X1 _16228_ ( .A1(_01964_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_03942_ ), .ZN(_00482_ ) );
OAI211_X1 _16229_ ( .A(_02006_ ), .B(_00482_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03943_ ), .ZN(_00483_ ) );
OAI21_X2 _16230_ ( .A(_00483_ ), .B1(\io_master_rdata [15] ), .B2(_02006_ ), .ZN(_00484_ ) );
NOR2_X1 _16231_ ( .A1(_00484_ ), .A2(_03911_ ), .ZN(\myifu.data_in [15] ) );
OR3_X1 _16232_ ( .A1(_02010_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00485_ ) );
OAI211_X1 _16233_ ( .A(_00461_ ), .B(_00485_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03944_ ), .ZN(_00486_ ) );
OAI21_X1 _16234_ ( .A(_00486_ ), .B1(\io_master_rdata [14] ), .B2(_02007_ ), .ZN(_00487_ ) );
NOR2_X1 _16235_ ( .A1(_00487_ ), .A2(_03911_ ), .ZN(\myifu.data_in [14] ) );
OR2_X1 _16236_ ( .A1(_02007_ ), .A2(\io_master_rdata [13] ), .ZN(_00488_ ) );
OR3_X1 _16237_ ( .A1(_02010_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00464_ ), .ZN(_00489_ ) );
OAI211_X1 _16238_ ( .A(_02007_ ), .B(_00489_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03945_ ), .ZN(_00490_ ) );
AND3_X1 _16239_ ( .A1(_00488_ ), .A2(_00490_ ), .A3(_03894_ ), .ZN(\myifu.data_in [13] ) );
OR2_X1 _16240_ ( .A1(_02008_ ), .A2(\io_master_rdata [12] ), .ZN(_00491_ ) );
OR3_X1 _16241_ ( .A1(_02012_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00492_ ) );
OAI211_X1 _16242_ ( .A(_02009_ ), .B(_00492_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00493_ ) );
AND3_X1 _16243_ ( .A1(_00491_ ), .A2(_00493_ ), .A3(_03894_ ), .ZN(\myifu.data_in [12] ) );
OR3_X1 _16244_ ( .A1(_02010_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00464_ ), .ZN(_00494_ ) );
OAI211_X1 _16245_ ( .A(_00461_ ), .B(_00494_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03944_ ), .ZN(_00495_ ) );
OAI21_X2 _16246_ ( .A(_00495_ ), .B1(\io_master_rdata [29] ), .B2(_02007_ ), .ZN(_00496_ ) );
BUF_X4 _16247_ ( .A(_03796_ ), .Z(_00497_ ) );
NOR2_X1 _16248_ ( .A1(_00496_ ), .A2(_00497_ ), .ZN(\myifu.data_in [29] ) );
OR2_X1 _16249_ ( .A1(_02007_ ), .A2(\io_master_rdata [11] ), .ZN(_00498_ ) );
OR3_X1 _16250_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00464_ ), .ZN(_00499_ ) );
OAI211_X1 _16251_ ( .A(_00475_ ), .B(_00499_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03945_ ), .ZN(_00500_ ) );
AND3_X1 _16252_ ( .A1(_00498_ ), .A2(_00500_ ), .A3(_03894_ ), .ZN(\myifu.data_in [11] ) );
OR2_X1 _16253_ ( .A1(_02007_ ), .A2(\io_master_rdata [10] ), .ZN(_00501_ ) );
OR3_X1 _16254_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00464_ ), .ZN(_00502_ ) );
OAI211_X1 _16255_ ( .A(_00475_ ), .B(_00502_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03945_ ), .ZN(_00503_ ) );
AND3_X1 _16256_ ( .A1(_00501_ ), .A2(_00503_ ), .A3(_02012_ ), .ZN(\myifu.data_in [10] ) );
OR2_X1 _16257_ ( .A1(_02007_ ), .A2(\io_master_rdata [9] ), .ZN(_00504_ ) );
OR3_X1 _16258_ ( .A1(_02010_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00464_ ), .ZN(_00505_ ) );
OAI211_X1 _16259_ ( .A(_00475_ ), .B(_00505_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03945_ ), .ZN(_00506_ ) );
AND3_X1 _16260_ ( .A1(_00504_ ), .A2(_00506_ ), .A3(_03894_ ), .ZN(\myifu.data_in [9] ) );
OR2_X1 _16261_ ( .A1(_02007_ ), .A2(\io_master_rdata [8] ), .ZN(_00507_ ) );
OR3_X1 _16262_ ( .A1(_02010_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00464_ ), .ZN(_00508_ ) );
OAI211_X1 _16263_ ( .A(_00475_ ), .B(_00508_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03945_ ), .ZN(_00509_ ) );
AND3_X1 _16264_ ( .A1(_00507_ ), .A2(_00509_ ), .A3(_03894_ ), .ZN(\myifu.data_in [8] ) );
OR2_X1 _16265_ ( .A1(_02006_ ), .A2(\io_master_rdata [7] ), .ZN(_00510_ ) );
OR3_X1 _16266_ ( .A1(_01964_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00511_ ) );
OAI211_X1 _16267_ ( .A(_02006_ ), .B(_00511_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03943_ ), .ZN(_00512_ ) );
AND3_X1 _16268_ ( .A1(_00510_ ), .A2(_00512_ ), .A3(_03894_ ), .ZN(\myifu.data_in [7] ) );
OR3_X1 _16269_ ( .A1(_02010_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00513_ ) );
OAI211_X1 _16270_ ( .A(_00461_ ), .B(_00513_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03944_ ), .ZN(_00514_ ) );
OAI21_X2 _16271_ ( .A(_00514_ ), .B1(\io_master_rdata [6] ), .B2(_00461_ ), .ZN(_00515_ ) );
NOR2_X1 _16272_ ( .A1(_00515_ ), .A2(_00497_ ), .ZN(\myifu.data_in [6] ) );
OR3_X1 _16273_ ( .A1(_01964_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00516_ ) );
OAI211_X1 _16274_ ( .A(_00461_ ), .B(_00516_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03944_ ), .ZN(_00517_ ) );
OAI21_X2 _16275_ ( .A(_00517_ ), .B1(\io_master_rdata [5] ), .B2(_00461_ ), .ZN(_00518_ ) );
NOR2_X1 _16276_ ( .A1(_00518_ ), .A2(_00497_ ), .ZN(\myifu.data_in [5] ) );
OR3_X1 _16277_ ( .A1(_02012_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00519_ ) );
OAI211_X1 _16278_ ( .A(_02009_ ), .B(_00519_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00520_ ) );
OAI21_X1 _16279_ ( .A(_00520_ ), .B1(\io_master_rdata [4] ), .B2(_02009_ ), .ZN(_00521_ ) );
NOR2_X1 _16280_ ( .A1(_00521_ ), .A2(_03911_ ), .ZN(\myifu.data_in [4] ) );
OR3_X1 _16281_ ( .A1(_02012_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00522_ ) );
OAI211_X1 _16282_ ( .A(_02009_ ), .B(_00522_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00523_ ) );
OAI21_X1 _16283_ ( .A(_00523_ ), .B1(\io_master_rdata [3] ), .B2(_02009_ ), .ZN(_00524_ ) );
NOR2_X1 _16284_ ( .A1(_00524_ ), .A2(_00497_ ), .ZN(\myifu.data_in [3] ) );
OR3_X1 _16285_ ( .A1(_02012_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00525_ ) );
OAI211_X1 _16286_ ( .A(_02009_ ), .B(_00525_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00526_ ) );
OAI21_X1 _16287_ ( .A(_00526_ ), .B1(\io_master_rdata [2] ), .B2(_02009_ ), .ZN(_00527_ ) );
NOR2_X1 _16288_ ( .A1(_00527_ ), .A2(_03911_ ), .ZN(\myifu.data_in [2] ) );
OR2_X1 _16289_ ( .A1(_00475_ ), .A2(\io_master_rdata [28] ), .ZN(_00528_ ) );
OR3_X1 _16290_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00464_ ), .ZN(_00529_ ) );
OAI211_X1 _16291_ ( .A(_00475_ ), .B(_00529_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03945_ ), .ZN(_00530_ ) );
AND3_X1 _16292_ ( .A1(_00528_ ), .A2(_00530_ ), .A3(_03894_ ), .ZN(\myifu.data_in [28] ) );
OR3_X1 _16293_ ( .A1(_02011_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00465_ ), .ZN(_00531_ ) );
OAI211_X1 _16294_ ( .A(_02008_ ), .B(_00531_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(\io_master_araddr [2] ), .ZN(_00532_ ) );
OAI21_X1 _16295_ ( .A(_00532_ ), .B1(\io_master_rdata [1] ), .B2(_02008_ ), .ZN(_00533_ ) );
NOR2_X1 _16296_ ( .A1(_00533_ ), .A2(_03911_ ), .ZN(\myifu.data_in [1] ) );
OR3_X1 _16297_ ( .A1(_02011_ ), .A2(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ), .A3(_00465_ ), .ZN(_00534_ ) );
OAI211_X1 _16298_ ( .A(_02008_ ), .B(_00534_ ), .C1(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ), .C2(\io_master_araddr [2] ), .ZN(_00535_ ) );
OAI21_X1 _16299_ ( .A(_00535_ ), .B1(\io_master_rdata [0] ), .B2(_02008_ ), .ZN(_00536_ ) );
NOR2_X1 _16300_ ( .A1(_00536_ ), .A2(_03911_ ), .ZN(\myifu.data_in [0] ) );
MUX2_X1 _16301_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03944_ ), .Z(_00537_ ) );
OR2_X1 _16302_ ( .A1(_02062_ ), .A2(_00537_ ), .ZN(_00538_ ) );
NAND2_X1 _16303_ ( .A1(_02062_ ), .A2(\io_master_rdata [27] ), .ZN(_00539_ ) );
AOI21_X1 _16304_ ( .A(_03911_ ), .B1(_00538_ ), .B2(_00539_ ), .ZN(\myifu.data_in [27] ) );
NAND2_X1 _16305_ ( .A1(_02062_ ), .A2(\io_master_rdata [26] ), .ZN(_00540_ ) );
OR3_X1 _16306_ ( .A1(_02010_ ), .A2(_01665_ ), .A3(_00464_ ), .ZN(_00541_ ) );
OAI211_X1 _16307_ ( .A(_02060_ ), .B(_00541_ ), .C1(_01651_ ), .C2(_03945_ ), .ZN(_00542_ ) );
AOI21_X1 _16308_ ( .A(_03910_ ), .B1(_00540_ ), .B2(_00542_ ), .ZN(\myifu.data_in [26] ) );
MUX2_X1 _16309_ ( .A(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ), .B(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ), .S(_03944_ ), .Z(_00543_ ) );
OR2_X1 _16310_ ( .A1(_02062_ ), .A2(_00543_ ), .ZN(_00544_ ) );
NAND2_X1 _16311_ ( .A1(_02062_ ), .A2(\io_master_rdata [25] ), .ZN(_00545_ ) );
AOI21_X1 _16312_ ( .A(_03910_ ), .B1(_00544_ ), .B2(_00545_ ), .ZN(\myifu.data_in [25] ) );
NAND2_X1 _16313_ ( .A1(_02062_ ), .A2(\io_master_rdata [24] ), .ZN(_00546_ ) );
OR3_X1 _16314_ ( .A1(_02010_ ), .A2(_01725_ ), .A3(_00464_ ), .ZN(_00547_ ) );
OAI211_X1 _16315_ ( .A(_02060_ ), .B(_00547_ ), .C1(_01657_ ), .C2(_03945_ ), .ZN(_00548_ ) );
AOI21_X1 _16316_ ( .A(_03911_ ), .B1(_00546_ ), .B2(_00548_ ), .ZN(\myifu.data_in [24] ) );
OR3_X1 _16317_ ( .A1(_01964_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00549_ ) );
OAI211_X1 _16318_ ( .A(_02006_ ), .B(_00549_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03943_ ), .ZN(_00550_ ) );
OAI21_X4 _16319_ ( .A(_00550_ ), .B1(\io_master_rdata [23] ), .B2(_00461_ ), .ZN(_00551_ ) );
NOR2_X1 _16320_ ( .A1(_00551_ ), .A2(_00497_ ), .ZN(\myifu.data_in [23] ) );
OR3_X1 _16321_ ( .A1(_02010_ ), .A2(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ), .A3(_00452_ ), .ZN(_00552_ ) );
OAI211_X1 _16322_ ( .A(_00461_ ), .B(_00552_ ), .C1(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ), .C2(_03944_ ), .ZN(_00553_ ) );
OAI21_X2 _16323_ ( .A(_00553_ ), .B1(\io_master_rdata [22] ), .B2(_00461_ ), .ZN(_00554_ ) );
NOR2_X1 _16324_ ( .A1(_00554_ ), .A2(_00497_ ), .ZN(\myifu.data_in [22] ) );
INV_X1 _16325_ ( .A(_00164_ ), .ZN(_00555_ ) );
NAND2_X1 _16326_ ( .A1(_00555_ ), .A2(_02049_ ), .ZN(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16327_ ( .A1(_03726_ ), .A2(fanout_net_12 ), .ZN(_00556_ ) );
INV_X1 _16328_ ( .A(\myifu.myicache.valid_data_in ), .ZN(_00557_ ) );
OAI21_X1 _16329_ ( .A(_02049_ ), .B1(_00556_ ), .B2(_00557_ ), .ZN(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16330_ ( .A1(_03737_ ), .A2(fanout_net_16 ), .ZN(_00558_ ) );
OAI21_X1 _16331_ ( .A(_02049_ ), .B1(_00558_ ), .B2(_00557_ ), .ZN(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ) );
NAND2_X1 _16332_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .ZN(_00559_ ) );
OAI21_X1 _16333_ ( .A(_02049_ ), .B1(_00559_ ), .B2(_00557_ ), .ZN(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ) );
NAND2_X1 _16334_ ( .A1(_00439_ ), .A2(\IF_ID_inst [8] ), .ZN(_00560_ ) );
AND2_X1 _16335_ ( .A1(_00437_ ), .A2(_03395_ ), .ZN(_00561_ ) );
NAND3_X1 _16336_ ( .A1(_03147_ ), .A2(_03129_ ), .A3(_03371_ ), .ZN(_00562_ ) );
AOI21_X1 _16337_ ( .A(_03113_ ), .B1(_03147_ ), .B2(_03148_ ), .ZN(_00563_ ) );
AND4_X1 _16338_ ( .A1(_03055_ ), .A2(_03390_ ), .A3(_00562_ ), .A4(_00563_ ), .ZN(_00564_ ) );
NOR4_X1 _16339_ ( .A1(_03380_ ), .A2(_03382_ ), .A3(_03159_ ), .A4(_03220_ ), .ZN(_00565_ ) );
NAND3_X1 _16340_ ( .A1(_00561_ ), .A2(_00564_ ), .A3(_00565_ ), .ZN(_00566_ ) );
AND2_X1 _16341_ ( .A1(_00566_ ), .A2(_03300_ ), .ZN(_00567_ ) );
OAI221_X1 _16342_ ( .A(_00560_ ), .B1(_03285_ ), .B2(_03056_ ), .C1(_00567_ ), .C2(_03064_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ) );
NOR2_X1 _16343_ ( .A1(_03340_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00568_ ) );
AND3_X1 _16344_ ( .A1(_03440_ ), .A2(_03112_ ), .A3(\IF_ID_inst [31] ), .ZN(_00569_ ) );
NOR2_X1 _16345_ ( .A1(_00568_ ), .A2(_00569_ ), .ZN(_00570_ ) );
BUF_X4 _16346_ ( .A(_00570_ ), .Z(_00571_ ) );
OAI21_X1 _16347_ ( .A(_00571_ ), .B1(_00561_ ), .B2(_03058_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ) );
BUF_X4 _16348_ ( .A(_03395_ ), .Z(_00572_ ) );
BUF_X4 _16349_ ( .A(_00438_ ), .Z(_00573_ ) );
OAI221_X1 _16350_ ( .A(_00571_ ), .B1(_03063_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00573_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ) );
OAI221_X1 _16351_ ( .A(_00571_ ), .B1(_03064_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00573_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ) );
OAI221_X1 _16352_ ( .A(_00571_ ), .B1(_03067_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00573_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ) );
INV_X1 _16353_ ( .A(_00568_ ), .ZN(_00574_ ) );
BUF_X4 _16354_ ( .A(_03057_ ), .Z(_00575_ ) );
BUF_X4 _16355_ ( .A(_00437_ ), .Z(_00576_ ) );
OAI221_X1 _16356_ ( .A(_00574_ ), .B1(_00575_ ), .B2(_00576_ ), .C1(_03162_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ) );
OAI221_X1 _16357_ ( .A(_00574_ ), .B1(_00575_ ), .B2(_00576_ ), .C1(_03163_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ) );
OAI221_X1 _16358_ ( .A(_00574_ ), .B1(_00575_ ), .B2(_00576_ ), .C1(_03164_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ) );
OAI221_X1 _16359_ ( .A(_00574_ ), .B1(_00575_ ), .B2(_00576_ ), .C1(_03285_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ) );
OAI221_X1 _16360_ ( .A(_00574_ ), .B1(_00575_ ), .B2(_00438_ ), .C1(_03080_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ) );
OAI221_X1 _16361_ ( .A(_00574_ ), .B1(_00575_ ), .B2(_00438_ ), .C1(_03178_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ) );
OAI221_X1 _16362_ ( .A(_00574_ ), .B1(_00575_ ), .B2(_00438_ ), .C1(_03117_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ) );
OAI221_X1 _16363_ ( .A(_00574_ ), .B1(_03057_ ), .B2(_00438_ ), .C1(_03078_ ), .C2(_03160_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ) );
OAI221_X1 _16364_ ( .A(_00571_ ), .B1(_03068_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00573_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ) );
OR2_X1 _16365_ ( .A1(_03124_ ), .A2(_03057_ ), .ZN(_00577_ ) );
OR2_X1 _16366_ ( .A1(_03368_ ), .A2(_03079_ ), .ZN(_00578_ ) );
NAND4_X1 _16367_ ( .A1(_00574_ ), .A2(_03451_ ), .A3(_00577_ ), .A4(_00578_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ) );
INV_X1 _16368_ ( .A(_03517_ ), .ZN(_00579_ ) );
OAI221_X1 _16369_ ( .A(_00579_ ), .B1(_03340_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .C1(_00573_ ), .C2(_03063_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ) );
INV_X1 _16370_ ( .A(_03455_ ), .ZN(_00580_ ) );
OAI221_X1 _16371_ ( .A(_00580_ ), .B1(_03340_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C1(_00573_ ), .C2(_03068_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ) );
OAI221_X1 _16372_ ( .A(_03509_ ), .B1(_03340_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .C1(_00573_ ), .C2(_03069_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ) );
OR2_X1 _16373_ ( .A1(_00438_ ), .A2(_03070_ ), .ZN(_00581_ ) );
OAI221_X1 _16374_ ( .A(_00581_ ), .B1(_03070_ ), .B2(_03300_ ), .C1(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .C2(_03340_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ) );
INV_X1 _16375_ ( .A(_03497_ ), .ZN(_00582_ ) );
OAI221_X1 _16376_ ( .A(_00582_ ), .B1(_03340_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .C1(_00573_ ), .C2(_03071_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ) );
INV_X1 _16377_ ( .A(_03488_ ), .ZN(_00583_ ) );
OAI221_X1 _16378_ ( .A(_00583_ ), .B1(_03340_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ), .C1(_00573_ ), .C2(_03072_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ) );
OAI221_X1 _16379_ ( .A(_00571_ ), .B1(_03069_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00573_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ) );
OAI221_X1 _16380_ ( .A(_00571_ ), .B1(_03070_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00576_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ) );
OAI221_X1 _16381_ ( .A(_00571_ ), .B1(_03071_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00576_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ) );
OAI221_X1 _16382_ ( .A(_00571_ ), .B1(_03072_ ), .B2(_00572_ ), .C1(_03058_ ), .C2(_00576_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ) );
OAI221_X1 _16383_ ( .A(_00571_ ), .B1(_03073_ ), .B2(_00572_ ), .C1(_00575_ ), .C2(_00576_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ) );
OAI221_X1 _16384_ ( .A(_00570_ ), .B1(_03075_ ), .B2(_00572_ ), .C1(_00575_ ), .C2(_00576_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ) );
OAI221_X1 _16385_ ( .A(_00570_ ), .B1(_03076_ ), .B2(_03395_ ), .C1(_00575_ ), .C2(_00576_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ) );
OAI21_X1 _16386_ ( .A(\IF_ID_inst [19] ), .B1(_03050_ ), .B2(_03054_ ), .ZN(_00584_ ) );
OAI221_X1 _16387_ ( .A(_00584_ ), .B1(_03085_ ), .B2(_00438_ ), .C1(_00567_ ), .C2(_03073_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ) );
OAI21_X1 _16388_ ( .A(\IF_ID_inst [18] ), .B1(_03050_ ), .B2(_03054_ ), .ZN(_00585_ ) );
OAI221_X1 _16389_ ( .A(_00585_ ), .B1(_03086_ ), .B2(_00438_ ), .C1(_00567_ ), .C2(_03075_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ) );
OAI21_X1 _16390_ ( .A(\IF_ID_inst [17] ), .B1(_03050_ ), .B2(_03054_ ), .ZN(_00586_ ) );
OAI221_X1 _16391_ ( .A(_00586_ ), .B1(_03087_ ), .B2(_00438_ ), .C1(_00567_ ), .C2(_03076_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ) );
OR2_X1 _16392_ ( .A1(_03124_ ), .A2(_03079_ ), .ZN(_00587_ ) );
OAI221_X1 _16393_ ( .A(_00587_ ), .B1(_03080_ ), .B2(_03055_ ), .C1(_00566_ ), .C2(_03067_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ) );
BUF_X4 _16394_ ( .A(_03802_ ), .Z(_00588_ ) );
AOI21_X1 _16395_ ( .A(\IF_ID_pc [1] ), .B1(_03792_ ), .B2(\IF_ID_pc [2] ), .ZN(_00589_ ) );
INV_X1 _16396_ ( .A(_00589_ ), .ZN(_00590_ ) );
OAI21_X1 _16397_ ( .A(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ), .B1(_03792_ ), .B2(\IF_ID_pc [2] ), .ZN(_00591_ ) );
NOR2_X1 _16398_ ( .A1(_00590_ ), .A2(_00591_ ), .ZN(_00592_ ) );
BUF_X4 _16399_ ( .A(_00592_ ), .Z(_00593_ ) );
NAND2_X1 _16400_ ( .A1(_00507_ ), .A2(_00509_ ), .ZN(_00594_ ) );
OAI211_X1 _16401_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00594_ ), .C2(_03910_ ), .ZN(_00595_ ) );
AND2_X2 _16402_ ( .A1(_03802_ ), .A2(_00592_ ), .ZN(_00596_ ) );
BUF_X4 _16403_ ( .A(_00596_ ), .Z(_00597_ ) );
OAI211_X1 _16404_ ( .A(_00595_ ), .B(\myifu.state [2] ), .C1(_00597_ ), .C2(_03477_ ), .ZN(_00598_ ) );
AND3_X1 _16405_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][8] ), .ZN(_00599_ ) );
AND3_X1 _16406_ ( .A1(_03725_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][8] ), .ZN(_00600_ ) );
AOI211_X1 _16407_ ( .A(_00599_ ), .B(_00600_ ), .C1(\myifu.myicache.data[0][8] ), .C2(_03893_ ), .ZN(_00601_ ) );
NAND2_X1 _16408_ ( .A1(_00557_ ), .A2(\IF_ID_pc [2] ), .ZN(_00602_ ) );
BUF_X2 _16409_ ( .A(_00602_ ), .Z(_00603_ ) );
NAND2_X2 _16410_ ( .A1(\myifu.tmp_offset [2] ), .A2(\myifu.myicache.valid_data_in ), .ZN(_00604_ ) );
BUF_X4 _16411_ ( .A(_00604_ ), .Z(_00605_ ) );
BUF_X4 _16412_ ( .A(_00605_ ), .Z(_00606_ ) );
NAND3_X1 _16413_ ( .A1(_03737_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][8] ), .ZN(_00607_ ) );
NAND4_X1 _16414_ ( .A1(_00601_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00607_ ), .ZN(_00608_ ) );
NOR2_X1 _16415_ ( .A1(\myifu.state [1] ), .A2(\myifu.state [2] ), .ZN(_00609_ ) );
BUF_X4 _16416_ ( .A(_00609_ ), .Z(_00610_ ) );
BUF_X4 _16417_ ( .A(_00610_ ), .Z(_00611_ ) );
BUF_X4 _16418_ ( .A(_03485_ ), .Z(_00612_ ) );
BUF_X4 _16419_ ( .A(_00612_ ), .Z(_00613_ ) );
NAND3_X1 _16420_ ( .A1(_00613_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][8] ), .ZN(_00614_ ) );
NAND3_X1 _16421_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][8] ), .ZN(_00615_ ) );
AND2_X1 _16422_ ( .A1(_00614_ ), .A2(_00615_ ), .ZN(_00616_ ) );
NAND2_X1 _16423_ ( .A1(_00602_ ), .A2(_00604_ ), .ZN(_00617_ ) );
BUF_X2 _16424_ ( .A(_00617_ ), .Z(_00618_ ) );
BUF_X4 _16425_ ( .A(_03736_ ), .Z(_00619_ ) );
NAND3_X1 _16426_ ( .A1(_00619_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][8] ), .ZN(_00620_ ) );
BUF_X4 _16427_ ( .A(_03736_ ), .Z(_00621_ ) );
NAND3_X1 _16428_ ( .A1(_03726_ ), .A2(_00621_ ), .A3(\myifu.myicache.data[1][8] ), .ZN(_00622_ ) );
NAND4_X1 _16429_ ( .A1(_00616_ ), .A2(_00618_ ), .A3(_00620_ ), .A4(_00622_ ), .ZN(_00623_ ) );
NAND3_X1 _16430_ ( .A1(_00608_ ), .A2(_00611_ ), .A3(_00623_ ), .ZN(_00624_ ) );
NAND2_X1 _16431_ ( .A1(_00598_ ), .A2(_00624_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ) );
AND3_X1 _16432_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][31] ), .ZN(_00625_ ) );
CLKBUF_X2 _16433_ ( .A(_03485_ ), .Z(_00626_ ) );
AND3_X1 _16434_ ( .A1(_00626_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][31] ), .ZN(_00627_ ) );
BUF_X4 _16435_ ( .A(_03892_ ), .Z(_00628_ ) );
AOI211_X1 _16436_ ( .A(_00625_ ), .B(_00627_ ), .C1(\myifu.myicache.data[0][31] ), .C2(_00628_ ), .ZN(_00629_ ) );
BUF_X4 _16437_ ( .A(_00602_ ), .Z(_00630_ ) );
BUF_X4 _16438_ ( .A(_03736_ ), .Z(_00631_ ) );
NAND3_X1 _16439_ ( .A1(_00631_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][31] ), .ZN(_00632_ ) );
NAND4_X1 _16440_ ( .A1(_00629_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_00632_ ), .ZN(_00633_ ) );
BUF_X4 _16441_ ( .A(_00612_ ), .Z(_00634_ ) );
NAND3_X1 _16442_ ( .A1(_00634_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][31] ), .ZN(_00635_ ) );
NAND3_X1 _16443_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][31] ), .ZN(_00636_ ) );
AND2_X1 _16444_ ( .A1(_00635_ ), .A2(_00636_ ), .ZN(_00637_ ) );
BUF_X4 _16445_ ( .A(_00617_ ), .Z(_00638_ ) );
BUF_X4 _16446_ ( .A(_00638_ ), .Z(_00639_ ) );
BUF_X4 _16447_ ( .A(_03735_ ), .Z(_00640_ ) );
BUF_X4 _16448_ ( .A(_00640_ ), .Z(_00641_ ) );
NAND3_X1 _16449_ ( .A1(_00641_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][31] ), .ZN(_00642_ ) );
BUF_X4 _16450_ ( .A(_03725_ ), .Z(_00643_ ) );
BUF_X4 _16451_ ( .A(_00640_ ), .Z(_00644_ ) );
NAND3_X1 _16452_ ( .A1(_00643_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][31] ), .ZN(_00645_ ) );
NAND4_X1 _16453_ ( .A1(_00637_ ), .A2(_00639_ ), .A3(_00642_ ), .A4(_00645_ ), .ZN(_00646_ ) );
NAND3_X1 _16454_ ( .A1(_00633_ ), .A2(_00610_ ), .A3(_00646_ ), .ZN(_00647_ ) );
OAI21_X1 _16455_ ( .A(\myifu.state [2] ), .B1(_00597_ ), .B2(_03294_ ), .ZN(_00648_ ) );
NOR4_X1 _16456_ ( .A1(_03803_ ), .A2(\myifu.data_in [31] ), .A3(_00591_ ), .A4(_00590_ ), .ZN(_00649_ ) );
OAI21_X1 _16457_ ( .A(_00647_ ), .B1(_00648_ ), .B2(_00649_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ) );
OR4_X1 _16458_ ( .A1(_03803_ ), .A2(\myifu.data_in [30] ), .A3(_00591_ ), .A4(_00590_ ), .ZN(_00650_ ) );
OAI211_X1 _16459_ ( .A(_00650_ ), .B(\myifu.state [2] ), .C1(_03518_ ), .C2(_00597_ ), .ZN(_00651_ ) );
AND3_X1 _16460_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][30] ), .ZN(_00652_ ) );
CLKBUF_X2 _16461_ ( .A(_03724_ ), .Z(_00653_ ) );
AND3_X1 _16462_ ( .A1(_00653_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][30] ), .ZN(_00654_ ) );
AOI211_X1 _16463_ ( .A(_00652_ ), .B(_00654_ ), .C1(\myifu.myicache.data[0][30] ), .C2(_03893_ ), .ZN(_00655_ ) );
NAND3_X1 _16464_ ( .A1(_03737_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][30] ), .ZN(_00656_ ) );
NAND4_X1 _16465_ ( .A1(_00655_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00656_ ), .ZN(_00657_ ) );
NAND3_X1 _16466_ ( .A1(_00613_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][30] ), .ZN(_00658_ ) );
NAND3_X1 _16467_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][30] ), .ZN(_00659_ ) );
AND2_X1 _16468_ ( .A1(_00658_ ), .A2(_00659_ ), .ZN(_00660_ ) );
NAND3_X1 _16469_ ( .A1(_00619_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][30] ), .ZN(_00661_ ) );
NAND3_X1 _16470_ ( .A1(_03726_ ), .A2(_00621_ ), .A3(\myifu.myicache.data[1][30] ), .ZN(_00662_ ) );
NAND4_X1 _16471_ ( .A1(_00660_ ), .A2(_00618_ ), .A3(_00661_ ), .A4(_00662_ ), .ZN(_00663_ ) );
NAND3_X1 _16472_ ( .A1(_00657_ ), .A2(_00611_ ), .A3(_00663_ ), .ZN(_00664_ ) );
NAND2_X1 _16473_ ( .A1(_00651_ ), .A2(_00664_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ) );
INV_X1 _16474_ ( .A(\myifu.state [2] ), .ZN(_00665_ ) );
BUF_X4 _16475_ ( .A(_00665_ ), .Z(_00666_ ) );
INV_X4 _16476_ ( .A(_00596_ ), .ZN(_00667_ ) );
BUF_X2 _16477_ ( .A(_00667_ ), .Z(_00668_ ) );
AOI21_X1 _16478_ ( .A(_00666_ ), .B1(_00668_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00669_ ) );
OAI211_X1 _16479_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00462_ ), .C2(_03910_ ), .ZN(_00670_ ) );
NAND2_X1 _16480_ ( .A1(_00669_ ), .A2(_00670_ ), .ZN(_00671_ ) );
AND3_X1 _16481_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][21] ), .ZN(_00672_ ) );
AND3_X1 _16482_ ( .A1(_00653_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][21] ), .ZN(_00673_ ) );
AOI211_X1 _16483_ ( .A(_00672_ ), .B(_00673_ ), .C1(\myifu.myicache.data[0][21] ), .C2(_03893_ ), .ZN(_00674_ ) );
NAND3_X1 _16484_ ( .A1(_03737_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][21] ), .ZN(_00675_ ) );
NAND4_X1 _16485_ ( .A1(_00674_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00675_ ), .ZN(_00676_ ) );
NAND3_X1 _16486_ ( .A1(_00613_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][21] ), .ZN(_00677_ ) );
NAND3_X1 _16487_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][21] ), .ZN(_00678_ ) );
AND2_X1 _16488_ ( .A1(_00677_ ), .A2(_00678_ ), .ZN(_00679_ ) );
NAND3_X1 _16489_ ( .A1(_00619_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][21] ), .ZN(_00680_ ) );
NAND3_X1 _16490_ ( .A1(_03726_ ), .A2(_00621_ ), .A3(\myifu.myicache.data[1][21] ), .ZN(_00681_ ) );
NAND4_X1 _16491_ ( .A1(_00679_ ), .A2(_00618_ ), .A3(_00680_ ), .A4(_00681_ ), .ZN(_00682_ ) );
NAND3_X1 _16492_ ( .A1(_00676_ ), .A2(_00611_ ), .A3(_00682_ ), .ZN(_00683_ ) );
NAND2_X1 _16493_ ( .A1(_00671_ ), .A2(_00683_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ) );
NAND2_X1 _16494_ ( .A1(_00463_ ), .A2(_00467_ ), .ZN(_00684_ ) );
OAI211_X1 _16495_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00684_ ), .C2(_03796_ ), .ZN(_00685_ ) );
NAND2_X1 _16496_ ( .A1(_00685_ ), .A2(\myifu.state [2] ), .ZN(_00686_ ) );
BUF_X4 _16497_ ( .A(_00667_ ), .Z(_00687_ ) );
AOI21_X1 _16498_ ( .A(_00686_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00687_ ), .ZN(_00688_ ) );
AND3_X1 _16499_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][20] ), .ZN(_00689_ ) );
AND3_X1 _16500_ ( .A1(_03724_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][20] ), .ZN(_00690_ ) );
AOI211_X1 _16501_ ( .A(_00689_ ), .B(_00690_ ), .C1(\myifu.myicache.data[0][20] ), .C2(_03892_ ), .ZN(_00691_ ) );
NAND3_X1 _16502_ ( .A1(_03736_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][20] ), .ZN(_00692_ ) );
NAND4_X1 _16503_ ( .A1(_00691_ ), .A2(_00602_ ), .A3(_00604_ ), .A4(_00692_ ), .ZN(_00693_ ) );
NAND3_X1 _16504_ ( .A1(_03724_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[3][20] ), .ZN(_00694_ ) );
NAND3_X1 _16505_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[7][20] ), .ZN(_00695_ ) );
AND2_X1 _16506_ ( .A1(_00694_ ), .A2(_00695_ ), .ZN(_00696_ ) );
NAND3_X1 _16507_ ( .A1(_00640_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[5][20] ), .ZN(_00697_ ) );
NAND3_X1 _16508_ ( .A1(_03725_ ), .A2(_00640_ ), .A3(\myifu.myicache.data[1][20] ), .ZN(_00698_ ) );
NAND4_X1 _16509_ ( .A1(_00696_ ), .A2(_00638_ ), .A3(_00697_ ), .A4(_00698_ ), .ZN(_00699_ ) );
AND3_X1 _16510_ ( .A1(_00693_ ), .A2(_00609_ ), .A3(_00699_ ), .ZN(_00700_ ) );
OR2_X1 _16511_ ( .A1(_00688_ ), .A2(_00700_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ) );
AOI21_X1 _16512_ ( .A(_00666_ ), .B1(_00668_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00701_ ) );
NAND2_X1 _16513_ ( .A1(_00468_ ), .A2(_00470_ ), .ZN(_00702_ ) );
OAI21_X1 _16514_ ( .A(_00597_ ), .B1(_03917_ ), .B2(_00702_ ), .ZN(_00703_ ) );
NAND2_X1 _16515_ ( .A1(_00701_ ), .A2(_00703_ ), .ZN(_00704_ ) );
AND3_X1 _16516_ ( .A1(fanout_net_16 ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[6][19] ), .ZN(_00705_ ) );
AND3_X1 _16517_ ( .A1(_00653_ ), .A2(fanout_net_12 ), .A3(\myifu.myicache.data[2][19] ), .ZN(_00706_ ) );
AOI211_X1 _16518_ ( .A(_00705_ ), .B(_00706_ ), .C1(\myifu.myicache.data[0][19] ), .C2(_03893_ ), .ZN(_00707_ ) );
NAND3_X1 _16519_ ( .A1(_03737_ ), .A2(fanout_net_16 ), .A3(\myifu.myicache.data[4][19] ), .ZN(_00708_ ) );
NAND4_X1 _16520_ ( .A1(_00707_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00708_ ), .ZN(_00709_ ) );
NAND3_X1 _16521_ ( .A1(_00613_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][19] ), .ZN(_00710_ ) );
NAND3_X1 _16522_ ( .A1(fanout_net_16 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][19] ), .ZN(_00711_ ) );
AND2_X1 _16523_ ( .A1(_00710_ ), .A2(_00711_ ), .ZN(_00712_ ) );
BUF_X4 _16524_ ( .A(_00638_ ), .Z(_00713_ ) );
NAND3_X1 _16525_ ( .A1(_00619_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][19] ), .ZN(_00714_ ) );
NAND3_X1 _16526_ ( .A1(_03726_ ), .A2(_00621_ ), .A3(\myifu.myicache.data[1][19] ), .ZN(_00715_ ) );
NAND4_X1 _16527_ ( .A1(_00712_ ), .A2(_00713_ ), .A3(_00714_ ), .A4(_00715_ ), .ZN(_00716_ ) );
NAND3_X1 _16528_ ( .A1(_00709_ ), .A2(_00611_ ), .A3(_00716_ ), .ZN(_00717_ ) );
NAND2_X1 _16529_ ( .A1(_00704_ ), .A2(_00717_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ) );
AND3_X1 _16530_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][18] ), .ZN(_00718_ ) );
AND3_X1 _16531_ ( .A1(_00612_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][18] ), .ZN(_00719_ ) );
AOI211_X1 _16532_ ( .A(_00718_ ), .B(_00719_ ), .C1(\myifu.myicache.data[0][18] ), .C2(_00628_ ), .ZN(_00720_ ) );
NAND3_X1 _16533_ ( .A1(_00631_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][18] ), .ZN(_00721_ ) );
NAND4_X1 _16534_ ( .A1(_00720_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_00721_ ), .ZN(_00722_ ) );
NAND3_X1 _16535_ ( .A1(_00634_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][18] ), .ZN(_00723_ ) );
NAND3_X1 _16536_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][18] ), .ZN(_00724_ ) );
AND2_X1 _16537_ ( .A1(_00723_ ), .A2(_00724_ ), .ZN(_00725_ ) );
NAND3_X1 _16538_ ( .A1(_00641_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][18] ), .ZN(_00726_ ) );
NAND3_X1 _16539_ ( .A1(_00643_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][18] ), .ZN(_00727_ ) );
NAND4_X1 _16540_ ( .A1(_00725_ ), .A2(_00639_ ), .A3(_00726_ ), .A4(_00727_ ), .ZN(_00728_ ) );
NAND3_X1 _16541_ ( .A1(_00722_ ), .A2(_00610_ ), .A3(_00728_ ), .ZN(_00729_ ) );
AND2_X1 _16542_ ( .A1(_00668_ ), .A2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00730_ ) );
OAI21_X1 _16543_ ( .A(\myifu.state [2] ), .B1(_00668_ ), .B2(\myifu.data_in [18] ), .ZN(_00731_ ) );
OAI21_X1 _16544_ ( .A(_00729_ ), .B1(_00730_ ), .B2(_00731_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ) );
NAND2_X1 _16545_ ( .A1(_00476_ ), .A2(_00478_ ), .ZN(_00732_ ) );
OAI211_X1 _16546_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00732_ ), .C2(_03796_ ), .ZN(_00733_ ) );
NAND2_X1 _16547_ ( .A1(_00733_ ), .A2(\myifu.state [2] ), .ZN(_00734_ ) );
AOI21_X1 _16548_ ( .A(_00734_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00687_ ), .ZN(_00735_ ) );
AND3_X1 _16549_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][17] ), .ZN(_00736_ ) );
AND3_X1 _16550_ ( .A1(_03724_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][17] ), .ZN(_00737_ ) );
AOI211_X1 _16551_ ( .A(_00736_ ), .B(_00737_ ), .C1(\myifu.myicache.data[0][17] ), .C2(_03892_ ), .ZN(_00738_ ) );
NAND3_X1 _16552_ ( .A1(_03736_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][17] ), .ZN(_00739_ ) );
NAND4_X1 _16553_ ( .A1(_00738_ ), .A2(_00602_ ), .A3(_00604_ ), .A4(_00739_ ), .ZN(_00740_ ) );
NAND3_X1 _16554_ ( .A1(_03724_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][17] ), .ZN(_00741_ ) );
NAND3_X1 _16555_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][17] ), .ZN(_00742_ ) );
AND2_X1 _16556_ ( .A1(_00741_ ), .A2(_00742_ ), .ZN(_00743_ ) );
NAND3_X1 _16557_ ( .A1(_00640_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][17] ), .ZN(_00744_ ) );
NAND3_X1 _16558_ ( .A1(_03725_ ), .A2(_00640_ ), .A3(\myifu.myicache.data[1][17] ), .ZN(_00745_ ) );
NAND4_X1 _16559_ ( .A1(_00743_ ), .A2(_00638_ ), .A3(_00744_ ), .A4(_00745_ ), .ZN(_00746_ ) );
AND3_X1 _16560_ ( .A1(_00740_ ), .A2(_00609_ ), .A3(_00746_ ), .ZN(_00747_ ) );
OR2_X1 _16561_ ( .A1(_00735_ ), .A2(_00747_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ) );
AOI21_X1 _16562_ ( .A(_00666_ ), .B1(_00668_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00748_ ) );
NAND2_X1 _16563_ ( .A1(_00479_ ), .A2(_00481_ ), .ZN(_00749_ ) );
OAI211_X1 _16564_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00749_ ), .C2(_03910_ ), .ZN(_00750_ ) );
NAND2_X1 _16565_ ( .A1(_00748_ ), .A2(_00750_ ), .ZN(_00751_ ) );
AND3_X1 _16566_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][16] ), .ZN(_00752_ ) );
AND3_X1 _16567_ ( .A1(_00653_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][16] ), .ZN(_00753_ ) );
AOI211_X1 _16568_ ( .A(_00752_ ), .B(_00753_ ), .C1(\myifu.myicache.data[0][16] ), .C2(_03893_ ), .ZN(_00754_ ) );
NAND3_X1 _16569_ ( .A1(_03737_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][16] ), .ZN(_00755_ ) );
NAND4_X1 _16570_ ( .A1(_00754_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00755_ ), .ZN(_00756_ ) );
NAND3_X1 _16571_ ( .A1(_00613_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][16] ), .ZN(_00757_ ) );
NAND3_X1 _16572_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][16] ), .ZN(_00758_ ) );
AND2_X1 _16573_ ( .A1(_00757_ ), .A2(_00758_ ), .ZN(_00759_ ) );
NAND3_X1 _16574_ ( .A1(_00619_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][16] ), .ZN(_00760_ ) );
BUF_X4 _16575_ ( .A(_03725_ ), .Z(_00761_ ) );
NAND3_X1 _16576_ ( .A1(_00761_ ), .A2(_00621_ ), .A3(\myifu.myicache.data[1][16] ), .ZN(_00762_ ) );
NAND4_X1 _16577_ ( .A1(_00759_ ), .A2(_00713_ ), .A3(_00760_ ), .A4(_00762_ ), .ZN(_00763_ ) );
NAND3_X1 _16578_ ( .A1(_00756_ ), .A2(_00611_ ), .A3(_00763_ ), .ZN(_00764_ ) );
NAND2_X1 _16579_ ( .A1(_00751_ ), .A2(_00764_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ) );
AOI21_X1 _16580_ ( .A(_00666_ ), .B1(_00668_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00765_ ) );
OAI21_X1 _16581_ ( .A(_00596_ ), .B1(_03917_ ), .B2(_00484_ ), .ZN(_00766_ ) );
NAND2_X1 _16582_ ( .A1(_00765_ ), .A2(_00766_ ), .ZN(_00767_ ) );
AND3_X1 _16583_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][15] ), .ZN(_00768_ ) );
AND3_X1 _16584_ ( .A1(_00653_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][15] ), .ZN(_00769_ ) );
AOI211_X1 _16585_ ( .A(_00768_ ), .B(_00769_ ), .C1(\myifu.myicache.data[0][15] ), .C2(_03893_ ), .ZN(_00770_ ) );
BUF_X4 _16586_ ( .A(_00644_ ), .Z(_00771_ ) );
NAND3_X1 _16587_ ( .A1(_00771_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][15] ), .ZN(_00772_ ) );
NAND4_X1 _16588_ ( .A1(_00770_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00772_ ), .ZN(_00773_ ) );
NAND3_X1 _16589_ ( .A1(_00613_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][15] ), .ZN(_00774_ ) );
NAND3_X1 _16590_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][15] ), .ZN(_00775_ ) );
AND2_X1 _16591_ ( .A1(_00774_ ), .A2(_00775_ ), .ZN(_00776_ ) );
BUF_X4 _16592_ ( .A(_03736_ ), .Z(_00777_ ) );
NAND3_X1 _16593_ ( .A1(_00777_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][15] ), .ZN(_00778_ ) );
NAND3_X1 _16594_ ( .A1(_00761_ ), .A2(_00621_ ), .A3(\myifu.myicache.data[1][15] ), .ZN(_00779_ ) );
NAND4_X1 _16595_ ( .A1(_00776_ ), .A2(_00713_ ), .A3(_00778_ ), .A4(_00779_ ), .ZN(_00780_ ) );
NAND3_X1 _16596_ ( .A1(_00773_ ), .A2(_00611_ ), .A3(_00780_ ), .ZN(_00781_ ) );
NAND2_X1 _16597_ ( .A1(_00767_ ), .A2(_00781_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ) );
AOI21_X1 _16598_ ( .A(_00666_ ), .B1(_00668_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00782_ ) );
OAI211_X1 _16599_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00487_ ), .C2(_03910_ ), .ZN(_00783_ ) );
NAND2_X1 _16600_ ( .A1(_00782_ ), .A2(_00783_ ), .ZN(_00784_ ) );
AND3_X1 _16601_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][14] ), .ZN(_00785_ ) );
AND3_X1 _16602_ ( .A1(_00653_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][14] ), .ZN(_00786_ ) );
BUF_X4 _16603_ ( .A(_03892_ ), .Z(_00787_ ) );
AOI211_X1 _16604_ ( .A(_00785_ ), .B(_00786_ ), .C1(\myifu.myicache.data[0][14] ), .C2(_00787_ ), .ZN(_00788_ ) );
NAND3_X1 _16605_ ( .A1(_00771_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][14] ), .ZN(_00789_ ) );
NAND4_X1 _16606_ ( .A1(_00788_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00789_ ), .ZN(_00790_ ) );
BUF_X4 _16607_ ( .A(_00612_ ), .Z(_00791_ ) );
NAND3_X1 _16608_ ( .A1(_00791_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][14] ), .ZN(_00792_ ) );
NAND3_X1 _16609_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][14] ), .ZN(_00793_ ) );
AND2_X1 _16610_ ( .A1(_00792_ ), .A2(_00793_ ), .ZN(_00794_ ) );
NAND3_X1 _16611_ ( .A1(_00777_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][14] ), .ZN(_00795_ ) );
NAND3_X1 _16612_ ( .A1(_00761_ ), .A2(_00621_ ), .A3(\myifu.myicache.data[1][14] ), .ZN(_00796_ ) );
NAND4_X1 _16613_ ( .A1(_00794_ ), .A2(_00713_ ), .A3(_00795_ ), .A4(_00796_ ), .ZN(_00797_ ) );
NAND3_X1 _16614_ ( .A1(_00790_ ), .A2(_00611_ ), .A3(_00797_ ), .ZN(_00798_ ) );
NAND2_X1 _16615_ ( .A1(_00784_ ), .A2(_00798_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ) );
AOI21_X1 _16616_ ( .A(_00666_ ), .B1(_00668_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00799_ ) );
NAND2_X1 _16617_ ( .A1(_00488_ ), .A2(_00490_ ), .ZN(_00800_ ) );
OAI21_X1 _16618_ ( .A(_00596_ ), .B1(_03917_ ), .B2(_00800_ ), .ZN(_00801_ ) );
NAND2_X1 _16619_ ( .A1(_00799_ ), .A2(_00801_ ), .ZN(_00802_ ) );
AND3_X1 _16620_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][13] ), .ZN(_00803_ ) );
AND3_X1 _16621_ ( .A1(_00653_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][13] ), .ZN(_00804_ ) );
AOI211_X1 _16622_ ( .A(_00803_ ), .B(_00804_ ), .C1(\myifu.myicache.data[0][13] ), .C2(_00787_ ), .ZN(_00805_ ) );
NAND3_X1 _16623_ ( .A1(_00771_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][13] ), .ZN(_00806_ ) );
NAND4_X1 _16624_ ( .A1(_00805_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00806_ ), .ZN(_00807_ ) );
NAND3_X1 _16625_ ( .A1(_00791_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][13] ), .ZN(_00808_ ) );
NAND3_X1 _16626_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][13] ), .ZN(_00809_ ) );
AND2_X1 _16627_ ( .A1(_00808_ ), .A2(_00809_ ), .ZN(_00810_ ) );
NAND3_X1 _16628_ ( .A1(_00777_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][13] ), .ZN(_00811_ ) );
BUF_X4 _16629_ ( .A(_03736_ ), .Z(_00812_ ) );
NAND3_X1 _16630_ ( .A1(_00761_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][13] ), .ZN(_00813_ ) );
NAND4_X1 _16631_ ( .A1(_00810_ ), .A2(_00713_ ), .A3(_00811_ ), .A4(_00813_ ), .ZN(_00814_ ) );
NAND3_X1 _16632_ ( .A1(_00807_ ), .A2(_00611_ ), .A3(_00814_ ), .ZN(_00815_ ) );
NAND2_X1 _16633_ ( .A1(_00802_ ), .A2(_00815_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ) );
AOI21_X1 _16634_ ( .A(_00666_ ), .B1(_00668_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00816_ ) );
NAND2_X1 _16635_ ( .A1(_00491_ ), .A2(_00493_ ), .ZN(_00817_ ) );
OAI211_X1 _16636_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00817_ ), .C2(_03910_ ), .ZN(_00818_ ) );
NAND2_X1 _16637_ ( .A1(_00816_ ), .A2(_00818_ ), .ZN(_00819_ ) );
AND3_X1 _16638_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[6][12] ), .ZN(_00820_ ) );
AND3_X1 _16639_ ( .A1(_00653_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[2][12] ), .ZN(_00821_ ) );
AOI211_X1 _16640_ ( .A(_00820_ ), .B(_00821_ ), .C1(\myifu.myicache.data[0][12] ), .C2(_00787_ ), .ZN(_00822_ ) );
NAND3_X1 _16641_ ( .A1(_00771_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[4][12] ), .ZN(_00823_ ) );
NAND4_X1 _16642_ ( .A1(_00822_ ), .A2(_00603_ ), .A3(_00606_ ), .A4(_00823_ ), .ZN(_00824_ ) );
NAND3_X1 _16643_ ( .A1(_00791_ ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[3][12] ), .ZN(_00825_ ) );
NAND3_X1 _16644_ ( .A1(fanout_net_17 ), .A2(fanout_net_13 ), .A3(\myifu.myicache.data[7][12] ), .ZN(_00826_ ) );
AND2_X1 _16645_ ( .A1(_00825_ ), .A2(_00826_ ), .ZN(_00827_ ) );
NAND3_X1 _16646_ ( .A1(_00777_ ), .A2(fanout_net_17 ), .A3(\myifu.myicache.data[5][12] ), .ZN(_00828_ ) );
NAND3_X1 _16647_ ( .A1(_00761_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][12] ), .ZN(_00829_ ) );
NAND4_X1 _16648_ ( .A1(_00827_ ), .A2(_00713_ ), .A3(_00828_ ), .A4(_00829_ ), .ZN(_00830_ ) );
NAND3_X1 _16649_ ( .A1(_00824_ ), .A2(_00611_ ), .A3(_00830_ ), .ZN(_00831_ ) );
NAND2_X1 _16650_ ( .A1(_00819_ ), .A2(_00831_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ) );
AND3_X1 _16651_ ( .A1(fanout_net_17 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][29] ), .ZN(_00832_ ) );
AND3_X1 _16652_ ( .A1(_00612_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][29] ), .ZN(_00833_ ) );
AOI211_X1 _16653_ ( .A(_00832_ ), .B(_00833_ ), .C1(\myifu.myicache.data[0][29] ), .C2(_00628_ ), .ZN(_00834_ ) );
NAND3_X1 _16654_ ( .A1(_00631_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][29] ), .ZN(_00835_ ) );
NAND4_X1 _16655_ ( .A1(_00834_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_00835_ ), .ZN(_00836_ ) );
NAND3_X1 _16656_ ( .A1(_00634_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][29] ), .ZN(_00837_ ) );
NAND3_X1 _16657_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][29] ), .ZN(_00838_ ) );
AND2_X1 _16658_ ( .A1(_00837_ ), .A2(_00838_ ), .ZN(_00839_ ) );
NAND3_X1 _16659_ ( .A1(_00641_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][29] ), .ZN(_00840_ ) );
NAND3_X1 _16660_ ( .A1(_00643_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][29] ), .ZN(_00841_ ) );
NAND4_X1 _16661_ ( .A1(_00839_ ), .A2(_00639_ ), .A3(_00840_ ), .A4(_00841_ ), .ZN(_00842_ ) );
NAND3_X1 _16662_ ( .A1(_00836_ ), .A2(_00610_ ), .A3(_00842_ ), .ZN(_00843_ ) );
BUF_X4 _16663_ ( .A(_00667_ ), .Z(_00844_ ) );
NOR2_X1 _16664_ ( .A1(_00844_ ), .A2(\myifu.data_in [29] ), .ZN(_00845_ ) );
OAI21_X1 _16665_ ( .A(\myifu.state [2] ), .B1(_00597_ ), .B2(_03456_ ), .ZN(_00846_ ) );
OAI21_X1 _16666_ ( .A(_00843_ ), .B1(_00845_ ), .B2(_00846_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ) );
AND3_X1 _16667_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][11] ), .ZN(_00847_ ) );
AND3_X1 _16668_ ( .A1(_00612_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][11] ), .ZN(_00848_ ) );
AOI211_X1 _16669_ ( .A(_00847_ ), .B(_00848_ ), .C1(\myifu.myicache.data[0][11] ), .C2(_00628_ ), .ZN(_00849_ ) );
NAND3_X1 _16670_ ( .A1(_00631_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][11] ), .ZN(_00850_ ) );
NAND4_X1 _16671_ ( .A1(_00849_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_00850_ ), .ZN(_00851_ ) );
NAND3_X1 _16672_ ( .A1(_00634_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][11] ), .ZN(_00852_ ) );
NAND3_X1 _16673_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][11] ), .ZN(_00853_ ) );
AND2_X1 _16674_ ( .A1(_00852_ ), .A2(_00853_ ), .ZN(_00854_ ) );
NAND3_X1 _16675_ ( .A1(_00641_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][11] ), .ZN(_00855_ ) );
NAND3_X1 _16676_ ( .A1(_00643_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][11] ), .ZN(_00856_ ) );
NAND4_X1 _16677_ ( .A1(_00854_ ), .A2(_00638_ ), .A3(_00855_ ), .A4(_00856_ ), .ZN(_00857_ ) );
NAND3_X1 _16678_ ( .A1(_00851_ ), .A2(_00610_ ), .A3(_00857_ ), .ZN(_00858_ ) );
NOR2_X1 _16679_ ( .A1(_00844_ ), .A2(\myifu.data_in [11] ), .ZN(_00859_ ) );
OAI21_X1 _16680_ ( .A(\myifu.state [2] ), .B1(_00597_ ), .B2(_03461_ ), .ZN(_00860_ ) );
OAI21_X1 _16681_ ( .A(_00858_ ), .B1(_00859_ ), .B2(_00860_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ) );
AND3_X1 _16682_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][10] ), .ZN(_00861_ ) );
AND3_X1 _16683_ ( .A1(_00612_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][10] ), .ZN(_00862_ ) );
AOI211_X1 _16684_ ( .A(_00861_ ), .B(_00862_ ), .C1(\myifu.myicache.data[0][10] ), .C2(_00628_ ), .ZN(_00863_ ) );
NAND3_X1 _16685_ ( .A1(_00631_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][10] ), .ZN(_00864_ ) );
NAND4_X1 _16686_ ( .A1(_00863_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_00864_ ), .ZN(_00865_ ) );
NAND3_X1 _16687_ ( .A1(_00634_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][10] ), .ZN(_00866_ ) );
NAND3_X1 _16688_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][10] ), .ZN(_00867_ ) );
AND2_X1 _16689_ ( .A1(_00866_ ), .A2(_00867_ ), .ZN(_00868_ ) );
NAND3_X1 _16690_ ( .A1(_00641_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][10] ), .ZN(_00869_ ) );
NAND3_X1 _16691_ ( .A1(_00613_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][10] ), .ZN(_00870_ ) );
NAND4_X1 _16692_ ( .A1(_00868_ ), .A2(_00638_ ), .A3(_00869_ ), .A4(_00870_ ), .ZN(_00871_ ) );
NAND3_X1 _16693_ ( .A1(_00865_ ), .A2(_00610_ ), .A3(_00871_ ), .ZN(_00872_ ) );
OAI21_X1 _16694_ ( .A(\myifu.state [2] ), .B1(_00668_ ), .B2(\myifu.data_in [10] ), .ZN(_00873_ ) );
AOI21_X1 _16695_ ( .A(_03466_ ), .B1(_00588_ ), .B2(_00593_ ), .ZN(_00874_ ) );
OAI21_X1 _16696_ ( .A(_00872_ ), .B1(_00873_ ), .B2(_00874_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ) );
NAND2_X1 _16697_ ( .A1(_00504_ ), .A2(_00506_ ), .ZN(_00875_ ) );
OAI211_X1 _16698_ ( .A(_03802_ ), .B(_00592_ ), .C1(_00875_ ), .C2(_03796_ ), .ZN(_00876_ ) );
NAND2_X1 _16699_ ( .A1(_00876_ ), .A2(\myifu.state [2] ), .ZN(_00877_ ) );
AOI21_X1 _16700_ ( .A(_00877_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ), .B2(_00687_ ), .ZN(_00878_ ) );
AND3_X1 _16701_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][9] ), .ZN(_00879_ ) );
AND3_X1 _16702_ ( .A1(_03724_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][9] ), .ZN(_00880_ ) );
AOI211_X1 _16703_ ( .A(_00879_ ), .B(_00880_ ), .C1(\myifu.myicache.data[0][9] ), .C2(_03892_ ), .ZN(_00881_ ) );
NAND3_X1 _16704_ ( .A1(_03736_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][9] ), .ZN(_00882_ ) );
NAND4_X1 _16705_ ( .A1(_00881_ ), .A2(_00602_ ), .A3(_00604_ ), .A4(_00882_ ), .ZN(_00883_ ) );
NAND3_X1 _16706_ ( .A1(_03724_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][9] ), .ZN(_00884_ ) );
NAND3_X1 _16707_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][9] ), .ZN(_00885_ ) );
AND2_X1 _16708_ ( .A1(_00884_ ), .A2(_00885_ ), .ZN(_00886_ ) );
NAND3_X1 _16709_ ( .A1(_00640_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][9] ), .ZN(_00887_ ) );
NAND3_X1 _16710_ ( .A1(_03725_ ), .A2(_00640_ ), .A3(\myifu.myicache.data[1][9] ), .ZN(_00888_ ) );
NAND4_X1 _16711_ ( .A1(_00886_ ), .A2(_00638_ ), .A3(_00887_ ), .A4(_00888_ ), .ZN(_00889_ ) );
AND3_X1 _16712_ ( .A1(_00883_ ), .A2(_00609_ ), .A3(_00889_ ), .ZN(_00890_ ) );
OR2_X1 _16713_ ( .A1(_00878_ ), .A2(_00890_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ) );
AOI21_X1 _16714_ ( .A(_00666_ ), .B1(_00687_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ), .ZN(_00891_ ) );
NAND2_X1 _16715_ ( .A1(_00510_ ), .A2(_00512_ ), .ZN(_00892_ ) );
OAI211_X1 _16716_ ( .A(_00588_ ), .B(_00593_ ), .C1(_00892_ ), .C2(_03910_ ), .ZN(_00893_ ) );
NAND2_X1 _16717_ ( .A1(_00891_ ), .A2(_00893_ ), .ZN(_00894_ ) );
AND3_X1 _16718_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][7] ), .ZN(_00895_ ) );
AND3_X1 _16719_ ( .A1(_00653_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][7] ), .ZN(_00896_ ) );
AOI211_X1 _16720_ ( .A(_00895_ ), .B(_00896_ ), .C1(\myifu.myicache.data[0][7] ), .C2(_00787_ ), .ZN(_00897_ ) );
BUF_X4 _16721_ ( .A(_00630_ ), .Z(_00898_ ) );
BUF_X4 _16722_ ( .A(_00604_ ), .Z(_00899_ ) );
NAND3_X1 _16723_ ( .A1(_00771_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][7] ), .ZN(_00900_ ) );
NAND4_X1 _16724_ ( .A1(_00897_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_00900_ ), .ZN(_00901_ ) );
NAND3_X1 _16725_ ( .A1(_00791_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][7] ), .ZN(_00902_ ) );
NAND3_X1 _16726_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][7] ), .ZN(_00903_ ) );
AND2_X1 _16727_ ( .A1(_00902_ ), .A2(_00903_ ), .ZN(_00904_ ) );
NAND3_X1 _16728_ ( .A1(_00777_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][7] ), .ZN(_00905_ ) );
NAND3_X1 _16729_ ( .A1(_00761_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][7] ), .ZN(_00906_ ) );
NAND4_X1 _16730_ ( .A1(_00904_ ), .A2(_00713_ ), .A3(_00905_ ), .A4(_00906_ ), .ZN(_00907_ ) );
NAND3_X1 _16731_ ( .A1(_00901_ ), .A2(_00611_ ), .A3(_00907_ ), .ZN(_00908_ ) );
NAND2_X1 _16732_ ( .A1(_00894_ ), .A2(_00908_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ) );
AND3_X1 _16733_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][6] ), .ZN(_00909_ ) );
AND3_X1 _16734_ ( .A1(_00612_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][6] ), .ZN(_00910_ ) );
AOI211_X1 _16735_ ( .A(_00909_ ), .B(_00910_ ), .C1(\myifu.myicache.data[0][6] ), .C2(_00628_ ), .ZN(_00911_ ) );
NAND3_X1 _16736_ ( .A1(_00621_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][6] ), .ZN(_00912_ ) );
NAND4_X1 _16737_ ( .A1(_00911_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_00912_ ), .ZN(_00913_ ) );
NAND3_X1 _16738_ ( .A1(_00634_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][6] ), .ZN(_00914_ ) );
NAND3_X1 _16739_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][6] ), .ZN(_00915_ ) );
AND2_X1 _16740_ ( .A1(_00914_ ), .A2(_00915_ ), .ZN(_00916_ ) );
NAND3_X1 _16741_ ( .A1(_00641_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][6] ), .ZN(_00917_ ) );
NAND3_X1 _16742_ ( .A1(_00613_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][6] ), .ZN(_00918_ ) );
NAND4_X1 _16743_ ( .A1(_00916_ ), .A2(_00638_ ), .A3(_00917_ ), .A4(_00918_ ), .ZN(_00919_ ) );
NAND3_X1 _16744_ ( .A1(_00913_ ), .A2(_00610_ ), .A3(_00919_ ), .ZN(_00920_ ) );
NOR2_X1 _16745_ ( .A1(_00844_ ), .A2(\myifu.data_in [6] ), .ZN(_00921_ ) );
OAI21_X1 _16746_ ( .A(\myifu.state [2] ), .B1(_00597_ ), .B2(_03156_ ), .ZN(_00922_ ) );
OAI21_X1 _16747_ ( .A(_00920_ ), .B1(_00921_ ), .B2(_00922_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ) );
AOI21_X2 _16748_ ( .A(_00665_ ), .B1(_00687_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00923_ ) );
OAI21_X1 _16749_ ( .A(_00923_ ), .B1(\myifu.data_in [5] ), .B2(_00844_ ), .ZN(_00924_ ) );
AND3_X1 _16750_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][5] ), .ZN(_00925_ ) );
AND3_X1 _16751_ ( .A1(_00653_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][5] ), .ZN(_00926_ ) );
AOI211_X1 _16752_ ( .A(_00925_ ), .B(_00926_ ), .C1(\myifu.myicache.data[0][5] ), .C2(_00787_ ), .ZN(_00927_ ) );
NAND3_X1 _16753_ ( .A1(_00771_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][5] ), .ZN(_00928_ ) );
NAND4_X1 _16754_ ( .A1(_00927_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_00928_ ), .ZN(_00929_ ) );
BUF_X4 _16755_ ( .A(_00610_ ), .Z(_00930_ ) );
NAND3_X1 _16756_ ( .A1(_00791_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[3][5] ), .ZN(_00931_ ) );
NAND3_X1 _16757_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[7][5] ), .ZN(_00932_ ) );
AND2_X1 _16758_ ( .A1(_00931_ ), .A2(_00932_ ), .ZN(_00933_ ) );
NAND3_X1 _16759_ ( .A1(_00777_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[5][5] ), .ZN(_00934_ ) );
NAND3_X1 _16760_ ( .A1(_00761_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][5] ), .ZN(_00935_ ) );
NAND4_X1 _16761_ ( .A1(_00933_ ), .A2(_00713_ ), .A3(_00934_ ), .A4(_00935_ ), .ZN(_00936_ ) );
NAND3_X1 _16762_ ( .A1(_00929_ ), .A2(_00930_ ), .A3(_00936_ ), .ZN(_00937_ ) );
NAND2_X1 _16763_ ( .A1(_00924_ ), .A2(_00937_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ) );
AOI21_X1 _16764_ ( .A(_00666_ ), .B1(_00687_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00938_ ) );
OAI21_X1 _16765_ ( .A(_00596_ ), .B1(_00497_ ), .B2(_00521_ ), .ZN(_00939_ ) );
NAND2_X1 _16766_ ( .A1(_00938_ ), .A2(_00939_ ), .ZN(_00940_ ) );
AND3_X1 _16767_ ( .A1(fanout_net_18 ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[6][4] ), .ZN(_00941_ ) );
AND3_X1 _16768_ ( .A1(_00626_ ), .A2(fanout_net_14 ), .A3(\myifu.myicache.data[2][4] ), .ZN(_00942_ ) );
AOI211_X1 _16769_ ( .A(_00941_ ), .B(_00942_ ), .C1(\myifu.myicache.data[0][4] ), .C2(_00787_ ), .ZN(_00943_ ) );
NAND3_X1 _16770_ ( .A1(_00771_ ), .A2(fanout_net_18 ), .A3(\myifu.myicache.data[4][4] ), .ZN(_00944_ ) );
NAND4_X1 _16771_ ( .A1(_00943_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_00944_ ), .ZN(_00945_ ) );
NAND3_X1 _16772_ ( .A1(_00791_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][4] ), .ZN(_00946_ ) );
NAND3_X1 _16773_ ( .A1(fanout_net_18 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][4] ), .ZN(_00947_ ) );
AND2_X1 _16774_ ( .A1(_00946_ ), .A2(_00947_ ), .ZN(_00948_ ) );
NAND3_X1 _16775_ ( .A1(_00777_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][4] ), .ZN(_00949_ ) );
NAND3_X1 _16776_ ( .A1(_00761_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][4] ), .ZN(_00950_ ) );
NAND4_X1 _16777_ ( .A1(_00948_ ), .A2(_00713_ ), .A3(_00949_ ), .A4(_00950_ ), .ZN(_00951_ ) );
NAND3_X1 _16778_ ( .A1(_00945_ ), .A2(_00930_ ), .A3(_00951_ ), .ZN(_00952_ ) );
NAND2_X1 _16779_ ( .A1(_00940_ ), .A2(_00952_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ) );
AOI21_X1 _16780_ ( .A(_00665_ ), .B1(_00667_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00953_ ) );
OAI21_X1 _16781_ ( .A(_00953_ ), .B1(\myifu.data_in [3] ), .B2(_00844_ ), .ZN(_00954_ ) );
AND3_X1 _16782_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][3] ), .ZN(_00955_ ) );
AND3_X1 _16783_ ( .A1(_00626_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][3] ), .ZN(_00956_ ) );
AOI211_X1 _16784_ ( .A(_00955_ ), .B(_00956_ ), .C1(\myifu.myicache.data[0][3] ), .C2(_00787_ ), .ZN(_00957_ ) );
NAND3_X1 _16785_ ( .A1(_00771_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][3] ), .ZN(_00958_ ) );
NAND4_X1 _16786_ ( .A1(_00957_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_00958_ ), .ZN(_00959_ ) );
NAND3_X1 _16787_ ( .A1(_00791_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][3] ), .ZN(_00960_ ) );
NAND3_X1 _16788_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][3] ), .ZN(_00961_ ) );
AND2_X1 _16789_ ( .A1(_00960_ ), .A2(_00961_ ), .ZN(_00962_ ) );
NAND3_X1 _16790_ ( .A1(_00777_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][3] ), .ZN(_00963_ ) );
NAND3_X1 _16791_ ( .A1(_00761_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][3] ), .ZN(_00964_ ) );
NAND4_X1 _16792_ ( .A1(_00962_ ), .A2(_00713_ ), .A3(_00963_ ), .A4(_00964_ ), .ZN(_00965_ ) );
NAND3_X1 _16793_ ( .A1(_00959_ ), .A2(_00930_ ), .A3(_00965_ ), .ZN(_00966_ ) );
NAND2_X1 _16794_ ( .A1(_00954_ ), .A2(_00966_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ) );
AOI21_X1 _16795_ ( .A(_00666_ ), .B1(_00687_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00967_ ) );
OAI21_X1 _16796_ ( .A(_00596_ ), .B1(_00497_ ), .B2(_00527_ ), .ZN(_00968_ ) );
NAND2_X1 _16797_ ( .A1(_00967_ ), .A2(_00968_ ), .ZN(_00969_ ) );
AND3_X1 _16798_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][2] ), .ZN(_00970_ ) );
AND3_X1 _16799_ ( .A1(_00626_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][2] ), .ZN(_00971_ ) );
AOI211_X1 _16800_ ( .A(_00970_ ), .B(_00971_ ), .C1(\myifu.myicache.data[0][2] ), .C2(_00787_ ), .ZN(_00972_ ) );
NAND3_X1 _16801_ ( .A1(_00771_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][2] ), .ZN(_00973_ ) );
NAND4_X1 _16802_ ( .A1(_00972_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_00973_ ), .ZN(_00974_ ) );
NAND3_X1 _16803_ ( .A1(_00791_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][2] ), .ZN(_00975_ ) );
NAND3_X1 _16804_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][2] ), .ZN(_00976_ ) );
AND2_X1 _16805_ ( .A1(_00975_ ), .A2(_00976_ ), .ZN(_00977_ ) );
NAND3_X1 _16806_ ( .A1(_00777_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][2] ), .ZN(_00978_ ) );
NAND3_X1 _16807_ ( .A1(_00761_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][2] ), .ZN(_00979_ ) );
NAND4_X1 _16808_ ( .A1(_00977_ ), .A2(_00639_ ), .A3(_00978_ ), .A4(_00979_ ), .ZN(_00980_ ) );
NAND3_X1 _16809_ ( .A1(_00974_ ), .A2(_00930_ ), .A3(_00980_ ), .ZN(_00981_ ) );
NAND2_X1 _16810_ ( .A1(_00969_ ), .A2(_00981_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ) );
AOI21_X1 _16811_ ( .A(_00665_ ), .B1(_00687_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_00982_ ) );
OAI21_X1 _16812_ ( .A(_00596_ ), .B1(_00497_ ), .B2(_00533_ ), .ZN(_00983_ ) );
NAND2_X1 _16813_ ( .A1(_00982_ ), .A2(_00983_ ), .ZN(_00984_ ) );
AND3_X1 _16814_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][1] ), .ZN(_00985_ ) );
AND3_X1 _16815_ ( .A1(_00626_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][1] ), .ZN(_00986_ ) );
AOI211_X1 _16816_ ( .A(_00985_ ), .B(_00986_ ), .C1(\myifu.myicache.data[0][1] ), .C2(_00787_ ), .ZN(_00987_ ) );
NAND3_X1 _16817_ ( .A1(_00771_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][1] ), .ZN(_00988_ ) );
NAND4_X1 _16818_ ( .A1(_00987_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_00988_ ), .ZN(_00989_ ) );
NAND3_X1 _16819_ ( .A1(_00791_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][1] ), .ZN(_00990_ ) );
NAND3_X1 _16820_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][1] ), .ZN(_00991_ ) );
AND2_X1 _16821_ ( .A1(_00990_ ), .A2(_00991_ ), .ZN(_00992_ ) );
NAND3_X1 _16822_ ( .A1(_00777_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][1] ), .ZN(_00993_ ) );
NAND3_X1 _16823_ ( .A1(_00643_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][1] ), .ZN(_00994_ ) );
NAND4_X1 _16824_ ( .A1(_00992_ ), .A2(_00639_ ), .A3(_00993_ ), .A4(_00994_ ), .ZN(_00995_ ) );
NAND3_X1 _16825_ ( .A1(_00989_ ), .A2(_00930_ ), .A3(_00995_ ), .ZN(_00996_ ) );
NAND2_X1 _16826_ ( .A1(_00984_ ), .A2(_00996_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ) );
AOI21_X1 _16827_ ( .A(_00665_ ), .B1(_00667_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ), .ZN(_00997_ ) );
OAI21_X1 _16828_ ( .A(_00997_ ), .B1(\myifu.data_in [28] ), .B2(_00844_ ), .ZN(_00998_ ) );
AND3_X1 _16829_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][28] ), .ZN(_00999_ ) );
AND3_X1 _16830_ ( .A1(_00626_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][28] ), .ZN(_01000_ ) );
AOI211_X1 _16831_ ( .A(_00999_ ), .B(_01000_ ), .C1(\myifu.myicache.data[0][28] ), .C2(_00787_ ), .ZN(_01001_ ) );
NAND3_X1 _16832_ ( .A1(_00619_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][28] ), .ZN(_01002_ ) );
NAND4_X1 _16833_ ( .A1(_01001_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_01002_ ), .ZN(_01003_ ) );
NAND3_X1 _16834_ ( .A1(_00791_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][28] ), .ZN(_01004_ ) );
NAND3_X1 _16835_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][28] ), .ZN(_01005_ ) );
AND2_X1 _16836_ ( .A1(_01004_ ), .A2(_01005_ ), .ZN(_01006_ ) );
NAND3_X1 _16837_ ( .A1(_00631_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][28] ), .ZN(_01007_ ) );
NAND3_X1 _16838_ ( .A1(_00643_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][28] ), .ZN(_01008_ ) );
NAND4_X1 _16839_ ( .A1(_01006_ ), .A2(_00639_ ), .A3(_01007_ ), .A4(_01008_ ), .ZN(_01009_ ) );
NAND3_X1 _16840_ ( .A1(_01003_ ), .A2(_00930_ ), .A3(_01009_ ), .ZN(_01010_ ) );
NAND2_X1 _16841_ ( .A1(_00998_ ), .A2(_01010_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ) );
AOI21_X1 _16842_ ( .A(_00665_ ), .B1(_00687_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01011_ ) );
OAI21_X1 _16843_ ( .A(_00596_ ), .B1(_00497_ ), .B2(_00536_ ), .ZN(_01012_ ) );
NAND2_X1 _16844_ ( .A1(_01011_ ), .A2(_01012_ ), .ZN(_01013_ ) );
AND3_X1 _16845_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][0] ), .ZN(_01014_ ) );
AND3_X1 _16846_ ( .A1(_00626_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][0] ), .ZN(_01015_ ) );
AOI211_X1 _16847_ ( .A(_01014_ ), .B(_01015_ ), .C1(\myifu.myicache.data[0][0] ), .C2(_00628_ ), .ZN(_01016_ ) );
NAND3_X1 _16848_ ( .A1(_00619_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][0] ), .ZN(_01017_ ) );
NAND4_X1 _16849_ ( .A1(_01016_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_01017_ ), .ZN(_01018_ ) );
NAND3_X1 _16850_ ( .A1(_00634_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][0] ), .ZN(_01019_ ) );
NAND3_X1 _16851_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][0] ), .ZN(_01020_ ) );
AND2_X1 _16852_ ( .A1(_01019_ ), .A2(_01020_ ), .ZN(_01021_ ) );
NAND3_X1 _16853_ ( .A1(_00631_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][0] ), .ZN(_01022_ ) );
NAND3_X1 _16854_ ( .A1(_00643_ ), .A2(_00812_ ), .A3(\myifu.myicache.data[1][0] ), .ZN(_01023_ ) );
NAND4_X1 _16855_ ( .A1(_01021_ ), .A2(_00639_ ), .A3(_01022_ ), .A4(_01023_ ), .ZN(_01024_ ) );
NAND3_X1 _16856_ ( .A1(_01018_ ), .A2(_00930_ ), .A3(_01024_ ), .ZN(_01025_ ) );
NAND2_X1 _16857_ ( .A1(_01013_ ), .A2(_01025_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ) );
AND2_X1 _16858_ ( .A1(_00538_ ), .A2(_00539_ ), .ZN(_01026_ ) );
OAI211_X1 _16859_ ( .A(_00588_ ), .B(_00593_ ), .C1(_03910_ ), .C2(_01026_ ), .ZN(_01027_ ) );
OAI211_X1 _16860_ ( .A(_01027_ ), .B(\myifu.state [2] ), .C1(_00597_ ), .C2(_03501_ ), .ZN(_01028_ ) );
AND3_X1 _16861_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][27] ), .ZN(_01029_ ) );
AND3_X1 _16862_ ( .A1(_00626_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][27] ), .ZN(_01030_ ) );
AOI211_X1 _16863_ ( .A(_01029_ ), .B(_01030_ ), .C1(\myifu.myicache.data[0][27] ), .C2(_00628_ ), .ZN(_01031_ ) );
NAND3_X1 _16864_ ( .A1(_00619_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][27] ), .ZN(_01032_ ) );
NAND4_X1 _16865_ ( .A1(_01031_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_01032_ ), .ZN(_01033_ ) );
NAND3_X1 _16866_ ( .A1(_00634_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][27] ), .ZN(_01034_ ) );
NAND3_X1 _16867_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][27] ), .ZN(_01035_ ) );
AND2_X1 _16868_ ( .A1(_01034_ ), .A2(_01035_ ), .ZN(_01036_ ) );
NAND3_X1 _16869_ ( .A1(_00631_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][27] ), .ZN(_01037_ ) );
NAND3_X1 _16870_ ( .A1(_00643_ ), .A2(_00641_ ), .A3(\myifu.myicache.data[1][27] ), .ZN(_01038_ ) );
NAND4_X1 _16871_ ( .A1(_01036_ ), .A2(_00639_ ), .A3(_01037_ ), .A4(_01038_ ), .ZN(_01039_ ) );
NAND3_X1 _16872_ ( .A1(_01033_ ), .A2(_00930_ ), .A3(_01039_ ), .ZN(_01040_ ) );
NAND2_X1 _16873_ ( .A1(_01028_ ), .A2(_01040_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ) );
AND3_X1 _16874_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[6][26] ), .ZN(_01041_ ) );
AND3_X1 _16875_ ( .A1(_00612_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[2][26] ), .ZN(_01042_ ) );
AOI211_X1 _16876_ ( .A(_01041_ ), .B(_01042_ ), .C1(\myifu.myicache.data[0][26] ), .C2(_03892_ ), .ZN(_01043_ ) );
NAND3_X1 _16877_ ( .A1(_00621_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[4][26] ), .ZN(_01044_ ) );
NAND4_X1 _16878_ ( .A1(_01043_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_01044_ ), .ZN(_01045_ ) );
NAND3_X1 _16879_ ( .A1(_03725_ ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[3][26] ), .ZN(_01046_ ) );
NAND3_X1 _16880_ ( .A1(fanout_net_19 ), .A2(fanout_net_15 ), .A3(\myifu.myicache.data[7][26] ), .ZN(_01047_ ) );
AND2_X1 _16881_ ( .A1(_01046_ ), .A2(_01047_ ), .ZN(_01048_ ) );
NAND3_X1 _16882_ ( .A1(_00641_ ), .A2(fanout_net_19 ), .A3(\myifu.myicache.data[5][26] ), .ZN(_01049_ ) );
NAND3_X1 _16883_ ( .A1(_00613_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][26] ), .ZN(_01050_ ) );
NAND4_X1 _16884_ ( .A1(_01048_ ), .A2(_00638_ ), .A3(_01049_ ), .A4(_01050_ ), .ZN(_01051_ ) );
NAND3_X1 _16885_ ( .A1(_01045_ ), .A2(_00610_ ), .A3(_01051_ ), .ZN(_01052_ ) );
NOR2_X1 _16886_ ( .A1(_00844_ ), .A2(\myifu.data_in [26] ), .ZN(_01053_ ) );
OAI21_X1 _16887_ ( .A(\myifu.state [2] ), .B1(_00597_ ), .B2(_03498_ ), .ZN(_01054_ ) );
OAI21_X1 _16888_ ( .A(_01052_ ), .B1(_01053_ ), .B2(_01054_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ) );
AND3_X1 _16889_ ( .A1(fanout_net_19 ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][25] ), .ZN(_01055_ ) );
AND3_X1 _16890_ ( .A1(_00612_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][25] ), .ZN(_01056_ ) );
AOI211_X1 _16891_ ( .A(_01055_ ), .B(_01056_ ), .C1(\myifu.myicache.data[0][25] ), .C2(_03892_ ), .ZN(_01057_ ) );
NAND3_X1 _16892_ ( .A1(_00621_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][25] ), .ZN(_01058_ ) );
NAND4_X1 _16893_ ( .A1(_01057_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_01058_ ), .ZN(_01059_ ) );
NAND3_X1 _16894_ ( .A1(_03725_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][25] ), .ZN(_01060_ ) );
NAND3_X1 _16895_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][25] ), .ZN(_01061_ ) );
AND2_X1 _16896_ ( .A1(_01060_ ), .A2(_01061_ ), .ZN(_01062_ ) );
NAND3_X1 _16897_ ( .A1(_00644_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][25] ), .ZN(_01063_ ) );
NAND3_X1 _16898_ ( .A1(_00613_ ), .A2(_00644_ ), .A3(\myifu.myicache.data[1][25] ), .ZN(_01064_ ) );
NAND4_X1 _16899_ ( .A1(_01062_ ), .A2(_00638_ ), .A3(_01063_ ), .A4(_01064_ ), .ZN(_01065_ ) );
NAND3_X1 _16900_ ( .A1(_01059_ ), .A2(_00610_ ), .A3(_01065_ ), .ZN(_01066_ ) );
NOR2_X1 _16901_ ( .A1(_00844_ ), .A2(\myifu.data_in [25] ), .ZN(_01067_ ) );
OAI21_X1 _16902_ ( .A(\myifu.state [2] ), .B1(_00597_ ), .B2(_03489_ ), .ZN(_01068_ ) );
OAI21_X1 _16903_ ( .A(_01066_ ), .B1(_01067_ ), .B2(_01068_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ) );
AND2_X1 _16904_ ( .A1(_00546_ ), .A2(_00548_ ), .ZN(_01069_ ) );
OAI211_X1 _16905_ ( .A(_03802_ ), .B(_00592_ ), .C1(_03796_ ), .C2(_01069_ ), .ZN(_01070_ ) );
NAND2_X1 _16906_ ( .A1(_01070_ ), .A2(\myifu.state [2] ), .ZN(_01071_ ) );
AOI21_X1 _16907_ ( .A(_01071_ ), .B1(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .B2(_00687_ ), .ZN(_01072_ ) );
AND3_X1 _16908_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][24] ), .ZN(_01073_ ) );
AND3_X1 _16909_ ( .A1(_03724_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][24] ), .ZN(_01074_ ) );
AOI211_X1 _16910_ ( .A(_01073_ ), .B(_01074_ ), .C1(\myifu.myicache.data[0][24] ), .C2(_03892_ ), .ZN(_01075_ ) );
NAND3_X1 _16911_ ( .A1(_03736_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][24] ), .ZN(_01076_ ) );
NAND4_X1 _16912_ ( .A1(_01075_ ), .A2(_00602_ ), .A3(_00604_ ), .A4(_01076_ ), .ZN(_01077_ ) );
NAND3_X1 _16913_ ( .A1(_03724_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][24] ), .ZN(_01078_ ) );
NAND3_X1 _16914_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][24] ), .ZN(_01079_ ) );
AND2_X1 _16915_ ( .A1(_01078_ ), .A2(_01079_ ), .ZN(_01080_ ) );
NAND3_X1 _16916_ ( .A1(_00640_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][24] ), .ZN(_01081_ ) );
NAND3_X1 _16917_ ( .A1(_03725_ ), .A2(_00640_ ), .A3(\myifu.myicache.data[1][24] ), .ZN(_01082_ ) );
NAND4_X1 _16918_ ( .A1(_01080_ ), .A2(_00617_ ), .A3(_01081_ ), .A4(_01082_ ), .ZN(_01083_ ) );
AND3_X1 _16919_ ( .A1(_01077_ ), .A2(_00609_ ), .A3(_01083_ ), .ZN(_01084_ ) );
OR2_X1 _16920_ ( .A1(_01072_ ), .A2(_01084_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ) );
AOI21_X1 _16921_ ( .A(_00665_ ), .B1(_00667_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ), .ZN(_01085_ ) );
OAI21_X1 _16922_ ( .A(_01085_ ), .B1(\myifu.data_in [23] ), .B2(_00844_ ), .ZN(_01086_ ) );
AND3_X1 _16923_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][23] ), .ZN(_01087_ ) );
AND3_X1 _16924_ ( .A1(_00626_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][23] ), .ZN(_01088_ ) );
AOI211_X1 _16925_ ( .A(_01087_ ), .B(_01088_ ), .C1(\myifu.myicache.data[0][23] ), .C2(_00628_ ), .ZN(_01089_ ) );
NAND3_X1 _16926_ ( .A1(_00619_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][23] ), .ZN(_01090_ ) );
NAND4_X1 _16927_ ( .A1(_01089_ ), .A2(_00898_ ), .A3(_00899_ ), .A4(_01090_ ), .ZN(_01091_ ) );
NAND3_X1 _16928_ ( .A1(_00634_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][23] ), .ZN(_01092_ ) );
NAND3_X1 _16929_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][23] ), .ZN(_01093_ ) );
AND2_X1 _16930_ ( .A1(_01092_ ), .A2(_01093_ ), .ZN(_01094_ ) );
NAND3_X1 _16931_ ( .A1(_00631_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][23] ), .ZN(_01095_ ) );
NAND3_X1 _16932_ ( .A1(_00643_ ), .A2(_00641_ ), .A3(\myifu.myicache.data[1][23] ), .ZN(_01096_ ) );
NAND4_X1 _16933_ ( .A1(_01094_ ), .A2(_00639_ ), .A3(_01095_ ), .A4(_01096_ ), .ZN(_01097_ ) );
NAND3_X1 _16934_ ( .A1(_01091_ ), .A2(_00930_ ), .A3(_01097_ ), .ZN(_01098_ ) );
NAND2_X1 _16935_ ( .A1(_01086_ ), .A2(_01098_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ) );
AOI21_X1 _16936_ ( .A(_00665_ ), .B1(_00667_ ), .B2(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ), .ZN(_01099_ ) );
OAI21_X1 _16937_ ( .A(_01099_ ), .B1(\myifu.data_in [22] ), .B2(_00844_ ), .ZN(_01100_ ) );
AND3_X1 _16938_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[6][22] ), .ZN(_01101_ ) );
AND3_X1 _16939_ ( .A1(_00626_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[2][22] ), .ZN(_01102_ ) );
AOI211_X1 _16940_ ( .A(_01101_ ), .B(_01102_ ), .C1(\myifu.myicache.data[0][22] ), .C2(_00628_ ), .ZN(_01103_ ) );
NAND3_X1 _16941_ ( .A1(_00619_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[4][22] ), .ZN(_01104_ ) );
NAND4_X1 _16942_ ( .A1(_01103_ ), .A2(_00630_ ), .A3(_00605_ ), .A4(_01104_ ), .ZN(_01105_ ) );
NAND3_X1 _16943_ ( .A1(_00634_ ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[3][22] ), .ZN(_01106_ ) );
NAND3_X1 _16944_ ( .A1(\IF_ID_pc [4] ), .A2(\IF_ID_pc [3] ), .A3(\myifu.myicache.data[7][22] ), .ZN(_01107_ ) );
AND2_X1 _16945_ ( .A1(_01106_ ), .A2(_01107_ ), .ZN(_01108_ ) );
NAND3_X1 _16946_ ( .A1(_00631_ ), .A2(\IF_ID_pc [4] ), .A3(\myifu.myicache.data[5][22] ), .ZN(_01109_ ) );
NAND3_X1 _16947_ ( .A1(_00643_ ), .A2(_00641_ ), .A3(\myifu.myicache.data[1][22] ), .ZN(_01110_ ) );
NAND4_X1 _16948_ ( .A1(_01108_ ), .A2(_00639_ ), .A3(_01109_ ), .A4(_01110_ ), .ZN(_01111_ ) );
NAND3_X1 _16949_ ( .A1(_01105_ ), .A2(_00930_ ), .A3(_01111_ ), .ZN(_01112_ ) );
NAND2_X1 _16950_ ( .A1(_01100_ ), .A2(_01112_ ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ) );
AOI211_X1 _16951_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_03275_ ), .C1(_03640_ ), .C2(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ), .ZN(\myifu.pc_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16952_ ( .A(_03804_ ), .ZN(_01113_ ) );
NAND4_X1 _16953_ ( .A1(_03795_ ), .A2(\myifu.state [2] ), .A3(_01113_ ), .A4(_03801_ ), .ZN(_01114_ ) );
AND2_X1 _16954_ ( .A1(_01928_ ), .A2(_01894_ ), .ZN(_01115_ ) );
AND3_X1 _16955_ ( .A1(_01115_ ), .A2(_01834_ ), .A3(\myifu.state [0] ), .ZN(_01116_ ) );
INV_X1 _16956_ ( .A(\myidu.stall_quest_fencei ), .ZN(_01117_ ) );
AOI21_X1 _16957_ ( .A(_00449_ ), .B1(_01116_ ), .B2(_01117_ ), .ZN(_01118_ ) );
AOI21_X1 _16958_ ( .A(reset ), .B1(_01114_ ), .B2(_01118_ ), .ZN(\myifu.state_$_DFF_P__Q_1_D ) );
NOR2_X1 _16959_ ( .A1(_03872_ ), .A2(_03796_ ), .ZN(_01119_ ) );
INV_X1 _16960_ ( .A(_01119_ ), .ZN(_01120_ ) );
AND3_X1 _16961_ ( .A1(_01120_ ), .A2(_01117_ ), .A3(_01930_ ), .ZN(_01121_ ) );
AND2_X1 _16962_ ( .A1(\myidu.stall_quest_fencei ), .A2(\myifu.state [0] ), .ZN(_01122_ ) );
OR4_X1 _16963_ ( .A1(reset ), .A2(_01121_ ), .A3(\myifu.pc_$_SDFFE_PP1P__Q_E ), .A4(_01122_ ), .ZN(\myifu.state_$_DFF_P__Q_2_D ) );
OAI211_X1 _16964_ ( .A(_01626_ ), .B(\myifu.state [2] ), .C1(_03803_ ), .C2(_03804_ ), .ZN(_01123_ ) );
NAND2_X1 _16965_ ( .A1(_01119_ ), .A2(_02050_ ), .ZN(_01124_ ) );
NAND2_X1 _16966_ ( .A1(_01123_ ), .A2(_01124_ ), .ZN(\myifu.state_$_DFF_P__Q_D ) );
AND3_X1 _16967_ ( .A1(_03795_ ), .A2(\myifu.state [2] ), .A3(_03801_ ), .ZN(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ) );
AOI21_X1 _16968_ ( .A(_02078_ ), .B1(_02047_ ), .B2(_02085_ ), .ZN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_B_$_MUX__Y_A_$_NOR__B_Y ) );
INV_X1 _16969_ ( .A(\myifu.wen_$_ANDNOT__A_Y ), .ZN(_01125_ ) );
NOR3_X1 _16970_ ( .A1(_01125_ ), .A2(_00559_ ), .A3(_00618_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND4_X1 _16971_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_03893_ ), .A3(_00603_ ), .A4(_00606_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ) );
AND4_X1 _16972_ ( .A1(_03726_ ), .A2(\myifu.wen_$_ANDNOT__A_Y ), .A3(\IF_ID_pc [3] ), .A4(_00618_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _16973_ ( .A1(\IF_ID_pc [4] ), .A2(_03891_ ), .A3(\IF_ID_pc [3] ), .A4(_00618_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ) );
NOR3_X1 _16974_ ( .A1(_01125_ ), .A2(_00558_ ), .A3(_00618_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ) );
NOR3_X1 _16975_ ( .A1(_01125_ ), .A2(_00556_ ), .A3(_00618_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ) );
AND3_X1 _16976_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_03893_ ), .A3(_00618_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _16977_ ( .A1(\IF_ID_pc [4] ), .A2(_03891_ ), .A3(_03737_ ), .A4(_00618_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ) );
AND3_X1 _16978_ ( .A1(_02049_ ), .A2(_03893_ ), .A3(\myifu.myicache.valid_data_in ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ) );
AND3_X1 _16979_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(_03726_ ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ) );
AND3_X1 _16980_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(\IF_ID_pc [3] ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ) );
AND3_X1 _16981_ ( .A1(\myifu.wen_$_ANDNOT__A_Y ), .A2(\IF_ID_pc [4] ), .A3(_03737_ ), .ZN(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ) );
NAND3_X1 _16982_ ( .A1(_01115_ ), .A2(_01834_ ), .A3(\myifu.state [0] ), .ZN(_01126_ ) );
AND2_X1 _16983_ ( .A1(_00451_ ), .A2(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ), .ZN(_01127_ ) );
NOR4_X1 _16984_ ( .A1(_01127_ ), .A2(_03276_ ), .A3(_00449_ ), .A4(_01122_ ), .ZN(_01128_ ) );
NAND2_X1 _16985_ ( .A1(_01126_ ), .A2(_01128_ ), .ZN(_01129_ ) );
AND2_X1 _16986_ ( .A1(_03802_ ), .A2(_01113_ ), .ZN(_01130_ ) );
INV_X1 _16987_ ( .A(_01130_ ), .ZN(_01131_ ) );
AOI221_X4 _16988_ ( .A(_01129_ ), .B1(\myifu.state [0] ), .B2(_01120_ ), .C1(_01131_ ), .C2(_01931_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E ) );
AOI211_X1 _16989_ ( .A(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ), .B(_03277_ ), .C1(_03273_ ), .C2(check_quest ), .ZN(\myidu.typ_$_SDFFE_PP0P__Q_E ) );
AOI211_X1 _16990_ ( .A(_00420_ ), .B(_00422_ ), .C1(_03056_ ), .C2(_03366_ ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ) );
OR4_X1 _16991_ ( .A1(reset ), .A2(_01127_ ), .A3(_00449_ ), .A4(_01122_ ), .ZN(_01132_ ) );
AOI211_X1 _16992_ ( .A(_03276_ ), .B(_01132_ ), .C1(_01929_ ), .C2(\myifu.state [0] ), .ZN(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
MUX2_X1 _16993_ ( .A(_03958_ ), .B(_01941_ ), .S(\mylsu.state [0] ), .Z(_01133_ ) );
NOR2_X1 _16994_ ( .A1(_03964_ ), .A2(_01133_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ) );
INV_X1 _16995_ ( .A(_03810_ ), .ZN(_01134_ ) );
NOR3_X1 _16996_ ( .A1(_03964_ ), .A2(_01134_ ), .A3(_01133_ ), .ZN(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ) );
NAND2_X1 _16997_ ( .A1(_03809_ ), .A2(_03884_ ), .ZN(_01135_ ) );
NOR2_X1 _16998_ ( .A1(_02074_ ), .A2(_01135_ ), .ZN(_01136_ ) );
NAND4_X1 _16999_ ( .A1(_03875_ ), .A2(_02017_ ), .A3(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A4(_01136_ ), .ZN(_01137_ ) );
AND2_X1 _17000_ ( .A1(_03795_ ), .A2(_03963_ ), .ZN(_01138_ ) );
OAI21_X1 _17001_ ( .A(_01137_ ), .B1(_01138_ ), .B2(_03886_ ), .ZN(\mylsu.state_$_DFF_P__Q_1_D ) );
AND2_X1 _17002_ ( .A1(io_master_awready ), .A2(io_master_wready ), .ZN(_01139_ ) );
AOI21_X1 _17003_ ( .A(_01139_ ), .B1(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .B2(_02152_ ), .ZN(_01140_ ) );
NAND4_X1 _17004_ ( .A1(_03857_ ), .A2(\mylsu.state [0] ), .A3(io_master_awready ), .A4(_01140_ ), .ZN(_01141_ ) );
NOR4_X1 _17005_ ( .A1(_02038_ ), .A2(_02037_ ), .A3(_02045_ ), .A4(_01141_ ), .ZN(_01142_ ) );
AND3_X1 _17006_ ( .A1(_03810_ ), .A2(\mylsu.state [2] ), .A3(_04017_ ), .ZN(_01143_ ) );
OR2_X1 _17007_ ( .A1(_01142_ ), .A2(_01143_ ), .ZN(\mylsu.state_$_DFF_P__Q_2_D ) );
AND4_X1 _17008_ ( .A1(EXU_valid_LSU ), .A2(_03884_ ), .A3(_02036_ ), .A4(_01139_ ), .ZN(_01144_ ) );
NAND4_X1 _17009_ ( .A1(_02046_ ), .A2(\mylsu.state [0] ), .A3(_03810_ ), .A4(_01144_ ), .ZN(_01145_ ) );
NAND4_X1 _17010_ ( .A1(fanout_net_5 ), .A2(_01458_ ), .A3(\mylsu.state [4] ), .A4(io_master_awready ), .ZN(_01146_ ) );
NAND4_X1 _17011_ ( .A1(fanout_net_5 ), .A2(_01457_ ), .A3(\mylsu.state [2] ), .A4(io_master_wready ), .ZN(_01147_ ) );
NAND3_X1 _17012_ ( .A1(_03969_ ), .A2(_03810_ ), .A3(\mylsu.state [1] ), .ZN(_01148_ ) );
NAND4_X1 _17013_ ( .A1(_01145_ ), .A2(_01146_ ), .A3(_01147_ ), .A4(_01148_ ), .ZN(\mylsu.state_$_DFF_P__Q_3_D ) );
NAND3_X1 _17014_ ( .A1(_03795_ ), .A2(_00205_ ), .A3(_03963_ ), .ZN(_01149_ ) );
AND3_X1 _17015_ ( .A1(_03966_ ), .A2(\mylsu.state [1] ), .A3(_03968_ ), .ZN(_01150_ ) );
NAND3_X1 _17016_ ( .A1(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .A2(_02152_ ), .A3(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_01151_ ) );
OAI211_X1 _17017_ ( .A(_03810_ ), .B(_01151_ ), .C1(_00418_ ), .C2(EXU_valid_LSU ), .ZN(_01152_ ) );
AND4_X1 _17018_ ( .A1(_02036_ ), .A2(_03810_ ), .A3(_03884_ ), .A4(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .ZN(_01153_ ) );
AOI211_X1 _17019_ ( .A(_01150_ ), .B(_01152_ ), .C1(_02045_ ), .C2(_01153_ ), .ZN(_01154_ ) );
OR4_X1 _17020_ ( .A1(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .A2(_00417_ ), .A3(_02074_ ), .A4(_01135_ ), .ZN(_01155_ ) );
INV_X1 _17021_ ( .A(_01155_ ), .ZN(_01156_ ) );
OR4_X1 _17022_ ( .A1(\EX_LS_dest_csreg_mem [28] ), .A2(_02032_ ), .A3(_02018_ ), .A4(_02015_ ), .ZN(_01157_ ) );
OAI21_X1 _17023_ ( .A(_01157_ ), .B1(_02017_ ), .B2(_02036_ ), .ZN(_01158_ ) );
AND3_X1 _17024_ ( .A1(_01158_ ), .A2(_03884_ ), .A3(_03857_ ), .ZN(_01159_ ) );
NAND3_X1 _17025_ ( .A1(_02032_ ), .A2(_03884_ ), .A3(_03857_ ), .ZN(_01160_ ) );
NOR4_X1 _17026_ ( .A1(_02016_ ), .A2(_01941_ ), .A3(_02037_ ), .A4(_01135_ ), .ZN(_01161_ ) );
NAND2_X1 _17027_ ( .A1(_01161_ ), .A2(_03883_ ), .ZN(_01162_ ) );
AND4_X1 _17028_ ( .A1(_04016_ ), .A2(_03811_ ), .A3(_04017_ ), .A4(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ), .ZN(_01163_ ) );
NAND4_X1 _17029_ ( .A1(_01163_ ), .A2(_03810_ ), .A3(_03856_ ), .A4(_01140_ ), .ZN(_01164_ ) );
OAI211_X1 _17030_ ( .A(_01160_ ), .B(_01162_ ), .C1(_02075_ ), .C2(_01164_ ), .ZN(_01165_ ) );
NOR3_X1 _17031_ ( .A1(_01156_ ), .A2(_01159_ ), .A3(_01165_ ), .ZN(_01166_ ) );
OAI211_X1 _17032_ ( .A(_01149_ ), .B(_01154_ ), .C1(_01166_ ), .C2(_00418_ ), .ZN(\mylsu.state_$_DFF_P__Q_4_D ) );
NAND4_X1 _17033_ ( .A1(_02046_ ), .A2(io_master_wready ), .A3(_03948_ ), .A4(_01140_ ), .ZN(_01167_ ) );
AOI211_X1 _17034_ ( .A(io_master_awready ), .B(_01134_ ), .C1(_01167_ ), .C2(_03954_ ), .ZN(\mylsu.state_$_DFF_P__Q_D ) );
NAND2_X1 _17035_ ( .A1(\EX_LS_flag [2] ), .A2(\EX_LS_result_csreg_mem [21] ), .ZN(_01168_ ) );
OAI21_X1 _17036_ ( .A(_01168_ ), .B1(_03824_ ), .B2(_02070_ ), .ZN(_01169_ ) );
MUX2_X1 _17037_ ( .A(_01169_ ), .B(\EX_LS_pc [21] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ) );
BUF_X4 _17038_ ( .A(_03817_ ), .Z(_01170_ ) );
AOI21_X1 _17039_ ( .A(\EX_LS_pc [20] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01171_ ) );
BUF_X4 _17040_ ( .A(_03823_ ), .Z(_01172_ ) );
MUX2_X1 _17041_ ( .A(\LS_WB_wdata_csreg [20] ), .B(\EX_LS_result_csreg_mem [20] ), .S(_01172_ ), .Z(_01173_ ) );
NOR3_X1 _17042_ ( .A1(_03813_ ), .A2(_03818_ ), .A3(_01173_ ), .ZN(_01174_ ) );
NOR2_X1 _17043_ ( .A1(_01171_ ), .A2(_01174_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ) );
MUX2_X1 _17044_ ( .A(\LS_WB_wdata_csreg [19] ), .B(\EX_LS_result_csreg_mem [19] ), .S(_03824_ ), .Z(_01175_ ) );
MUX2_X1 _17045_ ( .A(_01175_ ), .B(\EX_LS_pc [19] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ) );
MUX2_X1 _17046_ ( .A(\LS_WB_wdata_csreg [18] ), .B(\EX_LS_result_csreg_mem [18] ), .S(_03824_ ), .Z(_01176_ ) );
MUX2_X1 _17047_ ( .A(_01176_ ), .B(\EX_LS_pc [18] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ) );
AOI221_X4 _17048_ ( .A(_03819_ ), .B1(\LS_WB_wdata_csreg [17] ), .B2(_01945_ ), .C1(\EX_LS_result_csreg_mem [17] ), .C2(_03824_ ), .ZN(_01177_ ) );
AOI21_X1 _17049_ ( .A(\EX_LS_pc [17] ), .B1(_03868_ ), .B2(_01170_ ), .ZN(_01178_ ) );
NOR2_X1 _17050_ ( .A1(_01177_ ), .A2(_01178_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ) );
BUF_X4 _17051_ ( .A(_03823_ ), .Z(_01179_ ) );
MUX2_X1 _17052_ ( .A(\LS_WB_wdata_csreg [16] ), .B(\EX_LS_result_csreg_mem [16] ), .S(_01179_ ), .Z(_01180_ ) );
MUX2_X1 _17053_ ( .A(_01180_ ), .B(\EX_LS_pc [16] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ) );
MUX2_X1 _17054_ ( .A(\LS_WB_wdata_csreg [15] ), .B(\EX_LS_result_csreg_mem [15] ), .S(_01179_ ), .Z(_01181_ ) );
MUX2_X1 _17055_ ( .A(_01181_ ), .B(\EX_LS_pc [15] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ) );
AOI21_X1 _17056_ ( .A(\EX_LS_pc [14] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01182_ ) );
MUX2_X1 _17057_ ( .A(\LS_WB_wdata_csreg [14] ), .B(\EX_LS_result_csreg_mem [14] ), .S(_01172_ ), .Z(_01183_ ) );
NOR3_X1 _17058_ ( .A1(_03813_ ), .A2(_03818_ ), .A3(_01183_ ), .ZN(_01184_ ) );
NOR2_X1 _17059_ ( .A1(_01182_ ), .A2(_01184_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ) );
MUX2_X1 _17060_ ( .A(\LS_WB_wdata_csreg [13] ), .B(\EX_LS_result_csreg_mem [13] ), .S(_01179_ ), .Z(_01185_ ) );
MUX2_X1 _17061_ ( .A(_01185_ ), .B(\EX_LS_pc [13] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ) );
MUX2_X1 _17062_ ( .A(\LS_WB_wdata_csreg [12] ), .B(\EX_LS_result_csreg_mem [12] ), .S(_01179_ ), .Z(_01186_ ) );
MUX2_X1 _17063_ ( .A(_01186_ ), .B(\EX_LS_pc [12] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ) );
AOI21_X1 _17064_ ( .A(\EX_LS_pc [30] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01187_ ) );
MUX2_X1 _17065_ ( .A(\LS_WB_wdata_csreg [30] ), .B(\EX_LS_result_csreg_mem [30] ), .S(_01172_ ), .Z(_01188_ ) );
NOR3_X1 _17066_ ( .A1(_03813_ ), .A2(_03818_ ), .A3(_01188_ ), .ZN(_01189_ ) );
NOR2_X1 _17067_ ( .A1(_01187_ ), .A2(_01189_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ) );
MUX2_X1 _17068_ ( .A(\LS_WB_wdata_csreg [11] ), .B(\EX_LS_result_csreg_mem [11] ), .S(_01179_ ), .Z(_01190_ ) );
MUX2_X1 _17069_ ( .A(_01190_ ), .B(\EX_LS_pc [11] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ) );
MUX2_X1 _17070_ ( .A(\LS_WB_wdata_csreg [10] ), .B(\EX_LS_result_csreg_mem [10] ), .S(_01179_ ), .Z(_01191_ ) );
MUX2_X1 _17071_ ( .A(_01191_ ), .B(\EX_LS_pc [10] ), .S(_03820_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ) );
OAI22_X1 _17072_ ( .A1(_03824_ ), .A2(_02072_ ), .B1(_03829_ ), .B2(_05831_ ), .ZN(_01192_ ) );
BUF_X4 _17073_ ( .A(_03819_ ), .Z(_01193_ ) );
MUX2_X1 _17074_ ( .A(_01192_ ), .B(\EX_LS_pc [9] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ) );
AOI21_X1 _17075_ ( .A(\EX_LS_pc [8] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01194_ ) );
MUX2_X1 _17076_ ( .A(\LS_WB_wdata_csreg [8] ), .B(\EX_LS_result_csreg_mem [8] ), .S(_01172_ ), .Z(_01195_ ) );
NOR3_X1 _17077_ ( .A1(_03813_ ), .A2(_03818_ ), .A3(_01195_ ), .ZN(_01196_ ) );
NOR2_X1 _17078_ ( .A1(_01194_ ), .A2(_01196_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ) );
AOI21_X1 _17079_ ( .A(\EX_LS_pc [7] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01197_ ) );
INV_X1 _17080_ ( .A(_03823_ ), .ZN(_01198_ ) );
OAI21_X1 _17081_ ( .A(_03817_ ), .B1(_01198_ ), .B2(_03986_ ), .ZN(_01199_ ) );
AOI221_X4 _17082_ ( .A(_01199_ ), .B1(\LS_WB_wdata_csreg [7] ), .B2(_01198_ ), .C1(_02075_ ), .C2(_02036_ ), .ZN(_01200_ ) );
NOR2_X1 _17083_ ( .A1(_01197_ ), .A2(_01200_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ) );
OAI22_X1 _17084_ ( .A1(_03824_ ), .A2(_02073_ ), .B1(_03829_ ), .B2(_03987_ ), .ZN(_01201_ ) );
MUX2_X1 _17085_ ( .A(_01201_ ), .B(\EX_LS_pc [6] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ) );
MUX2_X1 _17086_ ( .A(\LS_WB_wdata_csreg [5] ), .B(\EX_LS_result_csreg_mem [5] ), .S(_01179_ ), .Z(_01202_ ) );
MUX2_X1 _17087_ ( .A(_01202_ ), .B(\EX_LS_pc [5] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ) );
OAI22_X1 _17088_ ( .A1(_03824_ ), .A2(_02069_ ), .B1(_03829_ ), .B2(_03975_ ), .ZN(_01203_ ) );
MUX2_X1 _17089_ ( .A(_01203_ ), .B(\EX_LS_pc [4] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ) );
MUX2_X1 _17090_ ( .A(\LS_WB_wdata_csreg [3] ), .B(\EX_LS_result_csreg_mem [3] ), .S(_01179_ ), .Z(_01204_ ) );
MUX2_X1 _17091_ ( .A(_01204_ ), .B(\EX_LS_pc [3] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ) );
AOI221_X4 _17092_ ( .A(_03819_ ), .B1(_01945_ ), .B2(\LS_WB_wdata_csreg [2] ), .C1(\EX_LS_result_csreg_mem [2] ), .C2(_03824_ ), .ZN(_01205_ ) );
AOI21_X1 _17093_ ( .A(\EX_LS_pc [2] ), .B1(_03868_ ), .B2(_03817_ ), .ZN(_01206_ ) );
NOR2_X1 _17094_ ( .A1(_01205_ ), .A2(_01206_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ) );
MUX2_X1 _17095_ ( .A(\LS_WB_wdata_csreg [29] ), .B(\EX_LS_result_csreg_mem [29] ), .S(_01179_ ), .Z(_01207_ ) );
MUX2_X1 _17096_ ( .A(_01207_ ), .B(\EX_LS_pc [29] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ) );
AOI21_X1 _17097_ ( .A(\EX_LS_pc [1] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01208_ ) );
OAI21_X1 _17098_ ( .A(_03817_ ), .B1(_01198_ ), .B2(_03978_ ), .ZN(_01209_ ) );
AOI221_X4 _17099_ ( .A(_01209_ ), .B1(\LS_WB_wdata_csreg [1] ), .B2(_01198_ ), .C1(_02075_ ), .C2(_02036_ ), .ZN(_01210_ ) );
NOR2_X1 _17100_ ( .A1(_01208_ ), .A2(_01210_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ) );
AOI21_X1 _17101_ ( .A(\EX_LS_pc [0] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01211_ ) );
OAI21_X1 _17102_ ( .A(_03817_ ), .B1(_01198_ ), .B2(_03979_ ), .ZN(_01212_ ) );
AOI221_X4 _17103_ ( .A(_01212_ ), .B1(\LS_WB_wdata_csreg [0] ), .B2(_01198_ ), .C1(_02075_ ), .C2(_02036_ ), .ZN(_01213_ ) );
NOR2_X1 _17104_ ( .A1(_01211_ ), .A2(_01213_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ) );
MUX2_X1 _17105_ ( .A(\LS_WB_wdata_csreg [28] ), .B(\EX_LS_result_csreg_mem [28] ), .S(_01179_ ), .Z(_01214_ ) );
MUX2_X1 _17106_ ( .A(_01214_ ), .B(\EX_LS_pc [28] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ) );
AOI21_X1 _17107_ ( .A(\EX_LS_pc [27] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01215_ ) );
MUX2_X1 _17108_ ( .A(\LS_WB_wdata_csreg [27] ), .B(\EX_LS_result_csreg_mem [27] ), .S(_01172_ ), .Z(_01216_ ) );
NOR3_X1 _17109_ ( .A1(_03813_ ), .A2(_03818_ ), .A3(_01216_ ), .ZN(_01217_ ) );
NOR2_X1 _17110_ ( .A1(_01215_ ), .A2(_01217_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ) );
MUX2_X1 _17111_ ( .A(\LS_WB_wdata_csreg [26] ), .B(\EX_LS_result_csreg_mem [26] ), .S(_01172_ ), .Z(_01218_ ) );
MUX2_X1 _17112_ ( .A(_01218_ ), .B(\EX_LS_pc [26] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ) );
AOI21_X1 _17113_ ( .A(\EX_LS_pc [25] ), .B1(_03869_ ), .B2(_01170_ ), .ZN(_01219_ ) );
MUX2_X1 _17114_ ( .A(\LS_WB_wdata_csreg [25] ), .B(\EX_LS_result_csreg_mem [25] ), .S(_03823_ ), .Z(_01220_ ) );
NOR3_X1 _17115_ ( .A1(_03813_ ), .A2(_03818_ ), .A3(_01220_ ), .ZN(_01221_ ) );
NOR2_X1 _17116_ ( .A1(_01219_ ), .A2(_01221_ ), .ZN(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ) );
MUX2_X1 _17117_ ( .A(\LS_WB_wdata_csreg [24] ), .B(\EX_LS_result_csreg_mem [24] ), .S(_01172_ ), .Z(_01222_ ) );
MUX2_X1 _17118_ ( .A(_01222_ ), .B(\EX_LS_pc [24] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ) );
MUX2_X1 _17119_ ( .A(\LS_WB_wdata_csreg [23] ), .B(\EX_LS_result_csreg_mem [23] ), .S(_01172_ ), .Z(_01223_ ) );
MUX2_X1 _17120_ ( .A(_01223_ ), .B(\EX_LS_pc [23] ), .S(_01193_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ) );
MUX2_X1 _17121_ ( .A(\LS_WB_wdata_csreg [22] ), .B(\EX_LS_result_csreg_mem [22] ), .S(_01172_ ), .Z(_01224_ ) );
MUX2_X1 _17122_ ( .A(_01224_ ), .B(\EX_LS_pc [22] ), .S(_03819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ) );
MUX2_X1 _17123_ ( .A(\LS_WB_wdata_csreg [31] ), .B(\EX_LS_result_csreg_mem [31] ), .S(_01172_ ), .Z(_01225_ ) );
MUX2_X1 _17124_ ( .A(_01225_ ), .B(\EX_LS_pc [31] ), .S(_03819_ ), .Z(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ) );
NOR2_X1 _17125_ ( .A1(\mylsu.araddr_tmp [0] ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01226_ ) );
INV_X1 _17126_ ( .A(_01226_ ), .ZN(_01227_ ) );
OR3_X2 _17127_ ( .A1(_00484_ ), .A2(_03873_ ), .A3(_01227_ ), .ZN(_01228_ ) );
NAND3_X1 _17128_ ( .A1(_00455_ ), .A2(_01979_ ), .A3(_01227_ ), .ZN(_01229_ ) );
NAND2_X1 _17129_ ( .A1(_01228_ ), .A2(_01229_ ), .ZN(_01230_ ) );
AND2_X1 _17130_ ( .A1(\mylsu.typ_tmp_$_NOT__A_Y ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01231_ ) );
INV_X1 _17131_ ( .A(\mylsu.typ_tmp [0] ), .ZN(_01232_ ) );
AND2_X1 _17132_ ( .A1(_01231_ ), .A2(_01232_ ), .ZN(_01233_ ) );
BUF_X4 _17133_ ( .A(_01233_ ), .Z(_01234_ ) );
INV_X1 _17134_ ( .A(_01234_ ), .ZN(_01235_ ) );
NOR2_X1 _17135_ ( .A1(_01230_ ), .A2(_01235_ ), .ZN(_01236_ ) );
OR2_X1 _17136_ ( .A1(_01232_ ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01237_ ) );
NOR2_X1 _17137_ ( .A1(_01237_ ), .A2(\mylsu.typ_tmp [2] ), .ZN(_01238_ ) );
NOR2_X1 _17138_ ( .A1(\mylsu.typ_tmp [0] ), .A2(\mylsu.typ_tmp [1] ), .ZN(_01239_ ) );
AND2_X2 _17139_ ( .A1(_01239_ ), .A2(\mylsu.typ_tmp_$_NOT__A_Y ), .ZN(_01240_ ) );
NOR2_X1 _17140_ ( .A1(_01238_ ), .A2(_01240_ ), .ZN(_01241_ ) );
INV_X1 _17141_ ( .A(_01241_ ), .ZN(_01242_ ) );
NOR2_X2 _17142_ ( .A1(_01236_ ), .A2(_01242_ ), .ZN(_01243_ ) );
BUF_X4 _17143_ ( .A(_01243_ ), .Z(_01244_ ) );
BUF_X4 _17144_ ( .A(_01234_ ), .Z(_01245_ ) );
AND2_X2 _17145_ ( .A1(_01231_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01246_ ) );
NOR3_X1 _17146_ ( .A1(_00462_ ), .A2(_03898_ ), .A3(_01246_ ), .ZN(_01247_ ) );
OAI21_X1 _17147_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01247_ ), .ZN(_01248_ ) );
BUF_X2 _17148_ ( .A(_03873_ ), .Z(_01249_ ) );
NAND2_X1 _17149_ ( .A1(_03903_ ), .A2(\mylsu.araddr_tmp [1] ), .ZN(_01250_ ) );
NOR3_X1 _17150_ ( .A1(_00551_ ), .A2(_01249_ ), .A3(_01250_ ), .ZN(_01251_ ) );
NOR3_X1 _17151_ ( .A1(_00484_ ), .A2(\mylsu.araddr_tmp [1] ), .A3(_01249_ ), .ZN(_01252_ ) );
OAI21_X2 _17152_ ( .A(_01227_ ), .B1(_01251_ ), .B2(_01252_ ), .ZN(_01253_ ) );
OR3_X1 _17153_ ( .A1(_00892_ ), .A2(_01249_ ), .A3(_01227_ ), .ZN(_01254_ ) );
NAND4_X1 _17154_ ( .A1(_00455_ ), .A2(\mylsu.araddr_tmp [0] ), .A3(\mylsu.araddr_tmp [1] ), .A4(_01979_ ), .ZN(_01255_ ) );
NAND3_X2 _17155_ ( .A1(_01253_ ), .A2(_01254_ ), .A3(_01255_ ), .ZN(_01256_ ) );
NAND2_X2 _17156_ ( .A1(_01256_ ), .A2(_01240_ ), .ZN(_01257_ ) );
BUF_X4 _17157_ ( .A(_01257_ ), .Z(_01258_ ) );
NAND2_X1 _17158_ ( .A1(_01248_ ), .A2(_01258_ ), .ZN(_01259_ ) );
MUX2_X1 _17159_ ( .A(\EX_LS_result_reg [21] ), .B(_01259_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ) );
NAND3_X1 _17160_ ( .A1(_00463_ ), .A2(_00467_ ), .A3(\io_master_arid [1] ), .ZN(_01260_ ) );
NOR2_X1 _17161_ ( .A1(_01260_ ), .A2(_01246_ ), .ZN(_01261_ ) );
OAI21_X1 _17162_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01261_ ), .ZN(_01262_ ) );
NAND2_X1 _17163_ ( .A1(_01262_ ), .A2(_01258_ ), .ZN(_01263_ ) );
MUX2_X1 _17164_ ( .A(\EX_LS_result_reg [20] ), .B(_01263_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ) );
NAND3_X1 _17165_ ( .A1(_00468_ ), .A2(_00470_ ), .A3(\io_master_arid [1] ), .ZN(_01264_ ) );
NOR2_X1 _17166_ ( .A1(_01264_ ), .A2(_01246_ ), .ZN(_01265_ ) );
OAI21_X1 _17167_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01265_ ), .ZN(_01266_ ) );
NAND2_X1 _17168_ ( .A1(_01266_ ), .A2(_01258_ ), .ZN(_01267_ ) );
MUX2_X1 _17169_ ( .A(\EX_LS_result_reg [19] ), .B(_01267_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ) );
AOI21_X1 _17170_ ( .A(_03874_ ), .B1(_00472_ ), .B2(_00474_ ), .ZN(_01268_ ) );
BUF_X4 _17171_ ( .A(_01231_ ), .Z(_01269_ ) );
NAND2_X1 _17172_ ( .A1(_01269_ ), .A2(\mylsu.typ_tmp [0] ), .ZN(_01270_ ) );
AOI21_X1 _17173_ ( .A(_01234_ ), .B1(_01268_ ), .B2(_01270_ ), .ZN(_01271_ ) );
OR3_X1 _17174_ ( .A1(_01236_ ), .A2(_01242_ ), .A3(_01271_ ), .ZN(_01272_ ) );
NAND2_X1 _17175_ ( .A1(_01272_ ), .A2(_01258_ ), .ZN(_01273_ ) );
MUX2_X1 _17176_ ( .A(\EX_LS_result_reg [18] ), .B(_01273_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ) );
AND4_X1 _17177_ ( .A1(\io_master_arid [1] ), .A2(_00476_ ), .A3(_00478_ ), .A4(_01270_ ), .ZN(_01274_ ) );
OAI21_X1 _17178_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01274_ ), .ZN(_01275_ ) );
NAND2_X1 _17179_ ( .A1(_01275_ ), .A2(_01258_ ), .ZN(_01276_ ) );
MUX2_X1 _17180_ ( .A(\EX_LS_result_reg [17] ), .B(_01276_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ) );
AND4_X1 _17181_ ( .A1(\io_master_arid [1] ), .A2(_00479_ ), .A3(_00481_ ), .A4(_01270_ ), .ZN(_01277_ ) );
OAI21_X1 _17182_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01277_ ), .ZN(_01278_ ) );
NAND2_X1 _17183_ ( .A1(_01278_ ), .A2(_01258_ ), .ZN(_01279_ ) );
MUX2_X1 _17184_ ( .A(\EX_LS_result_reg [16] ), .B(_01279_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ) );
AND2_X4 _17185_ ( .A1(_01256_ ), .A2(_01240_ ), .ZN(_01280_ ) );
NOR4_X1 _17186_ ( .A1(_00484_ ), .A2(_03897_ ), .A3(_01269_ ), .A4(_01242_ ), .ZN(_01281_ ) );
INV_X1 _17187_ ( .A(_01231_ ), .ZN(_01282_ ) );
AOI21_X1 _17188_ ( .A(_01282_ ), .B1(_01228_ ), .B2(_01229_ ), .ZN(_01283_ ) );
OR3_X2 _17189_ ( .A1(_01280_ ), .A2(_01281_ ), .A3(_01283_ ), .ZN(_01284_ ) );
MUX2_X2 _17190_ ( .A(\EX_LS_result_reg [15] ), .B(_01284_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ) );
NOR2_X1 _17191_ ( .A1(_00487_ ), .A2(_03874_ ), .ZN(_01285_ ) );
NOR2_X1 _17192_ ( .A1(_01282_ ), .A2(_01226_ ), .ZN(_01286_ ) );
OAI21_X1 _17193_ ( .A(_01241_ ), .B1(_01285_ ), .B2(_01286_ ), .ZN(_01287_ ) );
AND2_X1 _17194_ ( .A1(_00458_ ), .A2(_01979_ ), .ZN(_01288_ ) );
INV_X1 _17195_ ( .A(_01288_ ), .ZN(_01289_ ) );
AOI21_X1 _17196_ ( .A(_01287_ ), .B1(_01286_ ), .B2(_01289_ ), .ZN(_01290_ ) );
OR2_X1 _17197_ ( .A1(_01280_ ), .A2(_01290_ ), .ZN(_01291_ ) );
MUX2_X1 _17198_ ( .A(\EX_LS_result_reg [14] ), .B(_01291_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ) );
INV_X1 _17199_ ( .A(_01286_ ), .ZN(_01292_ ) );
NAND2_X1 _17200_ ( .A1(_01979_ ), .A2(_01292_ ), .ZN(_01293_ ) );
NOR2_X1 _17201_ ( .A1(_01293_ ), .A2(_01242_ ), .ZN(_01294_ ) );
NAND3_X1 _17202_ ( .A1(_00488_ ), .A2(_00490_ ), .A3(_01294_ ), .ZN(_01295_ ) );
NOR2_X1 _17203_ ( .A1(_00496_ ), .A2(_01249_ ), .ZN(_01296_ ) );
INV_X1 _17204_ ( .A(_01296_ ), .ZN(_01297_ ) );
OAI211_X1 _17205_ ( .A(_01257_ ), .B(_01295_ ), .C1(_01292_ ), .C2(_01297_ ), .ZN(_01298_ ) );
MUX2_X1 _17206_ ( .A(\EX_LS_result_reg [13] ), .B(_01298_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ) );
NAND3_X1 _17207_ ( .A1(_00491_ ), .A2(_00493_ ), .A3(_01294_ ), .ZN(_01299_ ) );
NAND4_X1 _17208_ ( .A1(_00528_ ), .A2(_00530_ ), .A3(\io_master_arid [1] ), .A4(_01286_ ), .ZN(_01300_ ) );
NAND3_X1 _17209_ ( .A1(_01257_ ), .A2(_01299_ ), .A3(_01300_ ), .ZN(_01301_ ) );
MUX2_X1 _17210_ ( .A(\EX_LS_result_reg [12] ), .B(_01301_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ) );
AND3_X1 _17211_ ( .A1(_00458_ ), .A2(\io_master_arid [1] ), .A3(_01282_ ), .ZN(_01302_ ) );
OAI21_X1 _17212_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01302_ ), .ZN(_01303_ ) );
NAND2_X1 _17213_ ( .A1(_01303_ ), .A2(_01258_ ), .ZN(_01304_ ) );
MUX2_X1 _17214_ ( .A(\EX_LS_result_reg [30] ), .B(_01304_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ) );
NOR3_X1 _17215_ ( .A1(_01026_ ), .A2(_03897_ ), .A3(_01292_ ), .ZN(_01305_ ) );
AND3_X1 _17216_ ( .A1(_00498_ ), .A2(_00500_ ), .A3(_01294_ ), .ZN(_01306_ ) );
OR3_X2 _17217_ ( .A1(_01280_ ), .A2(_01305_ ), .A3(_01306_ ), .ZN(_01307_ ) );
MUX2_X2 _17218_ ( .A(\EX_LS_result_reg [11] ), .B(_01307_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ) );
AND2_X1 _17219_ ( .A1(_00540_ ), .A2(_00542_ ), .ZN(_01308_ ) );
NOR3_X1 _17220_ ( .A1(_01308_ ), .A2(_03897_ ), .A3(_01292_ ), .ZN(_01309_ ) );
AND3_X1 _17221_ ( .A1(_00501_ ), .A2(_00503_ ), .A3(_01294_ ), .ZN(_01310_ ) );
OR3_X2 _17222_ ( .A1(_01280_ ), .A2(_01309_ ), .A3(_01310_ ), .ZN(_01311_ ) );
MUX2_X2 _17223_ ( .A(\EX_LS_result_reg [10] ), .B(_01311_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ) );
AND2_X1 _17224_ ( .A1(_00544_ ), .A2(_00545_ ), .ZN(_01312_ ) );
NOR3_X1 _17225_ ( .A1(_01312_ ), .A2(_03897_ ), .A3(_01292_ ), .ZN(_01313_ ) );
AND3_X1 _17226_ ( .A1(_00504_ ), .A2(_00506_ ), .A3(_01294_ ), .ZN(_01314_ ) );
OR3_X2 _17227_ ( .A1(_01280_ ), .A2(_01313_ ), .A3(_01314_ ), .ZN(_01315_ ) );
MUX2_X2 _17228_ ( .A(\EX_LS_result_reg [9] ), .B(_01315_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ) );
NOR3_X1 _17229_ ( .A1(_01069_ ), .A2(_03897_ ), .A3(_01292_ ), .ZN(_01316_ ) );
AND3_X1 _17230_ ( .A1(_00507_ ), .A2(_00509_ ), .A3(_01294_ ), .ZN(_01317_ ) );
OR3_X2 _17231_ ( .A1(_01280_ ), .A2(_01316_ ), .A3(_01317_ ), .ZN(_01318_ ) );
MUX2_X2 _17232_ ( .A(\EX_LS_result_reg [8] ), .B(_01318_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ) );
NOR3_X1 _17233_ ( .A1(_00551_ ), .A2(_03898_ ), .A3(_01292_ ), .ZN(_01319_ ) );
OAI21_X1 _17234_ ( .A(_01241_ ), .B1(_00892_ ), .B2(_01293_ ), .ZN(_01320_ ) );
OAI221_X1 _17235_ ( .A(\mylsu.state [3] ), .B1(_01319_ ), .B2(_01320_ ), .C1(_01256_ ), .C2(_01241_ ), .ZN(_01321_ ) );
NAND2_X1 _17236_ ( .A1(_03959_ ), .A2(\EX_LS_result_reg [7] ), .ZN(_01322_ ) );
NAND2_X1 _17237_ ( .A1(_01321_ ), .A2(_01322_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ) );
NAND2_X1 _17238_ ( .A1(_03900_ ), .A2(\mylsu.araddr_tmp [0] ), .ZN(_01323_ ) );
NOR3_X1 _17239_ ( .A1(_00554_ ), .A2(_03874_ ), .A3(_01250_ ), .ZN(_01324_ ) );
AND3_X1 _17240_ ( .A1(_00458_ ), .A2(_01979_ ), .A3(_01250_ ), .ZN(_01325_ ) );
OAI21_X1 _17241_ ( .A(_01323_ ), .B1(_01324_ ), .B2(_01325_ ), .ZN(_01326_ ) );
OR3_X1 _17242_ ( .A1(_00487_ ), .A2(_01249_ ), .A3(_01323_ ), .ZN(_01327_ ) );
AOI21_X1 _17243_ ( .A(_01226_ ), .B1(_01326_ ), .B2(_01327_ ), .ZN(_01328_ ) );
NOR3_X1 _17244_ ( .A1(_00515_ ), .A2(_01249_ ), .A3(_01227_ ), .ZN(_01329_ ) );
OAI21_X1 _17245_ ( .A(_01240_ ), .B1(_01328_ ), .B2(_01329_ ), .ZN(_01330_ ) );
NOR3_X1 _17246_ ( .A1(_00554_ ), .A2(_03874_ ), .A3(_01226_ ), .ZN(_01331_ ) );
OAI21_X1 _17247_ ( .A(_01246_ ), .B1(_01331_ ), .B2(_01329_ ), .ZN(_01332_ ) );
OR3_X1 _17248_ ( .A1(_00515_ ), .A2(_03874_ ), .A3(_01246_ ), .ZN(_01333_ ) );
AOI21_X1 _17249_ ( .A(_01234_ ), .B1(_01332_ ), .B2(_01333_ ), .ZN(_01334_ ) );
OR3_X1 _17250_ ( .A1(_00554_ ), .A2(_03874_ ), .A3(_01226_ ), .ZN(_01335_ ) );
OR3_X1 _17251_ ( .A1(_00515_ ), .A2(_01249_ ), .A3(_01227_ ), .ZN(_01336_ ) );
AOI21_X1 _17252_ ( .A(_01235_ ), .B1(_01335_ ), .B2(_01336_ ), .ZN(_01337_ ) );
OAI22_X1 _17253_ ( .A1(_01334_ ), .A2(_01337_ ), .B1(\mylsu.typ_tmp [2] ), .B2(_01237_ ), .ZN(_01338_ ) );
OAI21_X1 _17254_ ( .A(_01238_ ), .B1(_01328_ ), .B2(_01329_ ), .ZN(_01339_ ) );
AND2_X1 _17255_ ( .A1(_01338_ ), .A2(_01339_ ), .ZN(_01340_ ) );
OAI21_X1 _17256_ ( .A(_01330_ ), .B1(_01340_ ), .B2(_01240_ ), .ZN(_01341_ ) );
MUX2_X1 _17257_ ( .A(\EX_LS_result_reg [6] ), .B(_01341_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ) );
NAND2_X1 _17258_ ( .A1(_01296_ ), .A2(_01250_ ), .ZN(_01342_ ) );
OR3_X1 _17259_ ( .A1(_00462_ ), .A2(_01249_ ), .A3(_01250_ ), .ZN(_01343_ ) );
AOI22_X1 _17260_ ( .A1(_01342_ ), .A2(_01343_ ), .B1(\mylsu.araddr_tmp [0] ), .B2(_03900_ ), .ZN(_01344_ ) );
NOR3_X1 _17261_ ( .A1(_00800_ ), .A2(_03874_ ), .A3(_01323_ ), .ZN(_01345_ ) );
OAI21_X1 _17262_ ( .A(_01227_ ), .B1(_01344_ ), .B2(_01345_ ), .ZN(_01346_ ) );
NOR3_X1 _17263_ ( .A1(_00518_ ), .A2(_01249_ ), .A3(_01227_ ), .ZN(_01347_ ) );
INV_X1 _17264_ ( .A(_01347_ ), .ZN(_01348_ ) );
NAND2_X1 _17265_ ( .A1(_01346_ ), .A2(_01348_ ), .ZN(_01349_ ) );
NAND2_X1 _17266_ ( .A1(_01349_ ), .A2(_01240_ ), .ZN(_01350_ ) );
NOR3_X1 _17267_ ( .A1(_00462_ ), .A2(_01249_ ), .A3(_01226_ ), .ZN(_01351_ ) );
INV_X1 _17268_ ( .A(_01351_ ), .ZN(_01352_ ) );
AOI21_X1 _17269_ ( .A(_01270_ ), .B1(_01348_ ), .B2(_01352_ ), .ZN(_01353_ ) );
NOR3_X1 _17270_ ( .A1(_00518_ ), .A2(_03874_ ), .A3(_01246_ ), .ZN(_01354_ ) );
OAI21_X1 _17271_ ( .A(_01235_ ), .B1(_01353_ ), .B2(_01354_ ), .ZN(_01355_ ) );
OAI21_X1 _17272_ ( .A(_01234_ ), .B1(_01347_ ), .B2(_01351_ ), .ZN(_01356_ ) );
AOI21_X1 _17273_ ( .A(_01238_ ), .B1(_01355_ ), .B2(_01356_ ), .ZN(_01357_ ) );
AOI21_X1 _17274_ ( .A(_01357_ ), .B1(_01238_ ), .B2(_01349_ ), .ZN(_01358_ ) );
OAI21_X1 _17275_ ( .A(_01350_ ), .B1(_01358_ ), .B2(_01240_ ), .ZN(_01359_ ) );
MUX2_X1 _17276_ ( .A(\EX_LS_result_reg [5] ), .B(_01359_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ) );
NOR3_X1 _17277_ ( .A1(_01238_ ), .A2(_01269_ ), .A3(_01240_ ), .ZN(_01360_ ) );
NOR2_X1 _17278_ ( .A1(_01360_ ), .A2(_01226_ ), .ZN(_01361_ ) );
INV_X1 _17279_ ( .A(_01361_ ), .ZN(_01362_ ) );
AOI211_X1 _17280_ ( .A(_03958_ ), .B(_03899_ ), .C1(_00521_ ), .C2(_01362_ ), .ZN(_01363_ ) );
NOR2_X1 _17281_ ( .A1(_01241_ ), .A2(_03903_ ), .ZN(_01364_ ) );
NOR2_X1 _17282_ ( .A1(_01362_ ), .A2(_01364_ ), .ZN(_01365_ ) );
NAND2_X1 _17283_ ( .A1(_00684_ ), .A2(_01365_ ), .ZN(_01366_ ) );
AND3_X1 _17284_ ( .A1(_00528_ ), .A2(_00530_ ), .A3(\mylsu.araddr_tmp [1] ), .ZN(_01367_ ) );
OAI21_X1 _17285_ ( .A(_01364_ ), .B1(_00817_ ), .B2(\mylsu.araddr_tmp [1] ), .ZN(_01368_ ) );
OAI211_X1 _17286_ ( .A(_01363_ ), .B(_01366_ ), .C1(_01367_ ), .C2(_01368_ ), .ZN(_01369_ ) );
NAND2_X1 _17287_ ( .A1(_03959_ ), .A2(\EX_LS_result_reg [4] ), .ZN(_01370_ ) );
NAND2_X1 _17288_ ( .A1(_01369_ ), .A2(_01370_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ) );
NAND2_X1 _17289_ ( .A1(_03959_ ), .A2(\EX_LS_result_reg [3] ), .ZN(_01371_ ) );
AOI211_X1 _17290_ ( .A(_03959_ ), .B(_03899_ ), .C1(_00702_ ), .C2(_01365_ ), .ZN(_01372_ ) );
NAND2_X1 _17291_ ( .A1(_00524_ ), .A2(_01362_ ), .ZN(_01373_ ) );
NAND2_X1 _17292_ ( .A1(_01372_ ), .A2(_01373_ ), .ZN(_01374_ ) );
NAND3_X1 _17293_ ( .A1(_00498_ ), .A2(_00500_ ), .A3(_03900_ ), .ZN(_01375_ ) );
NAND2_X1 _17294_ ( .A1(_02009_ ), .A2(_00537_ ), .ZN(_01376_ ) );
OAI211_X1 _17295_ ( .A(_01376_ ), .B(\mylsu.araddr_tmp [1] ), .C1(\io_master_rdata [27] ), .C2(_02009_ ), .ZN(_01377_ ) );
AND3_X1 _17296_ ( .A1(_01375_ ), .A2(_01364_ ), .A3(_01377_ ), .ZN(_01378_ ) );
OAI21_X1 _17297_ ( .A(_01371_ ), .B1(_01374_ ), .B2(_01378_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ) );
NAND2_X1 _17298_ ( .A1(_03959_ ), .A2(\EX_LS_result_reg [2] ), .ZN(_01379_ ) );
NAND2_X1 _17299_ ( .A1(_00527_ ), .A2(_01362_ ), .ZN(_01380_ ) );
NAND3_X1 _17300_ ( .A1(_00472_ ), .A2(_00474_ ), .A3(_01365_ ), .ZN(_01381_ ) );
NAND4_X1 _17301_ ( .A1(_01380_ ), .A2(\mylsu.state [3] ), .A3(\io_master_arid [1] ), .A4(_01381_ ), .ZN(_01382_ ) );
NAND3_X1 _17302_ ( .A1(_00501_ ), .A2(_00503_ ), .A3(_03900_ ), .ZN(_01383_ ) );
OR2_X1 _17303_ ( .A1(_01308_ ), .A2(_03900_ ), .ZN(_01384_ ) );
AND3_X1 _17304_ ( .A1(_01383_ ), .A2(_01364_ ), .A3(_01384_ ), .ZN(_01385_ ) );
OAI21_X1 _17305_ ( .A(_01379_ ), .B1(_01382_ ), .B2(_01385_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ) );
NOR3_X1 _17306_ ( .A1(_00496_ ), .A2(_03898_ ), .A3(_01269_ ), .ZN(_01386_ ) );
OAI21_X1 _17307_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01386_ ), .ZN(_01387_ ) );
NAND2_X1 _17308_ ( .A1(_01387_ ), .A2(_01258_ ), .ZN(_01388_ ) );
MUX2_X1 _17309_ ( .A(\EX_LS_result_reg [29] ), .B(_01388_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ) );
AOI211_X1 _17310_ ( .A(_03958_ ), .B(_03898_ ), .C1(_00732_ ), .C2(_01365_ ), .ZN(_01389_ ) );
NAND2_X1 _17311_ ( .A1(_00533_ ), .A2(_01362_ ), .ZN(_01390_ ) );
NAND2_X1 _17312_ ( .A1(_01389_ ), .A2(_01390_ ), .ZN(_01391_ ) );
MUX2_X1 _17313_ ( .A(_01312_ ), .B(_00875_ ), .S(_03900_ ), .Z(_01392_ ) );
AOI21_X1 _17314_ ( .A(_01391_ ), .B1(_01364_ ), .B2(_01392_ ), .ZN(_01393_ ) );
AND2_X1 _17315_ ( .A1(_03959_ ), .A2(\EX_LS_result_reg [1] ), .ZN(_01394_ ) );
OR2_X1 _17316_ ( .A1(_01393_ ), .A2(_01394_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ) );
AOI211_X1 _17317_ ( .A(_03958_ ), .B(_03897_ ), .C1(_00749_ ), .C2(_01365_ ), .ZN(_01395_ ) );
NAND2_X1 _17318_ ( .A1(_00536_ ), .A2(_01362_ ), .ZN(_01396_ ) );
NAND2_X1 _17319_ ( .A1(_01395_ ), .A2(_01396_ ), .ZN(_01397_ ) );
MUX2_X1 _17320_ ( .A(_01069_ ), .B(_00594_ ), .S(_03900_ ), .Z(_01398_ ) );
AOI21_X1 _17321_ ( .A(_01397_ ), .B1(_01364_ ), .B2(_01398_ ), .ZN(_01399_ ) );
AND2_X1 _17322_ ( .A1(_03959_ ), .A2(\EX_LS_result_reg [0] ), .ZN(_01400_ ) );
OR2_X1 _17323_ ( .A1(_01399_ ), .A2(_01400_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ) );
AND4_X1 _17324_ ( .A1(_01979_ ), .A2(_00528_ ), .A3(_00530_ ), .A4(_01282_ ), .ZN(_01401_ ) );
OAI21_X1 _17325_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01401_ ), .ZN(_01402_ ) );
NAND2_X1 _17326_ ( .A1(_01402_ ), .A2(_01258_ ), .ZN(_01403_ ) );
MUX2_X1 _17327_ ( .A(\EX_LS_result_reg [28] ), .B(_01403_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ) );
AND2_X4 _17328_ ( .A1(_01258_ ), .A2(\mylsu.state [3] ), .ZN(_01404_ ) );
AOI211_X1 _17329_ ( .A(_03898_ ), .B(_01269_ ), .C1(_00538_ ), .C2(_00539_ ), .ZN(_01405_ ) );
OAI21_X1 _17330_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01405_ ), .ZN(_01406_ ) );
AOI22_X1 _17331_ ( .A1(_01404_ ), .A2(_01406_ ), .B1(_03959_ ), .B2(_04457_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ) );
AOI211_X1 _17332_ ( .A(_03897_ ), .B(_01269_ ), .C1(_00540_ ), .C2(_00542_ ), .ZN(_01407_ ) );
OAI21_X1 _17333_ ( .A(_01243_ ), .B1(_01234_ ), .B2(_01407_ ), .ZN(_01408_ ) );
NAND2_X1 _17334_ ( .A1(_01408_ ), .A2(_01257_ ), .ZN(_01409_ ) );
MUX2_X1 _17335_ ( .A(\EX_LS_result_reg [26] ), .B(_01409_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ) );
AOI211_X1 _17336_ ( .A(_03898_ ), .B(_01269_ ), .C1(_00544_ ), .C2(_00545_ ), .ZN(_01410_ ) );
OAI21_X1 _17337_ ( .A(_01244_ ), .B1(_01245_ ), .B2(_01410_ ), .ZN(_01411_ ) );
AOI22_X1 _17338_ ( .A1(_01404_ ), .A2(_01411_ ), .B1(_03959_ ), .B2(_04535_ ), .ZN(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ) );
AOI211_X1 _17339_ ( .A(_03897_ ), .B(_01269_ ), .C1(_00546_ ), .C2(_00548_ ), .ZN(_01412_ ) );
OAI21_X1 _17340_ ( .A(_01243_ ), .B1(_01234_ ), .B2(_01412_ ), .ZN(_01413_ ) );
NAND2_X1 _17341_ ( .A1(_01413_ ), .A2(_01257_ ), .ZN(_01414_ ) );
MUX2_X1 _17342_ ( .A(\EX_LS_result_reg [24] ), .B(_01414_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ) );
NOR3_X1 _17343_ ( .A1(_00551_ ), .A2(_03898_ ), .A3(_01269_ ), .ZN(_01415_ ) );
OAI21_X1 _17344_ ( .A(_01243_ ), .B1(_01234_ ), .B2(_01415_ ), .ZN(_01416_ ) );
NAND2_X1 _17345_ ( .A1(_01416_ ), .A2(_01257_ ), .ZN(_01417_ ) );
MUX2_X1 _17346_ ( .A(\EX_LS_result_reg [23] ), .B(_01417_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ) );
NOR3_X1 _17347_ ( .A1(_00554_ ), .A2(_03898_ ), .A3(_01269_ ), .ZN(_01418_ ) );
OAI21_X1 _17348_ ( .A(_01243_ ), .B1(_01234_ ), .B2(_01418_ ), .ZN(_01419_ ) );
NAND2_X1 _17349_ ( .A1(_01419_ ), .A2(_01257_ ), .ZN(_01420_ ) );
MUX2_X1 _17350_ ( .A(\EX_LS_result_reg [22] ), .B(_01420_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17351_ ( .A1(_00455_ ), .A2(\io_master_arid [1] ), .A3(_01282_ ), .ZN(_01421_ ) );
OAI21_X1 _17352_ ( .A(_01243_ ), .B1(_01234_ ), .B2(_01421_ ), .ZN(_01422_ ) );
NAND2_X1 _17353_ ( .A1(_01422_ ), .A2(_01257_ ), .ZN(_01423_ ) );
MUX2_X1 _17354_ ( .A(\EX_LS_result_reg [31] ), .B(_01423_ ), .S(\mylsu.state [3] ), .Z(\mylsu.wdata_reg_$_DFFE_PP__Q_D ) );
AND4_X1 _17355_ ( .A1(_01626_ ), .A2(fanout_net_5 ), .A3(IDU_valid_EXU ), .A4(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ), .ZN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ) );
AND4_X1 _17356_ ( .A1(_01458_ ), .A2(fanout_net_5 ), .A3(\mylsu.state [0] ), .A4(_03856_ ), .ZN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ) );
INV_X1 _17357_ ( .A(\LS_WB_waddr_reg [3] ), .ZN(_01424_ ) );
NOR2_X1 _17358_ ( .A1(\LS_WB_waddr_reg [3] ), .A2(\LS_WB_waddr_reg [0] ), .ZN(_01425_ ) );
INV_X1 _17359_ ( .A(\LS_WB_waddr_reg [2] ), .ZN(_01426_ ) );
INV_X1 _17360_ ( .A(\LS_WB_waddr_reg [1] ), .ZN(_01427_ ) );
NAND3_X1 _17361_ ( .A1(_01425_ ), .A2(_01426_ ), .A3(_01427_ ), .ZN(_01428_ ) );
AND2_X1 _17362_ ( .A1(_01456_ ), .A2(LS_WB_wen_reg ), .ZN(_01429_ ) );
NAND2_X1 _17363_ ( .A1(_01428_ ), .A2(_01429_ ), .ZN(_01430_ ) );
NOR2_X1 _17364_ ( .A1(_01430_ ), .A2(_01427_ ), .ZN(_01431_ ) );
BUF_X4 _17365_ ( .A(_01430_ ), .Z(_01432_ ) );
NOR2_X1 _17366_ ( .A1(_01432_ ), .A2(_01426_ ), .ZN(_01433_ ) );
INV_X1 _17367_ ( .A(\LS_WB_waddr_reg [0] ), .ZN(_01434_ ) );
AND4_X1 _17368_ ( .A1(_01424_ ), .A2(_01431_ ), .A3(_01433_ ), .A4(_01434_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ) );
AND4_X1 _17369_ ( .A1(_01424_ ), .A2(_01431_ ), .A3(_01433_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ) );
NOR2_X1 _17370_ ( .A1(_01430_ ), .A2(_01424_ ), .ZN(_01435_ ) );
AND4_X1 _17371_ ( .A1(_01426_ ), .A2(_01431_ ), .A3(_01435_ ), .A4(\LS_WB_waddr_reg [0] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ) );
AOI21_X1 _17372_ ( .A(_01432_ ), .B1(_01424_ ), .B2(_01426_ ), .ZN(_01436_ ) );
NOR4_X1 _17373_ ( .A1(_01436_ ), .A2(_01431_ ), .A3(_01434_ ), .A4(_01432_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ) );
NOR2_X1 _17374_ ( .A1(_01432_ ), .A2(_01434_ ), .ZN(_01437_ ) );
NOR4_X1 _17375_ ( .A1(_01436_ ), .A2(_01437_ ), .A3(_01427_ ), .A4(_01432_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ) );
NOR4_X1 _17376_ ( .A1(_01436_ ), .A2(_01427_ ), .A3(_01434_ ), .A4(_01432_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ) );
AOI21_X1 _17377_ ( .A(_01432_ ), .B1(_01427_ ), .B2(_01434_ ), .ZN(_01438_ ) );
NOR4_X1 _17378_ ( .A1(_01438_ ), .A2(_01435_ ), .A3(_01426_ ), .A4(_01432_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ) );
NOR4_X1 _17379_ ( .A1(_01438_ ), .A2(_01433_ ), .A3(_01424_ ), .A4(_01432_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ) );
AND4_X1 _17380_ ( .A1(_01426_ ), .A2(_01437_ ), .A3(_01435_ ), .A4(_01427_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ) );
NOR4_X1 _17381_ ( .A1(_01438_ ), .A2(_01424_ ), .A3(_01426_ ), .A4(_01432_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ) );
AND4_X1 _17382_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01437_ ), .A3(_01435_ ), .A4(_01427_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ) );
AND4_X1 _17383_ ( .A1(_01426_ ), .A2(_01431_ ), .A3(_01435_ ), .A4(_01434_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ) );
AND4_X1 _17384_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01431_ ), .A3(_01435_ ), .A4(_01434_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ) );
AND4_X1 _17385_ ( .A1(\LS_WB_waddr_reg [2] ), .A2(_01437_ ), .A3(_01435_ ), .A4(\LS_WB_waddr_reg [1] ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ) );
CLKBUF_X1 _17386_ ( .A(reset ), .Z(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ) );
AND4_X1 _17387_ ( .A1(_01424_ ), .A2(_01437_ ), .A3(_01433_ ), .A4(_01427_ ), .ZN(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ) );
NAND3_X1 _17388_ ( .A1(_01932_ ), .A2(_01564_ ), .A3(_01939_ ), .ZN(_01439_ ) );
NAND2_X1 _17389_ ( .A1(_01439_ ), .A2(_01735_ ), .ZN(\myminixbar.state_$_DFF_P__Q_1_D ) );
AOI211_X1 _17390_ ( .A(reset ), .B(_01932_ ), .C1(_01933_ ), .C2(_01961_ ), .ZN(\myminixbar.state_$_DFF_P__Q_D ) );
CLKBUF_X2 _17391_ ( .A(_01428_ ), .Z(_01440_ ) );
CLKBUF_X2 _17392_ ( .A(_01429_ ), .Z(_01441_ ) );
AND3_X1 _17393_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [21] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ) );
AND3_X1 _17394_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [20] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ) );
AND3_X1 _17395_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [19] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ) );
AND3_X1 _17396_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [18] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ) );
AND3_X1 _17397_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [17] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ) );
AND3_X1 _17398_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [16] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ) );
AND3_X1 _17399_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [15] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ) );
AND3_X1 _17400_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [14] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ) );
AND3_X1 _17401_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [13] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ) );
AND3_X1 _17402_ ( .A1(_01440_ ), .A2(\LS_WB_wdata_reg [12] ), .A3(_01441_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ) );
CLKBUF_X2 _17403_ ( .A(_01428_ ), .Z(_01442_ ) );
CLKBUF_X2 _17404_ ( .A(_01429_ ), .Z(_01443_ ) );
AND3_X1 _17405_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [30] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ) );
AND3_X1 _17406_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [11] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ) );
AND3_X1 _17407_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [10] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ) );
AND3_X1 _17408_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [9] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ) );
AND3_X1 _17409_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [8] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ) );
AND3_X1 _17410_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [7] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ) );
AND3_X1 _17411_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [6] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ) );
AND3_X1 _17412_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [5] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ) );
AND3_X1 _17413_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [4] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ) );
AND3_X1 _17414_ ( .A1(_01442_ ), .A2(\LS_WB_wdata_reg [3] ), .A3(_01443_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ) );
CLKBUF_X2 _17415_ ( .A(_01428_ ), .Z(_01444_ ) );
CLKBUF_X2 _17416_ ( .A(_01429_ ), .Z(_01445_ ) );
AND3_X1 _17417_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [2] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ) );
AND3_X1 _17418_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [29] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ) );
AND3_X1 _17419_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [1] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ) );
AND3_X1 _17420_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [0] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ) );
AND3_X1 _17421_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [28] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ) );
AND3_X1 _17422_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [27] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ) );
AND3_X1 _17423_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [26] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ) );
AND3_X1 _17424_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [25] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ) );
AND3_X1 _17425_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [24] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ) );
AND3_X1 _17426_ ( .A1(_01444_ ), .A2(\LS_WB_wdata_reg [23] ), .A3(_01445_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ) );
AND3_X1 _17427_ ( .A1(_01428_ ), .A2(\LS_WB_wdata_reg [22] ), .A3(_01429_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ) );
AND3_X1 _17428_ ( .A1(_01428_ ), .A2(\LS_WB_wdata_reg [31] ), .A3(_01429_ ), .ZN(\myreg.Reg[9]_$_DFFE_PP__Q_D ) );
AND3_X1 _17429_ ( .A1(_01564_ ), .A2(\mysc.state [2] ), .A3(\mylsu.previous_load_done ), .ZN(\mysc.state_$_DFF_P__Q_1_D ) );
NAND2_X1 _17430_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01446_ ) );
AND2_X1 _17431_ ( .A1(_01446_ ), .A2(\myidu.stall_quest_loaduse ), .ZN(_01447_ ) );
INV_X1 _17432_ ( .A(_01447_ ), .ZN(_01448_ ) );
NOR2_X1 _17433_ ( .A1(\ID_EX_pc [2] ), .A2(LS_WB_pc ), .ZN(_01449_ ) );
OAI211_X1 _17434_ ( .A(_01456_ ), .B(\mysc.state [0] ), .C1(_01448_ ), .C2(_01449_ ), .ZN(_01450_ ) );
INV_X1 _17435_ ( .A(_01450_ ), .ZN(_01451_ ) );
OR3_X1 _17436_ ( .A1(_01451_ ), .A2(reset ), .A3(\mysc.state [1] ), .ZN(\mysc.state_$_DFF_P__Q_2_D ) );
NOR3_X1 _17437_ ( .A1(_01448_ ), .A2(reset ), .A3(_01449_ ), .ZN(_01452_ ) );
NAND2_X1 _17438_ ( .A1(_01452_ ), .A2(\mysc.state [0] ), .ZN(_01453_ ) );
OR3_X1 _17439_ ( .A1(_03890_ ), .A2(reset ), .A3(\mylsu.previous_load_done ), .ZN(_01454_ ) );
NAND2_X1 _17440_ ( .A1(_01453_ ), .A2(_01454_ ), .ZN(\mysc.state_$_DFF_P__Q_D ) );
CLKGATE_X1 _17441_ ( .CK(clock ), .E(\mylsu.previous_load_done ), .GCK(_07921_ ) );
CLKGATE_X1 _17442_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07922_ ) );
CLKGATE_X1 _17443_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07923_ ) );
CLKGATE_X1 _17444_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07924_ ) );
CLKGATE_X1 _17445_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_Y ), .GCK(_07925_ ) );
CLKGATE_X1 _17446_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_AND__A_Y ), .GCK(_07926_ ) );
CLKGATE_X1 _17447_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_14_Y ), .GCK(_07927_ ) );
CLKGATE_X1 _17448_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_13_Y ), .GCK(_07928_ ) );
CLKGATE_X1 _17449_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_12_Y ), .GCK(_07929_ ) );
CLKGATE_X1 _17450_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_11_Y ), .GCK(_07930_ ) );
CLKGATE_X1 _17451_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_8_Y ), .GCK(_07931_ ) );
CLKGATE_X1 _17452_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07932_ ) );
CLKGATE_X1 _17453_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07933_ ) );
CLKGATE_X1 _17454_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07934_ ) );
CLKGATE_X1 _17455_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_10_Y ), .GCK(_07935_ ) );
CLKGATE_X1 _17456_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07936_ ) );
CLKGATE_X1 _17457_ ( .CK(clock ), .E(\mylsu.wen_reg_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__A_9_Y ), .GCK(_07937_ ) );
CLKGATE_X1 _17458_ ( .CK(clock ), .E(io_master_bvalid_$_ANDNOT__A_Y_$_ANDNOT__A_Y_$_ANDNOT__B_Y_$_NOR__A_Y_$_ANDNOT__A_Y ), .GCK(_07938_ ) );
CLKGATE_X1 _17459_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_ANDNOT__A_Y ), .GCK(_07939_ ) );
CLKGATE_X1 _17460_ ( .CK(clock ), .E(\mylsu.previous_load_done_$_SDFFE_PP0P__Q_E ), .GCK(_07940_ ) );
CLKGATE_X1 _17461_ ( .CK(clock ), .E(\mylsu.pc_out_$_SDFFE_PP0P__Q_E ), .GCK(_07941_ ) );
CLKGATE_X1 _17462_ ( .CK(clock ), .E(io_master_wready_$_NOR__B_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_Y ), .GCK(_07942_ ) );
CLKGATE_X1 _17463_ ( .CK(clock ), .E(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_OR__B_Y_$_ANDNOT__B_Y ), .GCK(_07943_ ) );
CLKGATE_X1 _17464_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E ), .GCK(_07944_ ) );
CLKGATE_X1 _17465_ ( .CK(clock ), .E(\myifu.tmp_offset_$_SDFFE_PP0P__Q_E ), .GCK(_07945_ ) );
CLKGATE_X1 _17466_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP1P__Q_E ), .GCK(_07946_ ) );
CLKGATE_X1 _17467_ ( .CK(clock ), .E(\myifu.pc_$_SDFFE_PP0P__Q_E ), .GCK(_07947_ ) );
CLKGATE_X1 _17468_ ( .CK(clock ), .E(\myifu.myicache.valid[3]_$_DFFE_PP__Q_E ), .GCK(_07948_ ) );
CLKGATE_X1 _17469_ ( .CK(clock ), .E(\myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q_E ), .GCK(_07949_ ) );
CLKGATE_X1 _17470_ ( .CK(clock ), .E(\myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q_E ), .GCK(_07950_ ) );
CLKGATE_X1 _17471_ ( .CK(clock ), .E(\myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q_E ), .GCK(_07951_ ) );
CLKGATE_X1 _17472_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_2_Y ), .GCK(_07952_ ) );
CLKGATE_X1 _17473_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_3_Y ), .GCK(_07953_ ) );
CLKGATE_X1 _17474_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_1_Y ), .GCK(_07954_ ) );
CLKGATE_X1 _17475_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_AND__B_Y ), .GCK(_07955_ ) );
CLKGATE_X1 _17476_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_3_Y ), .GCK(_07956_ ) );
CLKGATE_X1 _17477_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07957_ ) );
CLKGATE_X1 _17478_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_7_Y ), .GCK(_07958_ ) );
CLKGATE_X1 _17479_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_4_Y ), .GCK(_07959_ ) );
CLKGATE_X1 _17480_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_2_Y ), .GCK(_07960_ ) );
CLKGATE_X1 _17481_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_5_Y ), .GCK(_07961_ ) );
CLKGATE_X1 _17482_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_6_Y ), .GCK(_07962_ ) );
CLKGATE_X1 _17483_ ( .CK(clock ), .E(\myifu.wen_$_ANDNOT__A_Y_$_ANDNOT__A_1_Y ), .GCK(_07963_ ) );
CLKGATE_X1 _17484_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07964_ ) );
CLKGATE_X1 _17485_ ( .CK(clock ), .E(\myifu.check_assert_$_DFFE_PP__Q_E ), .GCK(_07965_ ) );
CLKGATE_X1 _17486_ ( .CK(clock ), .E(\myidu.typ_$_SDFFE_PP0P__Q_E ), .GCK(_07966_ ) );
CLKGATE_X1 _17487_ ( .CK(clock ), .E(\myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q_E ), .GCK(_07967_ ) );
CLKGATE_X1 _17488_ ( .CK(clock ), .E(\myidu.stall_quest_fencei_$_SDFFE_PP0P__Q_E ), .GCK(_07968_ ) );
CLKGATE_X1 _17489_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07969_ ) );
CLKGATE_X1 _17490_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_A_$_OR__Y_B_$_OR__Y_A_$_OR__Y_A_$_OR__Y_A_$_OR__A_Y_$_OR__B_Y_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07970_ ) );
CLKGATE_X1 _17491_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__B_Y_$_OR__A_Y_$_NOR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07971_ ) );
CLKGATE_X1 _17492_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_A_$_ANDNOT__A_Y ), .GCK(_07972_ ) );
CLKGATE_X1 _17493_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_NOR__B_Y_$_ANDNOT__B_Y_$_ANDNOT__Y_4_B_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_OR__Y_A_$_ORNOT__Y_A_$_ORNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07973_ ) );
CLKGATE_X1 _17494_ ( .CK(clock ), .E(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E ), .GCK(_07974_ ) );
CLKGATE_X1 _17495_ ( .CK(clock ), .E(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_E ), .GCK(_07975_ ) );
CLKGATE_X1 _17496_ ( .CK(clock ), .E(\myifu.wen_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_B_$_ORNOT__Y_A_$_ANDNOT__A_Y_$_NAND__B_Y_$_ANDNOT__B_Y ), .GCK(_07976_ ) );
CLKGATE_X1 _17497_ ( .CK(clock ), .E(\myifu.check_assert_$_ORNOT__A_Y_$_MUX__A_S_$_OR__A_Y_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07977_ ) );
CLKGATE_X1 _17498_ ( .CK(clock ), .E(\myifu.check_assert_$_ORNOT__A_Y_$_MUX__A_S_$_OR__A_Y_$_ANDNOT__A_B_$_NOR__B_Y ), .GCK(_07978_ ) );
CLKGATE_X1 _17499_ ( .CK(clock ), .E(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B_$_ANDNOT__A_Y_$_ANDNOT__A_Y ), .GCK(_07979_ ) );
CLKGATE_X1 _17500_ ( .CK(clock ), .E(\myec.state_$_SDFFE_PP0P__Q_E ), .GCK(_07980_ ) );
CLKGATE_X1 _17501_ ( .CK(clock ), .E(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_B_$_MUX__Y_A_$_NOR__B_Y ), .GCK(_07981_ ) );
CLKGATE_X1 _17502_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_B_$_OR__Y_B_$_OR__Y_A_$_OR__B_Y_$_OR__A_Y_$_ANDNOT__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07982_ ) );
CLKGATE_X1 _17503_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_1_Y ), .GCK(_07983_ ) );
CLKGATE_X1 _17504_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_Y ), .GCK(_07984_ ) );
CLKGATE_X1 _17505_ ( .CK(clock ), .E(\mycsreg.excp_written_$_SDFF_PN0__Q_R_$_ANDNOT__A_B_$_OR__Y_A_$_OR__Y_B_$_OR__A_Y_$_OR__A_Y_$_OR__A_Y_$_ANDNOT__B_Y ), .GCK(_07985_ ) );
LOGIC1_X1 _17506_ ( .Z(\io_master_awid [0] ) );
LOGIC0_X1 _17507_ ( .Z(\io_master_arburst [1] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q ( .D(_00001_ ), .CK(clock ), .Q(\myclint.mtime [63] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_1 ( .D(_00002_ ), .CK(clock ), .Q(\myclint.mtime [62] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_10 ( .D(_00003_ ), .CK(clock ), .Q(\myclint.mtime [53] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_11 ( .D(_00004_ ), .CK(clock ), .Q(\myclint.mtime [52] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_12 ( .D(_00005_ ), .CK(clock ), .Q(\myclint.mtime [51] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_13 ( .D(_00006_ ), .CK(clock ), .Q(\myclint.mtime [50] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_14 ( .D(_00007_ ), .CK(clock ), .Q(\myclint.mtime [49] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_15 ( .D(_00008_ ), .CK(clock ), .Q(\myclint.mtime [48] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_16 ( .D(_00009_ ), .CK(clock ), .Q(\myclint.mtime [47] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_17 ( .D(_00010_ ), .CK(clock ), .Q(\myclint.mtime [46] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_18 ( .D(_00011_ ), .CK(clock ), .Q(\myclint.mtime [45] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_19 ( .D(_00012_ ), .CK(clock ), .Q(\myclint.mtime [44] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_2 ( .D(_00013_ ), .CK(clock ), .Q(\myclint.mtime [61] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_20 ( .D(_00014_ ), .CK(clock ), .Q(\myclint.mtime [43] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_21 ( .D(_00015_ ), .CK(clock ), .Q(\myclint.mtime [42] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_22 ( .D(_00016_ ), .CK(clock ), .Q(\myclint.mtime [41] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_23 ( .D(_00017_ ), .CK(clock ), .Q(\myclint.mtime [40] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_24 ( .D(_00018_ ), .CK(clock ), .Q(\myclint.mtime [39] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_25 ( .D(_00019_ ), .CK(clock ), .Q(\myclint.mtime [38] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_26 ( .D(_00020_ ), .CK(clock ), .Q(\myclint.mtime [37] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_27 ( .D(_00021_ ), .CK(clock ), .Q(\myclint.mtime [36] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_28 ( .D(_00022_ ), .CK(clock ), .Q(\myclint.mtime [35] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_29 ( .D(_00023_ ), .CK(clock ), .Q(\myclint.mtime [34] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_3 ( .D(_00024_ ), .CK(clock ), .Q(\myclint.mtime [60] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_30 ( .D(_00025_ ), .CK(clock ), .Q(\myclint.mtime [33] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_31 ( .D(_00026_ ), .CK(clock ), .Q(\myclint.mtime [32] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D_$_MUX__A_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_32 ( .D(_00027_ ), .CK(clock ), .Q(\myclint.mtime [31] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_33 ( .D(_00028_ ), .CK(clock ), .Q(\myclint.mtime [30] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_1_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_34 ( .D(_00029_ ), .CK(clock ), .Q(\myclint.mtime [29] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_2_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_35 ( .D(_00030_ ), .CK(clock ), .Q(\myclint.mtime [28] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_3_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_36 ( .D(_00031_ ), .CK(clock ), .Q(\myclint.mtime [27] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_37 ( .D(_00032_ ), .CK(clock ), .Q(\myclint.mtime [26] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_38 ( .D(_00033_ ), .CK(clock ), .Q(\myclint.mtime [25] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_39 ( .D(_00034_ ), .CK(clock ), .Q(\myclint.mtime [24] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_4 ( .D(_00035_ ), .CK(clock ), .Q(\myclint.mtime [59] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_4_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_40 ( .D(_00036_ ), .CK(clock ), .Q(\myclint.mtime [23] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_41 ( .D(_00037_ ), .CK(clock ), .Q(\myclint.mtime [22] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_42 ( .D(_00038_ ), .CK(clock ), .Q(\myclint.mtime [21] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_10_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_43 ( .D(_00039_ ), .CK(clock ), .Q(\myclint.mtime [20] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_11_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_44 ( .D(_00040_ ), .CK(clock ), .Q(\myclint.mtime [19] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_12_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_45 ( .D(_00041_ ), .CK(clock ), .Q(\myclint.mtime [18] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_13_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_46 ( .D(_00042_ ), .CK(clock ), .Q(\myclint.mtime [17] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_14_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_47 ( .D(_00043_ ), .CK(clock ), .Q(\myclint.mtime [16] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_15_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_48 ( .D(_00044_ ), .CK(clock ), .Q(\myclint.mtime [15] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_16_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_49 ( .D(_00045_ ), .CK(clock ), .Q(\myclint.mtime [14] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_17_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_5 ( .D(_00046_ ), .CK(clock ), .Q(\myclint.mtime [58] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_5_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_50 ( .D(_00047_ ), .CK(clock ), .Q(\myclint.mtime [13] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_18_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_51 ( .D(_00048_ ), .CK(clock ), .Q(\myclint.mtime [12] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_19_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_52 ( .D(_00049_ ), .CK(clock ), .Q(\myclint.mtime [11] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_20_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_53 ( .D(_00050_ ), .CK(clock ), .Q(\myclint.mtime [10] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_21_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_54 ( .D(_00051_ ), .CK(clock ), .Q(\myclint.mtime [9] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_22_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_55 ( .D(_00052_ ), .CK(clock ), .Q(\myclint.mtime [8] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_23_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_56 ( .D(_00053_ ), .CK(clock ), .Q(\myclint.mtime [7] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_24_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_57 ( .D(_00054_ ), .CK(clock ), .Q(\myclint.mtime [6] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_25_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_58 ( .D(_00055_ ), .CK(clock ), .Q(\myclint.mtime [5] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_26_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_59 ( .D(_00056_ ), .CK(clock ), .Q(\myclint.mtime [4] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_27_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_6 ( .D(_00057_ ), .CK(clock ), .Q(\myclint.mtime [57] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_6_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_60 ( .D(_00058_ ), .CK(clock ), .Q(\myclint.mtime [3] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_28_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_61 ( .D(_00059_ ), .CK(clock ), .Q(\myclint.mtime [2] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_29_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_62 ( .D(_00060_ ), .CK(clock ), .Q(\myclint.mtime [1] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_30_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_63 ( .D(_00061_ ), .CK(clock ), .Q(\myclint.mtime [0] ), .QN(\myclint.mtime_$_SDFF_PP0__Q_63_D [0] ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_7 ( .D(_00062_ ), .CK(clock ), .Q(\myclint.mtime [56] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_7_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_8 ( .D(_00063_ ), .CK(clock ), .Q(\myclint.mtime [55] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_8_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.mtime_$_SDFF_PP0__Q_9 ( .D(_00064_ ), .CK(clock ), .Q(\myclint.mtime [54] ), .QN(\myifu.myicache.data_data_in_$_ANDNOT__Y_9_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myclint.state_r_$_SDFF_PP0__Q ( .D(_00065_ ), .CK(clock ), .Q(\myclint.rvalid ), .QN(\myclint.state_r_$_NOT__A_Y ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][31] ), .QN(_08215_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][30] ), .QN(_08216_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][21] ), .QN(_08217_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][20] ), .QN(_08218_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][19] ), .QN(_08219_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][18] ), .QN(_08220_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][17] ), .QN(_08221_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][16] ), .QN(_08222_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][15] ), .QN(_08223_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][14] ), .QN(_08224_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][13] ), .QN(_08225_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][12] ), .QN(_08226_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][29] ), .QN(_08227_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][11] ), .QN(_08228_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][10] ), .QN(_08229_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][9] ), .QN(_08230_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][8] ), .QN(_08231_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][7] ), .QN(_08232_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][6] ), .QN(_08233_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][5] ), .QN(_08234_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][4] ), .QN(_08235_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][3] ), .QN(_08236_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][2] ), .QN(_08237_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][28] ), .QN(_08238_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][1] ), .QN(_08239_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][0] ), .QN(_08240_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][27] ), .QN(_08241_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][26] ), .QN(_08242_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][25] ), .QN(_08243_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][24] ), .QN(_08244_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][23] ), .QN(_08245_ ) );
DFF_X1 \mycsreg.CSReg[0]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07985_ ), .Q(\mycsreg.CSReg[0][22] ), .QN(_08246_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07984_ ), .Q(\mtvec [31] ), .QN(_08247_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07984_ ), .Q(\mtvec [30] ), .QN(_08248_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07984_ ), .Q(\mtvec [21] ), .QN(_08249_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07984_ ), .Q(\mtvec [20] ), .QN(_08250_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07984_ ), .Q(\mtvec [19] ), .QN(_08251_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07984_ ), .Q(\mtvec [18] ), .QN(_08252_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07984_ ), .Q(\mtvec [17] ), .QN(_08253_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07984_ ), .Q(\mtvec [16] ), .QN(_08254_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07984_ ), .Q(\mtvec [15] ), .QN(_08255_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07984_ ), .Q(\mtvec [14] ), .QN(_08256_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07984_ ), .Q(\mtvec [13] ), .QN(_08257_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07984_ ), .Q(\mtvec [12] ), .QN(_08258_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07984_ ), .Q(\mtvec [29] ), .QN(_08259_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07984_ ), .Q(\mtvec [11] ), .QN(_08260_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07984_ ), .Q(\mtvec [10] ), .QN(_08261_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07984_ ), .Q(\mtvec [9] ), .QN(_08262_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07984_ ), .Q(\mtvec [8] ), .QN(_08263_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07984_ ), .Q(\mtvec [7] ), .QN(_08264_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07984_ ), .Q(\mtvec [6] ), .QN(_08265_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07984_ ), .Q(\mtvec [5] ), .QN(_08266_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07984_ ), .Q(\mtvec [4] ), .QN(_08267_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07984_ ), .Q(\mtvec [3] ), .QN(_08268_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07984_ ), .Q(\mtvec [2] ), .QN(_08269_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07984_ ), .Q(\mtvec [28] ), .QN(_08270_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07984_ ), .Q(\mtvec [1] ), .QN(_08271_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07984_ ), .Q(\mtvec [0] ), .QN(_08272_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07984_ ), .Q(\mtvec [27] ), .QN(_08273_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07984_ ), .Q(\mtvec [26] ), .QN(_08274_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07984_ ), .Q(\mtvec [25] ), .QN(_08275_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07984_ ), .Q(\mtvec [24] ), .QN(_08276_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07984_ ), .Q(\mtvec [23] ), .QN(_08277_ ) );
DFF_X1 \mycsreg.CSReg[1]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07984_ ), .Q(\mtvec [22] ), .QN(_08278_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q ( .D(\LS_WB_wdata_csreg [31] ), .CK(_07983_ ), .Q(\mepc [31] ), .QN(_08279_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_1 ( .D(\LS_WB_wdata_csreg [30] ), .CK(_07983_ ), .Q(\mepc [30] ), .QN(_08280_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_10 ( .D(\LS_WB_wdata_csreg [21] ), .CK(_07983_ ), .Q(\mepc [21] ), .QN(_08281_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_11 ( .D(\LS_WB_wdata_csreg [20] ), .CK(_07983_ ), .Q(\mepc [20] ), .QN(_08282_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_12 ( .D(\LS_WB_wdata_csreg [19] ), .CK(_07983_ ), .Q(\mepc [19] ), .QN(_08283_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_13 ( .D(\LS_WB_wdata_csreg [18] ), .CK(_07983_ ), .Q(\mepc [18] ), .QN(_08284_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_14 ( .D(\LS_WB_wdata_csreg [17] ), .CK(_07983_ ), .Q(\mepc [17] ), .QN(_08285_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_15 ( .D(\LS_WB_wdata_csreg [16] ), .CK(_07983_ ), .Q(\mepc [16] ), .QN(_08286_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_16 ( .D(\LS_WB_wdata_csreg [15] ), .CK(_07983_ ), .Q(\mepc [15] ), .QN(_08287_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_17 ( .D(\LS_WB_wdata_csreg [14] ), .CK(_07983_ ), .Q(\mepc [14] ), .QN(_08288_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_18 ( .D(\LS_WB_wdata_csreg [13] ), .CK(_07983_ ), .Q(\mepc [13] ), .QN(_08289_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_19 ( .D(\LS_WB_wdata_csreg [12] ), .CK(_07983_ ), .Q(\mepc [12] ), .QN(_08290_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_2 ( .D(\LS_WB_wdata_csreg [29] ), .CK(_07983_ ), .Q(\mepc [29] ), .QN(_08291_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_20 ( .D(\LS_WB_wdata_csreg [11] ), .CK(_07983_ ), .Q(\mepc [11] ), .QN(_08292_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_21 ( .D(\LS_WB_wdata_csreg [10] ), .CK(_07983_ ), .Q(\mepc [10] ), .QN(_08293_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_22 ( .D(\LS_WB_wdata_csreg [9] ), .CK(_07983_ ), .Q(\mepc [9] ), .QN(_08294_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_23 ( .D(\LS_WB_wdata_csreg [8] ), .CK(_07983_ ), .Q(\mepc [8] ), .QN(_08295_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_24 ( .D(\LS_WB_wdata_csreg [7] ), .CK(_07983_ ), .Q(\mepc [7] ), .QN(_08296_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_25 ( .D(\LS_WB_wdata_csreg [6] ), .CK(_07983_ ), .Q(\mepc [6] ), .QN(_08297_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_26 ( .D(\LS_WB_wdata_csreg [5] ), .CK(_07983_ ), .Q(\mepc [5] ), .QN(_08298_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_27 ( .D(\LS_WB_wdata_csreg [4] ), .CK(_07983_ ), .Q(\mepc [4] ), .QN(_08299_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_28 ( .D(\LS_WB_wdata_csreg [3] ), .CK(_07983_ ), .Q(\mepc [3] ), .QN(_08300_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_29 ( .D(\LS_WB_wdata_csreg [2] ), .CK(_07983_ ), .Q(\mepc [2] ), .QN(_08301_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_3 ( .D(\LS_WB_wdata_csreg [28] ), .CK(_07983_ ), .Q(\mepc [28] ), .QN(_08302_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_30 ( .D(\LS_WB_wdata_csreg [1] ), .CK(_07983_ ), .Q(\mepc [1] ), .QN(_08303_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_31 ( .D(\LS_WB_wdata_csreg [0] ), .CK(_07983_ ), .Q(\mepc [0] ), .QN(_08304_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_4 ( .D(\LS_WB_wdata_csreg [27] ), .CK(_07983_ ), .Q(\mepc [27] ), .QN(_08305_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_5 ( .D(\LS_WB_wdata_csreg [26] ), .CK(_07983_ ), .Q(\mepc [26] ), .QN(_08306_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_6 ( .D(\LS_WB_wdata_csreg [25] ), .CK(_07983_ ), .Q(\mepc [25] ), .QN(_08307_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_7 ( .D(\LS_WB_wdata_csreg [24] ), .CK(_07983_ ), .Q(\mepc [24] ), .QN(_08308_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_8 ( .D(\LS_WB_wdata_csreg [23] ), .CK(_07983_ ), .Q(\mepc [23] ), .QN(_08309_ ) );
DFF_X1 \mycsreg.CSReg[2]_$_DFFE_PP__Q_9 ( .D(\LS_WB_wdata_csreg [22] ), .CK(_07983_ ), .Q(\mepc [22] ), .QN(_08310_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_D ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][3] ), .QN(_08311_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_1 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_1_D ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][2] ), .QN(_08312_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_2 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_2_D ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][1] ), .QN(_08313_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_DFFE_PP__Q_3 ( .D(\mycsreg.CSReg[3]_$_DFFE_PP__Q_3_D ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][0] ), .QN(_08214_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q ( .D(_00066_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][5] ), .QN(_08213_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_1 ( .D(_00067_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][4] ), .QN(_08212_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_10 ( .D(_00068_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][23] ), .QN(_08211_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_11 ( .D(_00069_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][22] ), .QN(_08210_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_12 ( .D(_00070_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][21] ), .QN(_08209_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_13 ( .D(_00071_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][20] ), .QN(_08208_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_14 ( .D(_00072_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][19] ), .QN(_08207_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_15 ( .D(_00073_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][18] ), .QN(_08206_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_16 ( .D(_00074_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][17] ), .QN(_08205_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_17 ( .D(_00075_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][16] ), .QN(_08204_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_18 ( .D(_00076_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][15] ), .QN(_08203_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_19 ( .D(_00077_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][14] ), .QN(_08202_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_2 ( .D(_00078_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][31] ), .QN(_08201_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_20 ( .D(_00079_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][13] ), .QN(_08200_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_21 ( .D(_00080_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][12] ), .QN(_08199_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_22 ( .D(_00081_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][11] ), .QN(_08198_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_23 ( .D(_00082_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][10] ), .QN(_08197_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_24 ( .D(_00083_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][9] ), .QN(_08196_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_25 ( .D(_00084_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][8] ), .QN(_08195_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_26 ( .D(_00085_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][7] ), .QN(_08194_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_27 ( .D(_00086_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][6] ), .QN(_08193_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_3 ( .D(_00087_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][30] ), .QN(_08192_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_4 ( .D(_00088_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][29] ), .QN(_08191_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_5 ( .D(_00089_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][28] ), .QN(_08190_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_6 ( .D(_00090_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][27] ), .QN(_08189_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_7 ( .D(_00091_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][26] ), .QN(_08188_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_8 ( .D(_00092_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][25] ), .QN(_08187_ ) );
DFF_X1 \mycsreg.CSReg[3]_$_SDFFCE_PP0P__Q_9 ( .D(_00093_ ), .CK(_07982_ ), .Q(\mycsreg.CSReg[3][24] ), .QN(_08314_ ) );
DFF_X1 \mycsreg.excp_written_$_SDFF_PN0__Q ( .D(_00094_ ), .CK(clock ), .Q(excp_written ), .QN(_08315_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [31] ), .QN(_08186_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_1 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_1_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [30] ), .QN(_08316_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_10 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_10_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [21] ), .QN(_08317_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_11 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_11_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [20] ), .QN(_08318_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_12 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_12_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [19] ), .QN(_08319_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_13 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_13_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [18] ), .QN(_08320_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_14 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_14_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [17] ), .QN(_08321_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_15 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_15_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [16] ), .QN(_08322_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_16 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_16_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [15] ), .QN(_08323_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_17 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_17_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [14] ), .QN(_08324_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_18 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_18_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [13] ), .QN(_08325_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_19 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_19_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [12] ), .QN(_08326_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_2 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_2_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [29] ), .QN(_08327_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_20 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_20_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [11] ), .QN(_08328_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_21 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_21_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [10] ), .QN(_08329_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_22 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_22_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [9] ), .QN(_08330_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_23 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_23_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [8] ), .QN(_08331_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_24 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_24_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [7] ), .QN(_08332_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_25 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_25_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [6] ), .QN(_08333_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_26 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_26_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [5] ), .QN(_08334_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_27 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_27_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [4] ), .QN(_08335_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_28 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_28_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [3] ), .QN(_08336_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_29 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_29_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [2] ), .QN(_08337_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_3 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_3_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [28] ), .QN(_08338_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_30 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_30_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [1] ), .QN(_08339_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_31 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_31_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [0] ), .QN(_08340_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_4 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_4_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [27] ), .QN(_08341_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_5 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_5_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [26] ), .QN(_08342_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_6 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_6_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [25] ), .QN(_08343_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_7 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_7_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [24] ), .QN(_08344_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_8 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_8_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [23] ), .QN(_08345_ ) );
DFF_X1 \myec.mepc_tmp_$_DFFE_PP__Q_9 ( .D(\myec.mepc_tmp_$_DFFE_PP__Q_9_D ), .CK(_07981_ ), .Q(\myec.mepc_tmp [22] ), .QN(_08185_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q ( .D(_00095_ ), .CK(_07980_ ), .Q(\myec.state [1] ), .QN(_08184_ ) );
DFF_X1 \myec.state_$_SDFFE_PP0P__Q_1 ( .D(_00096_ ), .CK(_07980_ ), .Q(\myec.state [0] ), .QN(_08346_ ) );
DFFR_X1 \myexu.check_quest_$_DFF_PP0__Q ( .D(\myexu.check_quest_$_DFF_PP0__Q_D ), .RN(fanout_net_5 ), .CK(clock ), .Q(check_quest ), .QN(_08347_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [11] ), .QN(_08183_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [10] ), .QN(_08348_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [1] ), .QN(_08349_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [0] ), .QN(_08350_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [9] ), .QN(_08351_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [8] ), .QN(_08352_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [7] ), .QN(_08353_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [6] ), .QN(_08354_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [5] ), .QN(_08355_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [4] ), .QN(_08356_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [3] ), .QN(_08357_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.dest_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [2] ), .QN(_08182_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q ( .D(_00097_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [31] ), .QN(_08181_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_1 ( .D(_00098_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [30] ), .QN(_08180_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_10 ( .D(_00099_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [21] ), .QN(_08179_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_11 ( .D(_00100_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [20] ), .QN(_08178_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_12 ( .D(_00101_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [19] ), .QN(_08177_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_13 ( .D(_00102_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [18] ), .QN(_08176_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_14 ( .D(_00103_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [17] ), .QN(_08175_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_15 ( .D(_00104_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [16] ), .QN(_08174_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_16 ( .D(_00105_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [15] ), .QN(_08173_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_17 ( .D(_00106_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [14] ), .QN(_08172_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_18 ( .D(_00107_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [13] ), .QN(_08171_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_19 ( .D(_00108_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [12] ), .QN(_08170_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_2 ( .D(_00109_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [29] ), .QN(_08169_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_3 ( .D(_00110_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [28] ), .QN(_08168_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_4 ( .D(_00111_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [27] ), .QN(_08167_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_5 ( .D(_00112_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [26] ), .QN(_08166_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_6 ( .D(_00113_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [25] ), .QN(_08165_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_7 ( .D(_00114_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [24] ), .QN(_08164_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_8 ( .D(_00115_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [23] ), .QN(_08163_ ) );
DFF_X1 \myexu.dest_csreg_mem_$_SDFFCE_PP0P__Q_9 ( .D(_00116_ ), .CK(_07979_ ), .Q(\EX_LS_dest_csreg_mem [22] ), .QN(_08162_ ) );
DFFR_X1 \myexu.dest_reg_$_DFFE_PP0P__Q ( .D(\myexu.dest_reg_$_DFFE_PP0P__Q_D ), .RN(fanout_net_5 ), .CK(_07978_ ), .Q(\EX_LS_dest_reg [4] ), .QN(_08161_ ) );
DFFR_X1 \myexu.dest_reg_$_DFFE_PP0P__Q_1 ( .D(\myexu.dest_reg_$_DFFE_PP0P__Q_1_D ), .RN(fanout_net_5 ), .CK(_07978_ ), .Q(\EX_LS_dest_reg [3] ), .QN(_08160_ ) );
DFFR_X1 \myexu.dest_reg_$_DFFE_PP0P__Q_2 ( .D(\myexu.dest_reg_$_DFFE_PP0P__Q_2_D ), .RN(fanout_net_5 ), .CK(_07978_ ), .Q(\EX_LS_dest_reg [2] ), .QN(_08159_ ) );
DFFR_X1 \myexu.dest_reg_$_DFFE_PP0P__Q_3 ( .D(\myexu.dest_reg_$_DFFE_PP0P__Q_3_D ), .RN(fanout_net_5 ), .CK(_07978_ ), .Q(\EX_LS_dest_reg [1] ), .QN(_08158_ ) );
DFFR_X1 \myexu.dest_reg_$_DFFE_PP0P__Q_4 ( .D(\myexu.dest_reg_$_DFFE_PP0P__Q_4_D ), .RN(fanout_net_5 ), .CK(_07978_ ), .Q(\EX_LS_dest_reg [0] ), .QN(_08157_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [30] ), .QN(_08156_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_1 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_1_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [29] ), .QN(_08155_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_10 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_10_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [20] ), .QN(_08154_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_11 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_11_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [19] ), .QN(_08153_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_12 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_12_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [18] ), .QN(_08152_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_13 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_13_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [17] ), .QN(_08151_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_14 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_14_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [16] ), .QN(_08150_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_15 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_15_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [15] ), .QN(_08149_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_16 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_16_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [14] ), .QN(_08148_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_17 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_17_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [13] ), .QN(_08147_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_18 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_18_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [12] ), .QN(_08146_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_19 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_19_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [11] ), .QN(_08145_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_2 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_2_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [28] ), .QN(_08144_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_20 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_20_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [10] ), .QN(_08143_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_21 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_21_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [9] ), .QN(_08142_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_22 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_22_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [8] ), .QN(_08141_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_23 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_23_D ), .RN(fanout_net_5 ), .CK(_07977_ ), .Q(\myexu.pc_jump [7] ), .QN(_08140_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_24 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_24_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [6] ), .QN(_08139_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_25 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_25_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [5] ), .QN(_08138_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_26 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_26_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [4] ), .QN(_08137_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_27 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_27_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [3] ), .QN(_08136_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_28 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_28_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [2] ), .QN(_08135_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_29 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_29_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [1] ), .QN(_08134_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_3 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_3_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [27] ), .QN(_08133_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_30 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_30_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [0] ), .QN(_08132_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_4 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_4_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [26] ), .QN(_08131_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_5 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_5_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [25] ), .QN(_08130_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_6 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_6_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [24] ), .QN(_08129_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_7 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_7_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [23] ), .QN(_08128_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_8 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_8_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [22] ), .QN(_08127_ ) );
DFFR_X1 \myexu.pc_jump_$_DFFE_PP0P__Q_9 ( .D(\myexu.pc_jump_$_DFFE_PP0P__Q_9_D ), .RN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [21] ), .QN(_08126_ ) );
DFFS_X1 \myexu.pc_jump_$_DFFE_PP1P__Q ( .D(\myexu.pc_jump_$_DFFE_PP1P__Q_D ), .SN(fanout_net_6 ), .CK(_07977_ ), .Q(\myexu.pc_jump [31] ), .QN(_08125_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [31] ), .QN(_08124_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_1 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_1_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [30] ), .QN(_08123_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_10 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_10_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [21] ), .QN(_08122_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_11 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_11_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [20] ), .QN(_08121_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_12 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_12_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [19] ), .QN(_08120_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_13 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_13_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [18] ), .QN(_08119_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_14 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_14_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [17] ), .QN(_08118_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_15 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_15_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [16] ), .QN(_08117_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_16 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_16_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [15] ), .QN(_08116_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_17 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_17_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [14] ), .QN(_08115_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_18 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_18_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [13] ), .QN(_08114_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_19 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_19_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [12] ), .QN(_08113_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_2 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_2_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [29] ), .QN(_08112_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_20 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_20_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [11] ), .QN(_08111_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_21 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_21_D ), .RN(fanout_net_6 ), .CK(_07978_ ), .Q(\EX_LS_pc [10] ), .QN(_08110_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_22 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_22_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [9] ), .QN(_08109_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_23 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_23_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [8] ), .QN(_08108_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_24 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_24_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [7] ), .QN(_08107_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_25 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_25_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [6] ), .QN(_08106_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_26 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_26_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [5] ), .QN(_08105_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_27 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_27_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [4] ), .QN(_08104_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_28 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_28_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [3] ), .QN(_08103_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_29 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_29_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [2] ), .QN(_08102_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_3 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_3_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [28] ), .QN(_08101_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_30 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_30_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [1] ), .QN(_08100_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_31 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_31_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [0] ), .QN(_08099_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_4 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_4_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [27] ), .QN(_08098_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_5 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_5_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [26] ), .QN(_08097_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_6 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_6_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [25] ), .QN(_08096_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_7 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_7_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [24] ), .QN(_08095_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_8 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_8_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [23] ), .QN(_08094_ ) );
DFFR_X1 \myexu.pc_out_$_DFFE_PP0P__Q_9 ( .D(\myexu.pc_out_$_DFFE_PP0P__Q_9_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_pc [22] ), .QN(_08358_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [31] ), .QN(_08359_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_1 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_1_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [30] ), .QN(_08360_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_10 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_10_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [21] ), .QN(_08361_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_11 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_11_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [20] ), .QN(_08362_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_12 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_12_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [19] ), .QN(_08363_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_13 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_13_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [18] ), .QN(_08364_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_14 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_14_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [17] ), .QN(_08365_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_15 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_15_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [16] ), .QN(_08366_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_16 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_16_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [15] ), .QN(_08367_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_17 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_17_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [14] ), .QN(_08368_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_18 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_18_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [13] ), .QN(_08369_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_19 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_19_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [12] ), .QN(_08370_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_2 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [29] ), .QN(_08371_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_20 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_20_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [11] ), .QN(_08372_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_21 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [10] ), .QN(_08373_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_22 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_22_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [9] ), .QN(_08374_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_23 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_23_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [8] ), .QN(_08375_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_24 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [7] ), .QN(_08376_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_25 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [6] ), .QN(_08377_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_26 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [5] ), .QN(_08378_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_27 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [4] ), .QN(_08379_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_28 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [3] ), .QN(_08380_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_29 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [2] ), .QN(_08381_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_3 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [28] ), .QN(_08382_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_30 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_30_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [1] ), .QN(_08383_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_31 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_31_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [0] ), .QN(_08384_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_4 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [27] ), .QN(_08385_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_5 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [26] ), .QN(_08386_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_6 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [25] ), .QN(_08387_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_7 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [24] ), .QN(_08388_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_8 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_8_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [23] ), .QN(_08389_ ) );
DFF_X1 \myexu.result_csreg_mem_$_DFFE_PP__Q_9 ( .D(\myexu.result_csreg_mem_$_DFFE_PP__Q_9_D ), .CK(_07979_ ), .Q(\EX_LS_result_csreg_mem [22] ), .QN(_08390_ ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q ( .D(\myexu.result_reg_$_DFFE_PP__Q_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_1 ( .D(\myexu.result_reg_$_DFFE_PP__Q_1_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_10 ( .D(\myexu.result_reg_$_DFFE_PP__Q_10_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_11 ( .D(\myexu.result_reg_$_DFFE_PP__Q_11_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_12 ( .D(\myexu.result_reg_$_DFFE_PP__Q_12_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_13 ( .D(\myexu.result_reg_$_DFFE_PP__Q_13_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_14 ( .D(\myexu.result_reg_$_DFFE_PP__Q_14_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_15 ( .D(\myexu.result_reg_$_DFFE_PP__Q_15_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_16 ( .D(\myexu.result_reg_$_DFFE_PP__Q_16_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_17 ( .D(\myexu.result_reg_$_DFFE_PP__Q_17_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_18 ( .D(\myexu.result_reg_$_DFFE_PP__Q_18_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_19 ( .D(\myexu.result_reg_$_DFFE_PP__Q_19_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_2 ( .D(\myexu.result_reg_$_DFFE_PP__Q_2_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_20 ( .D(\myexu.result_reg_$_DFFE_PP__Q_20_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_21 ( .D(\myexu.result_reg_$_DFFE_PP__Q_21_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_22 ( .D(\myexu.result_reg_$_DFFE_PP__Q_22_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_23 ( .D(\myexu.result_reg_$_DFFE_PP__Q_23_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_24 ( .D(\myexu.result_reg_$_DFFE_PP__Q_24_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_25 ( .D(\myexu.result_reg_$_DFFE_PP__Q_25_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_26 ( .D(\myexu.result_reg_$_DFFE_PP__Q_26_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_27 ( .D(\myexu.result_reg_$_DFFE_PP__Q_27_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_28 ( .D(\myexu.result_reg_$_DFFE_PP__Q_28_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_29 ( .D(\myexu.result_reg_$_DFFE_PP__Q_29_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_3 ( .D(\myexu.result_reg_$_DFFE_PP__Q_3_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_30 ( .D(\myexu.result_reg_$_DFFE_PP__Q_30_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_31 ( .D(\myexu.result_reg_$_DFFE_PP__Q_31_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_4 ( .D(\myexu.result_reg_$_DFFE_PP__Q_4_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_5 ( .D(\myexu.result_reg_$_DFFE_PP__Q_5_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_6 ( .D(\myexu.result_reg_$_DFFE_PP__Q_6_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_7 ( .D(\myexu.result_reg_$_DFFE_PP__Q_7_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_Y_$_MUX__A_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_8 ( .D(\myexu.result_reg_$_DFFE_PP__Q_8_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myexu.result_reg_$_DFFE_PP__Q_9 ( .D(\myexu.result_reg_$_DFFE_PP__Q_9_D ), .CK(_07979_ ), .Q(\EX_LS_result_reg [22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_B ) );
DFFR_X1 \myexu.state_$_DFF_PP0__Q ( .D(\myexu.state_$_DFF_PP0__Q_D ), .RN(_00000_ ), .CK(clock ), .Q(EXU_valid_LSU ), .QN(\mylsu.wen_csreg_$_SDFFE_PP0P__Q_D_$_ANDNOT__Y_B_$_OR__Y_B ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_flag [2] ), .QN(\myidu.fc_disenable_$_NOT__A_Y_$_ANDNOT__A_B_$_OR__Y_B_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_B_$_ANDNOT__Y_A ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q_1 ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_1_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_flag [1] ), .QN(_08093_ ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q_2 ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_2_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_flag [0] ), .QN(_08092_ ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q_3 ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_3_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_typ [4] ), .QN(_08091_ ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q_4 ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_4_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_typ [3] ), .QN(_08090_ ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q_5 ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_5_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_typ [2] ), .QN(_08089_ ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q_6 ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_6_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_typ [1] ), .QN(_08088_ ) );
DFFR_X1 \myexu.typ_out_$_DFFE_PP0P__Q_7 ( .D(\myexu.typ_out_$_DFFE_PP0P__Q_7_D ), .RN(_00000_ ), .CK(_07978_ ), .Q(\EX_LS_typ [0] ), .QN(_08087_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q ( .D(_00117_ ), .CK(_07976_ ), .Q(\ID_EX_csr [11] ), .QN(_08086_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_1 ( .D(_00118_ ), .CK(_07976_ ), .Q(\ID_EX_csr [10] ), .QN(_08085_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_10 ( .D(_00119_ ), .CK(_07976_ ), .Q(\ID_EX_csr [1] ), .QN(_08084_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_11 ( .D(_00120_ ), .CK(_07976_ ), .Q(\ID_EX_csr [0] ), .QN(_08083_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_2 ( .D(_00121_ ), .CK(_07976_ ), .Q(\ID_EX_csr [9] ), .QN(_08082_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_3 ( .D(_00122_ ), .CK(_07976_ ), .Q(\ID_EX_csr [8] ), .QN(_08081_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_4 ( .D(_00123_ ), .CK(_07976_ ), .Q(\ID_EX_csr [7] ), .QN(_08080_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_5 ( .D(_00124_ ), .CK(_07976_ ), .Q(\ID_EX_csr [6] ), .QN(_08079_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_6 ( .D(_00125_ ), .CK(_07976_ ), .Q(\ID_EX_csr [5] ), .QN(_08078_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_7 ( .D(_00126_ ), .CK(_07976_ ), .Q(\ID_EX_csr [4] ), .QN(_08077_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_8 ( .D(_00127_ ), .CK(_07976_ ), .Q(\ID_EX_csr [3] ), .QN(_08076_ ) );
DFF_X1 \myidu.csr_$_SDFFE_PP0P__Q_9 ( .D(_00128_ ), .CK(_07976_ ), .Q(\ID_EX_csr [2] ), .QN(_08075_ ) );
DFF_X1 \myidu.exception_quest_IDU_$_SDFFE_PP0P__Q ( .D(_00129_ ), .CK(_07975_ ), .Q(exception_quest_IDU ), .QN(_08074_ ) );
DFF_X1 \myidu.fc_disenable_$_SDFFE_PP0P__Q ( .D(_00130_ ), .CK(_07974_ ), .Q(fc_disenable ), .QN(\myidu.fc_disenable_$_NOT__A_Y ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [31] ), .CK(_07973_ ), .Q(\ID_EX_imm [31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [30] ), .CK(_07973_ ), .Q(\ID_EX_imm [30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [21] ), .CK(_07973_ ), .Q(\ID_EX_imm [21] ), .QN(_08391_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [20] ), .CK(_07973_ ), .Q(\ID_EX_imm [20] ), .QN(_08392_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [19] ), .CK(_07973_ ), .Q(\ID_EX_imm [19] ), .QN(_08393_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [18] ), .CK(_07973_ ), .Q(\ID_EX_imm [18] ), .QN(_08394_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [17] ), .CK(_07973_ ), .Q(\ID_EX_imm [17] ), .QN(_08395_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [16] ), .CK(_07973_ ), .Q(\ID_EX_imm [16] ), .QN(_08396_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [15] ), .CK(_07973_ ), .Q(\ID_EX_imm [15] ), .QN(_08397_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [14] ), .CK(_07973_ ), .Q(\ID_EX_imm [14] ), .QN(_08398_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [13] ), .CK(_07973_ ), .Q(\ID_EX_imm [13] ), .QN(_08399_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [12] ), .CK(_07973_ ), .Q(\ID_EX_imm [12] ), .QN(_08400_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [29] ), .CK(_07973_ ), .Q(\ID_EX_imm [29] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [11] ), .CK(_07973_ ), .Q(\ID_EX_imm [11] ), .QN(_08401_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [10] ), .CK(_07973_ ), .Q(\ID_EX_imm [10] ), .QN(_08402_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [9] ), .CK(_07973_ ), .Q(\ID_EX_imm [9] ), .QN(_08403_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [8] ), .CK(_07973_ ), .Q(\ID_EX_imm [8] ), .QN(_08404_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [7] ), .CK(_07973_ ), .Q(\ID_EX_imm [7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [6] ), .CK(_07973_ ), .Q(\ID_EX_imm [6] ), .QN(_08405_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [5] ), .CK(_07973_ ), .Q(\ID_EX_imm [5] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [4] ), .CK(_07973_ ), .Q(\ID_EX_imm [4] ), .QN(_08406_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [3] ), .CK(_07973_ ), .Q(\ID_EX_imm [3] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_8_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [2] ), .CK(_07973_ ), .Q(\ID_EX_imm [2] ), .QN(_08407_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [28] ), .CK(_07973_ ), .Q(\ID_EX_imm [28] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_1_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [1] ), .CK(_07973_ ), .Q(\ID_EX_imm [1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_A_$_ANDNOT__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [0] ), .CK(_07973_ ), .Q(\ID_EX_imm [0] ), .QN(_08408_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [27] ), .CK(_07973_ ), .Q(\ID_EX_imm [27] ), .QN(_08409_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [26] ), .CK(_07973_ ), .Q(\ID_EX_imm [26] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_3_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [25] ), .CK(_07973_ ), .Q(\ID_EX_imm [25] ), .QN(_08410_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [24] ), .CK(_07973_ ), .Q(\ID_EX_imm [24] ), .QN(_08411_ ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [23] ), .CK(_07973_ ), .Q(\ID_EX_imm [23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_ANDNOT__B_A_$_OR__Y_B ) );
DFF_X1 \myidu.imm_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_OR__A_Y_$_OR__A_Y_$_OR__B_Y_$_MUX__B_Y [22] ), .CK(_07973_ ), .Q(\ID_EX_imm [22] ), .QN(_08412_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07972_ ), .Q(\ID_EX_pc [31] ), .QN(_08413_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07972_ ), .Q(\ID_EX_pc [30] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_1_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07972_ ), .Q(\ID_EX_pc [21] ), .QN(_08414_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07972_ ), .Q(\ID_EX_pc [20] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07972_ ), .Q(\ID_EX_pc [19] ), .QN(_08415_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07972_ ), .Q(\ID_EX_pc [18] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_13_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07972_ ), .Q(\ID_EX_pc [17] ), .QN(_08416_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07972_ ), .Q(\ID_EX_pc [16] ), .QN(_08417_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07972_ ), .Q(\ID_EX_pc [15] ), .QN(_08418_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07972_ ), .Q(\ID_EX_pc [14] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_17_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07972_ ), .Q(\ID_EX_pc [13] ), .QN(_08419_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07972_ ), .Q(\ID_EX_pc [12] ), .QN(_08420_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07972_ ), .Q(\ID_EX_pc [29] ), .QN(_08421_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07972_ ), .Q(\ID_EX_pc [11] ), .QN(_08422_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07972_ ), .Q(\ID_EX_pc [10] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_21_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07972_ ), .Q(\ID_EX_pc [9] ), .QN(_08423_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07972_ ), .Q(\ID_EX_pc [8] ), .QN(_08424_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07972_ ), .Q(\ID_EX_pc [7] ), .QN(_08425_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07972_ ), .Q(\ID_EX_pc [6] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_25_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07972_ ), .Q(\ID_EX_pc [5] ), .QN(_08426_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_27 ( .D(\IF_ID_pc [4] ), .CK(_07972_ ), .Q(\ID_EX_pc [4] ), .QN(_08427_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_28 ( .D(\IF_ID_pc [3] ), .CK(_07972_ ), .Q(\ID_EX_pc [3] ), .QN(_08428_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_29 ( .D(\IF_ID_pc [2] ), .CK(_07972_ ), .Q(\ID_EX_pc [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_29_D_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07972_ ), .Q(\ID_EX_pc [28] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_30 ( .D(\IF_ID_pc [1] ), .CK(_07972_ ), .Q(\ID_EX_pc [1] ), .QN(\myexu.pc_jump_$_DFFE_PP0P__Q_29_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_31 ( .D(\IF_ID_pc [0] ), .CK(_07972_ ), .Q(\ID_EX_pc [0] ), .QN(\myexu.pc_jump_$_DFFE_PP0P__Q_30_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07972_ ), .Q(\ID_EX_pc [27] ), .QN(_08429_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07972_ ), .Q(\ID_EX_pc [26] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07972_ ), .Q(\ID_EX_pc [25] ), .QN(_08430_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07972_ ), .Q(\ID_EX_pc [24] ), .QN(_08431_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07972_ ), .Q(\ID_EX_pc [23] ), .QN(_08432_ ) );
DFF_X1 \myidu.pc_out_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07972_ ), .Q(\ID_EX_pc [22] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_9_D_$_MUX__Y_A_$_MUX__Y_B_$_NOT__Y_A_$_XOR__Y_B ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q ( .D(_00131_ ), .CK(_07971_ ), .Q(\ID_EX_rd [4] ), .QN(_08073_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_1 ( .D(_00132_ ), .CK(_07971_ ), .Q(\ID_EX_rd [3] ), .QN(_08072_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_2 ( .D(_00133_ ), .CK(_07971_ ), .Q(\ID_EX_rd [2] ), .QN(_08071_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_3 ( .D(_00134_ ), .CK(_07971_ ), .Q(\ID_EX_rd [1] ), .QN(_08070_ ) );
DFF_X1 \myidu.rd_$_SDFFE_PP0P__Q_4 ( .D(_00135_ ), .CK(_07971_ ), .Q(\ID_EX_rd [0] ), .QN(_08069_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q ( .D(_00136_ ), .CK(_07970_ ), .Q(\ID_EX_rs1 [4] ), .QN(_08068_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1 ( .D(_00137_ ), .CK(_07970_ ), .Q(\ID_EX_rs1 [3] ), .QN(_08067_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00139_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08065_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2 ( .D(_00138_ ), .CK(_07970_ ), .Q(\ID_EX_rs1 [2] ), .QN(_08066_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00141_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08063_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3 ( .D(_00140_ ), .CK(_07970_ ), .Q(\ID_EX_rs1 [1] ), .QN(_08064_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00143_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08061_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4 ( .D(_00142_ ), .CK(_07970_ ), .Q(\ID_EX_rs1 [0] ), .QN(_08062_ ) );
DFF_X1 \myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00145_ ), .CK(clock ), .Q(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08059_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q ( .D(_00144_ ), .CK(_07969_ ), .Q(\ID_EX_rs2 [4] ), .QN(_08060_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1 ( .D(_00146_ ), .CK(_07969_ ), .Q(\ID_EX_rs2 [3] ), .QN(_08058_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_1_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00148_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .QN(_08056_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2 ( .D(_00147_ ), .CK(_07969_ ), .Q(\ID_EX_rs2 [2] ), .QN(_08057_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_2_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00150_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .QN(_08054_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3 ( .D(_00149_ ), .CK(_07969_ ), .Q(\ID_EX_rs2 [1] ), .QN(_08055_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_3_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00152_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08052_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4 ( .D(_00151_ ), .CK(_07969_ ), .Q(\ID_EX_rs2 [0] ), .QN(_08053_ ) );
DFF_X1 \myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00154_ ), .CK(clock ), .Q(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08050_ ) );
DFF_X1 \myidu.stall_quest_fencei_$_SDFFE_PP0P__Q ( .D(_00153_ ), .CK(_07968_ ), .Q(\myidu.stall_quest_fencei ), .QN(_08051_ ) );
DFF_X1 \myidu.stall_quest_loaduse_$_SDFFE_PP0P__Q ( .D(_00155_ ), .CK(_07967_ ), .Q(\myidu.stall_quest_loaduse ), .QN(_08049_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q ( .D(\myidu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myidu.state [2] ), .QN(_08434_ ) );
DFF_X1 \myidu.state_$_DFF_P__Q_1 ( .D(\myidu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(IDU_valid_EXU ), .QN(\myidu.exception_quest_IDU_$_SDFFE_PP0P__Q_D ) );
DFF_X1 \myidu.state_$_DFF_P__Q_2 ( .D(\myidu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(IDU_ready_IFU ), .QN(\myidu.fc_disenable_$_SDFFE_PP0P__Q_E_$_ANDNOT__Y_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q ( .D(_00156_ ), .CK(_07966_ ), .Q(\ID_EX_typ [7] ), .QN(_08433_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_1 ( .D(_00157_ ), .CK(_07966_ ), .Q(\ID_EX_typ [6] ), .QN(_08048_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_2 ( .D(_00158_ ), .CK(_07966_ ), .Q(\ID_EX_typ [5] ), .QN(_08047_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_3 ( .D(_00159_ ), .CK(_07966_ ), .Q(\ID_EX_typ [4] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_B_$_NOR__Y_B_$_OR__B_A_$_OR__A_Y_$_OR__A_B ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_4 ( .D(_00160_ ), .CK(_07966_ ), .Q(\ID_EX_typ [3] ), .QN(_08046_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_5 ( .D(_00161_ ), .CK(_07966_ ), .Q(\ID_EX_typ [2] ), .QN(\myexu.result_reg_$_DFFE_PP__Q_31_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_OR__Y_A_$_OR__Y_B_$_ANDNOT__Y_A_$_MUX__Y_A_$_NOR__Y_B_$_ANDNOT__B_1_A ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_6 ( .D(_00162_ ), .CK(_07966_ ), .Q(\ID_EX_typ [1] ), .QN(_08045_ ) );
DFF_X1 \myidu.typ_$_SDFFE_PP0P__Q_7 ( .D(_00163_ ), .CK(_07966_ ), .Q(\ID_EX_typ [0] ), .QN(\myexu.check_quest_$_DFF_PP0__Q_D_$_ANDNOT__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.check_assert_$_DFFE_PP__Q ( .D(\myifu.state [1] ), .CK(_07965_ ), .Q(check_assert ), .QN(_08435_ ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [31] ), .CK(_07964_ ), .Q(\IF_ID_inst [31] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_17_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_1 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [30] ), .CK(_07964_ ), .Q(\IF_ID_inst [30] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_20_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_10 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [21] ), .CK(_07964_ ), .Q(\IF_ID_inst [21] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_10_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_11 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [20] ), .CK(_07964_ ), .Q(\IF_ID_inst [20] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_11_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_12 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [19] ), .CK(_07964_ ), .Q(\IF_ID_inst [19] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_12_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_13 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [18] ), .CK(_07964_ ), .Q(\IF_ID_inst [18] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_13_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_14 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [17] ), .CK(_07964_ ), .Q(\IF_ID_inst [17] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_14_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_15 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [16] ), .CK(_07964_ ), .Q(\IF_ID_inst [16] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_15_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_16 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [15] ), .CK(_07964_ ), .Q(\IF_ID_inst [15] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_16_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_17 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [14] ), .CK(_07964_ ), .Q(\IF_ID_inst [14] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_17_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_18 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [13] ), .CK(_07964_ ), .Q(\IF_ID_inst [13] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_18_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_19 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [12] ), .CK(_07964_ ), .Q(\IF_ID_inst [12] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_19_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_2 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [29] ), .CK(_07964_ ), .Q(\IF_ID_inst [29] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_21_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_20 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [11] ), .CK(_07964_ ), .Q(\IF_ID_inst [11] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_NOR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_21 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [10] ), .CK(_07964_ ), .Q(\IF_ID_inst [10] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_22 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [9] ), .CK(_07964_ ), .Q(\IF_ID_inst [9] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_23 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [8] ), .CK(_07964_ ), .Q(\IF_ID_inst [8] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_24 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [7] ), .CK(_07964_ ), .Q(\IF_ID_inst [7] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_19_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_25 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [6] ), .CK(_07964_ ), .Q(\IF_ID_inst [6] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_24_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_26 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [5] ), .CK(_07964_ ), .Q(\IF_ID_inst [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_25_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_27 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [4] ), .CK(_07964_ ), .Q(\IF_ID_inst [4] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_26_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_28 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [3] ), .CK(_07964_ ), .Q(\IF_ID_inst [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_27_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_29 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [2] ), .CK(_07964_ ), .Q(\IF_ID_inst [2] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_28_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_3 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [28] ), .CK(_07964_ ), .Q(\IF_ID_inst [28] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__A_Y_$_OR__A_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_30 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [1] ), .CK(_07964_ ), .Q(\IF_ID_inst [1] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_29_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_31 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [0] ), .CK(_07964_ ), .Q(\IF_ID_inst [0] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_30_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_4 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [27] ), .CK(_07964_ ), .Q(\IF_ID_inst [27] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_23_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_ORNOT__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_5 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [26] ), .CK(_07964_ ), .Q(\IF_ID_inst [26] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_24_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_NOR__Y_B_$_ANDNOT__Y_B_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_6 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [25] ), .CK(_07964_ ), .Q(\IF_ID_inst [25] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_A_$_MUX__Y_B ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_7 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [24] ), .CK(_07964_ ), .Q(\IF_ID_inst [24] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_7_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_8 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [23] ), .CK(_07964_ ), .Q(\IF_ID_inst [23] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y_$_MUX__Y_8_A_$_ANDNOT__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myifu.inst_$_DFFE_PP__Q_9 ( .D(\myifu.pc_$_SDFFE_PP0P__Q_30_D_$_MUX__Y_A_$_MUX__Y_A_$_XNOR__Y_A_$_MUX__Y_B_$_MUX__A_Y_$_MUX__B_Y_$_ANDNOT__B_Y_$_MUX__A_Y [22] ), .CK(_07964_ ), .Q(\IF_ID_inst [22] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_29_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_B_$_XNOR__Y_A_$_MUX__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][31] ), .QN(_08436_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][30] ), .QN(_08437_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][21] ), .QN(_08438_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][20] ), .QN(_08439_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][19] ), .QN(_08440_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][18] ), .QN(_08441_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][17] ), .QN(_08442_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][16] ), .QN(_08443_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][15] ), .QN(_08444_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][14] ), .QN(_08445_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][13] ), .QN(_08446_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][12] ), .QN(_08447_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][29] ), .QN(_08448_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][11] ), .QN(_08449_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][10] ), .QN(_08450_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][9] ), .QN(_08451_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][8] ), .QN(_08452_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][7] ), .QN(_08453_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][6] ), .QN(_08454_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][5] ), .QN(_08455_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][4] ), .QN(_08456_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][3] ), .QN(_08457_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][2] ), .QN(_08458_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][28] ), .QN(_08459_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][1] ), .QN(_08460_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][0] ), .QN(_08461_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][27] ), .QN(_08462_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][26] ), .QN(_08463_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][25] ), .QN(_08464_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][24] ), .QN(_08465_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][23] ), .QN(_08466_ ) );
DFF_X1 \myifu.myicache.data[0]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07963_ ), .Q(\myifu.myicache.data[0][22] ), .QN(_08467_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][31] ), .QN(_08468_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][30] ), .QN(_08469_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][21] ), .QN(_08470_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][20] ), .QN(_08471_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][19] ), .QN(_08472_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][18] ), .QN(_08473_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][17] ), .QN(_08474_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][16] ), .QN(_08475_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][15] ), .QN(_08476_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][14] ), .QN(_08477_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][13] ), .QN(_08478_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][12] ), .QN(_08479_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][29] ), .QN(_08480_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][11] ), .QN(_08481_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][10] ), .QN(_08482_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][9] ), .QN(_08483_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][8] ), .QN(_08484_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][7] ), .QN(_08485_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][6] ), .QN(_08486_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][5] ), .QN(_08487_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][4] ), .QN(_08488_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][3] ), .QN(_08489_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][2] ), .QN(_08490_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][28] ), .QN(_08491_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][1] ), .QN(_08492_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][0] ), .QN(_08493_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][27] ), .QN(_08494_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][26] ), .QN(_08495_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][25] ), .QN(_08496_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][24] ), .QN(_08497_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][23] ), .QN(_08498_ ) );
DFF_X1 \myifu.myicache.data[1]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07962_ ), .Q(\myifu.myicache.data[1][22] ), .QN(_08499_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][31] ), .QN(_08500_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][30] ), .QN(_08501_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][21] ), .QN(_08502_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][20] ), .QN(_08503_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][19] ), .QN(_08504_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][18] ), .QN(_08505_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][17] ), .QN(_08506_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][16] ), .QN(_08507_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][15] ), .QN(_08508_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][14] ), .QN(_08509_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][13] ), .QN(_08510_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][12] ), .QN(_08511_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][29] ), .QN(_08512_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][11] ), .QN(_08513_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][10] ), .QN(_08514_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][9] ), .QN(_08515_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][8] ), .QN(_08516_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][7] ), .QN(_08517_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][6] ), .QN(_08518_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][5] ), .QN(_08519_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][4] ), .QN(_08520_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][3] ), .QN(_08521_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][2] ), .QN(_08522_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][28] ), .QN(_08523_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][1] ), .QN(_08524_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][0] ), .QN(_08525_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][27] ), .QN(_08526_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][26] ), .QN(_08527_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][25] ), .QN(_08528_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][24] ), .QN(_08529_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][23] ), .QN(_08530_ ) );
DFF_X1 \myifu.myicache.data[2]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07961_ ), .Q(\myifu.myicache.data[2][22] ), .QN(_08531_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][31] ), .QN(_08532_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][30] ), .QN(_08533_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][21] ), .QN(_08534_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][20] ), .QN(_08535_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][19] ), .QN(_08536_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][18] ), .QN(_08537_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][17] ), .QN(_08538_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][16] ), .QN(_08539_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][15] ), .QN(_08540_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][14] ), .QN(_08541_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][13] ), .QN(_08542_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][12] ), .QN(_08543_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][29] ), .QN(_08544_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][11] ), .QN(_08545_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][10] ), .QN(_08546_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][9] ), .QN(_08547_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][8] ), .QN(_08548_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][7] ), .QN(_08549_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][6] ), .QN(_08550_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][5] ), .QN(_08551_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][4] ), .QN(_08552_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][3] ), .QN(_08553_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][2] ), .QN(_08554_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][28] ), .QN(_08555_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][1] ), .QN(_08556_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][0] ), .QN(_08557_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][27] ), .QN(_08558_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][26] ), .QN(_08559_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][25] ), .QN(_08560_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][24] ), .QN(_08561_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][23] ), .QN(_08562_ ) );
DFF_X1 \myifu.myicache.data[3]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07960_ ), .Q(\myifu.myicache.data[3][22] ), .QN(_08563_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][31] ), .QN(_08564_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][30] ), .QN(_08565_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][21] ), .QN(_08566_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][20] ), .QN(_08567_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][19] ), .QN(_08568_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][18] ), .QN(_08569_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][17] ), .QN(_08570_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][16] ), .QN(_08571_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][15] ), .QN(_08572_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][14] ), .QN(_08573_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][13] ), .QN(_08574_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][12] ), .QN(_08575_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][29] ), .QN(_08576_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][11] ), .QN(_08577_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][10] ), .QN(_08578_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][9] ), .QN(_08579_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][8] ), .QN(_08580_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][7] ), .QN(_08581_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][6] ), .QN(_08582_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][5] ), .QN(_08583_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][4] ), .QN(_08584_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][3] ), .QN(_08585_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][2] ), .QN(_08586_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][28] ), .QN(_08587_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][1] ), .QN(_08588_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][0] ), .QN(_08589_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][27] ), .QN(_08590_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][26] ), .QN(_08591_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][25] ), .QN(_08592_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][24] ), .QN(_08593_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][23] ), .QN(_08594_ ) );
DFF_X1 \myifu.myicache.data[4]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07959_ ), .Q(\myifu.myicache.data[4][22] ), .QN(_08595_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][31] ), .QN(_08596_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][30] ), .QN(_08597_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][21] ), .QN(_08598_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][20] ), .QN(_08599_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][19] ), .QN(_08600_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][18] ), .QN(_08601_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][17] ), .QN(_08602_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][16] ), .QN(_08603_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][15] ), .QN(_08604_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][14] ), .QN(_08605_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][13] ), .QN(_08606_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][12] ), .QN(_08607_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][29] ), .QN(_08608_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][11] ), .QN(_08609_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][10] ), .QN(_08610_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][9] ), .QN(_08611_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][8] ), .QN(_08612_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][7] ), .QN(_08613_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][6] ), .QN(_08614_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][5] ), .QN(_08615_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][4] ), .QN(_08616_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][3] ), .QN(_08617_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][2] ), .QN(_08618_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][28] ), .QN(_08619_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][1] ), .QN(_08620_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][0] ), .QN(_08621_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][27] ), .QN(_08622_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][26] ), .QN(_08623_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][25] ), .QN(_08624_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][24] ), .QN(_08625_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][23] ), .QN(_08626_ ) );
DFF_X1 \myifu.myicache.data[5]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07958_ ), .Q(\myifu.myicache.data[5][22] ), .QN(_08627_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][31] ), .QN(_08628_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][30] ), .QN(_08629_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][21] ), .QN(_08630_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][20] ), .QN(_08631_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][19] ), .QN(_08632_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][18] ), .QN(_08633_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][17] ), .QN(_08634_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][16] ), .QN(_08635_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][15] ), .QN(_08636_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][14] ), .QN(_08637_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][13] ), .QN(_08638_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][12] ), .QN(_08639_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][29] ), .QN(_08640_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][11] ), .QN(_08641_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][10] ), .QN(_08642_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][9] ), .QN(_08643_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][8] ), .QN(_08644_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][7] ), .QN(_08645_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][6] ), .QN(_08646_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][5] ), .QN(_08647_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][4] ), .QN(_08648_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][3] ), .QN(_08649_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][2] ), .QN(_08650_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][28] ), .QN(_08651_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][1] ), .QN(_08652_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][0] ), .QN(_08653_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][27] ), .QN(_08654_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][26] ), .QN(_08655_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][25] ), .QN(_08656_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][24] ), .QN(_08657_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][23] ), .QN(_08658_ ) );
DFF_X1 \myifu.myicache.data[6]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07957_ ), .Q(\myifu.myicache.data[6][22] ), .QN(_08659_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q ( .D(\myifu.data_in [31] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][31] ), .QN(_08660_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_1 ( .D(\myifu.data_in [30] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][30] ), .QN(_08661_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_10 ( .D(\myifu.data_in [21] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][21] ), .QN(_08662_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_11 ( .D(\myifu.data_in [20] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][20] ), .QN(_08663_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_12 ( .D(\myifu.data_in [19] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][19] ), .QN(_08664_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_13 ( .D(\myifu.data_in [18] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][18] ), .QN(_08665_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_14 ( .D(\myifu.data_in [17] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][17] ), .QN(_08666_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_15 ( .D(\myifu.data_in [16] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][16] ), .QN(_08667_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_16 ( .D(\myifu.data_in [15] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][15] ), .QN(_08668_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_17 ( .D(\myifu.data_in [14] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][14] ), .QN(_08669_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_18 ( .D(\myifu.data_in [13] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][13] ), .QN(_08670_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_19 ( .D(\myifu.data_in [12] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][12] ), .QN(_08671_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_2 ( .D(\myifu.data_in [29] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][29] ), .QN(_08672_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_20 ( .D(\myifu.data_in [11] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][11] ), .QN(_08673_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_21 ( .D(\myifu.data_in [10] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][10] ), .QN(_08674_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_22 ( .D(\myifu.data_in [9] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][9] ), .QN(_08675_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_23 ( .D(\myifu.data_in [8] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][8] ), .QN(_08676_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_24 ( .D(\myifu.data_in [7] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][7] ), .QN(_08677_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_25 ( .D(\myifu.data_in [6] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][6] ), .QN(_08678_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_26 ( .D(\myifu.data_in [5] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][5] ), .QN(_08679_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_27 ( .D(\myifu.data_in [4] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][4] ), .QN(_08680_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_28 ( .D(\myifu.data_in [3] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][3] ), .QN(_08681_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_29 ( .D(\myifu.data_in [2] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][2] ), .QN(_08682_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_3 ( .D(\myifu.data_in [28] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][28] ), .QN(_08683_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_30 ( .D(\myifu.data_in [1] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][1] ), .QN(_08684_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_31 ( .D(\myifu.data_in [0] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][0] ), .QN(_08685_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_4 ( .D(\myifu.data_in [27] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][27] ), .QN(_08686_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_5 ( .D(\myifu.data_in [26] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][26] ), .QN(_08687_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_6 ( .D(\myifu.data_in [25] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][25] ), .QN(_08688_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_7 ( .D(\myifu.data_in [24] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][24] ), .QN(_08689_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_8 ( .D(\myifu.data_in [23] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][23] ), .QN(_08690_ ) );
DFF_X1 \myifu.myicache.data[7]_$_DFFE_PP__Q_9 ( .D(\myifu.data_in [22] ), .CK(_07956_ ), .Q(\myifu.myicache.data[7][22] ), .QN(_08691_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][26] ), .QN(_08692_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][25] ), .QN(_08693_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][16] ), .QN(_08694_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][15] ), .QN(_08695_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][14] ), .QN(_08696_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][13] ), .QN(_08697_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][12] ), .QN(_08698_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][11] ), .QN(_08699_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][10] ), .QN(_08700_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][9] ), .QN(_08701_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][8] ), .QN(_08702_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][7] ), .QN(_08703_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][24] ), .QN(_08704_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][6] ), .QN(_08705_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][5] ), .QN(_08706_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][4] ), .QN(_08707_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][3] ), .QN(_08708_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][2] ), .QN(_08709_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][1] ), .QN(_08710_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][0] ), .QN(_08711_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][23] ), .QN(_08712_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][22] ), .QN(_08713_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][21] ), .QN(_08714_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][20] ), .QN(_08715_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][19] ), .QN(_08716_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][18] ), .QN(_08717_ ) );
DFF_X1 \myifu.myicache.tag[0]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07955_ ), .Q(\myifu.myicache.tag[0][17] ), .QN(_08718_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][26] ), .QN(_08719_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][25] ), .QN(_08720_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][16] ), .QN(_08721_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][15] ), .QN(_08722_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][14] ), .QN(_08723_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][13] ), .QN(_08724_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][12] ), .QN(_08725_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][11] ), .QN(_08726_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][10] ), .QN(_08727_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][9] ), .QN(_08728_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][8] ), .QN(_08729_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][7] ), .QN(_08730_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][24] ), .QN(_08731_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][6] ), .QN(_08732_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][5] ), .QN(_08733_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][4] ), .QN(_08734_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][3] ), .QN(_08735_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][2] ), .QN(_08736_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][1] ), .QN(_08737_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][0] ), .QN(_08738_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][23] ), .QN(_08739_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][22] ), .QN(_08740_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][21] ), .QN(_08741_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][20] ), .QN(_08742_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][19] ), .QN(_08743_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][18] ), .QN(_08744_ ) );
DFF_X1 \myifu.myicache.tag[1]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07954_ ), .Q(\myifu.myicache.tag[1][17] ), .QN(_08745_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][26] ), .QN(_08746_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][25] ), .QN(_08747_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][16] ), .QN(_08748_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][15] ), .QN(_08749_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][14] ), .QN(_08750_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][13] ), .QN(_08751_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][12] ), .QN(_08752_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][11] ), .QN(_08753_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][10] ), .QN(_08754_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][9] ), .QN(_08755_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][8] ), .QN(_08756_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][7] ), .QN(_08757_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][24] ), .QN(_08758_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][6] ), .QN(_08759_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][5] ), .QN(_08760_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][4] ), .QN(_08761_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][3] ), .QN(_08762_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][2] ), .QN(_08763_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][1] ), .QN(_08764_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][0] ), .QN(_08765_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][23] ), .QN(_08766_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][22] ), .QN(_08767_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][21] ), .QN(_08768_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][20] ), .QN(_08769_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][19] ), .QN(_08770_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][18] ), .QN(_08771_ ) );
DFF_X1 \myifu.myicache.tag[2]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07953_ ), .Q(\myifu.myicache.tag[2][17] ), .QN(_08772_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q ( .D(\IF_ID_pc [31] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][26] ), .QN(_08773_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_1 ( .D(\IF_ID_pc [30] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][25] ), .QN(_08774_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_10 ( .D(\IF_ID_pc [21] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][16] ), .QN(_08775_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_11 ( .D(\IF_ID_pc [20] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][15] ), .QN(_08776_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_12 ( .D(\IF_ID_pc [19] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][14] ), .QN(_08777_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_13 ( .D(\IF_ID_pc [18] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][13] ), .QN(_08778_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_14 ( .D(\IF_ID_pc [17] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][12] ), .QN(_08779_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_15 ( .D(\IF_ID_pc [16] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][11] ), .QN(_08780_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_16 ( .D(\IF_ID_pc [15] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][10] ), .QN(_08781_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_17 ( .D(\IF_ID_pc [14] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][9] ), .QN(_08782_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_18 ( .D(\IF_ID_pc [13] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][8] ), .QN(_08783_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_19 ( .D(\IF_ID_pc [12] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][7] ), .QN(_08784_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_2 ( .D(\IF_ID_pc [29] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][24] ), .QN(_08785_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_20 ( .D(\IF_ID_pc [11] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][6] ), .QN(_08786_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_21 ( .D(\IF_ID_pc [10] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][5] ), .QN(_08787_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_22 ( .D(\IF_ID_pc [9] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][4] ), .QN(_08788_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_23 ( .D(\IF_ID_pc [8] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][3] ), .QN(_08789_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_24 ( .D(\IF_ID_pc [7] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][2] ), .QN(_08790_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_25 ( .D(\IF_ID_pc [6] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][1] ), .QN(_08791_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_26 ( .D(\IF_ID_pc [5] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][0] ), .QN(_08792_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_3 ( .D(\IF_ID_pc [28] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][23] ), .QN(_08793_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_4 ( .D(\IF_ID_pc [27] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][22] ), .QN(_08794_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_5 ( .D(\IF_ID_pc [26] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][21] ), .QN(_08795_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_6 ( .D(\IF_ID_pc [25] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][20] ), .QN(_08796_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_7 ( .D(\IF_ID_pc [24] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][19] ), .QN(_08797_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_8 ( .D(\IF_ID_pc [23] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][18] ), .QN(_08798_ ) );
DFF_X1 \myifu.myicache.tag[3]_$_DFFE_PP__Q_9 ( .D(\IF_ID_pc [22] ), .CK(_07952_ ), .Q(\myifu.myicache.tag[3][17] ), .QN(_08044_ ) );
DFF_X1 \myifu.myicache.valid[0]_$_SDFFCE_PN0P__Q ( .D(_00164_ ), .CK(_07951_ ), .Q(\myifu.myicache.valid [0] ), .QN(_08043_ ) );
DFF_X1 \myifu.myicache.valid[1]_$_SDFFCE_PN0P__Q ( .D(_00165_ ), .CK(_07950_ ), .Q(\myifu.myicache.valid [1] ), .QN(_08042_ ) );
DFF_X1 \myifu.myicache.valid[2]_$_SDFFCE_PN0P__Q ( .D(_00166_ ), .CK(_07949_ ), .Q(\myifu.myicache.valid [2] ), .QN(_08799_ ) );
DFF_X1 \myifu.myicache.valid[3]_$_DFFE_PP__Q ( .D(\myifu.wen_$_ANDNOT__A_Y ), .CK(_07948_ ), .Q(\myifu.myicache.valid [3] ), .QN(_08041_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q ( .D(_00167_ ), .CK(_07947_ ), .Q(\IF_ID_pc [0] ), .QN(\myifu.tmp_offset_$_XOR__B_Y_$_ANDNOT__B_A_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_1 ( .D(_00168_ ), .CK(_07946_ ), .Q(\IF_ID_pc [30] ), .QN(_08040_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_10 ( .D(_00169_ ), .CK(_07946_ ), .Q(\IF_ID_pc [21] ), .QN(_08039_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_11 ( .D(_00170_ ), .CK(_07946_ ), .Q(\IF_ID_pc [20] ), .QN(_08038_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_12 ( .D(_00171_ ), .CK(_07946_ ), .Q(\IF_ID_pc [19] ), .QN(_08037_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_13 ( .D(_00172_ ), .CK(_07946_ ), .Q(\IF_ID_pc [18] ), .QN(_08036_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_14 ( .D(_00173_ ), .CK(_07946_ ), .Q(\IF_ID_pc [17] ), .QN(_08035_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_15 ( .D(_00174_ ), .CK(_07946_ ), .Q(\IF_ID_pc [16] ), .QN(_08034_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_16 ( .D(_00175_ ), .CK(_07946_ ), .Q(\IF_ID_pc [15] ), .QN(_08033_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_17 ( .D(_00176_ ), .CK(_07946_ ), .Q(\IF_ID_pc [14] ), .QN(_08032_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_18 ( .D(_00177_ ), .CK(_07946_ ), .Q(\IF_ID_pc [13] ), .QN(_08031_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_19 ( .D(_00178_ ), .CK(_07946_ ), .Q(\IF_ID_pc [12] ), .QN(_08030_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_2 ( .D(_00179_ ), .CK(_07946_ ), .Q(\IF_ID_pc [29] ), .QN(_08029_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_20 ( .D(_00180_ ), .CK(_07946_ ), .Q(\IF_ID_pc [11] ), .QN(_08028_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_21 ( .D(_00181_ ), .CK(_07946_ ), .Q(\IF_ID_pc [10] ), .QN(_08027_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_22 ( .D(_00182_ ), .CK(_07946_ ), .Q(\IF_ID_pc [9] ), .QN(_08026_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_23 ( .D(_00183_ ), .CK(_07946_ ), .Q(\IF_ID_pc [8] ), .QN(_08025_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_24 ( .D(_00184_ ), .CK(_07946_ ), .Q(\IF_ID_pc [7] ), .QN(_08024_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_25 ( .D(_00185_ ), .CK(_07946_ ), .Q(\IF_ID_pc [6] ), .QN(_08023_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_26 ( .D(_00186_ ), .CK(_07946_ ), .Q(\IF_ID_pc [5] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_25_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27 ( .D(_00187_ ), .CK(_07946_ ), .Q(\IF_ID_pc [4] ), .QN(_08022_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00189_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .QN(_08021_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28 ( .D(_00188_ ), .CK(_07946_ ), .Q(\IF_ID_pc [3] ), .QN(\myifu.pc_$_SDFFE_PP0P__Q_27_D_$_MUX__Y_A_$_MUX__Y_A_$_XOR__Y_A_$_ANDNOT__Y_A_$_OR__Y_B ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D ( .D(_00191_ ), .CK(clock ), .Q(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .QN(_08019_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_29 ( .D(_00190_ ), .CK(_07946_ ), .Q(\IF_ID_pc [2] ), .QN(_08020_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_3 ( .D(_00192_ ), .CK(_07946_ ), .Q(\IF_ID_pc [28] ), .QN(_08018_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_30 ( .D(_00193_ ), .CK(_07946_ ), .Q(\IF_ID_pc [1] ), .QN(_08017_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_4 ( .D(_00194_ ), .CK(_07946_ ), .Q(\IF_ID_pc [27] ), .QN(_08016_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_5 ( .D(_00195_ ), .CK(_07946_ ), .Q(\IF_ID_pc [26] ), .QN(_08015_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_6 ( .D(_00196_ ), .CK(_07946_ ), .Q(\IF_ID_pc [25] ), .QN(_08014_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_7 ( .D(_00197_ ), .CK(_07946_ ), .Q(\IF_ID_pc [24] ), .QN(_08013_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_8 ( .D(_00198_ ), .CK(_07946_ ), .Q(\IF_ID_pc [23] ), .QN(_08012_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP0P__Q_9 ( .D(_00199_ ), .CK(_07946_ ), .Q(\IF_ID_pc [22] ), .QN(_08011_ ) );
DFF_X1 \myifu.pc_$_SDFFE_PP1P__Q ( .D(_00200_ ), .CK(_07946_ ), .Q(\IF_ID_pc [31] ), .QN(_08010_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q ( .D(\myifu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myifu.state [2] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_B_$_ANDNOT__Y_A ) );
DFF_X1 \myifu.state_$_DFF_P__Q_1 ( .D(\myifu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myifu.state [1] ), .QN(_08801_ ) );
DFF_X1 \myifu.state_$_DFF_P__Q_2 ( .D(\myifu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\myifu.state [0] ), .QN(_08009_ ) );
DFF_X1 \myifu.tmp_offset_$_SDFFE_PP0P__Q ( .D(_00201_ ), .CK(_07945_ ), .Q(\myifu.tmp_offset [2] ), .QN(_08800_ ) );
DFF_X1 \myifu.to_reset_$_SDFF_PP0__Q ( .D(_00203_ ), .CK(clock ), .Q(\myifu.to_reset ), .QN(\myifu.to_reset_$_SDFF_PP0__Q_D_$_MUX__Y_A_$_NAND__Y_B ) );
DFF_X1 \myifu.wen_$_SDFFE_PP0P__Q ( .D(_00202_ ), .CK(_07944_ ), .Q(\myifu.myicache.valid_data_in ), .QN(_08008_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [31] ), .QN(_08802_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [30] ), .QN(_08803_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [21] ), .QN(_08804_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [20] ), .QN(_08805_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [19] ), .QN(_08806_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [18] ), .QN(_08807_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [17] ), .QN(_08808_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [16] ), .QN(_08809_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [15] ), .QN(_08810_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [14] ), .QN(_08811_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [13] ), .QN(_08812_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [12] ), .QN(_08813_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [29] ), .QN(_08814_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [11] ), .QN(_08815_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [10] ), .QN(_08816_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [9] ), .QN(_08817_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [8] ), .QN(_08818_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [7] ), .QN(_08819_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [6] ), .QN(_08820_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [5] ), .QN(_08821_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [4] ), .QN(_08822_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [3] ), .QN(_08823_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [2] ), .QN(_08824_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [28] ), .QN(_08825_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [1] ), .QN(_08826_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [0] ), .QN(_08827_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [27] ), .QN(_08828_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [26] ), .QN(_08829_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [25] ), .QN(_08830_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [24] ), .QN(_08831_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [23] ), .QN(_08832_ ) );
DFF_X1 \mylsu.araddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07943_ ), .Q(\mylsu.araddr_tmp [22] ), .QN(_08833_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q ( .D(\EX_LS_dest_csreg_mem [31] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [31] ), .QN(_08834_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_csreg_mem [30] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [30] ), .QN(_08835_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_10 ( .D(\EX_LS_dest_csreg_mem [21] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [21] ), .QN(_08836_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_11 ( .D(\EX_LS_dest_csreg_mem [20] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [20] ), .QN(_08837_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_12 ( .D(\EX_LS_dest_csreg_mem [19] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [19] ), .QN(_08838_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_13 ( .D(\EX_LS_dest_csreg_mem [18] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [18] ), .QN(_08839_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_14 ( .D(\EX_LS_dest_csreg_mem [17] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [17] ), .QN(_08840_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_15 ( .D(\EX_LS_dest_csreg_mem [16] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [16] ), .QN(_08841_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_16 ( .D(\EX_LS_dest_csreg_mem [15] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [15] ), .QN(_08842_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_17 ( .D(\EX_LS_dest_csreg_mem [14] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [14] ), .QN(_08843_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_18 ( .D(\EX_LS_dest_csreg_mem [13] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [13] ), .QN(_08844_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_19 ( .D(\EX_LS_dest_csreg_mem [12] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [12] ), .QN(_08845_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_csreg_mem [29] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [29] ), .QN(_08846_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_20 ( .D(\EX_LS_dest_csreg_mem [11] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [11] ), .QN(_08847_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_21 ( .D(\EX_LS_dest_csreg_mem [10] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [10] ), .QN(_08848_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_22 ( .D(\EX_LS_dest_csreg_mem [9] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [9] ), .QN(_08849_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_23 ( .D(\EX_LS_dest_csreg_mem [8] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [8] ), .QN(_08850_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_24 ( .D(\EX_LS_dest_csreg_mem [7] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [7] ), .QN(_08851_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_25 ( .D(\EX_LS_dest_csreg_mem [6] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [6] ), .QN(_08852_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_26 ( .D(\EX_LS_dest_csreg_mem [5] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [5] ), .QN(_08853_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_27 ( .D(\EX_LS_dest_csreg_mem [4] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [4] ), .QN(_08854_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_28 ( .D(\EX_LS_dest_csreg_mem [3] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [3] ), .QN(_08855_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_29 ( .D(\EX_LS_dest_csreg_mem [2] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [2] ), .QN(_08856_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_csreg_mem [28] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [28] ), .QN(_08857_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_30 ( .D(\EX_LS_dest_csreg_mem [1] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [1] ), .QN(_08858_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_31 ( .D(\EX_LS_dest_csreg_mem [0] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [0] ), .QN(_08859_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_4 ( .D(\EX_LS_dest_csreg_mem [27] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [27] ), .QN(_08860_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_5 ( .D(\EX_LS_dest_csreg_mem [26] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [26] ), .QN(_08861_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_6 ( .D(\EX_LS_dest_csreg_mem [25] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [25] ), .QN(_08862_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_7 ( .D(\EX_LS_dest_csreg_mem [24] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [24] ), .QN(_08863_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_8 ( .D(\EX_LS_dest_csreg_mem [23] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [23] ), .QN(_08864_ ) );
DFF_X1 \mylsu.awaddr_tmp_$_DFFE_PP__Q_9 ( .D(\EX_LS_dest_csreg_mem [22] ), .CK(_07942_ ), .Q(\mylsu.awaddr_tmp [22] ), .QN(_08007_ ) );
DFF_X1 \mylsu.pc_out_$_SDFFE_PP0P__Q ( .D(_00204_ ), .CK(_07941_ ), .Q(LS_WB_pc ), .QN(_08006_ ) );
DFF_X1 \mylsu.previous_load_done_$_SDFFE_PP0P__Q ( .D(_00205_ ), .CK(_07940_ ), .Q(\mylsu.previous_load_done ), .QN(_08865_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q ( .D(\mylsu.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mylsu.state [4] ), .QN(_08866_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_1 ( .D(\mylsu.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mylsu.state [3] ), .QN(io_master_rready_$_ANDNOT__Y_B_$_MUX__Y_A_$_OR__Y_A_$_ANDNOT__Y_A ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_2 ( .D(\mylsu.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mylsu.state [2] ), .QN(_08867_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_3 ( .D(\mylsu.state_$_DFF_P__Q_3_D ), .CK(clock ), .Q(\mylsu.state [1] ), .QN(_08868_ ) );
DFF_X1 \mylsu.state_$_DFF_P__Q_4 ( .D(\mylsu.state_$_DFF_P__Q_4_D ), .CK(clock ), .Q(\mylsu.state [0] ), .QN(io_master_wready_$_NOR__B_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q ( .D(\EX_LS_typ [2] ), .CK(_07943_ ), .Q(\mylsu.typ_tmp [2] ), .QN(\mylsu.typ_tmp_$_NOT__A_Y ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_1 ( .D(\EX_LS_typ [1] ), .CK(_07943_ ), .Q(\mylsu.typ_tmp [1] ), .QN(_08869_ ) );
DFF_X1 \mylsu.typ_tmp_$_DFFE_PP__Q_2 ( .D(\EX_LS_typ [0] ), .CK(_07943_ ), .Q(\mylsu.typ_tmp [0] ), .QN(_08005_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q ( .D(_00206_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [11] ), .QN(_08004_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_1 ( .D(_00207_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [10] ), .QN(_08003_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_2 ( .D(_00208_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [7] ), .QN(_08002_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_3 ( .D(_00209_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [5] ), .QN(_08001_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_4 ( .D(_00210_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [4] ), .QN(_08000_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_5 ( .D(_00211_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [3] ), .QN(_07999_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_6 ( .D(_00212_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [2] ), .QN(_07998_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP0P__Q_7 ( .D(_00213_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [1] ), .QN(_07997_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q ( .D(_00214_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [9] ), .QN(_07996_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_1 ( .D(_00215_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [8] ), .QN(_07995_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_2 ( .D(_00216_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [6] ), .QN(_07994_ ) );
DFF_X1 \mylsu.waddr_csreg_$_SDFFCE_PP1P__Q_3 ( .D(_00217_ ), .CK(_07943_ ), .Q(\LS_WB_waddr_csreg [0] ), .QN(_08870_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q ( .D(\EX_LS_dest_reg [3] ), .CK(_07943_ ), .Q(\LS_WB_waddr_reg [3] ), .QN(_08871_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_1 ( .D(\EX_LS_dest_reg [2] ), .CK(_07943_ ), .Q(\LS_WB_waddr_reg [2] ), .QN(_08872_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_2 ( .D(\EX_LS_dest_reg [1] ), .CK(_07943_ ), .Q(\LS_WB_waddr_reg [1] ), .QN(_08873_ ) );
DFF_X1 \mylsu.waddr_reg_$_DFFE_PP__Q_3 ( .D(\EX_LS_dest_reg [0] ), .CK(_07943_ ), .Q(\LS_WB_waddr_reg [0] ), .QN(_08874_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [31] ), .QN(_08875_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_1_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [30] ), .QN(_08876_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_10_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [21] ), .QN(_08877_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_11_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [20] ), .QN(_08878_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_12_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [19] ), .QN(_08879_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_13_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [18] ), .QN(_08880_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_14_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [17] ), .QN(_08881_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_15_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [16] ), .QN(_08882_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_16_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [15] ), .QN(_08883_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_17_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [14] ), .QN(_08884_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_18_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [13] ), .QN(_08885_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_19_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [12] ), .QN(_08886_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_2_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [29] ), .QN(_08887_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_20_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [11] ), .QN(_08888_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_21_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [10] ), .QN(_08889_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_22_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [9] ), .QN(_08890_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_23_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [8] ), .QN(_08891_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_24_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [7] ), .QN(_08892_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_25_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [6] ), .QN(_08893_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_26_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [5] ), .QN(_08894_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_27_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [4] ), .QN(_08895_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_28_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [3] ), .QN(_08896_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_29_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [2] ), .QN(_08897_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_3_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [28] ), .QN(_08898_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_30_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [1] ), .QN(_08899_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_31_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [0] ), .QN(_08900_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_4_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [27] ), .QN(_08901_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_5_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [26] ), .QN(_08902_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_6_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [25] ), .QN(_08903_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_7_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [24] ), .QN(_08904_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_8_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [23] ), .QN(_08905_ ) );
DFF_X1 \mylsu.wdata_csreg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_csreg_$_DFFE_PP__Q_9_D ), .CK(_07943_ ), .Q(\LS_WB_wdata_csreg [22] ), .QN(_08906_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [31] ), .QN(_08907_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_1 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_1_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [30] ), .QN(_08908_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_10 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_10_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [21] ), .QN(_08909_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_11 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_11_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [20] ), .QN(_08910_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_12 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_12_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [19] ), .QN(_08911_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_13 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_13_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [18] ), .QN(_08912_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_14 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_14_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [17] ), .QN(_08913_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_15 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_15_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [16] ), .QN(_08914_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_16 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_16_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [15] ), .QN(_08915_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_17 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_17_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [14] ), .QN(_08916_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_18 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_18_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [13] ), .QN(_08917_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_19 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_19_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [12] ), .QN(_08918_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_2 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_2_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [29] ), .QN(_08919_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_20 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_20_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [11] ), .QN(_08920_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_21 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_21_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [10] ), .QN(_08921_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_22 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_22_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [9] ), .QN(_08922_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_23 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_23_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [8] ), .QN(_08923_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_24 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_24_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [7] ), .QN(_08924_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_25 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_25_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [6] ), .QN(_08925_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_26 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_26_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [5] ), .QN(_08926_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_27 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_27_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [4] ), .QN(_08927_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_28 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_28_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [3] ), .QN(_08928_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_29 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_29_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [2] ), .QN(_08929_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_3 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_3_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [28] ), .QN(_08930_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_30 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_30_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [1] ), .QN(_08931_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_31 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_31_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [0] ), .QN(_08932_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_4 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_4_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [27] ), .QN(_08933_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_5 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_5_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [26] ), .QN(_08934_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_6 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_6_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [25] ), .QN(_08935_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_7 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_7_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [24] ), .QN(_08936_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_8 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_8_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [23] ), .QN(_08937_ ) );
DFF_X1 \mylsu.wdata_reg_$_DFFE_PP__Q_9 ( .D(\mylsu.wdata_reg_$_DFFE_PP__Q_9_D ), .CK(_07939_ ), .Q(\LS_WB_wdata_reg [22] ), .QN(_07993_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q ( .D(_00218_ ), .CK(_07938_ ), .Q(\LS_WB_wen_csreg [7] ), .QN(_07992_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_1 ( .D(_00219_ ), .CK(_07938_ ), .Q(\LS_WB_wen_csreg [6] ), .QN(_07991_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_2 ( .D(_00220_ ), .CK(_07938_ ), .Q(\LS_WB_wen_csreg [3] ), .QN(_07990_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_3 ( .D(_00221_ ), .CK(_07938_ ), .Q(\LS_WB_wen_csreg [2] ), .QN(_07989_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_4 ( .D(_00222_ ), .CK(_07938_ ), .Q(\LS_WB_wen_csreg [1] ), .QN(_07988_ ) );
DFF_X1 \mylsu.wen_csreg_$_SDFFE_PP0P__Q_5 ( .D(_00223_ ), .CK(_07938_ ), .Q(\LS_WB_wen_csreg [0] ), .QN(_07987_ ) );
DFF_X1 \mylsu.wen_reg_$_SDFFE_PP0P__Q ( .D(_00224_ ), .CK(_07938_ ), .Q(LS_WB_wen_reg ), .QN(_08938_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q ( .D(\myminixbar.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\myminixbar.state [2] ), .QN(_08939_ ) );
DFF_X1 \myminixbar.state_$_DFF_P__Q_1 ( .D(\myminixbar.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\myminixbar.state [0] ), .QN(_08940_ ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[0]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07937_ ), .Q(\myreg.Reg[0][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[10]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07936_ ), .Q(\myreg.Reg[10][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[11]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07935_ ), .Q(\myreg.Reg[11][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[12]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07934_ ), .Q(\myreg.Reg[12][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[13]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07933_ ), .Q(\myreg.Reg[13][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[14]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07932_ ), .Q(\myreg.Reg[14][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[15]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07931_ ), .Q(\myreg.Reg[15][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[1]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07930_ ), .Q(\myreg.Reg[1][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[2]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07929_ ), .Q(\myreg.Reg[2][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[3]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07928_ ), .Q(\myreg.Reg[3][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[4]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07927_ ), .Q(\myreg.Reg[4][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[5]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07926_ ), .Q(\myreg.Reg[5][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[6]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07925_ ), .Q(\myreg.Reg[6][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[7]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07924_ ), .Q(\myreg.Reg[7][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[8]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07923_ ), .Q(\myreg.Reg[8][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][31] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_1 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_1_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][30] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_A_$_XOR__Y_B_$_XOR__Y_B_$_MUX__B_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_10 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_10_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][21] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_9_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_11 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_11_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][20] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_10_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_12 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_12_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][19] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_11_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_13 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_13_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][18] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_12_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_14 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_14_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][17] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_13_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_15 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_15_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][16] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_14_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_16 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_16_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][15] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_15_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_17 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_17_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][14] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_16_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_18 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_18_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][13] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_17_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_19 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_19_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][12] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_18_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_2 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_2_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][29] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_20 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_20_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][11] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_21 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_21_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][10] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_21_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_22 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_22_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][9] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_2_D_$_MUX__Y_A_$_NAND__Y_A_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_23 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_23_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][8] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_NAND__Y_A_$_XNOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_24 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_24_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][7] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_24_D_$_MUX__Y_B_$_MUX__Y_B_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_25 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_25_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][6] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_25_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_26 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_26_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][5] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_26_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_27 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_27_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][4] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_27_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_28 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_28_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][3] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_28_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_29 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_29_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][2] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_29_D_$_MUX__Y_B_$_MUX__Y_B_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_3 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_3_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][28] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_3_D_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_30 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_30_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][1] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_10_D_$_MUX__Y_A_$_ANDNOT__Y_B_$_XOR__Y_B_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_31 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_31_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][0] ), .QN(\myexu.dest_csreg_mem_$_DFFE_PP__Q_11_D_$_MUX__Y_A_$_OR__Y_A_$_XNOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_4 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_4_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][27] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_4_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_5 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_5_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][26] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_5_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_6 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_6_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][25] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_6_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_7 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_7_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][24] ), .QN(\myexu.result_csreg_mem_$_DFFE_PP__Q_7_D_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_A_$_NOT__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_8 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_8_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][23] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_7_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \myreg.Reg[9]_$_DFFE_PP__Q_9 ( .D(\myreg.Reg[9]_$_DFFE_PP__Q_9_D ), .CK(_07922_ ), .Q(\myreg.Reg[9][22] ), .QN(\myexu.src1_plus_imm_$_NOT__Y_8_A_$_XOR__Y_B_$_NOT__Y_A_$_XOR__Y_A_$_MUX__Y_A_$_MUX__Y_B_$_MUX__Y_A_$_MUX__Y_A_$_MUX__Y_B ) );
DFF_X1 \mysc.loaduse_clear_$_SDFFE_PP0P__Q ( .D(_00225_ ), .CK(_07921_ ), .Q(loaduse_clear ), .QN(_08941_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q ( .D(\mysc.state_$_DFF_P__Q_D ), .CK(clock ), .Q(\mysc.state [2] ), .QN(_08942_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_1 ( .D(\mysc.state_$_DFF_P__Q_1_D ), .CK(clock ), .Q(\mysc.state [1] ), .QN(_08943_ ) );
DFF_X1 \mysc.state_$_DFF_P__Q_2 ( .D(\mysc.state_$_DFF_P__Q_2_D ), .CK(clock ), .Q(\mysc.state [0] ), .QN(_07986_ ) );
BUF_X8 fanout_buf_1 ( .A(reset ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(reset ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(reset ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(reset ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(_00000_ ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(_00000_ ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\EX_LS_dest_csreg_mem [0] ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\ID_EX_typ [0] ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\ID_EX_typ [3] ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\ID_EX_typ [4] ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\IF_ID_pc [3] ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\IF_ID_pc [4] ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(io_master_wready_$_NOR__B_Y_$_OR__A_Y_$_ANDNOT__B_Y_$_ANDNOT__A_B_$_OR__Y_B ), .Z(fanout_net_20 ) );
BUF_X8 fanout_buf_21 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_21 ) );
BUF_X8 fanout_buf_22 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_22 ) );
BUF_X8 fanout_buf_23 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_23 ) );
BUF_X8 fanout_buf_24 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_24 ) );
BUF_X8 fanout_buf_25 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_25 ) );
BUF_X8 fanout_buf_26 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_26 ) );
BUF_X8 fanout_buf_27 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_27 ) );
BUF_X8 fanout_buf_28 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_28 ) );
BUF_X8 fanout_buf_29 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_29 ) );
BUF_X8 fanout_buf_30 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_30 ) );
BUF_X8 fanout_buf_31 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_31 ) );
BUF_X8 fanout_buf_32 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_32 ) );
BUF_X8 fanout_buf_33 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_33 ) );
BUF_X8 fanout_buf_34 ( .A(\myidu.rs1_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_34 ) );
BUF_X8 fanout_buf_35 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_35 ) );
BUF_X8 fanout_buf_36 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_36 ) );
BUF_X8 fanout_buf_37 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_37 ) );
BUF_X8 fanout_buf_38 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_38 ) );
BUF_X8 fanout_buf_39 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_39 ) );
BUF_X8 fanout_buf_40 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_40 ) );
BUF_X8 fanout_buf_41 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_41 ) );
BUF_X8 fanout_buf_42 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_42 ) );
BUF_X8 fanout_buf_43 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_43 ) );
BUF_X8 fanout_buf_44 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_44 ) );
BUF_X8 fanout_buf_45 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [1] ), .Z(fanout_net_45 ) );
BUF_X8 fanout_buf_46 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [2] ), .Z(fanout_net_46 ) );
BUF_X8 fanout_buf_47 ( .A(\myidu.rs2_$_SDFFE_PP0P__Q_4_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [3] ), .Z(fanout_net_47 ) );
BUF_X8 fanout_buf_48 ( .A(\myifu.pc_$_SDFFE_PP0P__Q_28_D_$_MUX__B_Y_$_SDFF_PP0__D_Q [0] ), .Z(fanout_net_48 ) );
BUF_X8 fanout_buf_49 ( .A(\myifu.to_reset ), .Z(fanout_net_49 ) );

endmodule
